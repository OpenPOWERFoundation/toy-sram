VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO 10T_toy_magic
  CLASS BLOCK ;
  FOREIGN 10T_toy_magic ;
  ORIGIN 0.500 0.095 ;
  SIZE 2.760 BY 1.350 ;
  PIN RWL
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.031500 ;
    PORT
      LAYER li1 ;
        RECT 1.895 0.415 2.045 0.585 ;
    END
  END RWL
  PIN RWL
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.031500 ;
    PORT
      LAYER li1 ;
        RECT -0.285 0.415 -0.135 0.585 ;
    END
  END RWL
  PIN WBL
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.024175 ;
    PORT
      LAYER li1 ;
        RECT 1.820 0.825 1.895 0.970 ;
    END
  END WBL
  PIN WBLb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.023100 ;
    PORT
      LAYER li1 ;
        RECT -0.130 0.825 -0.055 0.965 ;
    END
  END WBLb
  PIN RBL0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.045150 ;
    PORT
      LAYER li1 ;
        RECT 2.185 0.095 2.260 0.305 ;
    END
  END RBL0
  PIN RBL1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.045150 ;
    PORT
      LAYER li1 ;
        RECT -0.500 0.095 -0.425 0.305 ;
    END
  END RBL1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER nwell ;
        RECT 0.490 0.625 1.255 1.105 ;
      LAYER li1 ;
        RECT 0.800 1.035 0.960 1.105 ;
        RECT 0.810 1.025 0.950 1.035 ;
      LAYER met1 ;
        RECT -0.500 1.035 2.260 1.105 ;
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER pwell ;
        RECT -0.500 0.395 0.350 1.255 ;
        RECT 1.410 0.395 2.260 1.255 ;
        RECT -0.500 -0.095 2.260 0.395 ;
      LAYER li1 ;
        RECT 0.810 -0.025 0.950 -0.015 ;
        RECT 0.800 -0.095 0.960 -0.025 ;
      LAYER met1 ;
        RECT -0.500 -0.095 2.260 -0.025 ;
    END
  END GND
  OBS
      LAYER li1 ;
        RECT 0.275 0.825 0.350 0.965 ;
        RECT 0.490 0.775 0.565 0.915 ;
        RECT 1.195 0.835 1.255 0.915 ;
        POLYGON 1.195 0.835 1.255 0.835 1.255 0.775 ;
        RECT 1.410 0.825 1.485 0.965 ;
        RECT 0.220 0.305 0.370 0.475 ;
        RECT 0.610 0.440 0.760 0.610 ;
        RECT 1.000 0.440 1.150 0.610 ;
        RECT 1.390 0.305 1.540 0.475 ;
        RECT 0.485 0.220 0.535 0.255 ;
        POLYGON 0.535 0.255 0.570 0.220 0.535 0.220 ;
        RECT 0.485 0.095 0.570 0.220 ;
        RECT 1.190 0.095 1.275 0.255 ;
  END
END 10T_toy_magic
END LIBRARY

