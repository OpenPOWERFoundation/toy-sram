magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< obsli1 >>
rect 126 1532 1598 1598
rect 126 192 192 1532
rect 528 1130 1196 1196
rect 528 594 594 1130
rect 761 761 963 963
rect 1130 594 1196 1130
rect 528 528 1196 594
rect 1532 192 1598 1532
rect 126 126 1598 192
<< obsm1 >>
rect 130 1536 1594 1594
rect 130 188 188 1536
rect 532 1134 1192 1192
rect 532 590 590 1134
rect 761 761 963 963
rect 1134 590 1192 1134
rect 532 532 1192 590
rect 1536 188 1594 1536
rect 130 130 1594 188
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 1724 1724
string LEFview TRUE
string gencell sky130_fd_pr__rf_npn_05v5_W1p00L1p00
string library sky130
string parameter m=1
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 8602464
string GDS_START 8580692
<< end >>
