* NGSPICE file created from 10T_32x32_magic_flattened.ext - technology: sky130A

.subckt x10T_32x32_magic_flattened RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3
+ RBL0_3 RBL1_4 RBL0_4 RBL1_5 RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 RBL1_8 RBL0_8 RBL1_9
+ RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL0_11 RBL1_12 RBL0_12 RBL1_13 RBL0_13 RBL1_14 RBL0_14
+ RBL1_15 RBL0_15 WWL_0 RWL_0 WWL_1 RWL_1 WWL_2 RWL_2 WWL_3 RWL_3 WWL_4 RWL_4 WWL_5
+ RWL_5 WWL_6 RWL_6 WWL_7 RWL_7 WWL_8 RWL_8 WWL_9 RWL_9 WWL_10 RWL_10 WWL_11 RWL_11
+ WWL_12 RWL_12 WWL_13 RWL_13 WWL_14 RWL_14 WWL_15 RWL_15 WWL_16 RWL_16 WWL_17 RWL_17
+ WWL_18 RWL_18 WWL_19 RWL_19 WWL_20 RWL_20 WWL_21 RWL_21 WWL_22 RWL_22 WWL_23 RWL_23
+ WWL_24 RWL_24 WWL_25 RWL_25 WWL_26 RWL_26 WWL_27 RWL_27 WWL_28 RWL_28 WWL_29 RWL_29
+ WWL_30 RWL_30 WWL_31 RWL_31 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19
+ RBL0_19 RBL1_20 RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 RBL1_24
+ RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL0_27 RBL1_28 RBL0_28 RBL1_29
+ RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 WBL_0 WBLb_0 WBL_1 WBLb_1 WBL_2 WBLb_2 WBL_3
+ WBLb_19 WBL_4 WBLb_4 WBL_5 WBLb_5 WBL_22 WBLb_6 WBL_23 WBLb_7 WBL_24 WBLb_8 WBL_25
+ WBLb_9 WBL_26 WBLb_10 WBL_11 WBLb_11 WBL_12 WBLb_12 WBL_13 WBLb_13 WBL_14 WBLb_30
+ WBL_15 WBLb_31 VDD GND

M1000 GND a_12309_826# a_12253_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1001 a_2163_3818# a_1962_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1002 a_10569_2446# WWL_22 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1003 a_16313_4088# RWL_16 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1004 a_4483_4898# a_4282_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1005 a_12889_3526# WWL_18 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1006 a_4133_8138# RWL_1 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1007 RBL0_13 RWL_2 a_7963_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1008 WBL_14 WWL_12 a_8342_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1009 a_16083_6518# a_15882_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1010 WBL_5 WWL_20 a_3122_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1011 a_11242_1906# a_11149_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1012 a_7762_826# a_7669_826# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1013 a_18403_7598# a_18202_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1014 a_11242_5686# a_11149_5686# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1015 GND a_11242_7846# a_11149_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1016 a_4862_2986# a_4769_2986# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1017 GND a_9409_3526# a_9353_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1018 VDD a_2542_7846# a_2449_7846# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1019 GND a_10569_7846# a_10513_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1020 GND a_709_5416# a_653_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1021 GND a_4862_5146# a_4769_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1022 a_2973_7598# RWL_3 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1023 a_7383_309# a_7182_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1024 a_9703_578# a_9502_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1025 a_14923_5978# a_14722_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1026 a_423_2468# a_222_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1027 a_1382_286# a_1289_286# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1028 GND a_6602_1906# a_6509_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1029 a_802_3796# a_709_3796# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1030 VDD a_7182_6766# a_7089_6766# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1031 VDD a_6602_5686# a_6509_5686# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1032 a_5349_3256# WWL_19 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1033 RBL0_22 RWL_6 a_13183_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1034 GND a_5929_1906# a_5873_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1035 WBL_23 WWL_16 a_13562_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1036 RBL0_7 RWL_20 a_4483_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1037 GND a_18109_4066# a_18053_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1038 a_9502_8116# a_9409_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1039 RBL0_11 RWL_16 a_6803_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1040 a_423_308# a_222_286# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1041 GND a_15302_2446# a_15209_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1042 RBL0_15 RWL_24 a_9123_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1043 a_6022_2716# a_5929_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1044 RBL0_0 RWL_17 a_423_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1045 VDD a_15302_6226# a_15209_6226# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1046 a_1869_1636# WWL_25 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1047 a_6022_6496# a_5929_6496# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1048 GND a_14629_2446# a_14573_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1049 a_7613_3278# RWL_19 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1050 a_7383_5708# a_7182_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1052 a_653_1928# RWL_24 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1053 a_2163_3548# a_1962_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1054 a_15789_4336# WWL_15 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1055 VDD a_1962_826# a_1869_826# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1056 GND a_12309_556# a_12253_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1057 a_10569_2176# WWL_23 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1058 VDD a_11822_4606# a_11729_4606# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1059 a_9703_6788# a_9502_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1060 a_2449_826# WWL_28 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1061 RBL0_1 RWL_30 a_1003_308# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1062 a_13183_848# a_12982_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1063 a_1289_8386# WWL_0 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1064 RBL0_13 a_4683_7576# a_7963_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1065 WBL_14 WWL_13 a_8342_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1066 a_16083_6248# a_15882_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1067 a_10513_1118# RWL_27 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1068 a_16462_3796# a_16369_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1069 a_5442_287# a_5349_287# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1070 a_11242_1636# a_11149_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1071 a_16462_7576# a_16369_7576# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1072 a_11242_5416# a_11149_5416# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1073 WBL_31 WWL_29 a_18202_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1074 RBL0_11 RWL_31 a_6803_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1075 a_5873_8408# RWL_0 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1076 GND a_11242_7576# a_11149_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1077 a_1962_7846# a_1869_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1078 RBL0_7 RWL_9 a_4483_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1079 GND a_9409_3256# a_9353_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1080 GND a_10569_7576# a_10513_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1081 GND a_709_5146# a_653_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1082 a_12603_4628# a_12402_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1083 a_423_2198# a_222_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1084 GND a_6602_1636# a_6509_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1085 GND a_7182_2716# a_7089_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1086 a_15789_287# WWL_30 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1087 a_9502_1636# a_9409_1636# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1088 a_802_3526# a_709_3526# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1089 VDD a_7182_6496# a_7089_6496# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1090 VDD a_6602_5416# a_6509_5416# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1091 a_5349_2986# WWL_20 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1092 GND a_5929_1636# a_5873_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1093 WBL_27 WWL_25 a_15882_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1094 GND a_12309_1096# a_12253_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1095 GND a_15302_2176# a_15209_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1096 WBL_31 WWL_21 a_18202_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1097 a_9933_3008# RWL_20 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1098 RBL0_15 RWL_25 a_9123_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1099 a_6022_2446# a_5929_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1100 a_11822_7846# a_11729_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1101 a_1869_1366# WWL_26 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1102 RBL0_0 RWL_18 a_423_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1103 GND a_14629_2176# a_14573_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1104 WBL_10 WWL_6 a_6022_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1105 a_6022_6226# a_5929_6226# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1106 GND a_3029_7306# a_2973_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1107 a_11242_826# a_11149_826# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1108 a_7383_5438# a_7182_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1109 a_653_1658# RWL_25 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1110 a_15789_4066# WWL_16 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1111 a_10569_1906# WWL_24 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1112 a_2163_3278# a_1962_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1113 VDD a_11822_4336# a_11729_4336# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1114 a_7762_6766# a_7669_6766# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1115 a_2542_4606# a_2449_4606# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1116 a_3553_38# RWL_31 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1117 GND a_2542_6766# a_2449_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1118 a_13183_578# a_12982_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1119 a_1289_8116# WWL_1 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1120 VDD a_17622_826# a_17529_826# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1121 GND a_1869_6766# a_1813_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1122 a_16462_3526# a_16369_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1123 a_3903_3818# a_3702_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1124 GND a_14142_8386# a_14049_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1125 a_5442_17# a_5349_17# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1126 a_11242_1366# a_11149_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1127 a_16462_7306# a_16369_7306# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1128 WBL_19 WWL_10 a_11242_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1129 GND a_13469_8386# a_13413_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1130 RBL0_3 RWL_14 a_2163_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1131 a_5873_8138# RWL_1 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1132 RBL0_16 RWL_2 a_9703_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1133 a_1962_7576# a_1869_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1134 a_17823_6518# a_17622_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1135 a_12603_4358# a_12402_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1136 RBL0_27 RWL_4 a_16083_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1137 GND a_12982_7846# a_12889_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1138 a_9933_5978# RWL_9 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1139 GND a_7182_2446# a_7089_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1140 a_15789_17# WWL_31 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1141 GND a_6602_1366# a_6509_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1142 a_5293_4898# RWL_13 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1143 VDD a_7182_6226# a_7089_6226# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1144 WBL_1 WWL_17 a_802_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1145 GND a_5929_1366# a_5873_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1146 GND a_18202_2986# a_18109_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1147 WBL_27 WWL_26 a_15882_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1148 RBL0_21 RWL_10 a_12603_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1149 a_653_38# RWL_31 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1150 GND a_17529_2986# a_17473_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1151 a_3702_556# a_3609_556# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1152 RBL0_15 RWL_26 a_9123_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1153 a_11822_7576# a_11729_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1154 RBL0_25 RWL_6 a_14923_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1155 a_1869_1096# WWL_27 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1156 a_6022_2176# a_5929_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1157 RBL0_0 RWL_19 a_423_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1158 WBL_10 WWL_7 a_6022_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1159 GND a_3029_7036# a_2973_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1160 a_12833_3818# RWL_17 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1161 VDD a_14722_5146# a_14629_5146# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1162 RBL0_14 RWL_28 a_8543_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1163 VDD a_10082_4066# a_9989_4066# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1164 a_653_1388# RWL_26 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1165 a_7383_5168# a_7182_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1166 a_7762_2716# a_7669_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1167 a_7762_6496# a_7669_6496# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1168 a_2542_4336# a_2449_4336# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1169 a_18109_1636# WWL_25 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1170 VDD a_15302_287# a_15209_287# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1171 a_14142_5956# a_14049_5956# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1172 a_16462_3256# a_16369_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1173 a_3903_3548# a_3702_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1174 GND a_14142_8116# a_14049_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1175 a_16462_7036# a_16369_7036# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1176 a_8249_6766# WWL_6 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1177 WBL_28 WWL_3 a_16462_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1178 RBL0_12 RWL_7 a_7383_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1179 a_3029_4606# WWL_14 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1180 GND a_13469_8116# a_13413_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1181 WBL_19 WWL_11 a_11242_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1182 RBL0_3 RWL_15 a_2163_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1183 RBL0_16 a_4683_7576# a_9703_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1184 a_6602_287# a_6509_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1185 a_10283_3008# a_10082_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1186 a_17823_6248# a_17622_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1187 GND a_18202_5956# a_18109_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1188 a_12603_4088# a_12402_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1189 GND a_10662_6496# a_10569_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1190 a_8193_5708# RWL_10 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1191 VDD a_802_7846# a_709_7846# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1192 RBL0_27 RWL_5 a_16083_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1193 VDD a_9502_5956# a_9409_5956# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1194 GND a_17529_5956# a_17473_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1195 GND a_4189_1096# a_4133_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1196 GND a_7182_2176# a_7089_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1197 GND a_12982_7576# a_12889_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1198 a_3702_7846# a_3609_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1199 WBL_1 WWL_18 a_802_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1200 a_8193_309# RWL_30 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1201 a_13469_5686# WWL_10 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1202 a_8922_2986# a_8829_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1203 VDD a_222_4606# a_129_4606# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1204 a_14722_8386# a_14629_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1205 a_10082_7306# a_9989_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1206 WBL_27 WWL_27 a_15882_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1207 VDD a_1382_3256# a_1289_3256# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1208 RBL0_21 RWL_11 a_12603_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1209 a_3702_286# a_3609_286# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1210 WBL_10 WWL_8 a_6022_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1211 a_1233_38# RWL_31 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1212 GND a_14722_1096# a_14629_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1213 a_13413_4628# RWL_14 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1214 RBL0_10 RWL_30 a_6223_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1215 a_12833_3548# RWL_18 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1216 RBL0_14 RWL_29 a_8543_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1217 VDD a_14722_4876# a_14629_4876# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1218 a_5442_5146# a_5349_5146# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1219 a_8922_826# a_8829_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1220 a_7762_2446# a_7669_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1221 GND a_5442_7306# a_5349_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1222 WBL_13 WWL_6 a_7762_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1223 a_7762_6226# a_7669_6226# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1224 a_12402_826# a_12309_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1225 WBL_4 WWL_14 a_2542_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1226 GND a_4769_7306# a_4713_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1227 a_18109_1366# WWL_26 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1228 a_10283_5978# a_10082_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1229 VDD a_14142_1636# a_14049_1636# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1230 RBL0_29 RWL_27 a_17243_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1231 VDD a_15302_17# a_15209_17# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1232 a_709_826# WWL_28 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1233 a_3903_3278# a_3702_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1234 GND a_1962_5686# a_1869_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1235 a_8249_6496# WWL_7 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1236 WBL_28 WWL_4 a_16462_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1237 RBL0_12 RWL_8 a_7383_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1238 RBL0_3 RWL_16 a_2163_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1239 a_10662_4066# a_10569_4066# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1240 GND a_15882_8386# a_15789_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1241 GND a_15209_4606# a_15153_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1242 a_8193_5438# RWL_11 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1243 a_222_7846# a_129_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1244 GND a_10662_6226# a_10569_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1245 a_8922_5956# a_8829_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1246 a_1382_6496# a_1289_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1247 RBL0_6 RWL_14 a_3903_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1248 a_3702_7576# a_3609_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1249 RBL0_20 RWL_28 a_12023_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1250 VDD a_12402_6766# a_12309_6766# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1251 a_11149_4336# WWL_15 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1252 VDD a_13562_556# a_13469_556# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1253 GND a_9989_287# a_9933_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1254 a_4713_3818# RWL_17 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1255 a_5063_6788# a_4862_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1256 a_14049_556# WWL_29 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1257 a_14722_8116# a_14629_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1258 RBL0_30 RWL_4 a_17823_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1259 a_13469_5416# WWL_11 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1260 VDD a_222_4336# a_129_4336# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1261 a_10082_7036# a_9989_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1262 RBL0_21 RWL_12 a_12603_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1263 VDD a_1382_2986# a_1289_2986# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1264 WBL_15 WWL_5 a_8922_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1265 GND a_3122_826# a_3029_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1266 a_3702_16# a_3609_16# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1268 a_13413_4358# RWL_15 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1269 a_709_2446# WWL_22 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1270 a_12833_3278# RWL_19 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1271 a_14142_4876# a_14049_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1272 a_5442_1096# a_5349_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1273 a_1233_8408# RWL_0 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1274 a_5442_4876# a_5349_4876# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1275 a_8922_556# a_8829_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1276 a_13413_39# RWL_31 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1277 a_7762_2176# a_7669_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1278 GND a_5442_7036# a_5349_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1279 a_10082_287# a_9989_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1280 VDD a_17042_2446# a_16949_2446# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1281 a_12402_556# a_12309_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1282 WBL_13 WWL_7 a_7762_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1283 a_15503_7868# a_15302_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1284 GND a_4769_7036# a_4713_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1285 a_18109_1096# WWL_27 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1286 GND a_802_6766# a_709_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1287 WBL_24 WWL_9 a_14142_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1288 GND a_6509_3796# a_6453_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1289 GND a_9502_4876# a_9409_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1290 GND a_1962_5416# a_1869_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1291 a_8249_6226# WWL_8 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1292 GND a_16462_287# a_16369_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1293 GND a_8829_4876# a_8773_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1294 GND a_15789_826# a_15733_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1295 a_15882_5956# a_15789_5956# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1296 GND a_15209_4336# a_15153_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1297 WBL_18 WWL_15 a_10662_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1298 GND a_15882_8116# a_15789_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1299 a_9989_6766# WWL_6 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1300 a_8193_5168# RWL_12 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1301 a_6602_8386# a_6509_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1302 a_222_7576# a_129_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1303 a_4769_4606# WWL_14 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1304 a_1382_6226# a_1289_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1305 RBL0_6 RWL_15 a_3903_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1306 a_12023_3008# a_11822_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1307 GND a_12402_2716# a_12309_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1308 RBL0_20 RWL_29 a_12023_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1309 a_14722_1636# a_14629_1636# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1310 a_15302_2716# a_15209_2716# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1311 VDD a_12402_6496# a_12309_6496# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1312 a_11149_4066# WWL_16 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1313 GND a_11729_2716# a_11673_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1314 a_3122_6766# a_3029_6766# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1315 a_4713_3548# RWL_18 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1316 RBL0_30 RWL_5 a_17823_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1317 GND a_3122_556# a_3029_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1318 VDD a_222_826# a_129_826# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1319 a_17042_5686# a_16949_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1320 a_11093_3008# RWL_20 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1321 a_709_2176# WWL_23 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1322 a_13413_4088# RWL_16 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1323 a_1583_4898# a_1382_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1324 a_15733_309# RWL_30 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1325 a_1233_8138# RWL_1 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1326 RBL0_8 RWL_2 a_5063_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1327 WBL_9 WWL_12 a_5442_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1328 a_13183_6518# a_12982_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1329 VDD a_17042_2176# a_16949_2176# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1330 WBL_13 WWL_8 a_7762_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1331 a_15503_7598# a_15302_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1332 RBL0_23 RWL_30 a_13763_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1333 GND a_7089_4606# a_7033_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1334 GND a_6509_3526# a_6453_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1335 GND a_1962_5146# a_1869_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1336 a_12023_5978# a_11822_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1337 GND a_13469_287# a_13413_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1338 VDD a_15882_1636# a_15789_1636# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1339 GND a_15789_556# a_15733_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1340 GND a_3702_1906# a_3609_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1341 VDD a_4282_6766# a_4189_6766# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1342 VDD a_3702_5686# a_3609_5686# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1343 a_2449_3256# WWL_19 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1344 RBL0_17 RWL_6 a_10283_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1345 GND a_15209_4066# a_15153_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1346 WBL_18 WWL_16 a_10662_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1347 a_9989_6496# WWL_7 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1348 a_17243_1118# a_17042_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1349 RBL0_2 RWL_20 a_1583_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1350 a_6602_8116# a_6509_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1351 a_17622_2446# a_17529_2446# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1352 a_12982_1366# a_12889_1366# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1353 RBL0_6 RWL_16 a_3903_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1354 GND a_17622_4606# a_17529_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1355 GND a_12402_2446# a_12309_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1356 a_11093_5978# RWL_9 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1357 VDD a_17622_8386# a_17529_8386# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1358 a_16369_5956# WWL_9 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1359 RBL0_10 RWL_24 a_6223_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1360 a_3122_2716# a_3029_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1361 GND a_16949_4606# a_16893_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1362 VDD a_12402_6226# a_12309_6226# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1363 a_3122_6496# a_3029_6496# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1364 GND a_11729_2446# a_11673_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1365 a_4713_3278# RWL_19 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1366 a_11093_39# RWL_31 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1367 a_4483_5708# a_4282_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1368 a_17042_5416# a_16949_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1369 VDD a_8342_1366# a_8249_1366# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1370 a_12889_4336# WWL_15 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1371 a_6803_6788# a_6602_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1372 WBL_20 WWL_3 a_11822_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1373 a_709_1906# WWL_24 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1374 WBL_30 WWL_28 a_17622_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1375 a_18403_8408# a_18202_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1376 RBL0_8 a_4683_7576# a_5063_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1377 WBL_9 WWL_13 a_5442_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1378 a_13183_6248# a_12982_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1379 a_13562_3796# a_13469_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1380 VDD a_17042_1906# a_16949_1906# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1381 a_13562_7576# a_13469_7576# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1382 a_15882_4876# a_15789_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1383 a_2973_8408# RWL_0 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1384 RBL0_2 RWL_9 a_1583_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1385 GND a_6509_3256# a_6453_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1386 GND a_7089_4336# a_7033_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1387 GND a_8922_3796# a_8829_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1388 GND a_3702_1636# a_3609_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1389 GND a_4282_2716# a_4189_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1390 VDD a_8922_7576# a_8829_7576# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1391 a_7669_5146# WWL_12 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1392 a_6602_1636# a_6509_1636# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1393 VDD a_4282_6496# a_4189_6496# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1394 VDD a_3702_5416# a_3609_5416# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1395 a_2449_2986# WWL_20 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1396 a_9989_6226# WWL_8 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1397 a_17622_2176# a_17529_2176# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1398 a_18202_3256# a_18109_3256# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1399 a_12982_1096# a_12889_1096# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1400 WBL_22 WWL_25 a_12982_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1401 a_16313_7868# RWL_2 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1402 a_15733_6788# RWL_6 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1403 GND a_17622_4336# a_17529_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1404 GND a_12402_2176# a_12309_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1405 WBL_26 WWL_21 a_15302_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1406 a_8342_4606# a_8249_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1407 VDD a_17622_8116# a_17529_8116# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1408 RBL0_10 RWL_25 a_6223_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1409 a_3122_2446# a_3029_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1410 a_8342_8386# a_8249_8386# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1411 GND a_16949_4336# a_16893_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1412 GND a_11729_2176# a_11673_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1413 WBL_5 WWL_6 a_3122_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1414 a_3122_6226# a_3029_6226# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1415 a_4483_5438# a_4282_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1416 VDD a_8342_1096# a_8249_1096# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1417 a_12889_4066# WWL_16 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1418 a_17042_5146# a_16949_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1419 a_4862_6766# a_4769_6766# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1420 RBL0_13 RWL_0 a_7963_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1421 WBL_20 WWL_4 a_11822_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1422 VDD a_5442_826# a_5349_826# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1423 a_18403_8138# a_18202_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1424 a_13562_3526# a_13469_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1425 GND a_11242_8386# a_11149_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1426 a_13562_7306# a_13469_7306# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1427 GND a_18109_7846# a_18053_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1428 GND a_10569_8386# a_10513_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1429 a_2973_8138# RWL_1 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1430 RBL0_11 RWL_2 a_6803_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1431 a_9123_1118# a_8922_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1432 a_8922_287# a_8829_287# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1433 GND a_7089_4066# a_7033_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1434 a_14923_6518# a_14722_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1435 a_12402_287# a_12309_287# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1436 a_423_3008# a_222_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1437 a_9502_2446# a_9409_2446# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1438 a_14049_7576# WWL_3 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1439 RBL0_22 RWL_4 a_13183_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1440 GND a_129_2716# a_73_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1441 GND a_8922_3526# a_8829_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1442 GND a_4282_2446# a_4189_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1443 GND a_3702_1366# a_3609_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1444 a_2393_4898# RWL_13 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1445 VDD a_8922_7306# a_8829_7306# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1446 VDD a_4282_6226# a_4189_6226# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1447 a_7669_4876# WWL_13 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1448 GND a_15302_2986# a_15209_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1449 a_18202_2986# a_18109_2986# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1450 WBL_22 WWL_26 a_12982_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1451 a_17622_1906# a_17529_1906# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1452 WBL_30 WWL_22 a_17622_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1453 a_16313_7598# a_13963_7576# RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1454 a_653_848# RWL_28 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1455 GND a_14629_2986# a_14573_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1456 GND a_17622_4066# a_17529_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1457 a_8342_4336# a_8249_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1458 RBL0_10 RWL_26 a_6223_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1459 a_3122_2176# a_3029_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1460 GND a_16949_4066# a_16893_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1461 a_8342_8116# a_8249_8116# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1462 WBL_5 WWL_7 a_3122_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1463 VDD a_11822_5146# a_11729_5146# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1464 a_9703_7328# a_9502_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1465 a_4862_2716# a_4769_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1466 a_4483_5168# a_4282_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1467 a_4862_6496# a_4769_6496# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1468 RBL0_13 RWL_1 a_7963_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1469 a_18053_1118# RWL_27 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1470 a_15209_1636# WWL_25 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1471 a_423_5978# a_222_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1472 a_11242_5956# a_11149_5956# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1473 a_13562_3256# a_13469_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1474 GND a_11242_8116# a_11149_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1475 WBL_23 WWL_3 a_13562_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1476 a_13562_7036# a_13469_7036# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1477 a_5349_6766# WWL_6 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1478 a_1962_8386# a_1869_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1479 GND a_18109_7576# a_18053_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1480 RBL0_7 RWL_7 a_4483_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1481 GND a_10569_8116# a_10513_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1482 RBL0_11 a_4683_7576# a_6803_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1483 a_8922_17# a_8829_17# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1484 a_14923_6248# a_14722_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1485 GND a_15302_5956# a_15209_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1486 a_12402_17# a_12309_17# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1487 a_5293_5708# RWL_10 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1488 a_9502_2176# a_9409_2176# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1489 a_802_4066# a_709_4066# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1490 a_14049_7306# WWL_4 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1491 RBL0_22 RWL_5 a_13183_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1492 VDD a_6602_5956# a_6509_5956# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1493 GND a_14629_5956# a_14573_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1494 GND a_129_2446# a_73_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1495 a_7613_6788# RWL_6 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1496 GND a_1289_1096# a_1233_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1497 GND a_4282_2176# a_4189_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1498 GND a_8922_3256# a_8829_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1499 VDD a_8922_7036# a_8829_7036# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1500 WBL_23 WWL_29 a_13562_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1501 WBL_31 WWL_19 a_18202_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1502 a_10569_5686# WWL_10 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1503 WBL_30 WWL_23 a_17622_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1504 VDD a_6022_2716# a_5929_2716# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1505 a_6022_2986# a_5929_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1506 a_11822_8386# a_11729_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1507 WBL_22 WWL_27 a_12982_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1508 a_653_578# RWL_29 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1509 a_8342_4066# a_8249_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1510 WBL_14 WWL_0 a_8342_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1511 RBL0_29 RWL_31 a_17243_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1512 WBL_5 WWL_8 a_3122_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1513 GND a_11822_1096# a_11729_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1514 a_10513_4628# RWL_14 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1515 a_7182_556# a_7089_556# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1516 VDD a_11822_4876# a_11729_4876# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1517 a_9703_7058# a_9502_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1518 a_2542_5146# a_2449_5146# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1519 a_4862_2446# a_4769_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1520 GND a_2542_7306# a_2449_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1521 a_4862_6226# a_4769_6226# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1522 GND a_9409_6766# a_9353_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1523 GND a_1869_7306# a_1813_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1524 a_15209_1366# WWL_26 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1525 VDD a_16462_3796# a_16369_3796# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1526 RBL0_24 RWL_27 a_14343_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1527 VDD a_11242_1636# a_11149_1636# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1528 a_16462_7846# a_16369_7846# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1529 RBL0_16 RWL_0 a_9703_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1530 a_5349_6496# WWL_7 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1531 a_1962_8116# a_1869_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1532 WBL_23 WWL_4 a_13562_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1533 RBL0_7 RWL_8 a_4483_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1534 GND a_12982_8386# a_12889_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1535 a_9933_6518# RWL_7 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1536 GND a_7182_2986# a_7089_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1537 GND a_12309_4606# a_12253_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1538 a_5293_5438# RWL_11 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1539 a_9502_1906# a_9409_1906# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1540 WBL_16 WWL_22 a_9502_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1541 a_6022_5956# a_5929_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1542 WBL_1 WWL_15 a_802_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1543 GND a_129_2176# a_73_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1544 a_16663_2738# a_16462_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1545 VDD a_1382_556# a_1289_556# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1546 a_15789_7576# WWL_3 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1547 a_1813_3818# RWL_17 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1548 a_2163_6788# a_1962_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1549 a_10569_5416# WWL_11 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1550 WBL_30 WWL_24 a_17622_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1551 WBL_31 WWL_20 a_18202_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1552 a_11822_8116# a_11729_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1553 RBL0_25 RWL_4 a_14923_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1554 WBL_0 WWL_28 a_222_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1555 WBL_10 WWL_5 a_6022_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1556 WBL_14 WWL_1 a_8342_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1557 a_10513_4358# RWL_15 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1558 a_11242_4876# a_11149_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1559 a_2542_1096# a_2449_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1560 a_5873_848# RWL_28 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1561 a_2542_4876# a_2449_4876# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1562 a_4862_2176# a_4769_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1563 GND a_2542_7036# a_2449_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1564 VDD a_14142_2446# a_14049_2446# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1565 a_12603_7868# a_12402_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1566 GND a_1869_7036# a_1813_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1567 a_15209_1096# WWL_27 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1568 VDD a_16462_3526# a_16369_3526# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1569 a_7182_3796# a_7089_3796# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1570 a_1962_1636# a_1869_1636# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1571 GND a_7182_5956# a_7089_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1572 a_3029_5146# WWL_12 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1573 RBL0_6 RWL_28 a_3903_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1574 WBL_19 WWL_9 a_11242_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1575 GND a_3609_3796# a_3553_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1576 GND a_6602_4876# a_6509_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1577 RBL0_16 RWL_1 a_9703_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1578 a_5349_6226# WWL_8 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1579 a_7963_1928# a_7762_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1580 GND a_5929_4876# a_5873_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1581 a_5929_556# WWL_29 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1582 GND a_18202_6496# a_18109_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1583 GND a_17529_6496# a_17473_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1584 a_9933_6248# RWL_8 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1585 GND a_12309_4336# a_12253_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1586 GND a_12982_8116# a_12889_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1587 a_5293_5168# RWL_12 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1588 WBL_16 WWL_23 a_9502_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1589 RBL0_15 RWL_13 a_9123_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1590 a_3702_8386# a_3609_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1591 RBL0_0 RWL_6 a_423_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1592 WBL_1 WWL_16 a_802_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1593 a_1869_4606# WWL_14 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1594 a_16663_2468# a_16462_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1595 a_7033_1928# RWL_24 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1596 GND a_10082_3796# a_9989_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1597 VDD a_222_5146# a_129_5146# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1598 a_11822_1636# a_11729_1636# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1599 a_12402_2716# a_12309_2716# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1600 VDD a_10082_7576# a_9989_7576# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1601 VDD a_1382_286# a_1289_286# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1602 a_653_4898# RWL_13 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1603 a_15789_7306# WWL_4 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1604 a_1813_3548# RWL_18 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1605 RBL0_25 RWL_5 a_14923_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1606 VDD a_17042_556# a_16949_556# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1607 a_14142_5686# a_14049_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1608 RBL0_28 RWL_17 a_16663_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1609 RBL0_20 RWL_21 a_12023_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1610 a_16462_6766# a_16369_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1611 VDD a_7762_2716# a_7669_2716# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1612 a_7762_2986# a_7669_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1613 a_10513_4088# RWL_16 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1614 GND a_10082_826# a_9989_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1615 a_5873_578# RWL_29 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1616 RBL0_3 RWL_2 a_2163_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1617 WBL_4 WWL_12 a_2542_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1618 a_10283_6518# a_10082_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1619 VDD a_14142_2176# a_14049_2176# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1620 a_12603_7598# a_12402_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1621 GND a_9502_5686# a_9409_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1622 a_7182_3526# a_7089_3526# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1623 a_8249_7036# WWL_5 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1624 a_14722_556# a_14629_556# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1625 WBL_28 WWL_2 a_16462_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1626 GND a_8829_5686# a_8773_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1627 GND a_4189_4606# a_4133_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1628 a_3029_4876# WWL_13 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1629 RBL0_6 RWL_29 a_3903_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1630 GND a_3609_3526# a_3553_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1631 a_7963_1658# a_7762_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1632 GND a_18202_6226# a_18109_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1633 VDD a_12982_1636# a_12889_1636# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1634 a_222_8386# a_129_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1635 a_8922_6496# a_8829_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1636 WBL_27 WWL_14 a_15882_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1637 VDD a_1382_6766# a_1289_6766# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1638 GND a_17529_6226# a_17473_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1639 GND a_12309_4066# a_12253_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1640 a_14343_1118# a_14142_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1641 a_3702_8116# a_3609_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1642 WBL_16 WWL_24 a_9502_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1643 a_14722_2446# a_14629_2446# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1644 a_10082_1366# a_9989_1366# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1645 a_16663_2198# a_16462_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1646 GND a_222_1096# a_129_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1647 GND a_14722_4606# a_14629_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1648 a_7033_1658# RWL_25 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1649 GND a_10082_3526# a_9989_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1650 VDD a_14722_8386# a_14629_8386# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1651 a_5063_7328# a_4862_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1652 a_13469_5956# WWL_9 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1653 VDD a_10082_7306# a_9989_7306# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1654 RBL0_5 RWL_24 a_3323_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1655 VDD a_222_4876# a_129_4876# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1656 a_7762_5956# a_7669_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1657 VDD a_1382_16# a_1289_16# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1658 a_1813_3278# RWL_19 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1659 a_17622_287# a_17529_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1660 a_17529_3796# WWL_17 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1661 a_1583_5708# a_1382_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1662 a_14142_5416# a_14049_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1663 VDD a_5442_1366# a_5349_1366# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1664 RBL0_28 RWL_18 a_16663_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1665 RBL0_29 RWL_14 a_17243_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1666 RBL0_20 RWL_22 a_12023_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1667 a_16462_17# a_16369_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1668 a_3903_6788# a_3702_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1669 WBL_9 WWL_28 a_5442_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1670 GND a_10082_556# a_9989_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1671 WBL_13 WWL_5 a_7762_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1672 a_17473_2738# RWL_21 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1673 a_15503_8408# a_15302_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1674 RBL0_3 RWL_3 a_2163_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1675 WBL_4 WWL_13 a_2542_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1676 a_10283_6248# a_10082_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1677 a_10662_3796# a_10569_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1678 VDD a_14142_1906# a_14049_1906# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1680 a_10662_7576# a_10569_7576# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1681 GND a_802_7306# a_709_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1682 GND a_9502_5416# a_9409_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1683 WBL_12 WWL_17 a_7182_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1684 GND a_8829_5416# a_8773_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1685 a_9353_39# RWL_31 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1686 GND a_3609_3256# a_3553_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1687 GND a_4189_4336# a_4133_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1688 a_17823_39# a_17622_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1689 VDD a_15882_2446# a_15789_2446# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1690 a_7963_1388# a_7762_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1691 GND a_1382_2716# a_1289_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1692 a_222_8116# a_129_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1693 a_8922_6226# a_8829_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1694 a_4769_5146# WWL_12 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1695 a_3702_1636# a_3609_1636# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1696 VDD a_1382_6496# a_1289_6496# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1697 a_14722_2176# a_14629_2176# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1698 a_15302_3256# a_15209_3256# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1699 GND a_11822_287# a_11729_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1700 a_10082_1096# a_9989_1096# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1701 WBL_17 WWL_25 a_10082_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1702 a_9409_826# WWL_28 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1703 GND a_14722_4336# a_14629_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1704 a_13413_7868# RWL_2 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1705 a_12833_6788# RWL_6 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1706 a_7033_1388# RWL_26 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1707 GND a_10082_3256# a_9989_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1708 a_5063_7058# a_4862_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1709 WBL_21 WWL_21 a_12402_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1710 RBL0_14 RWL_17 a_8543_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1711 a_5442_4606# a_5349_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1712 VDD a_14722_8116# a_14629_8116# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1713 VDD a_10082_7036# a_9989_7036# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1714 RBL0_5 RWL_25 a_3323_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1715 a_5442_8386# a_5349_8386# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1716 a_8773_1928# RWL_24 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1717 a_17529_3526# WWL_18 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1718 a_18109_4606# WWL_14 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1719 a_1583_5438# a_1382_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1720 a_14142_5146# a_14049_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1721 VDD a_5442_1096# a_5349_1096# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1722 RBL0_29 RWL_15 a_17243_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1723 RBL0_20 RWL_23 a_12023_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1724 RBL0_28 RWL_19 a_16663_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1725 RBL0_8 RWL_0 a_5063_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1726 a_17473_2468# RWL_22 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1727 a_15503_8138# a_15302_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1728 a_15882_5686# a_15789_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1729 a_10662_3526# a_10569_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1730 GND a_15209_7846# a_15153_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1731 a_10662_7306# a_10569_7306# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1732 WBL_8 WWL_22 a_4862_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1733 GND a_9502_5146# a_9409_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1734 GND a_802_7036# a_709_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1735 WBL_12 WWL_18 a_7182_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1736 RBL0_6 RWL_2 a_3903_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1737 GND a_8829_5146# a_8773_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1738 a_6223_1118# a_6022_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1739 GND a_4189_4066# a_4133_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1740 a_12023_6518# a_11822_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1741 VDD a_15882_2176# a_15789_2176# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1742 a_6602_2446# a_6509_2446# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1743 a_222_1636# a_129_1636# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1744 a_73_3818# RWL_17 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1745 a_11149_7576# WWL_3 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1746 RBL0_17 RWL_4 a_10283_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1747 a_9989_7036# WWL_5 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1748 GND a_1382_2446# a_1289_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1749 VDD a_1382_6226# a_1289_6226# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1750 a_18202_826# a_18109_826# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1751 a_4769_4876# WWL_13 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1752 a_1813_308# RWL_30 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1753 GND a_12402_2986# a_12309_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1754 a_11093_6518# RWL_7 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1755 a_7089_287# WWL_30 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1756 a_14722_1906# a_14629_1906# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1757 a_15302_2986# a_15209_2986# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1758 WBL_17 WWL_26 a_10082_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1759 WBL_25 WWL_22 a_14722_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1760 a_13413_7598# a_4683_7576# RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1761 a_709_5686# WWL_10 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1762 a_8829_2716# WWL_21 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1763 GND a_11729_2986# a_11673_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1764 a_9409_3796# WWL_17 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1765 GND a_14722_4066# a_14629_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1767 RBL0_14 RWL_18 a_8543_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1768 a_5442_4336# a_5349_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1769 a_14142_17# a_14049_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1770 RBL0_5 RWL_26 a_3323_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1771 a_5442_8116# a_5349_8116# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1772 GND a_17042_1906# a_16949_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1773 VDD a_17042_5686# a_16949_5686# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1774 a_8543_848# a_8342_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1775 GND a_16369_1906# a_16313_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1776 a_12023_848# a_11822_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1777 a_8773_1658# RWL_25 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1778 a_6803_7328# a_6602_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1779 a_1583_5168# a_1382_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1780 RBL0_29 RWL_16 a_17243_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1781 RBL0_8 RWL_1 a_5063_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1782 a_15153_1118# RWL_27 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1783 a_12309_1636# WWL_25 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1784 a_7033_39# RWL_31 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1785 a_17473_2198# RWL_23 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1786 a_15882_5416# a_15789_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1787 a_15503_39# a_15302_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1788 a_10662_3256# a_10569_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1789 a_2449_6766# WWL_6 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1790 WBL_18 WWL_3 a_10662_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1791 a_10662_7036# a_10569_7036# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1792 WBL_8 WWL_23 a_4862_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1793 GND a_15209_7576# a_15153_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1794 RBL0_2 RWL_7 a_1583_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1795 a_17243_4628# a_17042_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1796 RBL0_6 RWL_3 a_3903_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1797 a_12023_6248# a_11822_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1798 VDD a_15882_1906# a_15789_1906# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1799 GND a_12402_5956# a_12309_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1800 a_2393_5708# RWL_10 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1801 a_6602_2176# a_6509_2176# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1802 a_73_3548# RWL_18 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1803 a_11149_7306# WWL_4 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1804 VDD a_3702_5956# a_3609_5956# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1805 RBL0_17 RWL_5 a_10283_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1806 GND a_11729_5956# a_11673_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1807 a_4713_6788# RWL_6 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1808 GND a_1382_2176# a_1289_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1809 WBL_2 WWL_29 a_1382_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1810 a_16313_8408# RWL_0 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1811 a_15733_7328# RWL_4 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1812 a_7089_2446# WWL_22 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1813 a_11093_6248# RWL_8 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1814 WBL_26 WWL_19 a_15302_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1815 a_7089_17# WWL_31 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1816 WBL_17 WWL_27 a_10082_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1817 WBL_25 WWL_23 a_14722_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1818 VDD a_3122_2716# a_3029_2716# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1819 a_3122_2986# a_3029_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1820 a_709_5416# WWL_11 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1821 a_9409_3526# WWL_18 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1822 RBL0_14 RWL_19 a_8543_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1823 a_5442_4066# a_5349_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1824 WBL_9 WWL_0 a_5442_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1825 GND a_17042_1636# a_16949_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1826 VDD a_17042_5416# a_16949_5416# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1827 a_8543_578# a_8342_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1828 GND a_16369_1636# a_16313_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1829 a_12023_578# a_11822_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1830 a_8773_1388# RWL_26 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1831 a_6803_7058# a_6602_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1832 WBL_20 WWL_2 a_11822_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1833 a_16949_826# WWL_28 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1834 GND a_7089_7846# a_7033_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1835 GND a_6509_6766# a_6453_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1836 a_16949_2446# WWL_22 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1837 a_8543_3818# a_8342_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1838 a_12309_1366# WWL_26 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1839 VDD a_13562_3796# a_13469_3796# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1840 RBL0_19 RWL_27 a_11443_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1841 GND a_18109_8386# a_18053_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1842 a_13562_7846# a_13469_7846# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1843 a_15882_5146# a_15789_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1844 RBL0_11 RWL_0 a_6803_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1845 a_2449_6496# WWL_7 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1846 WBL_8 WWL_24 a_4862_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1847 WBL_18 WWL_4 a_10662_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1848 RBL0_2 RWL_8 a_1583_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1849 a_17622_1906# a_17529_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1850 a_17243_4358# a_17042_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1851 VDD a_10082_287# a_9989_287# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1852 a_18202_6766# a_18109_6766# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1853 a_17622_5686# a_17529_5686# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1854 GND a_17622_17# a_17529_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1855 a_12982_4606# a_12889_4606# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1856 GND a_17622_7846# a_17529_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1857 GND a_4282_2986# a_4189_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1858 a_3122_5956# a_3029_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1859 a_2393_5438# RWL_11 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1860 a_6602_1906# a_6509_1906# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1861 WBL_11 WWL_22 a_6602_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1862 a_73_3278# RWL_19 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1863 VDD a_8922_7846# a_8829_7846# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1864 GND a_16949_7846# a_16893_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1865 a_13763_2738# a_13562_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1866 WBL_2 WWL_30 a_1382_286# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1867 a_16313_8138# RWL_1 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1868 a_12889_7576# WWL_3 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1869 a_15733_7058# RWL_5 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1870 a_7089_2176# WWL_23 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1871 VDD a_8342_4606# a_8249_4606# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1872 WBL_25 WWL_24 a_14722_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1873 WBL_26 WWL_20 a_15302_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1874 WBL_29 WWL_29 a_17042_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1875 WBL_5 WWL_5 a_3122_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1876 WBL_9 WWL_1 a_5442_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1877 GND a_17042_1366# a_16949_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1878 GND a_16369_1366# a_16313_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1879 a_14629_287# WWL_30 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1880 a_13183_39# a_12982_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1881 VDD a_11242_2446# a_11149_2446# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1882 GND a_7089_7576# a_7033_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1883 a_9123_4628# a_8922_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1884 a_423_6518# a_222_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1885 a_8543_3548# a_8342_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1886 a_12309_1096# WWL_27 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1887 a_16949_2176# WWL_23 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1888 VDD a_13562_3526# a_13469_3526# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1889 a_4282_3796# a_4189_3796# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1890 GND a_18109_8116# a_18053_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1891 GND a_4282_5956# a_4189_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1892 GND a_3702_4876# a_3609_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1893 a_7669_8386# WWL_0 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1894 RBL0_11 RWL_1 a_6803_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1895 a_2449_6226# WWL_8 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1896 GND a_3609_286# a_3553_308# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1897 a_16893_1118# RWL_27 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1898 a_17622_1636# a_17529_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1899 a_18202_2716# a_18109_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1900 a_17243_4088# a_17042_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1901 VDD a_10082_17# a_9989_17# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1902 a_18202_6496# a_18109_6496# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1903 GND a_15302_6496# a_15209_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1904 a_17622_5416# a_17529_5416# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1905 a_12982_4336# a_12889_4336# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1906 a_14049_7846# WWL_2 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1907 GND a_17622_7576# a_17529_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1908 GND a_14629_6496# a_14573_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1909 GND a_129_2986# a_73_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1910 a_7613_7328# RWL_4 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1911 a_8342_7846# a_8249_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1912 a_2393_5168# RWL_12 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1913 WBL_11 WWL_23 a_6602_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1914 RBL0_10 RWL_13 a_6223_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1915 GND a_16949_7576# a_16893_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1916 GND a_4862_17# a_4769_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1917 a_13763_2468# a_13562_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1918 a_4133_1928# RWL_24 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1919 WBL_2 WWL_31 a_1382_16# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1920 VDD a_6022_3256# a_5929_3256# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1921 a_12889_7306# WWL_4 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1922 a_7089_1906# WWL_24 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1923 VDD a_8342_4336# a_8249_4336# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1924 a_18053_4628# RWL_14 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1925 a_7762_826# a_7669_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1926 a_11242_5686# a_11149_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1927 RBL0_23 RWL_17 a_13763_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1928 a_13562_6766# a_13469_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1929 VDD a_4862_2716# a_4769_2716# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1930 a_4862_2986# a_4769_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1931 a_14629_17# WWL_31 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1932 GND a_9409_7306# a_9353_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1933 VDD a_11242_2176# a_11149_2176# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1934 a_423_6248# a_222_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1935 a_9353_848# RWL_28 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1936 a_9502_1906# a_9409_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1937 a_1962_2446# a_1869_2446# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1938 a_8543_3278# a_8342_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1939 a_802_3796# a_709_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1940 a_9123_4358# a_8922_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1941 GND a_15302_17# a_15209_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1942 a_16949_1906# WWL_24 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1943 a_9502_5686# a_9409_5686# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1944 GND a_6602_5686# a_6509_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1945 a_802_7576# a_709_7576# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1946 a_4282_3526# a_4189_3526# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1947 a_5349_7036# WWL_5 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1948 GND a_129_5956# a_73_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1949 a_2542_556# a_2449_556# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1950 WBL_23 WWL_2 a_13562_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1951 GND a_8922_6766# a_8829_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1952 GND a_5929_5686# a_5873_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1953 GND a_1289_4606# a_1233_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1954 a_7669_8116# WWL_1 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1955 a_18202_2446# a_18109_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1956 a_17622_1366# a_17529_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1957 a_18202_6226# a_18109_6226# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1958 GND a_15302_6226# a_15209_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1959 RBL0_12 RWL_28 a_7383_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1960 WBL_31 WWL_6 a_18202_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1961 WBL_30 WWL_10 a_17622_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1962 RBL0_15 RWL_10 a_9123_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1963 a_6022_6496# a_5929_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1964 a_4483_308# a_4282_286# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1965 WBL_22 WWL_14 a_12982_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1966 GND a_14629_6226# a_14573_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1967 VDD a_8922_556# a_8829_556# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1968 a_7613_7058# RWL_5 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1969 a_8342_7576# a_8249_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1970 a_11443_1118# a_11242_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1971 GND a_7089_826# a_7033_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1972 a_12889_556# WWL_29 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1973 WBL_11 WWL_24 a_6602_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1974 a_11822_2446# a_11729_2446# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1975 a_13763_2198# a_13562_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1976 a_9353_3818# RWL_17 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1977 a_653_5708# RWL_10 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1978 GND a_1962_826# a_1869_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1979 GND a_11822_4606# a_11729_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1980 a_4133_1658# RWL_25 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1981 VDD a_11822_8386# a_11729_8386# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1982 a_2163_7328# a_1962_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1983 a_10569_5956# WWL_9 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1984 VDD a_6022_2986# a_5929_2986# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1985 a_4862_5956# a_4769_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1986 a_5442_287# a_5349_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1987 a_18053_4358# RWL_15 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1988 a_14629_3796# WWL_17 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1989 a_11242_5416# a_11149_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1990 a_7762_556# a_7669_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1991 VDD a_2542_1366# a_2449_1366# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1992 RBL0_23 RWL_18 a_13763_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1993 RBL0_24 RWL_14 a_14343_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1994 GND a_9409_7036# a_9353_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1995 a_14573_2738# RWL_21 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1996 a_12603_8408# a_12402_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1997 VDD a_16462_4066# a_16369_4066# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1998 a_7033_309# RWL_30 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1999 VDD a_11242_1906# a_11149_1906# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2000 a_9353_578# RWL_29 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2001 a_9502_1636# a_9409_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2002 a_1962_2176# a_1869_2176# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2003 a_9123_4088# a_8922_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2004 GND a_7182_6496# a_7089_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2005 a_10513_309# RWL_30 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2006 a_802_3526# a_709_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2007 a_9502_5416# a_9409_5416# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2008 GND a_6602_5416# a_6509_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2009 a_802_7306# a_709_7306# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2010 a_2542_286# a_2449_286# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2011 WBL_7 WWL_17 a_4282_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2012 GND a_5929_5416# a_5873_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2013 GND a_1289_4336# a_1233_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2014 VDD a_12982_2446# a_12889_2446# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2015 a_18202_2176# a_18109_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2016 RBL0_8 RWL_30 a_5063_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2017 RBL0_12 RWL_29 a_7383_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2018 WBL_31 WWL_7 a_18202_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2019 WBL_30 WWL_11 a_17622_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2020 RBL0_15 RWL_11 a_9123_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2021 RBL0_0 RWL_4 a_423_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2022 a_6022_6226# a_5929_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2023 a_1869_5146# WWL_12 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2024 WBL_11 WWL_30 a_6602_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2025 a_16663_3008# a_16462_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2026 a_11242_826# a_11149_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2027 GND a_7089_556# a_7033_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2028 a_12402_3256# a_12309_3256# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2029 a_11822_2176# a_11729_2176# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2030 a_653_5438# RWL_11 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2031 GND a_1962_556# a_1869_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2032 a_9353_3548# RWL_18 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2033 GND a_11822_4336# a_11729_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2034 a_15789_7846# WWL_2 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2035 a_10513_7868# RWL_2 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2036 a_4133_1388# RWL_26 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2037 RBL0_9 RWL_17 a_5643_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2038 a_2163_7058# a_1962_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2039 a_2542_4606# a_2449_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2040 VDD a_11822_8116# a_11729_8116# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2041 a_2542_8386# a_2449_8386# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2042 a_4282_16# a_4189_16# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2043 GND a_17622_826# a_17529_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2044 a_5873_1928# RWL_24 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2045 a_18053_4088# RWL_16 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2046 a_16462_7306# a_16369_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2047 VDD a_7762_3256# a_7669_3256# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2048 a_14629_3526# WWL_18 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2049 a_15209_4606# WWL_14 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2050 a_11242_5146# a_11149_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2051 VDD a_2542_1096# a_2449_1096# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2052 RBL0_23 RWL_19 a_13763_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2053 RBL0_24 RWL_15 a_14343_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2054 RBL0_3 RWL_0 a_2163_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2055 a_14573_2468# RWL_22 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2056 a_12603_8138# a_12402_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2057 WBL_15 WWL_28 a_8922_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2058 a_7182_4066# a_7089_4066# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2059 VDD a_12402_556# a_12309_556# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2060 GND a_8829_287# a_8773_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2061 a_9502_1366# a_9409_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2062 a_1962_1906# a_1869_1906# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2063 GND a_12309_7846# a_12253_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2064 GND a_7182_6226# a_7089_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2065 WBL_21 WWL_28 a_12402_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2066 WBL_3 WWL_22 a_1962_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2067 a_802_3256# a_709_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2068 GND a_6602_5146# a_6509_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2069 WBL_1 WWL_3 a_802_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2070 a_802_7036# a_709_7036# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2071 WBL_16 WWL_10 a_9502_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2072 a_2542_16# a_2449_16# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2073 WBL_7 WWL_18 a_4282_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2074 a_16663_5978# a_16462_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2075 GND a_5929_5146# a_5873_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2076 a_3323_1118# a_3122_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2077 GND a_1289_4066# a_1233_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2079 VDD a_12982_2176# a_12889_2176# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2080 a_3702_2446# a_3609_2446# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2081 WBL_27 WWL_12 a_15882_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2082 WBL_31 WWL_8 a_18202_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2083 RBL0_0 RWL_5 a_423_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2084 RBL0_15 RWL_12 a_9123_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2085 a_1869_4876# WWL_13 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2086 WBL_11 WWL_31 a_6602_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2087 a_11242_556# a_11149_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2088 a_11822_1906# a_11729_1906# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2089 a_12402_2986# a_12309_2986# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2090 VDD a_10082_7846# a_9989_7846# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2091 a_653_5168# RWL_12 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2092 a_9353_3278# RWL_19 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2093 a_6509_3796# WWL_17 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2094 a_10513_7598# a_4683_7576# RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2095 a_7762_6496# a_7669_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2096 a_5929_2716# WWL_21 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2097 GND a_11822_4066# a_11729_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2098 RBL0_9 RWL_18 a_5643_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2099 a_2542_4336# a_2449_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2100 a_2542_8116# a_2449_8116# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2101 GND a_14142_1906# a_14049_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2102 GND a_15302_287# a_15209_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2103 GND a_17622_556# a_17529_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2104 a_17529_4336# WWL_15 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2105 VDD a_14142_5686# a_14049_5686# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2106 GND a_13469_1906# a_13413_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2107 RBL0_20 RWL_20 a_12023_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2108 GND a_14629_826# a_14573_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2109 a_5873_1658# RWL_25 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2110 a_3903_7328# a_3702_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2111 a_16462_7036# a_16369_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2112 VDD a_7762_2986# a_7669_2986# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2113 RBL0_24 RWL_16 a_14343_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2114 a_3029_8386# WWL_0 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2115 RBL0_3 RWL_1 a_2163_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2116 a_12253_1118# RWL_27 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2117 a_14573_2198# RWL_23 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2118 WBL_17 WWL_30 a_10082_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2119 WBL_12 WWL_15 a_7182_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2120 WBL_3 WWL_23 a_1962_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2121 GND a_12309_7576# a_12253_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2122 a_14343_4628# a_14142_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2123 WBL_1 WWL_4 a_802_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2124 WBL_16 WWL_11 a_9502_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2125 a_222_2446# a_129_2446# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2126 a_9703_309# a_9502_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2127 VDD a_12982_1906# a_12889_1906# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2128 GND a_222_4606# a_129_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2129 VDD a_222_8386# a_129_8386# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2130 a_3702_286# a_3609_286# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2131 a_3702_2176# a_3609_2176# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2132 GND a_8249_2716# a_8193_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2133 WBL_27 WWL_13 a_15882_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2134 a_802_556# a_709_556# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2135 a_1813_6788# RWL_6 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2136 a_1962_16# a_1869_16# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2137 a_13413_8408# RWL_0 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2138 a_12833_7328# RWL_4 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2139 a_4189_2446# WWL_22 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2140 RBL0_20 RWL_9 a_12023_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2141 WBL_21 WWL_19 a_12402_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2142 a_7762_6226# a_7669_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2143 a_6509_3526# WWL_18 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2144 RBL0_9 RWL_19 a_5643_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2145 a_2542_4066# a_2449_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2146 WBL_4 WWL_0 a_2542_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2147 GND a_14142_1636# a_14049_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2148 a_18109_5146# WWL_12 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2149 a_17529_4066# WWL_16 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2150 VDD a_14142_5416# a_14049_5416# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2151 GND a_12309_287# a_12253_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2152 GND a_13469_1636# a_13413_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2153 GND a_14629_556# a_14573_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2154 a_5873_1388# RWL_26 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2155 a_3903_7058# a_3702_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2156 a_4769_826# WWL_28 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2157 RBL0_5 RWL_30 a_3323_308# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2158 a_3323_38# a_3122_16# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2159 a_3029_8116# WWL_1 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2160 GND a_4189_7846# a_4133_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2161 GND a_3609_6766# a_3553_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2162 a_17473_3008# RWL_20 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2163 a_15503_848# a_15302_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2164 a_5643_3818# a_5442_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2165 VDD a_802_1366# a_709_1366# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2166 VDD a_10662_3796# a_10569_3796# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2167 a_7963_4898# a_7762_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2168 GND a_15209_8386# a_15153_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2169 a_10662_7846# a_10569_7846# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2170 a_7762_287# a_7669_287# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2171 WBL_17 WWL_31 a_10082_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2172 WBL_12 WWL_16 a_7182_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2173 RBL0_6 RWL_0 a_3903_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2174 WBL_3 WWL_24 a_1962_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2175 a_14722_1906# a_14629_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2176 a_14343_4358# a_14142_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2177 a_15302_6766# a_15209_6766# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2178 a_14722_5686# a_14629_5686# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2179 a_222_2176# a_129_2176# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2180 a_10082_4606# a_9989_4606# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2181 GND a_14722_7846# a_14629_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2182 GND a_10082_6766# a_9989_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2183 GND a_222_4336# a_129_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2184 a_7033_4898# RWL_13 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2185 GND a_1382_2986# a_1289_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2186 VDD a_222_8116# a_129_8116# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2187 a_3702_1906# a_3609_1906# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2188 GND a_8249_2446# a_8193_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2189 WBL_6 WWL_22 a_3702_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2190 a_802_286# a_709_286# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2191 a_10863_2738# a_10662_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2192 a_9409_4336# WWL_15 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2193 a_13413_8138# RWL_1 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2194 RBL0_29 RWL_2 a_17243_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2195 a_12833_7058# RWL_5 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2196 a_423_38# a_222_16# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2197 a_8829_3256# WWL_19 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2198 RBL0_28 RWL_6 a_16663_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2199 a_4189_2176# WWL_23 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2200 WBL_21 WWL_20 a_12402_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2201 VDD a_5442_4606# a_5349_4606# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2202 WBL_8 WWL_29 a_4862_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2203 a_17473_5978# RWL_9 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2204 WBL_4 WWL_1 a_2542_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2205 GND a_14142_1366# a_14049_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2206 a_13562_826# a_13469_826# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2207 a_18109_4876# WWL_13 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2208 GND a_13469_1366# a_13413_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2209 a_13183_309# a_12982_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2210 GND a_15882_1906# a_15789_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2211 GND a_4189_7576# a_4133_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2212 a_6223_4628# a_6022_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2213 VDD a_15882_5686# a_15789_5686# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2214 a_15503_578# a_15302_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2215 a_5643_3548# a_5442_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2216 VDD a_802_1096# a_709_1096# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2217 VDD a_10662_3526# a_10569_3526# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2218 a_1382_3796# a_1289_3796# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2219 a_7762_17# a_7669_17# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2220 GND a_15209_8116# a_15153_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2221 GND a_1382_5956# a_1289_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2222 GND a_17529_17# a_17473_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2223 a_4769_8386# WWL_0 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2224 RBL0_6 RWL_1 a_3903_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2225 a_13993_1118# RWL_27 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2226 a_14722_1636# a_14629_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2227 a_15302_2716# a_15209_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2228 a_14343_4088# a_14142_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2229 a_15302_6496# a_15209_6496# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2230 GND a_12402_6496# a_12309_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2231 a_14722_5416# a_14629_5416# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2232 a_222_1906# a_129_1906# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2233 WBL_0 WWL_22 a_222_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2234 a_10082_4336# a_9989_4336# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2235 a_11149_7846# WWL_2 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2236 RBL0_1 RWL_17 a_1003_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2237 GND a_14722_7576# a_14629_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2238 GND a_11729_6496# a_11673_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2239 GND a_222_4066# a_129_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2240 a_5442_7846# a_5349_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2241 a_4713_7328# RWL_4 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2242 WBL_6 WWL_23 a_3702_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2243 RBL0_5 RWL_13 a_3323_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2244 GND a_222_826# a_129_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2245 GND a_8249_2176# a_8193_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2246 a_802_16# a_709_16# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2247 a_10863_2468# a_10662_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2248 a_1233_1928# RWL_24 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2249 VDD a_3122_3256# a_3029_3256# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2250 RBL0_29 a_13963_7576# a_17243_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2251 a_709_5956# WWL_9 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2252 a_8829_2986# WWL_20 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2253 a_9409_4066# WWL_16 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2254 a_4189_1906# WWL_24 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2255 GND a_9989_2716# a_9933_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2256 VDD a_5442_4336# a_5349_4336# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2257 a_15153_4628# RWL_14 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2258 VDD a_17042_5956# a_16949_5956# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2259 a_11242_287# a_11149_287# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2260 RBL0_18 RWL_17 a_10863_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2261 a_10662_6766# a_10569_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2262 VDD a_1962_2716# a_1869_2716# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2263 WBL_8 WWL_10 a_4862_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2264 GND a_7089_8386# a_7033_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2265 GND a_6509_7306# a_6453_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2266 GND a_15882_1636# a_15789_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2267 VDD a_15882_5416# a_15789_5416# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2268 VDD a_17622_287# a_17529_287# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2269 a_6602_1906# a_6509_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2270 a_5643_3278# a_5442_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2271 a_6223_4358# a_6022_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2272 GND a_3702_5686# a_3609_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2273 a_6602_5686# a_6509_5686# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2274 a_1382_3526# a_1289_3526# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2275 WBL_18 WWL_2 a_10662_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2276 a_2449_7036# WWL_5 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2277 a_4769_8116# WWL_1 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2278 a_12982_5146# a_12889_5146# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2279 a_15302_2446# a_15209_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2280 GND a_17622_8386# a_17529_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2281 a_14722_1366# a_14629_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2282 WBL_26 WWL_6 a_15302_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2283 a_15302_6226# a_15209_6226# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2284 GND a_12402_6226# a_12309_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2285 a_3122_6496# a_3029_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2286 WBL_25 WWL_10 a_14722_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2287 RBL0_10 RWL_10 a_6223_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2288 WBL_0 WWL_23 a_222_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2289 GND a_16949_8386# a_16893_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2290 RBL0_1 RWL_18 a_1003_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2291 WBL_17 WWL_14 a_10082_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2292 GND a_11729_6226# a_11673_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2293 GND a_4769_17# a_4713_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2294 a_4713_7058# RWL_5 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2295 RBL0_14 RWL_6 a_8543_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2296 a_5442_7576# a_5349_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2297 WBL_6 WWL_24 a_3702_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2298 GND a_222_556# a_129_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2299 a_10863_2198# a_10662_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2300 a_6453_3818# RWL_17 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2301 a_1233_1658# RWL_25 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2302 VDD a_8342_5146# a_8249_5146# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2303 VDD a_3122_2986# a_3029_2986# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2304 a_8773_4898# RWL_13 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2305 GND a_9989_2446# a_9933_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2306 a_15153_4358# RWL_15 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2307 a_11729_3796# WWL_17 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2308 RBL0_18 RWL_18 a_10863_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2309 RBL0_19 RWL_14 a_11443_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2310 RBL0_14 RWL_30 a_8543_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2311 a_11242_17# a_11149_17# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2312 GND a_3122_16# a_3029_16# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2313 WBL_8 WWL_11 a_4862_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2314 GND a_7089_8116# a_7033_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2315 a_17243_7868# a_17042_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2316 GND a_6509_7036# a_6453_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2317 GND a_15209_17# a_15153_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2318 a_11673_2738# RWL_21 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2319 VDD a_13562_4066# a_13469_4066# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2320 GND a_15882_1366# a_15789_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2321 VDD a_17622_17# a_17529_17# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2322 a_6602_1636# a_6509_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2323 a_6223_4088# a_6022_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2324 GND a_4282_6496# a_4189_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2325 a_6602_5416# a_6509_5416# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2326 GND a_3702_5416# a_3609_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2327 a_73_6788# RWL_6 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2328 WBL_2 WWL_17 a_1382_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2329 a_12982_1096# a_12889_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2330 a_17622_5956# a_17529_5956# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2331 a_16313_848# RWL_28 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2332 a_12982_4876# a_12889_4876# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2333 a_15302_2176# a_15209_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2334 GND a_17622_8116# a_17529_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2335 a_6022_556# a_5929_556# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2336 a_8342_8386# a_8249_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2337 a_7089_5686# WWL_10 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2338 WBL_26 WWL_7 a_15302_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2339 WBL_25 WWL_11 a_14722_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2340 RBL0_10 RWL_11 a_6223_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2341 WBL_0 WWL_24 a_222_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2342 GND a_16949_8116# a_16893_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2343 a_3122_6226# a_3029_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2344 RBL0_1 RWL_19 a_1003_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2345 a_13763_3008# a_13562_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2346 a_17042_2716# a_16949_2716# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2347 GND a_14049_3796# a_13993_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2348 GND a_17042_4876# a_16949_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2349 GND a_8342_1096# a_8249_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2350 RBL0_24 RWL_28 a_14343_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2351 a_6453_3548# RWL_18 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2352 a_12889_7846# WWL_2 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2353 GND a_222_16# a_129_16# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2354 a_1233_1388# RWL_26 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2355 RBL0_4 RWL_17 a_2743_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2356 GND a_16369_4876# a_16313_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2357 VDD a_8342_4876# a_8249_4876# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2358 GND a_7669_1096# a_7613_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2359 VDD a_15882_556# a_15789_556# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2360 a_18403_1928# a_18202_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2361 a_16369_556# WWL_29 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2362 GND a_9989_2176# a_9933_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2363 GND a_5442_826# a_5349_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2364 a_16949_5686# WWL_10 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2365 a_2973_1928# RWL_24 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2366 a_15153_4088# RWL_16 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2367 a_12309_4606# WWL_14 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2368 a_13562_7306# a_13469_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2369 VDD a_4862_3256# a_4769_3256# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2370 a_11729_3526# WWL_18 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2371 RBL0_18 RWL_19 a_10863_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2372 RBL0_19 RWL_15 a_11443_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2373 a_8922_287# a_8829_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2374 a_12402_287# a_12309_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2375 a_16893_4628# RWL_14 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2376 a_17243_7598# a_17042_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2377 a_11673_2468# RWL_22 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2378 a_4282_4066# a_4189_4066# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2379 GND a_129_6496# a_73_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2380 a_6602_1366# a_6509_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2381 GND a_8922_7306# a_8829_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2382 GND a_4282_6226# a_4189_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2383 GND a_3702_5146# a_3609_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2384 WBL_11 WWL_10 a_6602_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2385 WBL_2 WWL_18 a_1382_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2386 a_13763_5978# a_13562_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2387 VDD a_17622_1636# a_17529_1636# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2388 a_18202_2986# a_18109_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2389 VDD a_6022_6766# a_5929_6766# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2390 a_16313_578# RWL_29 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2391 WBL_22 WWL_12 a_12982_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2392 a_7089_5416# WWL_11 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2393 a_8342_8116# a_8249_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2394 WBL_26 WWL_8 a_15302_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2395 RBL0_10 RWL_12 a_6223_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2396 RBL0_20 RWL_30 a_12023_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2397 RBL0_13 RWL_24 a_7963_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2398 GND a_14049_3526# a_13993_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2399 RBL0_24 RWL_29 a_14343_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2400 a_6453_3278# RWL_19 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2401 a_3609_3796# WWL_17 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2402 a_4862_6496# a_4769_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2403 a_13993_39# RWL_31 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2404 a_18403_1658# a_18202_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2405 RBL0_4 RWL_18 a_2743_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2406 GND a_11242_1906# a_11149_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2407 VDD a_11242_5686# a_11149_5686# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2408 GND a_5442_556# a_5349_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2409 a_14629_4336# WWL_15 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2410 GND a_10569_1906# a_10513_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2411 a_9123_7868# a_8922_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2412 a_8543_6788# a_8342_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2413 a_16949_5416# WWL_11 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2414 GND a_2449_826# a_2393_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2415 a_2973_1658# RWL_25 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2416 a_13562_7036# a_13469_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2417 VDD a_4862_2986# a_4769_2986# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2418 RBL0_19 RWL_16 a_11443_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2419 a_18202_5956# a_18109_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2420 a_16893_4358# RWL_15 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2421 a_11673_2198# RWL_23 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2422 a_17622_4876# a_17529_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2423 a_9502_5956# a_9409_5956# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2424 a_802_7846# a_709_7846# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2425 GND a_129_6226# a_73_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2426 WBL_7 WWL_15 a_4282_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2427 GND a_8922_7036# a_8829_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2428 a_11443_4628# a_11242_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2429 WBL_11 WWL_11 a_6602_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2430 GND a_6022_2716# a_5929_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2431 WBL_27 WWL_28 a_15882_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2432 a_8342_1636# a_8249_1636# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2433 WBL_31 WWL_5 a_18202_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2434 VDD a_6022_6496# a_5929_6496# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2435 WBL_30 WWL_9 a_17622_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2436 GND a_15789_287# a_15733_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2437 GND a_5349_2716# a_5293_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2438 WBL_22 WWL_13 a_12982_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2440 a_1003_2738# a_802_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2441 a_18053_7868# RWL_2 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2442 a_10513_8408# RWL_0 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2443 a_129_3796# WWL_17 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2444 RBL0_13 RWL_25 a_7963_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2445 a_1289_2446# WWL_22 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2446 WBL_29 WWL_21 a_17042_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2447 GND a_14049_3256# a_13993_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2448 a_4862_6226# a_4769_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2449 a_3609_3526# WWL_18 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2450 a_18403_1388# a_18202_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2451 RBL0_4 RWL_19 a_2743_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2452 GND a_16462_3796# a_16369_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2453 GND a_11242_1636# a_11149_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2454 VDD a_16462_7576# a_16369_7576# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2455 a_15209_5146# WWL_12 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2456 a_1962_1906# a_1869_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2457 GND a_15789_3796# a_15733_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2458 a_14629_4066# WWL_16 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2459 VDD a_11242_5416# a_11149_5416# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2461 a_9123_7598# a_8922_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2462 a_1962_5686# a_1869_5686# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2463 GND a_10569_1636# a_10513_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2464 GND a_2449_556# a_2393_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2465 a_2973_1388# RWL_26 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2466 GND a_1289_7846# a_1233_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2467 a_3323_848# a_3122_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2468 RBL0_31 RWL_21 a_18403_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2469 a_14573_3008# RWL_20 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2470 GND a_18109_826# a_18053_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2471 a_2743_3818# a_2542_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2472 a_16893_4088# RWL_16 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2473 GND a_12309_8386# a_12253_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2474 WBL_7 WWL_16 a_4282_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2475 a_16663_6518# a_16462_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2476 a_11822_1906# a_11729_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2477 a_11443_4358# a_11242_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2478 a_12402_6766# a_12309_6766# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2479 a_11822_5686# a_11729_5686# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2480 GND a_11822_7846# a_11729_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2481 GND a_6022_2446# a_5929_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2482 a_4133_4898# RWL_13 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2483 VDD a_6022_6226# a_5929_6226# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2484 GND a_5349_2446# a_5293_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2485 a_11673_39# RWL_31 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2486 a_1003_2468# a_802_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2487 a_18053_7598# a_13963_7576# RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2488 VDD a_7762_6766# a_7669_6766# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2489 a_6509_4336# WWL_15 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2490 a_10513_8138# RWL_1 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2491 RBL0_24 RWL_2 a_14343_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2492 RBL0_13 RWL_26 a_7963_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2493 a_5929_3256# WWL_19 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2494 a_129_3526# WWL_18 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2495 VDD a_2542_4606# a_2449_4606# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2496 RBL0_23 RWL_6 a_13763_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2497 a_1289_2176# WWL_23 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2498 a_16462_1366# a_16369_1366# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2499 GND a_16462_3526# a_16369_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2500 a_14573_5978# RWL_9 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2501 a_1382_826# a_1289_826# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2502 GND a_11242_1366# a_11149_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2503 RBL0_16 RWL_24 a_9703_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2504 a_7182_3796# a_7089_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2505 VDD a_16462_7306# a_16369_7306# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2506 a_1962_1636# a_1869_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2507 a_15209_4876# WWL_13 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2508 a_7182_7576# a_7089_7576# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2509 GND a_15789_3526# a_15733_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2510 a_1962_5416# a_1869_5416# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2511 GND a_10569_1366# a_10513_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2512 a_9502_4876# a_9409_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2513 a_802_6766# a_709_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2514 WBL_30 WWL_30 a_17622_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2515 GND a_12982_1906# a_12889_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2516 GND a_1289_7576# a_1233_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2517 a_7963_5708# a_7762_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2518 a_3323_578# a_3122_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2519 a_3323_4628# a_3122_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2520 VDD a_12982_5686# a_12889_5686# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2521 VDD a_7762_826# a_7669_826# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2522 GND a_18109_556# a_18053_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2523 RBL0_31 RWL_22 a_18403_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2524 a_2743_3548# a_2542_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2525 a_8249_826# WWL_28 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2526 GND a_12309_8116# a_12253_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2527 WBL_1 WWL_2 a_802_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2528 WBL_16 WWL_9 a_9502_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2529 a_1869_8386# WWL_0 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2530 a_16663_6248# a_16462_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2531 a_11822_1636# a_11729_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2532 a_12402_2716# a_12309_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2533 a_11443_4088# a_11242_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2534 a_7033_5708# RWL_10 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2535 a_12402_6496# a_12309_6496# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2536 a_11822_5416# a_11729_5416# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2537 GND a_1382_286# a_1289_286# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2538 a_9353_6788# RWL_6 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2539 GND a_3029_1096# a_2973_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2540 GND a_6022_2176# a_5929_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2541 GND a_11822_7576# a_11729_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2542 a_2542_7846# a_2449_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2543 a_1813_7328# RWL_4 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2544 GND a_5349_2176# a_5293_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2545 RBL0_20 RWL_7 a_12023_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2546 a_1003_2198# a_802_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2547 GND a_7762_2716# a_7669_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2548 RBL0_24 a_13963_7576# a_14343_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2549 VDD a_7762_6496# a_7669_6496# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2550 a_5929_2986# WWL_20 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2551 a_6509_4066# WWL_16 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2552 a_1289_1906# WWL_24 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2553 VDD a_2542_4336# a_2449_4336# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2554 a_16462_1096# a_16369_1096# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2555 a_12253_4628# RWL_14 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2556 WBL_28 WWL_25 a_16462_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2557 VDD a_14142_5956# a_14049_5956# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2558 GND a_16462_3256# a_16369_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2559 RBL0_16 RWL_25 a_9703_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2560 a_7182_3526# a_7089_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2561 VDD a_16462_7036# a_16369_7036# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2562 a_1962_1366# a_1869_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2563 GND a_15789_3256# a_15733_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2564 a_7182_7306# a_7089_7306# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2565 WBL_3 WWL_10 a_1962_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2566 GND a_4189_8386# a_4133_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2567 GND a_3609_7306# a_3553_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2568 VDD a_18202_3796# a_18109_3796# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2569 a_17042_826# a_16949_826# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2570 RBL0_27 RWL_27 a_16083_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2571 WBL_30 WWL_31 a_17622_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2572 GND a_12982_1636# a_12889_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2573 a_7963_5438# a_7762_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2574 VDD a_5442_287# a_5349_287# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2575 a_3702_1906# a_3609_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2576 a_3323_4358# a_3122_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2577 VDD a_12982_5416# a_12889_5416# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2578 RBL0_31 RWL_23 a_18403_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2579 a_2743_3278# a_2542_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2580 WBL_27 WWL_0 a_15882_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2581 a_3702_5686# a_3609_5686# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2582 a_1869_8116# WWL_1 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2583 a_10082_5146# a_9989_5146# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2584 a_11822_1366# a_11729_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2585 a_12402_2446# a_12309_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2586 GND a_14722_8386# a_14629_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2587 GND a_10082_7306# a_9989_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2588 a_7033_5438# RWL_11 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2589 WBL_21 WWL_6 a_12402_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2590 a_12402_6226# a_12309_6226# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2591 a_10863_848# a_10662_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2592 RBL0_5 RWL_10 a_3323_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2593 GND a_8249_2986# a_8193_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2594 a_1813_7058# RWL_5 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2595 RBL0_9 RWL_6 a_5643_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2596 a_2542_7576# a_2449_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2597 a_17529_7576# WWL_3 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2598 a_3553_3818# RWL_17 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2599 RBL0_29 RWL_0 a_17243_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2600 RBL0_28 RWL_4 a_16663_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2601 RBL0_20 RWL_8 a_12023_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2602 VDD a_5442_5146# a_5349_5146# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2603 GND a_7762_2446# a_7669_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2604 a_5873_4898# RWL_13 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2605 VDD a_7762_6226# a_7669_6226# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2606 a_17473_6518# RWL_7 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2607 VDD a_11242_826# a_11149_826# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2608 WBL_28 WWL_26 a_16462_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2609 a_12253_4358# RWL_15 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2610 a_9502_556# a_9409_556# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2611 RBL0_16 RWL_26 a_9703_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2612 a_7182_3256# a_7089_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2613 WBL_12 WWL_3 a_7182_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2614 a_7182_7036# a_7089_7036# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2615 WBL_3 WWL_11 a_1962_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2616 GND a_4189_8116# a_4133_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2617 a_14343_7868# a_14142_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2618 a_222_1906# a_129_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2619 GND a_3609_7036# a_3553_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2620 VDD a_18202_3526# a_18109_3526# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2621 a_8922_3796# a_8829_3796# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2622 VDD a_10662_4066# a_10569_4066# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2623 a_222_5686# a_129_5686# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2624 GND a_12982_1366# a_12889_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2625 a_7963_5168# a_7762_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2626 VDD a_5442_17# a_5349_17# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2627 GND a_222_7846# a_129_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2628 a_3702_1636# a_3609_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2629 a_3323_4088# a_3122_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2630 GND a_1382_6496# a_1289_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2631 WBL_27 WWL_1 a_15882_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2632 a_3702_5416# a_3609_5416# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2633 GND a_8249_5956# a_8193_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2634 a_10082_1096# a_9989_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2635 a_14722_5956# a_14629_5956# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2636 a_10082_4876# a_9989_4876# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2637 a_12402_2176# a_12309_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2638 GND a_14722_8116# a_14629_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2639 GND a_10082_7036# a_9989_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2640 a_8829_6766# WWL_6 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2641 a_7033_5168# RWL_12 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2642 a_5442_8386# a_5349_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2643 a_4189_5686# WWL_10 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2644 a_10863_578# a_10662_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2645 WBL_21 WWL_7 a_12402_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2646 RBL0_5 RWL_11 a_3323_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2647 a_10863_3008# a_10662_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2648 RBL0_30 RWL_31 a_17823_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2649 a_14142_2716# a_14049_2716# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2650 a_8773_5708# RWL_10 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2651 GND a_11149_3796# a_11093_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2652 GND a_14142_4876# a_14049_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2653 a_18109_8386# WWL_0 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2654 GND a_5442_1096# a_5349_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2655 a_3553_3548# RWL_18 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2656 RBL0_29 RWL_1 a_17243_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2657 a_17529_7306# WWL_4 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2658 RBL0_28 RWL_5 a_16663_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2659 a_15503_1928# a_15302_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2660 GND a_13469_4876# a_13413_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2661 VDD a_5442_4876# a_5349_4876# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2662 GND a_4769_1096# a_4713_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2663 a_4189_556# WWL_29 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2664 GND a_7762_2176# a_7669_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2665 a_17473_6248# RWL_8 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2666 VDD a_9502_2716# a_9409_2716# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2667 WBL_28 WWL_27 a_16462_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2668 a_12253_4088# RWL_16 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2669 VDD a_802_4606# a_709_4606# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2670 a_10662_7306# a_10569_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2671 GND a_3029_16# a_2973_38# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2672 VDD a_1962_3256# a_1869_3256# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2673 WBL_12 WWL_4 a_7182_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2674 a_13993_4628# RWL_14 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2675 a_14343_7598# a_14142_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2676 VDD a_15882_5956# a_15789_5956# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2677 a_222_1636# a_129_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2678 a_8922_3526# a_8829_3526# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2679 a_222_5416# a_129_5416# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2680 a_1382_4066# a_1289_4066# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2681 GND a_222_7576# a_129_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2682 a_3702_1366# a_3609_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2683 GND a_1382_6226# a_1289_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2684 WBL_6 WWL_10 a_3702_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2685 a_18202_826# a_18109_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2686 a_10863_5978# a_10662_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2687 RBL0_30 RWL_27 a_17823_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2688 VDD a_14722_1636# a_14629_1636# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2689 a_15302_2986# a_15209_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2690 VDD a_3122_6766# a_3029_6766# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2691 WBL_17 WWL_12 a_10082_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2692 a_9409_7576# WWL_3 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2693 a_8829_6496# WWL_7 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2694 RBL0_14 RWL_4 a_8543_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2695 a_4189_5416# WWL_11 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2696 a_5442_8116# a_5349_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2697 WBL_21 WWL_8 a_12402_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2698 RBL0_5 RWL_12 a_3323_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2699 GND a_17042_5686# a_16949_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2700 GND a_129_16# a_73_38# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2701 GND a_16369_5686# a_16313_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2702 a_12982_556# a_12889_556# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2703 RBL0_8 RWL_24 a_5063_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2704 a_8773_5438# RWL_11 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2705 GND a_11149_3526# a_11093_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2706 a_18109_8116# WWL_1 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2707 a_3553_3278# RWL_19 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2708 GND a_9989_2986# a_9933_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2709 a_4189_286# WWL_30 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2710 a_15503_1658# a_15302_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2711 a_11729_4336# WWL_15 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2712 a_6223_7868# a_6022_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2713 a_5643_6788# a_5442_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2714 VDD a_802_4336# a_709_4336# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2715 a_10662_7036# a_10569_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2716 VDD a_1962_2986# a_1869_2986# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2717 WBL_8 WWL_9 a_4862_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2718 a_5873_309# RWL_30 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2719 a_17243_8408# a_17042_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2720 a_15302_5956# a_15209_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2721 a_13993_4358# RWL_15 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2722 a_222_1366# a_129_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2723 a_14722_4876# a_14629_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2724 a_6602_5956# a_6509_5956# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2725 WBL_0 WWL_10 a_222_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2726 WBL_15 WWL_17 a_8922_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2727 a_73_7328# RWL_4 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2728 WBL_2 WWL_15 a_1382_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2729 a_9123_39# a_8922_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2730 VDD a_17622_2446# a_17529_2446# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2731 a_18202_556# a_18109_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2732 WBL_6 WWL_11 a_3702_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2733 RBL0_26 RWL_31 a_15503_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2734 GND a_3122_2716# a_3029_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2735 a_5442_1636# a_5349_1636# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2736 WBL_26 WWL_5 a_15302_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2737 VDD a_3122_6496# a_3029_6496# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2738 WBL_25 WWL_9 a_14722_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2739 GND a_2449_2716# a_2393_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2740 WBL_17 WWL_13 a_10082_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2741 a_9409_7306# WWL_4 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2742 RBL0_14 RWL_5 a_8543_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2743 a_8829_6226# WWL_8 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2744 GND a_9989_5956# a_9933_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2745 a_17042_3256# a_16949_3256# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2746 a_1813_38# RWL_31 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2747 WBL_20 WWL_25 a_11822_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2748 GND a_17042_5416# a_16949_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2749 a_15153_7868# RWL_2 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2750 WBL_24 WWL_21 a_14142_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2751 GND a_16369_5416# a_16313_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2752 RBL0_8 RWL_25 a_5063_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2753 GND a_11149_3256# a_11093_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2754 a_8773_5168# RWL_12 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2755 a_11673_848# RWL_28 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2756 a_15503_1388# a_15302_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2757 a_4189_16# WWL_31 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2758 GND a_13562_3796# a_13469_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2759 a_15882_2716# a_15789_2716# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2760 VDD a_13562_7576# a_13469_7576# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2761 a_12309_5146# WWL_12 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2762 GND a_12889_3796# a_12833_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2763 a_11729_4066# WWL_16 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2764 GND a_15882_4876# a_15789_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2765 a_6223_7598# a_6022_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2766 WBL_13 WWL_28 a_7762_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2767 GND a_10082_287# a_9989_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2768 a_17243_8138# a_17042_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2769 a_17622_5686# a_17529_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2770 a_11729_556# WWL_29 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2771 RBL0_26 RWL_21 a_15503_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2772 a_11673_3008# RWL_20 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2773 a_12982_4606# a_12889_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2774 a_12982_8386# a_12889_8386# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2775 a_13993_4088# RWL_16 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2776 WBL_15 WWL_18 a_8922_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2777 a_73_7058# RWL_5 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2778 WBL_0 WWL_11 a_222_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2779 a_16313_1928# RWL_24 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2780 RBL0_1 RWL_6 a_1003_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2781 WBL_2 WWL_16 a_1382_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2782 a_13763_6518# a_13562_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2783 VDD a_17622_2176# a_17529_2176# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2784 a_8342_2446# a_8249_2446# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2785 GND a_8342_4606# a_8249_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2786 GND a_3122_2446# a_3029_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2787 VDD a_8342_8386# a_8249_8386# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2788 a_7089_5956# WWL_9 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2789 a_1233_4898# RWL_13 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2790 VDD a_3122_6226# a_3029_6226# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2791 GND a_7669_4606# a_7613_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2792 GND a_2449_2446# a_2393_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2793 a_17042_2986# a_16949_2986# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2794 WBL_20 WWL_26 a_11822_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2795 GND a_17042_5146# a_16949_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2796 a_15153_7598# a_13963_7576# RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2797 VDD a_4862_6766# a_4769_6766# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2798 a_3609_4336# WWL_15 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2799 RBL0_19 RWL_2 a_11443_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2800 GND a_16369_5146# a_16313_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2801 RBL0_8 RWL_26 a_5063_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2802 RBL0_18 RWL_6 a_10863_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2803 a_11673_578# RWL_29 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2804 a_13562_1366# a_13469_1366# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2805 GND a_18109_1906# a_18053_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2806 GND a_13562_3526# a_13469_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2807 a_9123_8408# a_8922_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2808 a_8543_7328# a_8342_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2809 a_11673_5978# RWL_9 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2810 a_16949_5956# WWL_9 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2811 RBL0_11 RWL_24 a_6803_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2812 a_4282_3796# a_4189_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2813 VDD a_13562_7306# a_13469_7306# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2814 a_12309_4876# WWL_13 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2815 a_4282_7576# a_4189_7576# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2816 GND a_12889_3526# a_12833_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2817 a_6602_4876# a_6509_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2818 a_9933_39# RWL_31 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2819 a_14049_1636# WWL_25 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2820 WBL_9 WWL_30 a_5442_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2821 a_18202_6496# a_18109_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2822 a_16369_2716# WWL_21 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2823 a_17622_5416# a_17529_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2824 VDD a_8922_1366# a_8829_1366# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2825 a_12982_4336# a_12889_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2826 RBL0_26 RWL_22 a_15503_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2827 a_12982_8116# a_12889_8116# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2828 RBL0_22 RWL_31 a_13183_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2829 WBL_11 WWL_9 a_6602_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2830 a_16313_1658# RWL_25 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2831 a_13763_6248# a_13562_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2832 VDD a_17622_1906# a_17529_1906# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2833 a_4133_5708# RWL_10 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2834 a_8342_2176# a_8249_2176# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2835 GND a_8342_4336# a_8249_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2836 a_6453_6788# RWL_6 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2837 GND a_3122_2176# a_3029_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2838 VDD a_8342_8116# a_8249_8116# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2839 GND a_7669_4336# a_7613_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2840 GND a_2449_2176# a_2393_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2841 a_18053_8408# RWL_0 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2842 WBL_29 WWL_19 a_17042_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2843 a_129_4336# WWL_15 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2844 WBL_20 WWL_27 a_11822_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2845 GND a_4862_2716# a_4769_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2846 a_9409_287# WWL_30 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2847 VDD a_4862_6496# a_4769_6496# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2848 a_3609_4066# WWL_16 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2849 RBL0_19 a_4683_7576# a_11443_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2850 WBL_19 WWL_28 a_11242_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2851 a_13562_1096# a_13469_1096# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2852 GND a_18109_1636# a_18053_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2853 WBL_23 WWL_25 a_13562_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2854 a_16893_7868# RWL_2 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2855 VDD a_11242_5956# a_11149_5956# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2856 a_9123_8138# a_8922_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2857 a_9502_5686# a_9409_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2859 GND a_13562_3256# a_13469_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2860 a_8543_7058# a_8342_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2861 RBL0_11 RWL_25 a_6803_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2862 a_4282_3526# a_4189_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2863 VDD a_13562_7036# a_13469_7036# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2864 a_4282_7306# a_4189_7306# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2865 GND a_12889_3256# a_12833_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2866 GND a_1289_8386# a_1233_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2867 a_14049_1366# WWL_26 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2868 VDD a_15302_3796# a_15209_3796# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2869 GND a_709_286# a_653_308# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2870 WBL_9 WWL_31 a_5442_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2871 RBL0_22 RWL_27 a_13183_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2872 a_18202_6226# a_18109_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2873 VDD a_8922_1096# a_8829_1096# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2874 a_17622_5146# a_17529_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2875 RBL0_26 RWL_23 a_15503_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2876 a_12982_4066# a_12889_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2877 WBL_22 WWL_0 a_12982_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2878 a_16313_1388# RWL_26 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2879 GND a_11822_8386# a_11729_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2880 a_15209_826# WWL_28 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2881 GND a_6022_2986# a_5929_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2882 a_4133_5438# RWL_11 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2883 a_8342_1906# a_8249_1906# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2884 WBL_14 WWL_22 a_8342_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2885 GND a_14049_6766# a_13993_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2886 GND a_5349_2986# a_5293_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2887 a_16083_3818# a_15882_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2888 GND a_8342_4066# a_8249_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2889 a_14722_17# a_14629_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2890 RBL0_4 RWL_6 a_2743_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2891 GND a_7669_4066# a_7613_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2892 a_18403_4898# a_18202_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2893 a_9703_1118# a_9502_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2894 a_1003_3008# a_802_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2895 a_18202_287# a_18109_287# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2896 a_18053_8138# RWL_1 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2897 WBL_6 WWL_29 a_3702_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2898 a_14629_7576# WWL_3 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2899 a_129_4066# WWL_16 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2900 RBL0_24 RWL_0 a_14343_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2901 VDD a_2542_5146# a_2449_5146# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2902 GND a_709_2716# a_653_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2903 WBL_29 WWL_20 a_17042_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2904 RBL0_23 RWL_4 a_13763_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2905 GND a_4862_2446# a_4769_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2906 a_9409_17# WWL_31 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2907 a_2973_4898# RWL_13 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2908 VDD a_4862_6226# a_4769_6226# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2909 a_14573_6518# RWL_7 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2910 VDD a_16462_7846# a_16369_7846# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2911 GND a_18109_1366# a_18053_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2912 WBL_23 WWL_26 a_13562_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2913 a_8543_309# a_8342_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2914 a_16893_7598# a_13963_7576# RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2915 a_1962_5956# a_1869_5956# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2916 a_9502_5416# a_9409_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2917 a_12023_309# a_11822_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2918 a_802_7306# a_709_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2919 a_4282_3256# a_4189_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2920 a_2542_286# a_2449_286# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2921 RBL0_11 RWL_26 a_6803_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2922 WBL_7 WWL_3 a_4282_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2923 a_4282_7036# a_4189_7036# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2924 GND a_1289_8116# a_1233_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2925 a_11443_7868# a_11242_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2926 a_14049_1096# WWL_27 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2927 VDD a_15302_3526# a_15209_3526# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2928 RBL0_31 RWL_20 a_18403_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2929 a_6022_3796# a_5929_3796# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2930 GND a_6022_5956# a_5929_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2931 WBL_22 WWL_1 a_12982_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2932 GND a_5349_5956# a_5293_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2933 a_4133_308# RWL_30 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2934 a_15789_1636# WWL_25 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2935 a_73_38# RWL_31 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2936 a_11822_5956# a_11729_5956# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2937 a_1003_5978# a_802_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2938 a_9353_7328# RWL_4 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2939 GND a_11822_8116# a_11729_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2940 a_5929_6766# WWL_6 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2941 a_4133_5168# RWL_12 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2942 RBL0_13 RWL_13 a_7963_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2943 a_2542_8386# a_2449_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2944 a_1289_5686# WWL_10 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2945 WBL_14 WWL_23 a_8342_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2946 a_16083_3548# a_15882_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2947 RBL0_3 RWL_30 a_2163_308# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2948 a_11242_2716# a_11149_2716# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2949 a_14343_848# a_14142_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2950 a_18202_17# a_18109_17# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2951 a_5873_5708# RWL_10 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2952 GND a_2542_1096# a_2449_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2953 WBL_6 WWL_30 a_3702_286# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2954 GND a_11242_4876# a_11149_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2955 a_15209_8386# WWL_0 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2956 RBL0_24 RWL_1 a_14343_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2957 a_14629_7306# WWL_4 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2958 RBL0_23 RWL_5 a_13763_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2959 a_12603_1928# a_12402_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2960 GND a_709_2446# a_653_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2961 GND a_10569_4876# a_10513_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2962 VDD a_2542_4876# a_2449_4876# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2963 GND a_1869_1096# a_1813_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2964 GND a_4862_2176# a_4769_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2965 a_14573_6248# RWL_8 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2966 RBL0_31 RWL_9 a_18403_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2967 VDD a_6602_2716# a_6509_2716# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2968 VDD a_7182_3796# a_7089_3796# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2969 WBL_23 WWL_27 a_13562_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2970 a_7182_7846# a_7089_7846# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2971 a_9502_5146# a_9409_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2972 a_802_7036# a_709_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2973 a_16949_287# WWL_30 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2974 WBL_7 WWL_4 a_4282_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2975 a_11443_7598# a_11242_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2976 VDD a_12982_5956# a_12889_5956# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2977 a_6022_3526# a_5929_3526# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2978 GND a_3029_4606# a_2973_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2979 a_7383_2738# a_7182_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2980 a_15789_1366# WWL_26 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2981 RBL0_25 RWL_27 a_14923_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2982 VDD a_11822_1636# a_11729_1636# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2983 a_12402_2986# a_12309_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2984 a_9353_7058# RWL_5 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2985 a_6509_7576# WWL_3 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2986 a_5929_6496# WWL_7 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2987 a_2542_8116# a_2449_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2988 RBL0_9 RWL_4 a_5643_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2989 a_1289_5416# WWL_11 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2990 WBL_14 WWL_24 a_8342_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2991 a_16083_3278# a_15882_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2992 GND a_14142_5686# a_14049_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2993 a_16462_4606# a_16369_4606# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2994 GND a_16462_6766# a_16369_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2995 GND a_13469_5686# a_13413_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2996 a_14343_578# a_14142_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2997 RBL0_3 RWL_24 a_2163_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2998 a_5873_5438# RWL_11 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2999 WBL_6 WWL_31 a_3702_16# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3000 GND a_7762_2986# a_7669_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3001 a_15209_8116# WWL_1 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3002 GND a_15789_6766# a_15733_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3003 a_17823_3818# a_17622_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3004 a_1962_4876# a_1869_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3005 a_13763_39# a_13562_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3006 GND a_709_2176# a_653_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3007 a_12603_1658# a_12402_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3008 RBL0_27 RWL_14 a_16083_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3009 VDD a_7182_556# a_7089_556# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3010 a_3323_7868# a_3122_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3011 a_2743_6788# a_2542_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3012 VDD a_7182_3526# a_7089_3526# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3013 WBL_3 WWL_9 a_1962_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3014 a_14343_8408# a_14142_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3015 a_16949_17# WWL_31 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3016 VDD a_18202_4066# a_18109_4066# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3017 a_12402_5956# a_12309_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3018 GND a_222_8386# a_129_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3019 a_11822_4876# a_11729_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3020 GND a_8249_6496# a_8193_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3021 a_3702_5956# a_3609_5956# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3022 WBL_10 WWL_17 a_6022_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3023 GND a_3029_4336# a_2973_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3024 a_4862_556# a_4769_556# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3025 VDD a_10082_1366# a_9989_1366# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3026 VDD a_14722_2446# a_14629_2446# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3027 a_7383_2468# a_7182_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3028 a_15789_1096# WWL_27 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3029 a_7762_3796# a_7669_3796# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3030 a_2542_1636# a_2449_1636# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3031 WBL_21 WWL_5 a_12402_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3032 GND a_7762_5956# a_7669_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3033 RBL0_16 RWL_28 a_9703_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3034 a_6509_7306# WWL_4 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3035 RBL0_9 RWL_5 a_5643_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3036 a_5929_6226# WWL_8 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3037 a_14142_3256# a_14049_3256# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3038 GND a_14142_5416# a_14049_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3039 a_12253_7868# RWL_2 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3040 a_16462_4336# a_16369_4336# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3041 a_17529_7846# WWL_2 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3042 WBL_19 WWL_21 a_11242_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3043 RBL0_12 RWL_17 a_7383_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3044 GND a_13469_5416# a_13413_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3045 RBL0_3 RWL_25 a_2163_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3046 a_7182_6766# a_7089_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3047 a_5873_5168# RWL_12 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3048 RBL0_16 RWL_13 a_9703_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3049 a_17823_3548# a_17622_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3050 a_12603_1388# a_12402_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3051 GND a_10662_3796# a_10569_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3052 VDD a_9502_3256# a_9409_3256# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3053 VDD a_10662_7576# a_10569_7576# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3054 VDD a_802_5146# a_709_5146# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3055 RBL0_27 RWL_15 a_16083_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3056 a_7762_287# a_7669_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3057 GND a_12982_4876# a_12889_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3058 a_3323_7598# a_3122_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3059 WBL_12 WWL_2 a_7182_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3060 a_14343_8138# a_14142_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3061 a_14722_5686# a_14629_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3062 RBL0_21 RWL_21 a_12603_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3063 a_10082_4606# a_9989_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3064 a_8922_4066# a_8829_4066# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3065 a_10082_8386# a_9989_8386# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3066 a_222_5956# a_129_5956# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3067 GND a_222_8116# a_129_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3068 a_9353_309# RWL_30 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3069 RBL0_5 RWL_31 a_3323_38# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3070 a_802_286# a_709_286# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3071 WBL_10 WWL_18 a_6022_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3072 GND a_8249_6226# a_8193_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3073 a_13413_1928# RWL_24 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3074 a_5063_1118# a_4862_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3075 GND a_3029_4066# a_2973_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3076 a_10863_6518# a_10662_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3077 VDD a_10082_1096# a_9989_1096# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3078 VDD a_14722_2176# a_14629_2176# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3079 a_5442_2446# a_5349_2446# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3080 a_7383_2198# a_7182_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3081 GND a_5442_4606# a_5349_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3082 a_8829_7036# WWL_5 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3083 a_7762_3526# a_7669_3526# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3084 VDD a_5442_8386# a_5349_8386# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3085 a_4189_5956# WWL_9 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3086 RBL0_12 RWL_30 a_7383_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3087 RBL0_16 RWL_29 a_9703_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3088 GND a_4769_4606# a_4713_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3089 a_11443_39# a_11242_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3090 a_14142_2986# a_14049_2986# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3091 a_13562_826# a_13469_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3092 GND a_7089_287# a_7033_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3093 GND a_14142_5146# a_14049_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3094 a_12253_7598# a_4683_7576# RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3095 a_8249_3796# WWL_17 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3096 WBL_28 WWL_14 a_16462_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3097 VDD a_1962_6766# a_1869_6766# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3098 RBL0_12 RWL_18 a_7383_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3099 GND a_13469_5146# a_13413_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3100 RBL0_3 RWL_26 a_2163_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3101 RBL0_0 RWL_30 a_423_308# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3102 a_10662_1366# a_10569_1366# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3103 a_17823_3278# a_17622_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3104 GND a_15882_5686# a_15789_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3105 GND a_15209_1906# a_15153_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3106 GND a_802_1096# a_709_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3107 a_8193_2738# RWL_21 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3108 GND a_10662_3526# a_10569_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3109 a_6223_8408# a_6022_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3110 a_5643_7328# a_5442_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3111 a_15153_848# RWL_28 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3112 RBL0_0 RWL_31 a_423_38# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3113 RBL0_6 RWL_24 a_3903_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3114 VDD a_9502_2986# a_9409_2986# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3115 a_1382_3796# a_1289_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3116 RBL0_27 RWL_16 a_16083_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3117 VDD a_802_4876# a_709_4876# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3118 VDD a_10662_7306# a_10569_7306# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3119 a_1382_7576# a_1289_7576# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3120 a_3702_4876# a_3609_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3121 a_11149_1636# WWL_25 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3122 a_15302_6496# a_15209_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3123 VDD a_222_1636# a_129_1636# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3124 a_13469_2716# WWL_21 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3125 RBL0_30 RWL_14 a_17823_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3126 a_14722_5416# a_14629_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3127 RBL0_21 RWL_22 a_12603_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3128 a_10082_4336# a_9989_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3129 RBL0_22 RWL_28 a_13183_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3130 WBL_15 WWL_15 a_8922_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3131 a_10082_8116# a_9989_8116# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3132 VDD a_14722_556# a_14629_556# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3133 WBL_6 WWL_9 a_3702_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3134 a_13413_1658# RWL_25 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3135 a_10863_6248# a_10662_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3136 VDD a_14722_1906# a_14629_1906# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3137 a_1233_5708# RWL_10 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3138 a_5442_2176# a_5349_2176# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3139 GND a_5442_4336# a_5349_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3140 a_9409_7846# WWL_2 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3141 a_3553_6788# RWL_6 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3142 WBL_13 WWL_17 a_7762_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3143 VDD a_5442_8116# a_5349_8116# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3144 GND a_9989_6496# a_9933_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3145 GND a_4769_4336# a_4713_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3146 a_15153_8408# RWL_0 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3147 a_11242_287# a_11149_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3148 WBL_24 WWL_19 a_14142_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3149 a_13562_556# a_13469_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3150 GND a_1962_2716# a_1869_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3151 a_8249_3526# WWL_18 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3152 VDD a_1962_6496# a_1869_6496# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3153 RBL0_12 RWL_19 a_7383_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3154 a_15882_3256# a_15789_3256# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3155 a_10662_1096# a_10569_1096# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3156 GND a_15882_5416# a_15789_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3157 GND a_17622_287# a_17529_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3158 GND a_15209_1636# a_15153_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3159 WBL_18 WWL_25 a_10662_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3160 a_13993_7868# RWL_2 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3161 a_8193_2468# RWL_22 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3162 a_6223_8138# a_6022_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3163 a_6602_5686# a_6509_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3164 GND a_10662_3256# a_10569_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3165 a_222_4876# a_129_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3166 a_5643_7058# a_5442_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3167 a_15153_578# RWL_29 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3168 RBL0_6 RWL_25 a_3903_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3169 a_1382_3526# a_1289_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3170 VDD a_10662_7036# a_10569_7036# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3171 GND a_16949_826# a_16893_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3172 a_1382_7306# a_1289_7306# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3173 RBL0_1 RWL_31 a_1003_38# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3174 a_11149_1366# WWL_26 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3175 VDD a_12402_3796# a_12309_3796# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3176 RBL0_17 RWL_27 a_10283_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3177 a_15302_6226# a_15209_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3178 a_14722_5146# a_14629_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3179 a_10082_4066# a_9989_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3180 RBL0_30 RWL_15 a_17823_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3181 RBL0_21 RWL_23 a_12603_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3182 RBL0_22 RWL_29 a_13183_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3183 WBL_15 WWL_16 a_8922_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3184 WBL_17 WWL_0 a_10082_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3185 RBL0_1 RWL_4 a_1003_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3186 WBL_0 WWL_9 a_222_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3187 WBL_15 WWL_30 a_8922_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3188 WBL_21 WWL_30 a_12402_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3189 a_17042_6766# a_16949_6766# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3190 a_13413_1388# RWL_26 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3191 GND a_3122_2986# a_3029_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3192 a_1233_5438# RWL_11 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3193 a_5442_1906# a_5349_1906# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3194 WBL_9 WWL_22 a_5442_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3195 GND a_11149_6766# a_11093_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3196 GND a_2449_2986# a_2393_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3197 a_13183_3818# a_12982_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3198 GND a_5442_4066# a_5349_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3199 WBL_13 WWL_18 a_7762_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3200 GND a_9989_6226# a_9933_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3201 GND a_4769_4066# a_4713_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3202 a_15503_4898# a_15302_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3203 a_6803_1118# a_6602_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3204 a_15153_8138# RWL_1 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3205 a_11729_7576# WWL_3 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3206 GND a_7089_1906# a_7033_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3207 RBL0_19 RWL_0 a_11443_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3208 RBL0_18 RWL_4 a_10863_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3209 WBL_24 WWL_20 a_14142_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3210 GND a_1962_2446# a_1869_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3211 VDD a_1962_6226# a_1869_6226# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3212 a_11673_6518# RWL_7 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3213 a_15882_2986# a_15789_2986# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3214 VDD a_13562_7846# a_13469_7846# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3215 GND a_15209_1366# a_15153_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3216 WBL_18 WWL_26 a_10662_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3217 a_13993_7598# a_13963_7576# RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3218 GND a_15882_5146# a_15789_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3219 a_8193_2198# RWL_23 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3220 a_9989_3796# WWL_17 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3221 a_6602_5416# a_6509_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3222 GND a_14629_287# a_14573_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3223 RBL0_6 RWL_26 a_3903_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3224 a_1382_3256# a_1289_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3225 GND a_16949_556# a_16893_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3226 GND a_17622_1906# a_17529_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3227 WBL_2 WWL_3 a_1382_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3228 a_1382_7036# a_1289_7036# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3229 VDD a_17622_5686# a_17529_5686# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3230 a_16369_3256# WWL_19 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3231 a_11149_1096# WWL_27 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3232 GND a_16949_1906# a_16893_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3233 VDD a_12402_3526# a_12309_3526# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3234 a_17823_848# a_17622_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3235 RBL0_26 RWL_20 a_15503_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3236 a_3122_3796# a_3029_3796# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3237 GND a_3122_5956# a_3029_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3238 RBL0_30 RWL_16 a_17823_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3239 WBL_17 WWL_1 a_10082_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3240 GND a_2449_5956# a_2393_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3241 WBL_15 WWL_31 a_8922_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3242 RBL0_1 RWL_5 a_1003_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3243 a_15733_1118# RWL_27 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3244 a_12889_1636# WWL_25 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3245 a_17042_2716# a_16949_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3246 WBL_21 WWL_31 a_12402_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3247 a_17042_6496# a_16949_6496# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3248 a_2542_16# a_2449_16# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3249 a_6453_7328# RWL_4 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3250 a_1233_5168# RWL_12 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3251 WBL_9 WWL_23 a_5442_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3252 RBL0_8 RWL_13 a_5063_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3253 a_18403_5708# a_18202_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3254 a_13183_3548# a_12982_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3255 a_2163_848# a_1962_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3256 a_2973_5708# RWL_10 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3257 a_12309_8386# WWL_0 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3258 a_11729_7306# WWL_4 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3259 GND a_7089_1636# a_7033_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3260 RBL0_19 RWL_1 a_11443_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3261 RBL0_18 RWL_5 a_10863_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3262 a_3903_38# a_3702_16# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3263 GND a_1962_2176# a_1869_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3264 WBL_12 WWL_29 a_7182_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3265 a_16893_8408# RWL_0 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3266 a_11673_6248# RWL_8 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3267 a_7669_2446# WWL_22 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3268 a_12982_7846# a_12889_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3269 RBL0_26 RWL_9 a_15503_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3270 VDD a_3702_2716# a_3609_2716# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3271 VDD a_4282_3796# a_4189_3796# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3272 WBL_18 WWL_27 a_10662_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3273 a_4282_7846# a_4189_7846# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3274 a_15882_826# a_15789_826# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3275 a_9989_3526# WWL_18 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3276 a_6602_5146# a_6509_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3277 a_4769_287# WWL_30 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3278 GND a_17622_1636# a_17529_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3279 WBL_2 WWL_4 a_1382_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3280 VDD a_17622_5416# a_17529_5416# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3281 a_8342_1906# a_8249_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3282 a_16369_2986# WWL_20 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3283 a_15503_309# a_15302_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3284 GND a_16949_1636# a_16893_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3285 a_8342_5686# a_8249_5686# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3286 a_17823_578# a_17622_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3287 a_3122_3526# a_3029_3526# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3288 GND a_8342_7846# a_8249_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3289 GND a_7669_7846# a_7613_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3290 a_17042_2446# a_16949_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3291 a_4483_2738# a_4282_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3292 a_12889_1366# WWL_26 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3293 a_17042_6226# a_16949_6226# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3294 WBL_29 WWL_6 a_17042_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3295 RBL0_13 RWL_10 a_7963_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3296 a_1003_38# a_802_16# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3297 WBL_20 WWL_14 a_11822_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3298 GND a_14049_7306# a_13993_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3299 a_6453_7058# RWL_5 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3300 a_3609_7576# WWL_3 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3301 RBL0_4 RWL_4 a_2743_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3302 a_18403_5438# a_18202_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3303 WBL_9 WWL_24 a_5442_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3304 a_13183_3278# a_12982_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3305 GND a_11242_5686# a_11149_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3306 a_13562_4606# a_13469_4606# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3307 a_2163_578# a_1962_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3308 GND a_13562_6766# a_13469_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3309 GND a_10569_5686# a_10513_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3310 VDD a_6602_826# a_6509_826# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3311 GND a_4862_2986# a_4769_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3312 a_2973_5438# RWL_11 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3313 a_12309_8116# WWL_1 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3314 GND a_12889_6766# a_12833_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3315 GND a_7089_1366# a_7033_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3316 a_14923_3818# a_14722_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3317 a_10569_826# WWL_28 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3318 a_7613_39# RWL_31 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3319 RBL0_22 RWL_14 a_13183_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3320 a_16893_8138# RWL_1 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3321 a_7669_2176# WWL_23 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3322 VDD a_8922_4606# a_8829_4606# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3323 a_12982_7576# a_12889_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3324 a_13562_287# a_13469_287# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3325 VDD a_4282_3526# a_4189_3526# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3326 a_11443_8408# a_11242_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3327 VDD a_15302_4066# a_15209_4066# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3328 a_4769_17# WWL_31 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3329 GND a_17622_1366# a_17529_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3330 a_7613_1118# RWL_27 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3331 a_16313_4898# RWL_13 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3332 a_8342_1636# a_8249_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3333 GND a_6022_6496# a_5929_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3334 a_8342_5416# a_8249_5416# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3335 GND a_16949_1366# a_16893_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3336 GND a_8342_7576# a_8249_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3337 GND a_5349_6496# a_5293_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3338 WBL_5 WWL_17 a_3122_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3339 VDD a_11822_2446# a_11729_2446# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3340 GND a_7669_7576# a_7613_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3341 a_9703_4628# a_9502_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3342 a_1003_6518# a_802_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3343 a_17042_2176# a_16949_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3344 a_4483_2468# a_4282_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3345 a_12889_1096# WWL_27 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3346 a_4862_3796# a_4769_3796# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3347 a_129_7576# WWL_3 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3348 WBL_29 WWL_7 a_17042_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3349 RBL0_13 RWL_11 a_7963_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3350 a_18053_39# RWL_31 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3351 GND a_14049_7036# a_13993_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3352 GND a_4862_5956# a_4769_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3353 a_3609_7306# WWL_4 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3354 RBL0_4 RWL_5 a_2743_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3355 a_18403_5168# a_18202_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3356 a_1583_38# a_1382_16# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3357 a_11242_3256# a_11149_3256# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3358 GND a_11242_5416# a_11149_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3359 a_14629_7846# WWL_2 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3360 a_1962_5686# a_1869_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3361 a_13562_4336# a_13469_4336# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3362 GND a_18109_4876# a_18053_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3363 GND a_9409_1096# a_9353_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3364 RBL0_7 RWL_17 a_4483_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3365 GND a_10569_5416# a_10513_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3366 GND a_709_2986# a_653_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3367 a_2973_5168# RWL_12 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3368 a_4282_6766# a_4189_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3369 RBL0_11 RWL_13 a_6803_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3370 a_14923_3548# a_14722_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3371 a_802_1366# a_709_1366# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3372 RBL0_31 RWL_7 a_18403_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3373 VDD a_6602_3256# a_6509_3256# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3374 a_14049_4606# WWL_14 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3375 RBL0_22 RWL_15 a_13183_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3376 a_7669_1906# WWL_24 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3377 VDD a_8922_4336# a_8829_4336# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3378 a_13562_17# a_13469_17# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3379 WBL_7 WWL_2 a_4282_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3380 a_11443_8138# a_11242_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3381 a_11822_5686# a_11729_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3382 a_6022_4066# a_5929_4066# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3383 WBL_25 WWL_29 a_14722_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3384 a_8342_1366# a_8249_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3385 GND a_6022_6226# a_5929_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3386 WBL_14 WWL_10 a_8342_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3387 WBL_5 WWL_18 a_3122_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3388 GND a_5349_6226# a_5293_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3389 a_10513_1928# RWL_24 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3390 a_2163_1118# a_1962_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3391 a_12402_17# a_12309_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3392 VDD a_11822_2176# a_11729_2176# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3393 a_2542_2446# a_2449_2446# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3394 a_9703_4358# a_9502_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3395 a_1003_6248# a_802_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3396 a_4483_2198# a_4282_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3397 GND a_2542_4606# a_2449_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3398 a_129_7306# WWL_4 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3399 a_5929_7036# WWL_5 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3400 WBL_29 WWL_8 a_17042_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3401 a_8342_556# a_8249_556# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3402 a_4862_3526# a_4769_3526# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3403 VDD a_2542_8386# a_2449_8386# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3404 a_1289_5956# WWL_9 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3405 GND a_709_5956# a_653_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3406 RBL0_13 RWL_12 a_7963_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3407 GND a_1869_4606# a_1813_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3408 a_16462_5146# a_16369_5146# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3409 a_1382_826# a_1289_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3410 a_11242_2986# a_11149_2986# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3411 GND a_16462_7306# a_16369_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3412 GND a_11242_5146# a_11149_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3413 a_5349_3796# WWL_17 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3414 RBL0_16 RWL_10 a_9703_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3415 a_5293_39# RWL_31 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3416 WBL_23 WWL_14 a_13562_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3417 GND a_15789_7306# a_15733_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3418 a_1962_5416# a_1869_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3419 RBL0_7 RWL_18 a_4483_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3420 GND a_10569_5146# a_10513_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3421 GND a_3702_16# a_3609_16# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3422 GND a_12309_1906# a_12253_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3423 a_14923_3278# a_14722_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3424 GND a_12982_5686# a_12889_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3425 a_423_848# a_222_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3426 GND a_7762_826# a_7669_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3427 a_5293_2738# RWL_21 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3428 a_9933_3818# RWL_17 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3429 a_802_1096# a_709_1096# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3430 WBL_1 WWL_25 a_802_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3431 a_3323_8408# a_3122_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3432 a_2743_7328# a_2542_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3433 RBL0_31 RWL_8 a_18403_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3434 VDD a_6602_2986# a_6509_2986# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3435 VDD a_7182_4066# a_7089_4066# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3436 RBL0_22 RWL_16 a_13183_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3437 a_12402_6496# a_12309_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3438 RBL0_0 RWL_27 a_423_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3439 a_10569_2716# WWL_21 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3440 RBL0_25 RWL_14 a_14923_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3441 a_11822_5416# a_11729_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3442 RBL0_1 RWL_28 a_1003_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3443 WBL_10 WWL_15 a_6022_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3444 VDD a_2542_556# a_2449_556# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3445 WBL_14 WWL_11 a_8342_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3446 a_3029_556# WWL_29 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3447 a_16083_6788# a_15882_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3448 a_10513_1658# RWL_25 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3449 a_7383_3008# a_7182_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3450 VDD a_11822_1906# a_11729_1906# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3451 a_9703_4088# a_9502_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3452 GND a_802_16# a_709_16# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3453 a_16313_309# RWL_30 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3454 a_2542_2176# a_2449_2176# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3455 GND a_7762_6496# a_7669_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3456 GND a_2542_4336# a_2449_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3457 a_6509_7846# WWL_2 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3458 VDD a_2542_8116# a_2449_8116# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3459 GND a_1869_4336# a_1813_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3460 a_16462_1096# a_16369_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3461 a_12253_8408# RWL_0 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3462 a_3029_2446# WWL_22 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3463 a_16462_4876# a_16369_4876# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3464 WBL_19 WWL_19 a_11242_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3465 GND a_16462_7036# a_16369_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3466 a_1382_556# a_1289_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3467 RBL0_24 RWL_30 a_14343_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3468 a_7182_7306# a_7089_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3469 RBL0_16 RWL_11 a_9703_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3470 a_5349_3526# WWL_18 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3471 GND a_15789_7036# a_15733_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3472 a_1962_5146# a_1869_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3473 RBL0_7 RWL_19 a_4483_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3474 GND a_18202_3796# a_18109_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3475 a_17042_826# a_16949_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3476 VDD a_18202_7576# a_18109_7576# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3477 GND a_5442_287# a_5349_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3478 GND a_17529_3796# a_17473_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3479 GND a_12982_5416# a_12889_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3480 GND a_12309_1636# a_12253_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3481 a_9933_3548# RWL_18 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3482 a_423_578# a_222_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3483 GND a_7762_556# a_7669_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3484 GND a_15882_17# a_15789_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3485 a_5293_2468# RWL_22 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3486 a_3323_8138# a_3122_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3487 a_2743_7058# a_2542_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3488 a_3702_5686# a_3609_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3489 WBL_1 WWL_26 a_802_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3490 GND a_4769_826# a_4713_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3491 GND a_3029_7846# a_2973_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3492 VDD a_222_2446# a_129_2446# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3493 a_7383_5978# a_7182_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3494 a_15789_4606# WWL_14 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3495 a_12402_6226# a_12309_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3496 RBL0_25 RWL_15 a_14923_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3497 a_11822_5146# a_11729_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3498 a_10082_17# a_9989_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3499 RBL0_1 RWL_29 a_1003_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3500 WBL_10 WWL_16 a_6022_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3501 VDD a_2542_286# a_2449_286# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3502 a_14142_6766# a_14049_6766# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3503 a_3029_286# WWL_30 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3504 a_10513_1388# RWL_26 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3505 VDD a_18202_556# a_18109_556# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3506 a_7762_4066# a_7669_4066# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3507 a_2542_1906# a_2449_1906# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3508 WBL_4 WWL_22 a_2542_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3509 GND a_7762_6226# a_7669_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3510 WBL_31 WWL_28 a_18202_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3511 a_10283_3818# a_10082_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3512 GND a_2542_4066# a_2449_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3513 GND a_11242_826# a_11149_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3514 GND a_1869_4066# a_1813_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3515 a_12603_4898# a_12402_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3516 a_3903_1118# a_3702_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3517 VDD a_9502_6766# a_9409_6766# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3519 a_12253_8138# RWL_1 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3520 RBL0_27 RWL_2 a_16083_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3521 WBL_28 WWL_12 a_16462_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3522 a_8249_4336# WWL_15 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3523 GND a_4189_1906# a_4133_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3524 a_3029_2176# WWL_23 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3525 WBL_19 WWL_20 a_11242_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3526 a_7182_7036# a_7089_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3527 RBL0_16 RWL_12 a_9703_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3528 GND a_18202_3526# a_18109_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3529 a_17042_556# a_16949_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3530 a_8922_3796# a_8829_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3531 VDD a_18202_7306# a_18109_7306# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3532 a_222_5686# a_129_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3533 VDD a_10662_7846# a_10569_7846# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3534 a_8922_7576# a_8829_7576# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3535 GND a_17529_3526# a_17473_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3536 GND a_12982_5146# a_12889_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3537 GND a_12309_1366# a_12253_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3538 a_9933_3278# RWL_19 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3539 a_5293_2198# RWL_23 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3540 a_3702_5416# a_3609_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3542 WBL_1 WWL_27 a_802_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3543 GND a_4769_556# a_4713_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3544 GND a_14722_1906# a_14629_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3545 GND a_3029_7576# a_2973_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3546 a_5063_4628# a_4862_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3547 VDD a_14722_5686# a_14629_5686# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3548 VDD a_222_2176# a_129_2176# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3549 a_13469_3256# WWL_19 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3550 RBL0_21 RWL_20 a_12603_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3551 VDD a_10082_4606# a_9989_4606# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3552 RBL0_25 RWL_16 a_14923_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3553 RBL0_29 RWL_24 a_17243_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3554 a_12833_1118# RWL_27 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3555 VDD a_2542_16# a_2449_16# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3556 a_14142_2716# a_14049_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3557 a_14142_6496# a_14049_6496# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3558 a_3029_16# WWL_31 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3559 a_3553_7328# RWL_4 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3560 WBL_27 WWL_30 a_15882_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3561 WBL_13 WWL_15 a_7762_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3562 WBL_4 WWL_23 a_2542_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3563 RBL0_3 RWL_13 a_2163_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3564 a_15503_5708# a_15302_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3565 a_10283_3548# a_10082_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3566 a_17823_6788# a_17622_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3567 GND a_11242_556# a_11149_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3568 GND a_9502_2716# a_9409_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3569 GND a_802_4606# a_709_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3570 VDD a_802_8386# a_709_8386# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3571 RBL0_27 a_13963_7576# a_16083_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3572 VDD a_9502_6496# a_9409_6496# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3573 a_8249_4066# WWL_16 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3574 GND a_4189_1636# a_4133_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3575 a_3029_1906# WWL_24 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3576 GND a_8829_2716# a_8773_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3577 WBL_28 WWL_13 a_16462_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3578 GND a_13562_17# a_13469_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3579 GND a_18202_3256# a_18109_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3580 a_13993_8408# RWL_0 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3581 a_8193_3008# RWL_20 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3582 a_8922_3526# a_8829_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3583 a_10082_7846# a_9989_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3584 VDD a_18202_7036# a_18109_7036# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3585 a_222_5416# a_129_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3586 a_4769_2446# WWL_22 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3587 VDD a_1382_3796# a_1289_3796# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3588 RBL0_21 RWL_9 a_12603_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3589 GND a_17529_3256# a_17473_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3590 a_8922_7306# a_8829_7306# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3591 a_3702_826# a_3609_826# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3592 a_1382_7846# a_1289_7846# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3593 a_3702_5146# a_3609_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3594 GND a_14722_1636# a_14629_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3595 VDD a_14722_5416# a_14629_5416# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3596 a_5442_1906# a_5349_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3597 VDD a_222_1906# a_129_1906# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3598 a_13469_2986# WWL_20 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3599 a_5063_4358# a_4862_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3600 GND a_18109_287# a_18053_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3601 VDD a_10082_4336# a_9989_4336# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3602 a_5442_5686# a_5349_5686# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3603 GND a_5442_7846# a_5349_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3604 GND a_4769_7846# a_4713_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3605 RBL0_29 RWL_25 a_17243_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3606 a_14142_2446# a_14049_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3607 a_1583_2738# a_1382_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3608 a_14142_6226# a_14049_6226# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3609 WBL_24 WWL_6 a_14142_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3610 RBL0_8 RWL_10 a_5063_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3611 GND a_11149_7306# a_11093_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3612 a_3553_7058# RWL_5 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3613 RBL0_12 RWL_6 a_7383_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3614 WBL_27 WWL_31 a_15882_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3615 WBL_13 WWL_16 a_7762_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3616 a_15503_5438# a_15302_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3617 WBL_4 WWL_24 a_2542_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3618 a_10283_3278# a_10082_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3619 a_15882_6766# a_15789_6766# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3620 a_10662_4606# a_10569_4606# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3621 a_8193_5978# RWL_9 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3622 GND a_9502_2446# a_9409_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3623 GND a_802_4336# a_709_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3624 GND a_10662_6766# a_10569_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3626 GND a_1962_2986# a_1869_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3627 VDD a_9502_6226# a_9409_6226# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3628 VDD a_802_8116# a_709_8116# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3629 GND a_4189_1366# a_4133_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3630 GND a_8829_2446# a_8773_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3631 a_12023_3818# a_11822_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3632 RBL0_17 RWL_14 a_10283_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3633 a_13993_8138# RWL_1 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3634 a_9989_4336# WWL_15 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3635 RBL0_30 RWL_2 a_17823_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3636 a_222_5146# a_129_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3637 a_4769_2176# WWL_23 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3638 a_8922_3256# a_8829_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3639 a_10082_7576# a_9989_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3640 VDD a_1382_3526# a_1289_3526# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3641 WBL_15 WWL_3 a_8922_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3642 a_8922_7036# a_8829_7036# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3643 a_11093_3818# RWL_17 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3644 VDD a_12402_4066# a_12309_4066# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3645 GND a_14722_1366# a_14629_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3646 a_13413_4898# RWL_13 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3647 a_4713_1118# RWL_27 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3648 a_2973_308# RWL_30 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3649 a_5442_1636# a_5349_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3650 a_5063_4088# a_4862_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3651 GND a_3122_6496# a_3029_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3652 a_5442_5416# a_5349_5416# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3653 VDD a_7762_287# a_7669_287# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3654 a_8249_287# WWL_30 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3655 GND a_5442_7576# a_5349_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3656 GND a_2449_6496# a_2393_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3657 GND a_4769_7576# a_4713_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3658 a_6803_4628# a_6602_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3659 RBL0_29 RWL_26 a_17243_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3660 a_14142_2176# a_14049_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3661 a_1583_2468# a_1382_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3662 WBL_24 WWL_7 a_14142_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3663 RBL0_8 RWL_11 a_5063_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3664 GND a_1962_5956# a_1869_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3665 GND a_11149_7036# a_11093_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3666 RBL0_15 RWL_31 a_9123_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3667 a_15503_5168# a_15302_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3668 a_15882_2716# a_15789_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3669 GND a_11242_17# a_11149_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3670 a_15882_6496# a_15789_6496# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3671 a_11729_7846# WWL_2 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3672 RBL0_2 RWL_17 a_1583_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3673 a_10662_4336# a_10569_4336# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3674 GND a_15209_4876# a_15153_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3675 GND a_6509_1096# a_6453_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3676 a_17243_1928# a_17042_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3677 GND a_9502_2176# a_9409_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3678 GND a_802_4066# a_709_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3679 a_1382_6766# a_1289_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3680 GND a_8829_2176# a_8773_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3681 RBL0_6 RWL_13 a_3903_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3682 a_12023_3548# a_11822_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3683 a_16369_6766# WWL_6 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3684 a_12982_8386# a_12889_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3685 RBL0_26 RWL_7 a_15503_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3686 VDD a_3702_3256# a_3609_3256# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3687 a_11149_4606# WWL_14 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3688 VDD a_13562_826# a_13469_826# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3689 RBL0_17 RWL_15 a_10283_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3690 a_14049_826# WWL_28 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3691 a_9989_4066# WWL_16 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3692 RBL0_30 a_13963_7576# a_17823_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3693 a_4769_1906# WWL_24 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3694 WBL_15 WWL_4 a_8922_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3695 a_16313_5708# RWL_10 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3696 WBL_2 WWL_2 a_1382_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3697 a_11093_3548# RWL_18 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3698 a_15733_4628# RWL_14 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3699 VDD a_17622_5956# a_17529_5956# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3700 a_17042_287# a_16949_287# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3701 WBL_4 WWL_29 a_2542_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3702 a_709_2716# WWL_21 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3703 a_3122_4066# a_3029_4066# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3704 GND a_8342_8386# a_8249_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3705 a_5442_1366# a_5349_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3706 GND a_3122_6226# a_3029_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3707 VDD a_7762_17# a_7669_17# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3708 GND a_7669_8386# a_7613_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3709 WBL_9 WWL_10 a_5442_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3710 a_8249_17# WWL_31 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3711 GND a_2449_6226# a_2393_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3712 VDD a_17042_2716# a_16949_2716# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3713 a_17042_2986# a_16949_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3714 a_6803_4358# a_6602_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3715 WBL_20 WWL_12 a_11822_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3716 a_1583_2198# a_1382_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3717 WBL_24 WWL_8 a_14142_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3718 RBL0_8 RWL_12 a_5063_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3719 a_10863_309# a_10662_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3720 GND a_18109_5686# a_18053_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3721 a_13562_5146# a_13469_5146# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3722 a_15882_2446# a_15789_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3723 GND a_13562_7306# a_13469_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3724 a_15882_6226# a_15789_6226# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3725 RBL0_11 RWL_10 a_6803_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3726 a_2449_3796# WWL_17 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3727 WBL_18 WWL_14 a_10662_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3728 GND a_12889_7306# a_12833_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3729 a_17243_1658# a_17042_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3730 RBL0_2 RWL_18 a_1583_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3731 a_6509_556# WWL_29 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3732 a_12023_3278# a_11822_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3733 a_2393_2738# RWL_21 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3734 a_16369_6496# WWL_7 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3735 VDD a_8922_5146# a_8829_5146# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3736 a_12982_8116# a_12889_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3737 RBL0_26 RWL_8 a_15503_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3738 VDD a_11242_287# a_11149_287# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3739 VDD a_3702_2986# a_3609_2986# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3740 VDD a_4282_4066# a_4189_4066# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3741 RBL0_17 RWL_16 a_10283_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3742 a_17042_5956# a_16949_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3743 a_16313_5438# RWL_11 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3744 a_15733_4358# RWL_15 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3745 a_11093_3278# RWL_19 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3746 a_8342_5956# a_8249_5956# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3747 a_17042_17# a_16949_17# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3748 WBL_4 WWL_30 a_2542_286# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3749 GND a_8342_8116# a_8249_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3750 WBL_5 WWL_15 a_3122_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3751 WBL_9 WWL_11 a_5442_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3752 GND a_7669_8116# a_7613_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3753 a_13183_6788# a_12982_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3754 a_4483_3008# a_4282_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3755 WBL_29 WWL_5 a_17042_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3756 a_6803_4088# a_6602_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3757 WBL_20 WWL_13 a_11822_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3758 GND a_4862_6496# a_4769_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3759 a_3609_7846# WWL_2 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3760 a_9123_1928# a_8922_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3761 GND a_7089_4876# a_7033_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3762 a_423_3818# a_222_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3763 a_13562_1096# a_13469_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3764 GND a_18109_5416# a_18053_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3765 a_13562_4876# a_13469_4876# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3766 a_15882_2176# a_15789_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3767 GND a_13562_7036# a_13469_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3768 a_7669_5686# WWL_10 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3769 GND a_3609_16# a_3553_38# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3770 a_15302_556# a_15209_556# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3771 a_4282_7306# a_4189_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3772 RBL0_11 RWL_11 a_6803_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3773 a_2449_3526# WWL_18 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3774 GND a_12889_7036# a_12833_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3775 a_17243_1388# a_17042_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3776 RBL0_2 RWL_19 a_1583_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3777 GND a_15302_3796# a_15209_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3778 a_17622_2716# a_17529_2716# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3779 a_18202_3796# a_18109_3796# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3780 a_12982_1636# a_12889_1636# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3781 VDD a_15302_7576# a_15209_7576# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3782 a_14049_5146# WWL_12 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3783 GND a_14629_3796# a_14573_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3784 GND a_8922_1096# a_8829_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3785 a_7613_4628# RWL_14 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3786 GND a_17622_4876# a_17529_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3787 a_16369_6226# WWL_8 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3788 a_2393_2468# RWL_22 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3789 VDD a_8922_4876# a_8829_4876# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3790 VDD a_11242_17# a_11149_17# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3791 GND a_16949_4876# a_16893_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3792 a_4483_5978# a_4282_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3793 a_16313_5168# RWL_12 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3794 a_15733_4088# RWL_16 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3795 VDD a_8342_1636# a_8249_1636# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3796 a_12889_4606# WWL_14 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3797 WBL_4 WWL_31 a_2542_16# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3798 a_18053_1928# RWL_24 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3799 WBL_5 WWL_16 a_3122_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3800 a_18202_287# a_18109_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3801 a_11242_6766# a_11149_6766# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3802 GND a_709_16# a_653_38# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3803 a_129_7846# WWL_2 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3804 VDD a_6022_556# a_5929_556# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3805 a_4862_4066# a_4769_4066# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3806 GND a_9409_4606# a_9353_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3807 GND a_709_6496# a_653_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3808 GND a_4862_6226# a_4769_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3809 a_9123_1658# a_8922_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3810 a_423_3548# a_222_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3812 a_8342_17# a_8249_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3813 VDD a_6602_6766# a_6509_6766# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3814 a_5349_4336# WWL_15 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3815 RBL0_22 RWL_2 a_13183_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3816 WBL_23 WWL_12 a_13562_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3817 GND a_1289_1906# a_1233_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3818 GND a_18109_5146# a_18053_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3819 a_7669_5416# WWL_11 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3820 a_4282_7036# a_4189_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3821 RBL0_11 RWL_12 a_6803_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3822 a_13993_848# RWL_28 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3823 GND a_15302_3526# a_15209_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3824 a_18202_3526# a_18109_3526# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3825 GND a_15789_17# a_15733_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3826 a_6022_3796# a_5929_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3827 VDD a_15302_7306# a_15209_7306# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3828 a_14049_4876# WWL_13 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3829 a_6022_7576# a_5929_7576# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3830 GND a_14629_3526# a_14573_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3831 a_7613_4358# RWL_15 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3832 a_8342_4876# a_8249_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3833 a_2393_2198# RWL_23 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3834 a_9703_39# a_9502_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3835 GND a_11822_1906# a_11729_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3836 a_2163_4628# a_1962_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3837 VDD a_11822_5686# a_11729_5686# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3838 a_10569_3256# WWL_19 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3839 a_9703_7868# a_9502_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3840 GND a_8249_826# a_8193_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3841 WBL_14 WWL_9 a_8342_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3842 a_18053_1658# RWL_25 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3843 a_16083_7328# a_15882_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3844 RBL0_24 RWL_24 a_14343_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3845 a_11242_2716# a_11149_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3846 a_11242_6496# a_11149_6496# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3847 WBL_1 WWL_29 a_802_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3848 GND a_9409_4336# a_9353_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3849 GND a_709_6226# a_653_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3850 a_12603_5708# a_12402_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3851 VDD a_16462_1366# a_16369_1366# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3852 a_14923_6788# a_14722_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3853 a_9123_1388# a_8922_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3854 a_423_3278# a_222_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3855 GND a_6602_2716# a_6509_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3856 GND a_7182_3796# a_7089_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3857 a_9502_2716# a_9409_2716# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3858 a_802_4606# a_709_4606# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3859 VDD a_7182_7576# a_7089_7576# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3860 RBL0_22 a_4683_7576# a_13183_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3861 VDD a_6602_6496# a_6509_6496# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3862 a_5349_4066# WWL_16 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3863 WBL_23 WWL_13 a_13562_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3864 GND a_1289_1636# a_1233_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3865 GND a_5929_2716# a_5873_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3866 a_11673_309# RWL_30 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3867 a_13993_578# RWL_29 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3868 GND a_15302_3256# a_15209_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3869 WBL_31 WWL_17 a_18202_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3870 RBL0_15 RWL_21 a_9123_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3871 WBL_30 WWL_21 a_17622_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3872 a_5293_3008# RWL_20 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3873 a_6022_3526# a_5929_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3874 VDD a_15302_7036# a_15209_7036# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3875 a_1869_2446# WWL_22 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3876 RBL0_0 RWL_14 a_423_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3877 GND a_14629_3256# a_14573_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3878 a_6022_7306# a_5929_7306# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3879 a_7613_4088# RWL_16 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3880 GND a_3029_8386# a_2973_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3881 a_7383_6518# a_7182_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3882 GND a_11822_1636# a_11729_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3883 a_653_2738# RWL_21 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3884 a_15789_5146# WWL_12 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3885 WBL_13 WWL_30 a_7762_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3886 VDD a_11822_5416# a_11729_5416# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3887 a_2542_1906# a_2449_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3888 a_10569_2986# WWL_20 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3889 a_2163_4358# a_1962_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3890 a_9703_7598# a_9502_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3891 a_2542_5686# a_2449_5686# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3892 GND a_8249_556# a_8193_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3893 GND a_2542_7846# a_2449_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3894 GND a_1869_7846# a_1813_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3895 a_18053_1388# RWL_26 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3896 a_16083_7058# a_15882_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3897 a_9123_848# a_8922_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3898 a_16462_4606# a_16369_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3899 RBL0_24 RWL_25 a_14343_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3900 a_11242_2446# a_11149_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3901 a_16462_8386# a_16369_8386# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3902 WBL_19 WWL_6 a_11242_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3903 a_11242_6226# a_11149_6226# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3904 RBL0_3 RWL_10 a_2163_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3905 WBL_1 WWL_30 a_802_286# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3906 a_6022_17# a_5929_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3907 RBL0_7 RWL_6 a_4483_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3908 GND a_9409_4066# a_9353_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3909 a_12603_5438# a_12402_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3910 VDD a_16462_1096# a_16369_1096# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3911 GND a_1382_16# a_1289_16# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3912 a_7182_1366# a_7089_1366# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3913 RBL0_27 RWL_0 a_16083_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3914 GND a_7182_3526# a_7089_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3915 a_5293_5978# RWL_9 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3916 GND a_13469_17# a_13413_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3917 GND a_6602_2446# a_6509_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3918 VDD a_7182_7306# a_7089_7306# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3919 a_802_4336# a_709_4336# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3920 VDD a_6602_6226# a_6509_6226# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3921 GND a_1289_1366# a_1233_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3922 GND a_5929_2446# a_5873_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3923 WBL_23 WWL_28 a_13562_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3924 WBL_27 WWL_22 a_15882_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3925 VDD a_18202_7846# a_18109_7846# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3926 a_7383_39# a_7182_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3927 RBL0_15 RWL_22 a_9123_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3928 WBL_31 WWL_18 a_18202_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3929 RBL0_25 RWL_2 a_14923_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3930 a_1869_2176# WWL_23 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3931 a_6022_3256# a_5929_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3932 RBL0_0 RWL_15 a_423_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3934 RBL0_23 RWL_31 a_13763_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3935 WBL_10 WWL_3 a_6022_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3936 a_6022_7036# a_5929_7036# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3937 GND a_3029_8116# a_2973_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3938 VDD a_10082_5146# a_9989_5146# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3939 GND a_11822_1366# a_11729_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3940 a_653_2468# RWL_22 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3941 a_10513_4898# RWL_13 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3942 a_7383_6248# a_7182_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3943 a_1813_1118# RWL_27 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3944 a_7182_826# a_7089_826# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3945 WBL_13 WWL_31 a_7762_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3946 a_7762_3796# a_7669_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3947 a_15789_4876# WWL_13 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3948 a_2542_1636# a_2449_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3949 a_2163_4088# a_1962_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3950 a_7762_7576# a_7669_7576# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3951 a_2542_5416# a_2449_5416# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3952 GND a_2542_7576# a_2449_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3953 a_17529_1636# WWL_25 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3955 GND a_1869_7576# a_1813_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3956 a_9123_578# a_8922_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3957 a_16462_4336# a_16369_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3958 a_3903_4628# a_3702_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3959 RBL0_24 RWL_26 a_14343_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3960 a_11242_2176# a_11149_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3961 a_16462_8116# a_16369_8116# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3962 a_3029_5686# WWL_10 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3963 WBL_19 WWL_7 a_11242_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3964 RBL0_3 RWL_11 a_2163_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3965 WBL_1 WWL_31 a_802_16# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3966 a_17823_7328# a_17622_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3967 a_12603_5168# a_12402_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3968 a_7182_1096# a_7089_1096# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3969 WBL_12 WWL_25 a_7182_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3970 RBL0_27 RWL_1 a_16083_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3971 a_9933_6788# RWL_6 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3972 GND a_7182_3256# a_7089_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3973 GND a_12309_4876# a_12253_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3974 GND a_3609_1096# a_3553_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3975 a_14343_1928# a_14142_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3976 GND a_6602_2176# a_6509_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3977 WBL_16 WWL_21 a_9502_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3978 VDD a_7182_7036# a_7089_7036# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3979 WBL_1 WWL_14 a_802_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3980 GND a_5929_2176# a_5873_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3981 GND a_222_1906# a_129_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3982 WBL_19 WWL_30 a_11242_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3983 a_13469_6766# WWL_6 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3984 VDD a_222_5686# a_129_5686# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3985 a_10082_8386# a_9989_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3986 WBL_27 WWL_23 a_15882_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3987 RBL0_21 RWL_7 a_12603_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3988 VDD a_1382_826# a_1289_826# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3989 a_8922_7846# a_8829_7846# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3990 RBL0_15 RWL_23 a_9123_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3991 RBL0_25 a_13963_7576# a_14923_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3992 a_1869_1906# WWL_24 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3993 RBL0_0 RWL_16 a_423_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3994 WBL_10 WWL_4 a_6022_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3995 GND a_9502_17# a_9409_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3996 a_13413_5708# RWL_10 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3997 GND a_10082_1096# a_9989_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3998 a_12833_4628# RWL_14 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3999 VDD a_14722_5956# a_14629_5956# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4000 VDD a_10082_4876# a_9989_4876# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4001 a_653_2198# RWL_23 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4002 a_7762_3526# a_7669_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4003 GND a_5442_8386# a_5349_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4004 a_2542_1366# a_2449_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4005 a_7762_7306# a_7669_7306# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4006 WBL_4 WWL_10 a_2542_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4007 GND a_4769_8386# a_4713_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4008 a_18109_2446# WWL_22 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4009 a_17529_1366# WWL_26 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4010 VDD a_14142_2716# a_14049_2716# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4011 RBL0_28 RWL_27 a_16663_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4012 a_14142_2986# a_14049_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4013 a_16462_4066# a_16369_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4014 a_3903_4358# a_3702_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4015 a_8249_7576# WWL_3 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4016 WBL_28 WWL_0 a_16462_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4017 RBL0_12 RWL_4 a_7383_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4018 a_3029_5416# WWL_11 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4019 a_15209_287# WWL_30 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4020 WBL_19 WWL_8 a_11242_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4021 RBL0_3 RWL_12 a_2163_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4022 GND a_11149_17# a_11093_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4023 a_17823_7058# a_17622_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4024 a_10662_5146# a_10569_5146# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4025 a_5929_826# WWL_28 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4026 GND a_18202_6766# a_18109_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4027 GND a_15209_5686# a_15153_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4028 RBL0_7 RWL_30 a_4483_308# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4029 a_8193_6518# RWL_7 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4030 GND a_9502_2986# a_9409_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4031 GND a_10662_7306# a_10569_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4032 WBL_12 WWL_26 a_7182_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4033 GND a_17529_6766# a_17473_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4034 RBL0_6 RWL_10 a_3903_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4035 a_16663_848# a_16462_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4036 a_5063_39# a_4862_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4037 GND a_8829_2986# a_8773_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4038 a_14343_1658# a_14142_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4039 GND a_4189_286# a_4133_308# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4040 GND a_222_1636# a_129_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4041 WBL_19 WWL_31 a_11242_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4042 a_5063_7868# a_4862_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4043 a_13469_6496# WWL_7 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4044 RBL0_30 RWL_0 a_17823_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4045 VDD a_222_5416# a_129_5416# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4046 WBL_27 WWL_24 a_15882_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4047 a_10082_8116# a_9989_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4048 RBL0_21 RWL_8 a_12603_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4049 VDD a_1382_4066# a_1289_4066# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4050 a_13413_5438# RWL_11 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4051 a_9409_1636# WWL_25 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4052 a_14142_5956# a_14049_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4053 VDD a_17042_826# a_16949_826# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4054 a_12833_4358# RWL_15 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4055 a_5442_5956# a_5349_5956# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4056 a_7762_3256# a_7669_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4057 GND a_5442_8116# a_5349_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4058 a_7762_7036# a_7669_7036# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4059 WBL_13 WWL_3 a_7762_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4060 GND a_4769_8116# a_4713_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4061 WBL_4 WWL_11 a_2542_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4062 a_18109_2176# WWL_23 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4063 a_10283_6788# a_10082_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4064 a_17529_1096# WWL_27 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4065 WBL_10 WWL_29 a_6022_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4066 a_1583_3008# a_1382_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4067 GND a_802_7846# a_709_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4068 WBL_24 WWL_5 a_14142_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4069 GND a_9502_5956# a_9409_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4070 a_3903_4088# a_3702_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4071 GND a_1962_6496# a_1869_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4072 a_8249_7306# WWL_4 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4073 WBL_28 WWL_1 a_16462_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4074 RBL0_12 RWL_5 a_7383_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4075 GND a_8829_5956# a_8773_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4076 a_14722_826# a_14629_826# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4077 a_15209_17# WWL_31 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4078 a_6223_1928# a_6022_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4079 GND a_4189_4876# a_4133_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4080 a_10662_1096# a_10569_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4081 GND a_15209_5416# a_15153_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4082 a_10662_4876# a_10569_4876# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4083 a_8193_6248# RWL_8 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4084 a_14343_309# a_14142_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4085 GND a_10662_7036# a_10569_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4086 a_8922_6766# a_8829_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4087 a_4769_5686# WWL_10 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4088 a_1382_7306# a_1289_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4089 a_16663_578# a_16462_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4090 WBL_12 WWL_27 a_7182_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4091 RBL0_6 RWL_11 a_3903_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4092 a_14343_1388# a_14142_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4093 GND a_12402_3796# a_12309_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4094 a_14722_2716# a_14629_2716# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4095 a_15302_3796# a_15209_3796# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4096 VDD a_12402_7576# a_12309_7576# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4097 a_11149_5146# WWL_12 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4098 a_10082_1636# a_9989_1636# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4099 GND a_11729_3796# a_11673_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4100 GND a_14722_4876# a_14629_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4101 GND a_222_1366# a_129_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4102 a_4713_4628# RWL_14 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4103 a_5063_7598# a_4862_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4104 RBL0_30 RWL_1 a_17823_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4105 a_13469_6226# WWL_8 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4106 WBL_15 WWL_2 a_8922_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4107 a_9409_1366# WWL_26 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4108 a_1583_5978# a_1382_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4109 a_13413_5168# RWL_12 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4110 VDD a_5442_1636# a_5349_1636# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4111 a_709_3256# WWL_19 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4112 a_12833_4088# RWL_16 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4113 RBL0_29 RWL_13 a_17243_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4114 RBL0_14 RWL_27 a_8543_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4115 a_15153_1928# RWL_24 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4116 VDD a_17042_3256# a_16949_3256# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4117 WBL_13 WWL_4 a_7762_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4118 a_18109_1906# WWL_24 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4119 GND a_7089_5686# a_7033_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4120 GND a_6509_4606# a_6453_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4121 GND a_802_7576# a_709_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4122 GND a_1962_6226# a_1869_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4123 a_6223_1658# a_6022_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4124 VDD a_15882_2716# a_15789_2716# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4125 a_15882_2986# a_15789_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4126 VDD a_3702_6766# a_3609_6766# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4127 a_2449_4336# WWL_15 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4128 RBL0_17 RWL_2 a_10283_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4129 WBL_18 WWL_12 a_10662_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4130 GND a_15209_5146# a_15153_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4131 a_9989_7576# WWL_3 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4132 a_4769_5416# WWL_11 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4133 a_1382_7036# a_1289_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4134 RBL0_6 RWL_12 a_3903_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4135 a_1813_848# RWL_28 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4136 a_12982_2446# a_12889_2446# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4137 GND a_17622_5686# a_17529_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4138 GND a_12402_3526# a_12309_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4139 a_15302_3526# a_15209_3526# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4140 a_16369_7036# WWL_5 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4141 GND a_16949_5686# a_16893_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4142 a_73_1118# RWL_27 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4143 a_3122_3796# a_3029_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4144 VDD a_12402_7306# a_12309_7306# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4145 a_11149_4876# WWL_13 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4146 a_3122_7576# a_3029_7576# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4147 GND a_11729_3526# a_11673_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4148 a_4713_4358# RWL_15 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4149 a_5442_4876# a_5349_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4150 a_17042_6496# a_16949_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4151 VDD a_8342_2446# a_8249_2446# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4152 a_6803_7868# a_6602_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4153 a_1869_556# WWL_29 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4154 a_9409_1096# WWL_27 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4155 a_709_2986# WWL_20 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4156 WBL_9 WWL_9 a_5442_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4157 a_15153_1658# RWL_25 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4158 a_13183_7328# a_12982_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4159 RBL0_19 RWL_24 a_11443_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4160 VDD a_17042_2986# a_16949_2986# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4161 a_15882_5956# a_15789_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4162 WBL_8 WWL_21 a_4862_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4163 GND a_7089_5416# a_7033_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4164 GND a_6509_4336# a_6453_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4165 RBL0_16 RWL_30 a_9703_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4166 VDD a_13562_1366# a_13469_1366# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4167 a_6223_1388# a_6022_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4168 a_12023_6788# a_11822_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4169 GND a_3702_2716# a_3609_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4170 GND a_4282_3796# a_4189_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4171 a_6602_2716# a_6509_2716# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4172 VDD a_4282_7576# a_4189_7576# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4173 a_15882_826# a_15789_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4174 RBL0_17 a_4683_7576# a_10283_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4175 VDD a_3702_6496# a_3609_6496# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4176 a_2449_4066# WWL_16 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4177 WBL_18 WWL_13 a_10662_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4178 a_9989_7306# WWL_4 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4179 a_17622_3256# a_17529_3256# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4180 a_12982_2176# a_12889_2176# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4181 a_1813_578# RWL_29 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4182 a_15733_7868# RWL_2 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4183 GND a_17622_5416# a_17529_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4184 a_11093_6788# RWL_6 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4185 a_8342_5686# a_8249_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4186 GND a_12402_3256# a_12309_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4187 WBL_26 WWL_17 a_15302_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4188 RBL0_10 RWL_21 a_6223_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4189 WBL_25 WWL_21 a_14722_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4190 a_2393_3008# RWL_20 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4191 a_3122_3526# a_3029_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4192 VDD a_12402_7036# a_12309_7036# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4193 GND a_16949_5416# a_16893_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4194 a_3122_7306# a_3029_7306# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4195 GND a_11729_3256# a_11673_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4196 a_17473_848# RWL_28 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4197 RBL0_6 RWL_31 a_3903_38# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4198 a_4713_4088# RWL_16 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4199 a_10662_556# a_10569_556# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4200 a_4483_6518# a_4282_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4201 a_17042_6226# a_16949_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4202 a_12889_5146# WWL_12 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4203 VDD a_8342_2176# a_8249_2176# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4204 a_6803_7598# a_6602_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4205 WBL_20 WWL_0 a_11822_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4206 a_1869_286# WWL_30 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4207 RBL0_26 RWL_28 a_15503_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4208 a_15153_1388# RWL_26 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4209 a_13183_7058# a_12982_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4210 a_17529_556# WWL_29 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4211 RBL0_19 RWL_25 a_11443_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4212 a_13562_4606# a_13469_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4213 a_13562_8386# a_13469_8386# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4214 GND a_6602_826# a_6509_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4215 a_16893_1928# RWL_24 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4216 RBL0_2 RWL_6 a_1583_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4217 GND a_7089_5146# a_7033_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4218 GND a_6509_4066# a_6453_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4219 a_17243_4898# a_17042_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4220 a_8543_1118# a_8342_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4221 VDD a_13562_1096# a_13469_1096# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4222 a_4282_1366# a_4189_1366# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4223 RBL0_22 RWL_0 a_13183_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4224 GND a_129_3796# a_73_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4225 GND a_8922_4606# a_8829_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4226 a_13562_287# a_13469_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4227 GND a_3702_2446# a_3609_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4228 GND a_4282_3526# a_4189_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4229 a_2393_5978# RWL_9 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4230 VDD a_8922_8386# a_8829_8386# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4231 VDD a_4282_7306# a_4189_7306# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4232 a_7669_5956# WWL_9 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4233 a_15882_556# a_15789_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4234 VDD a_3702_6226# a_3609_6226# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4235 WBL_2 WWL_28 a_1382_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4236 a_18202_4066# a_18109_4066# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4237 a_12982_1906# a_12889_1906# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4238 WBL_22 WWL_22 a_12982_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4239 a_17622_2986# a_17529_2986# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4240 VDD a_15302_7846# a_15209_7846# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4241 GND a_17622_5146# a_17529_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4242 a_15733_7598# a_13963_7576# RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4243 a_8342_5416# a_8249_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4244 a_7089_2716# WWL_21 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4245 RBL0_10 RWL_22 a_6223_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4246 a_3122_3256# a_3029_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4247 WBL_26 WWL_18 a_15302_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4248 GND a_16949_5146# a_16893_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4249 a_15153_309# RWL_30 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4250 WBL_5 WWL_3 a_3122_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4251 a_3122_7036# a_3029_7036# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4252 a_17473_578# RWL_29 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4253 a_9703_8408# a_9502_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4254 a_4483_6248# a_4282_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4255 a_4862_3796# a_4769_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4256 VDD a_8342_1906# a_8249_1906# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4257 a_12889_4876# WWL_13 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4258 a_4862_7576# a_4769_7576# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4259 WBL_20 WWL_1 a_11822_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4260 a_1869_16# WWL_31 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4261 RBL0_22 RWL_30 a_13183_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4262 RBL0_26 RWL_29 a_15503_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4263 a_14629_1636# WWL_25 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4264 a_16949_2716# WWL_21 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4265 a_13562_4336# a_13469_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4266 RBL0_19 RWL_26 a_11443_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4267 a_13562_8116# a_13469_8116# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4268 GND a_6602_556# a_6509_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4269 GND a_3609_826# a_3553_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4270 GND a_1289_16# a_1233_38# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4271 a_16893_1658# RWL_25 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4272 a_14923_7328# a_14722_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4273 a_802_5146# a_709_5146# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4274 a_9502_3256# a_9409_3256# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4275 a_14049_8386# WWL_0 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4276 a_4282_1096# a_4189_1096# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4277 WBL_7 WWL_25 a_4282_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4278 RBL0_22 RWL_1 a_13183_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4279 GND a_129_3526# a_73_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4280 a_7613_7868# RWL_2 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4281 a_11443_1928# a_11242_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4282 GND a_4282_3256# a_4189_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4283 GND a_8922_4336# a_8829_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4284 GND a_3702_2176# a_3609_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4285 WBL_11 WWL_21 a_6602_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4286 VDD a_8922_8116# a_8829_8116# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4287 VDD a_4282_7036# a_4189_7036# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4288 RBL0_2 RWL_31 a_1583_38# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4289 WBL_31 WWL_15 a_18202_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4290 a_10569_6766# WWL_6 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4291 WBL_30 WWL_19 a_17622_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4292 VDD a_6022_3796# a_5929_3796# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4293 WBL_22 WWL_23 a_12982_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4294 a_6022_7846# a_5929_7846# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4295 a_8342_5146# a_8249_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4296 RBL0_10 RWL_23 a_6223_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4297 WBL_29 WWL_28 a_17042_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4298 WBL_5 WWL_4 a_3122_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4299 GND a_16949_287# a_16893_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4300 a_10513_5708# RWL_10 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4301 VDD a_11822_5956# a_11729_5956# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4302 a_9703_8138# a_9502_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4304 a_4862_3526# a_4769_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4305 GND a_2542_8386# a_2449_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4306 a_4862_7306# a_4769_7306# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4307 GND a_9409_7846# a_9353_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4308 GND a_1869_8386# a_1813_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4309 a_15209_2446# WWL_22 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4310 a_14629_1366# WWL_26 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4311 VDD a_11242_2716# a_11149_2716# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4312 RBL0_23 RWL_27 a_13763_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4313 a_11242_2986# a_11149_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4314 a_423_6788# a_222_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4315 a_9123_4898# a_8922_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4316 a_13562_4066# a_13469_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4317 a_5349_7576# WWL_3 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4318 WBL_23 WWL_0 a_13562_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4319 RBL0_7 RWL_4 a_4483_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4321 GND a_3609_556# a_3553_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4323 a_16893_1388# RWL_26 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4324 a_14923_7058# a_14722_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4325 a_802_1096# a_709_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4326 GND a_15302_6766# a_15209_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4327 GND a_12309_5686# a_12253_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4328 a_5293_6518# RWL_7 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4329 GND a_6602_2986# a_6509_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4330 a_9502_2986# a_9409_2986# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4331 a_14049_8116# WWL_1 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4332 VDD a_7182_7846# a_7089_7846# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4333 a_4483_848# a_4282_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4334 WBL_7 WWL_26 a_4282_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4335 a_802_4876# a_709_4876# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4336 GND a_14629_6766# a_14573_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4337 GND a_129_3256# a_73_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4338 a_16663_3818# a_16462_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4339 a_7613_7598# a_4683_7576# RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4340 GND a_5929_2986# a_5873_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4341 GND a_8922_4066# a_8829_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4342 a_11443_1658# a_11242_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4343 WBL_16 WWL_29 a_9502_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4344 a_2163_7868# a_1962_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4345 a_10569_6496# WWL_7 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4346 RBL0_15 RWL_20 a_9123_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4347 WBL_30 WWL_20 a_17622_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4348 VDD a_6022_3526# a_5929_3526# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4349 WBL_31 WWL_16 a_18202_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4350 RBL0_25 RWL_0 a_14923_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4351 WBL_22 WWL_24 a_12982_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4352 GND a_9409_17# a_9353_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4353 a_9353_1118# RWL_27 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4354 a_18053_4898# RWL_13 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4355 a_10513_5438# RWL_11 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4356 a_6509_1636# WWL_25 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4357 a_653_3008# RWL_20 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4358 a_11242_5956# a_11149_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4359 a_2542_5956# a_2449_5956# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4360 a_17823_309# a_17622_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4361 a_4862_3256# a_4769_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4362 GND a_2542_8116# a_2449_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4363 a_4862_7036# a_4769_7036# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4364 GND a_9409_7576# a_9353_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4365 GND a_1869_8116# a_1813_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4366 a_15209_2176# WWL_23 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4367 VDD a_16462_4606# a_16369_4606# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4368 a_14629_1096# WWL_27 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4369 a_1962_2716# a_1869_2716# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4370 WBL_19 WWL_5 a_11242_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4371 GND a_6602_5956# a_6509_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4372 a_5349_7306# WWL_4 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4373 a_2542_826# a_2449_826# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4374 WBL_23 WWL_1 a_13562_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4375 RBL0_7 RWL_5 a_4483_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4376 GND a_5929_5956# a_5873_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4377 GND a_1289_4876# a_1233_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4378 a_3323_1928# a_3122_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4379 a_9933_7328# RWL_4 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4380 GND a_12309_5416# a_12253_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4381 a_5293_6248# RWL_8 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4382 RBL0_15 RWL_9 a_9123_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4383 WBL_16 WWL_19 a_9502_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4384 RBL0_0 RWL_2 a_423_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4385 a_6022_6766# a_5929_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4386 a_1869_5686# WWL_10 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4387 WBL_1 WWL_12 a_802_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4388 a_4483_578# a_4282_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4389 VDD a_8922_826# a_8829_826# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4390 WBL_7 WWL_27 a_4282_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4391 a_16663_3548# a_16462_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4392 a_11443_1388# a_11242_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4393 a_12889_826# WWL_28 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4394 a_11822_2716# a_11729_2716# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4395 a_12402_3796# a_12309_3796# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4396 a_653_5978# RWL_9 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4397 GND a_11822_4876# a_11729_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4398 a_15789_8386# WWL_0 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4399 a_1813_4628# RWL_14 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4400 a_2163_7598# a_1962_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4401 RBL0_25 RWL_1 a_14923_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4402 a_10569_6226# WWL_8 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4403 WBL_10 WWL_2 a_6022_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4404 a_15882_287# a_15789_287# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4405 GND a_2542_286# a_2449_286# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4406 a_129_556# WWL_29 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4407 RBL0_20 RWL_17 a_12023_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4408 a_16462_7846# a_16369_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4409 a_6509_1366# WWL_26 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4410 VDD a_7762_3796# a_7669_3796# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4411 a_10513_5168# RWL_12 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4412 VDD a_2542_1636# a_2449_1636# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4413 RBL0_24 RWL_13 a_14343_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4414 RBL0_9 RWL_27 a_5643_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4415 a_7762_7846# a_7669_7846# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4416 a_12253_1928# RWL_24 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4417 VDD a_14142_3256# a_14049_3256# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4418 a_15209_1906# WWL_24 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4419 VDD a_16462_4336# a_16369_4336# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4420 a_7182_4606# a_7089_4606# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4421 GND a_7182_6766# a_7089_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4422 a_3029_5956# WWL_9 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4423 GND a_4189_5686# a_4133_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4424 GND a_3609_4606# a_3553_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4425 WBL_22 WWL_29 a_12982_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4426 a_3323_1658# a_3122_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4427 a_7963_2738# a_7762_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4428 GND a_18202_7306# a_18109_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4429 VDD a_12982_2716# a_12889_2716# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4430 WBL_27 WWL_10 a_15882_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4431 GND a_17529_7306# a_17473_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4432 GND a_12309_5146# a_12253_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4433 a_9933_7058# RWL_5 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4434 RBL0_0 RWL_3 a_423_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4435 a_1869_5416# WWL_11 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4436 VDD a_6602_287# a_6509_287# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4437 WBL_16 WWL_20 a_9502_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4438 WBL_1 WWL_13 a_802_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4439 a_10082_2446# a_9989_2446# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4440 a_16663_3278# a_16462_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4441 GND a_14722_5686# a_14629_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4442 a_10569_287# WWL_30 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4443 RBL0_19 RWL_31 a_11443_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4444 a_7033_2738# RWL_21 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4445 GND a_10082_4606# a_9989_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4446 a_5063_8408# a_4862_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4447 a_13469_7036# WWL_5 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4448 a_12402_3526# a_12309_3526# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4449 VDD a_10082_8386# a_9989_8386# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4450 VDD a_222_5956# a_129_5956# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4451 a_1813_4358# RWL_15 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4452 a_15789_8116# WWL_1 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4453 a_2542_4876# a_2449_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4454 a_15882_17# a_15789_17# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4455 a_14142_6496# a_14049_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4456 RBL0_29 RWL_10 a_17243_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4457 VDD a_5442_2446# a_5349_2446# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4458 RBL0_28 RWL_14 a_16663_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4459 a_129_286# WWL_30 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4460 RBL0_20 RWL_18 a_12023_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4461 a_3903_7868# a_3702_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4462 a_16462_7576# a_16369_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4463 a_6509_1096# WWL_27 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4464 VDD a_7762_3526# a_7669_3526# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4465 a_17473_3818# RWL_17 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4466 WBL_4 WWL_9 a_2542_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4467 a_12253_1658# RWL_25 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4468 a_10283_7328# a_10082_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4469 VDD a_14142_2986# a_14049_2986# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4470 GND a_802_8386# a_709_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4471 GND a_9502_6496# a_9409_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4472 a_7182_4336# a_7089_4336# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4473 a_8249_7846# WWL_2 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4474 VDD a_12402_826# a_12309_826# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4475 GND a_8829_6496# a_8773_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4476 WBL_3 WWL_21 a_1962_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4477 GND a_4189_5416# a_4133_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4478 GND a_3609_4336# a_3553_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4479 VDD a_10662_1366# a_10569_1366# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4480 a_3323_1388# a_3122_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4481 a_7963_2468# a_7762_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4482 GND a_18202_7036# a_18109_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4483 GND a_1382_3796# a_1289_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4484 a_8922_7306# a_8829_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4485 WBL_27 WWL_11 a_15882_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4486 a_3702_826# a_3609_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4487 a_3702_2716# a_3609_2716# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4488 VDD a_1382_7576# a_1289_7576# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4489 GND a_17529_7036# a_17473_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4490 VDD a_6602_17# a_6509_17# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4491 a_14722_3256# a_14629_3256# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4492 a_10082_2176# a_9989_2176# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4493 GND a_14722_5416# a_14629_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4494 a_10569_17# WWL_31 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4495 a_12833_7868# RWL_2 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4496 GND a_7182_17# a_7089_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4497 a_7033_2468# RWL_22 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4498 GND a_10082_4336# a_9989_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4499 a_5063_8138# a_4862_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4500 a_5442_5686# a_5349_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4501 WBL_21 WWL_17 a_12402_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4502 VDD a_10082_8116# a_9989_8116# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4503 RBL0_5 RWL_21 a_3323_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4504 a_7762_6766# a_7669_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4505 a_5293_848# RWL_28 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4506 a_1813_4088# RWL_16 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4507 a_18109_5686# WWL_10 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4508 a_17529_4606# WWL_14 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4509 a_1583_6518# a_1382_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4510 a_14142_6226# a_14049_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4511 RBL0_29 RWL_11 a_17243_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4512 VDD a_5442_2176# a_5349_2176# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4513 a_129_16# WWL_31 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4514 RBL0_20 RWL_19 a_12023_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4515 RBL0_28 RWL_15 a_16663_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4516 a_3903_7598# a_3702_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4517 RBL0_5 RWL_28 a_3323_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4518 WBL_13 WWL_2 a_7762_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4519 a_17473_3548# RWL_18 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4520 VDD a_4862_556# a_4769_556# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4521 a_12253_1388# RWL_26 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4522 a_5349_556# WWL_29 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4523 a_10283_7058# a_10082_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4524 a_10662_4606# a_10569_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4525 a_10662_8386# a_10569_8386# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4526 GND a_9502_6226# a_9409_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4527 a_5873_39# RWL_31 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4528 GND a_802_8116# a_709_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4529 WBL_12 WWL_14 a_7182_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4530 GND a_8829_6226# a_8773_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4531 a_13993_1928# RWL_24 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4532 GND a_4189_5146# a_4133_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4533 GND a_3609_4066# a_3553_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4534 a_14343_4898# a_14142_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4535 a_5643_1118# a_5442_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4536 VDD a_15882_3256# a_15789_3256# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4537 VDD a_10662_1096# a_10569_1096# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4538 a_222_2716# a_129_2716# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4539 a_1382_1366# a_1289_1366# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4540 a_7963_2198# a_7762_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4541 RBL0_17 RWL_0 a_10283_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4542 GND a_222_4876# a_129_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4543 GND a_1382_3526# a_1289_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4544 a_8922_7036# a_8829_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4545 a_4769_5956# WWL_9 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4546 a_3702_556# a_3609_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4547 VDD a_1382_7306# a_1289_7306# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4548 a_802_826# a_709_826# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4549 a_14722_2986# a_14629_2986# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4550 a_15302_4066# a_15209_4066# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4551 a_10082_1906# a_9989_1906# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4552 WBL_17 WWL_22 a_10082_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4553 VDD a_12402_7846# a_12309_7846# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4554 a_12833_7598# a_4683_7576# RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4555 a_709_6766# WWL_6 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4556 GND a_14722_5146# a_14629_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4557 a_7033_2198# RWL_23 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4558 a_8829_3796# WWL_17 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4559 GND a_10082_4066# a_9989_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4560 a_5442_5416# a_5349_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4561 GND a_7762_287# a_7669_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4562 a_4189_2716# WWL_21 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4563 WBL_21 WWL_18 a_12402_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4564 RBL0_14 RWL_14 a_8543_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4565 RBL0_5 RWL_22 a_3323_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4566 a_5293_578# RWL_29 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4567 VDD a_17042_6766# a_16949_6766# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4568 a_8773_2738# RWL_21 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4569 a_6803_8408# a_6602_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4570 a_18109_5416# WWL_11 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4571 a_1583_6248# a_1382_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4572 RBL0_29 RWL_12 a_17243_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4573 VDD a_5442_1906# a_5349_1906# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4574 RBL0_28 RWL_16 a_16663_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4575 a_14142_556# a_14049_556# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4576 RBL0_5 RWL_29 a_3323_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4577 a_11729_1636# WWL_25 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4578 a_17473_3278# RWL_19 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4579 a_15882_6496# a_15789_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4580 VDD a_802_1636# a_709_1636# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4581 a_10662_4336# a_10569_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4582 a_10662_8116# a_10569_8116# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4583 WBL_8 WWL_19 a_4862_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4584 a_17243_5708# a_17042_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4585 a_13993_1658# RWL_25 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4586 a_12023_7328# a_11822_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4587 VDD a_15882_2986# a_15789_2986# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4588 GND a_13562_826# a_13469_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4589 a_6602_3256# a_6509_3256# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4590 a_73_4628# RWL_14 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4591 a_11149_8386# WWL_0 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4592 a_1382_1096# a_1289_1096# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4593 WBL_2 WWL_25 a_1382_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4594 RBL0_17 RWL_1 a_10283_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4595 a_4713_7868# RWL_2 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4596 GND a_1382_3256# a_1289_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4597 a_9989_7846# WWL_2 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4598 WBL_6 WWL_21 a_3702_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4599 VDD a_1382_7036# a_1289_7036# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4600 a_15733_8408# RWL_0 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4601 a_11093_7328# RWL_4 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4602 a_17042_287# a_16949_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4603 WBL_26 WWL_15 a_15302_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4604 WBL_17 WWL_23 a_10082_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4605 WBL_25 WWL_19 a_14722_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4606 VDD a_3122_3796# a_3029_3796# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4607 RBL0_1 RWL_27 a_1003_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4608 a_3122_7846# a_3029_7846# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4609 a_709_6496# WWL_7 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4610 a_10662_17# a_10569_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4611 a_8829_3526# WWL_18 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4612 a_9409_4606# WWL_14 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4613 a_5442_5146# a_5349_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4614 RBL0_14 RWL_15 a_8543_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4615 RBL0_5 RWL_23 a_3323_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4616 WBL_8 WWL_28 a_4862_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4617 GND a_4769_287# a_4713_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4618 GND a_17042_2716# a_16949_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4619 VDD a_17042_6496# a_16949_6496# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4620 GND a_16369_2716# a_16313_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4621 a_8773_2468# RWL_22 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4622 a_6803_8138# a_6602_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4623 GND a_6509_7846# a_6453_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4624 a_12309_2446# WWL_22 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4625 a_12833_848# RWL_28 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4626 a_11729_1366# WWL_26 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4627 RBL0_18 RWL_27 a_10863_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4628 a_12023_39# a_11822_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4629 a_6223_4898# a_6022_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4630 a_15882_6226# a_15789_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4631 a_10662_4066# a_10569_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4632 WBL_18 WWL_0 a_10662_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4633 a_2449_7576# WWL_3 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4634 WBL_8 WWL_20 a_4862_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4635 RBL0_2 RWL_4 a_1583_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4636 a_17243_5438# a_17042_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4637 WBL_31 WWL_30 a_18202_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4638 a_12982_1906# a_12889_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4639 a_17622_6766# a_17529_6766# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4640 a_12982_5686# a_12889_5686# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4641 RBL0_18 RWL_28 a_10863_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4642 a_13993_1388# RWL_26 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4643 a_12023_7058# a_11822_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4644 GND a_12402_6766# a_12309_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4645 GND a_11242_287# a_11149_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4646 GND a_3702_2986# a_3609_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4647 a_2393_6518# RWL_7 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4648 GND a_13562_556# a_13469_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4649 WBL_0 WWL_21 a_222_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4650 a_6602_2986# a_6509_2986# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4651 a_73_4358# RWL_15 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4652 a_11149_8116# WWL_1 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4653 VDD a_4282_7846# a_4189_7846# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4654 WBL_2 WWL_26 a_1382_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4655 GND a_11729_6766# a_11673_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4656 a_13763_3818# a_13562_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4657 a_4713_7598# a_4683_7576# RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4658 GND a_10569_826# a_10513_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4659 GND a_8342_1906# a_8249_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4660 a_15733_8138# RWL_1 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4661 a_11093_7058# RWL_5 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4662 VDD a_8342_5686# a_8249_5686# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4663 a_7089_3256# WWL_19 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4664 GND a_7669_1906# a_7613_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4665 RBL0_10 RWL_20 a_6223_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4666 WBL_25 WWL_20 a_14722_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4667 VDD a_3122_3526# a_3029_3526# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4668 WBL_26 WWL_16 a_15302_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4669 WBL_17 WWL_24 a_10082_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4670 a_709_6226# WWL_8 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4671 RBL0_14 RWL_16 a_8543_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4672 GND a_17042_2446# a_16949_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4673 a_6453_1118# RWL_27 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4674 a_15153_4898# RWL_13 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4675 VDD a_17042_6226# a_16949_6226# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4676 a_3609_1636# WWL_25 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4677 GND a_16369_2446# a_16313_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4678 a_8773_2198# RWL_23 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4679 a_9123_5708# a_8922_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4680 GND a_6509_7576# a_6453_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4681 a_8543_4628# a_8342_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4682 a_12309_2176# WWL_23 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4683 a_16949_3256# WWL_19 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4684 VDD a_13562_4606# a_13469_4606# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4685 a_12833_578# RWL_29 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4686 a_11729_1096# WWL_27 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4687 GND a_3702_5956# a_3609_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4688 a_2449_7306# WWL_4 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4689 WBL_18 WWL_1 a_10662_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4690 RBL0_2 RWL_5 a_1583_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4691 a_17622_2716# a_17529_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4692 a_18202_3796# a_18109_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4693 a_17243_5168# a_17042_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4694 WBL_31 WWL_31 a_18202_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4695 a_12982_1636# a_12889_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4696 a_18202_7576# a_18109_7576# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4697 a_17622_6496# a_17529_6496# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4698 a_12982_5416# a_12889_5416# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4699 RBL0_18 RWL_29 a_10863_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4700 a_7613_8408# RWL_0 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4701 a_2393_6248# RWL_8 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4702 RBL0_10 RWL_9 a_6223_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4703 WBL_11 WWL_19 a_6602_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4704 a_3122_6766# a_3029_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4705 WBL_2 WWL_27 a_1382_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4706 a_73_4088# RWL_16 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4708 GND a_10569_556# a_10513_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4709 a_13763_3548# a_13562_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4710 GND a_8342_1636# a_8249_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4711 a_12889_8386# WWL_0 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4712 VDD a_8342_5416# a_8249_5416# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4713 a_7089_2986# WWL_20 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4714 GND a_7669_1636# a_7613_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4715 WBL_5 WWL_2 a_3122_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4716 a_18053_5708# RWL_10 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4717 a_129_1636# WWL_25 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4718 GND a_14049_1096# a_13993_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4719 GND a_17042_2176# a_16949_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4720 a_13562_7846# a_13469_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4721 a_3609_1366# WWL_26 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4722 VDD a_4862_3796# a_4769_3796# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4723 RBL0_4 RWL_27 a_2743_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4724 GND a_16369_2176# a_16313_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4725 RBL0_19 RWL_13 a_11443_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4726 GND a_9409_8386# a_9353_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4727 a_4862_7846# a_4769_7846# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4728 VDD a_11242_3256# a_11149_3256# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4729 a_423_7328# a_222_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4730 a_9123_5438# a_8922_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4731 a_8543_4358# a_8342_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4732 a_12309_1906# WWL_24 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4733 a_16949_2986# WWL_20 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4734 VDD a_13562_4336# a_13469_4336# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4735 a_9502_6766# a_9409_6766# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4736 a_4282_4606# a_4189_4606# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4737 GND a_8922_7846# a_8829_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4738 GND a_4282_6766# a_4189_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4739 GND a_1289_5686# a_1233_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4740 a_18202_3526# a_18109_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4741 a_12982_1366# a_12889_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4742 a_17622_2446# a_17529_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4743 a_18202_7306# a_18109_7306# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4744 GND a_15302_7306# a_15209_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4745 WBL_30 WWL_6 a_17622_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4746 a_17622_6226# a_17529_6226# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4747 WBL_22 WWL_10 a_12982_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4748 GND a_14629_7306# a_14573_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4749 a_6022_826# a_5929_826# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4750 a_7613_8138# RWL_1 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4751 WBL_11 WWL_20 a_6602_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4752 a_13763_3278# a_13562_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4753 GND a_11822_5686# a_11729_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4754 a_4133_2738# RWL_21 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4755 a_2163_8408# a_1962_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4756 a_10569_7036# WWL_5 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4757 VDD a_6022_4066# a_5929_4066# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4758 GND a_8342_1366# a_8249_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4759 a_12889_8116# WWL_1 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4760 VDD a_15882_826# a_15789_826# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4761 GND a_7669_1366# a_7613_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4762 a_16369_826# WWL_28 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4763 a_18053_5438# RWL_11 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4764 a_129_1366# WWL_26 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4765 a_11242_6496# a_11149_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4766 RBL0_24 RWL_10 a_14343_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4767 VDD a_2542_2446# a_2449_2446# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4768 RBL0_23 RWL_14 a_13763_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4769 a_13562_7576# a_13469_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4770 a_3609_1096# WWL_27 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4771 VDD a_4862_3526# a_4769_3526# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4772 RBL0_16 RWL_31 a_9703_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4773 GND a_9409_8116# a_9353_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4774 a_14573_3818# RWL_17 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4775 VDD a_16462_5146# a_16369_5146# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4776 VDD a_11242_2986# a_11149_2986# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4777 GND a_11822_17# a_11729_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4778 a_16893_4898# RWL_13 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4779 a_423_7058# a_222_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4780 a_9123_5168# a_8922_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4781 a_9502_2716# a_9409_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4782 a_1962_3256# a_1869_3256# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4783 a_8543_4088# a_8342_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4784 a_802_4606# a_709_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4785 a_9502_6496# a_9409_6496# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4786 GND a_6602_6496# a_6509_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4787 a_802_8386# a_709_8386# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4788 a_4282_4336# a_4189_4336# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4789 a_5349_7846# WWL_2 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4790 GND a_129_6766# a_73_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4791 GND a_8922_7576# a_8829_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4792 GND a_5929_6496# a_5873_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4793 GND a_1289_5416# a_1233_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4794 a_18202_3256# a_18109_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4795 a_17622_2176# a_17529_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4796 GND a_15302_7036# a_15209_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4797 WBL_31 WWL_3 a_18202_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4798 a_18202_7036# a_18109_7036# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4799 WBL_30 WWL_7 a_17622_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4800 RBL0_15 RWL_7 a_9123_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4801 RBL0_0 RWL_0 a_423_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4802 a_6022_7306# a_5929_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4803 WBL_22 WWL_11 a_12982_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4804 GND a_14629_7036# a_14573_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4805 a_11822_3256# a_11729_3256# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4806 a_653_6518# RWL_7 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4807 GND a_11822_5416# a_11729_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4808 a_9353_4628# RWL_14 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4809 a_4133_2468# RWL_22 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4810 a_2163_8138# a_1962_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4811 a_2542_5686# a_2449_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4812 VDD a_13562_287# a_13469_287# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4813 a_4862_6766# a_4769_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4814 a_14049_287# WWL_30 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4815 a_18053_5168# RWL_12 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4816 a_16462_8386# a_16369_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4817 a_15209_5686# WWL_10 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4818 a_129_1096# WWL_27 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4819 a_14629_4606# WWL_14 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4820 a_11242_6226# a_11149_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4821 RBL0_24 RWL_11 a_14343_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4822 VDD a_2542_2176# a_2449_2176# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4823 RBL0_23 RWL_15 a_13763_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4824 GND a_16462_1096# a_16369_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4825 GND a_3029_286# a_2973_308# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4826 a_14573_3548# RWL_18 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4827 GND a_15789_1096# a_15733_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4828 VDD a_16462_4876# a_16369_4876# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4829 a_7182_5146# a_7089_5146# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4830 a_9502_2446# a_9409_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4831 a_1962_2986# a_1869_2986# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4832 GND a_7182_7306# a_7089_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4833 a_802_4336# a_709_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4834 a_9502_6226# a_9409_6226# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4835 GND a_6602_6226# a_6509_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4836 a_802_8116# a_709_8116# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4837 WBL_16 WWL_6 a_9502_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4838 WBL_7 WWL_14 a_4282_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4839 GND a_5929_6226# a_5873_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4840 GND a_1289_5146# a_1233_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4841 a_11443_4898# a_11242_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4842 a_2743_1118# a_2542_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4843 VDD a_12982_3256# a_12889_3256# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4844 GND a_3029_1906# a_2973_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4845 WBL_31 WWL_4 a_18202_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4846 RBL0_0 RWL_1 a_423_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4847 a_6022_7036# a_5929_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4848 WBL_30 WWL_8 a_17622_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4849 RBL0_15 RWL_8 a_9123_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4850 a_1869_5956# WWL_9 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4851 GND a_7089_17# a_7033_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4852 a_11822_2986# a_11729_2986# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4853 a_12402_4066# a_12309_4066# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4854 a_7182_826# a_7089_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4855 a_653_6248# RWL_8 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4856 a_9353_4358# RWL_15 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4857 GND a_11822_5146# a_11729_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4858 a_4133_2198# RWL_23 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4859 a_5929_3796# WWL_17 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4860 a_2542_5416# a_2449_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4861 a_1289_2716# WWL_21 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4862 RBL0_9 RWL_14 a_5643_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4863 VDD a_13562_17# a_13469_17# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4864 a_14049_17# WWL_31 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4865 VDD a_14142_6766# a_14049_6766# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4866 RBL0_12 RWL_31 a_7383_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4867 a_5873_2738# RWL_21 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4868 a_3903_8408# a_3702_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4869 a_16462_8116# a_16369_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4870 a_15209_5416# WWL_11 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4871 VDD a_7762_4066# a_7669_4066# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4872 RBL0_24 RWL_12 a_14343_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4873 VDD a_2542_1906# a_2449_1906# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4874 RBL0_23 RWL_16 a_13763_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4875 a_1962_556# a_1869_556# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4876 RBL0_27 RWL_24 a_16083_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4877 a_14573_3278# RWL_19 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4878 a_7182_1096# a_7089_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4879 a_7182_4876# a_7089_4876# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4880 a_9502_2176# a_9409_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4881 WBL_3 WWL_19 a_1962_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4882 a_802_4066# a_709_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4883 GND a_7182_7036# a_7089_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4884 a_14343_5708# a_14142_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4885 VDD a_18202_1366# a_18109_1366# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4886 WBL_1 WWL_0 a_802_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4887 WBL_16 WWL_7 a_9502_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4888 VDD a_8342_556# a_8249_556# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4889 a_16663_6788# a_16462_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4890 a_12309_556# WWL_29 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4891 a_7963_3008# a_7762_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4892 GND a_222_5686# a_129_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4893 VDD a_12982_2986# a_12889_2986# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4894 GND a_1382_826# a_1289_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4895 WBL_27 WWL_9 a_15882_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4896 a_3702_3256# a_3609_3256# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4897 GND a_8249_3796# a_8193_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4898 GND a_3029_1636# a_2973_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4899 a_1813_7868# RWL_2 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4900 a_12833_8408# RWL_0 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4901 a_7033_3008# RWL_20 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4902 a_4133_38# RWL_31 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4903 WBL_21 WWL_15 a_12402_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4904 a_7182_556# a_7089_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4905 a_9353_4088# RWL_16 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4906 a_7762_7306# a_7669_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4907 a_5929_3526# WWL_18 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4908 a_6509_4606# WWL_14 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4909 a_2542_5146# a_2449_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4910 RBL0_9 RWL_15 a_5643_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4911 GND a_14142_2716# a_14049_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4912 a_17529_5146# WWL_12 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4913 a_16462_1636# a_16369_1636# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4914 VDD a_14142_6496# a_14049_6496# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4915 GND a_13469_2716# a_13413_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4916 a_5873_2468# RWL_22 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4917 a_3903_8138# a_3702_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4918 GND a_3609_7846# a_3553_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4919 a_1962_286# a_1869_286# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4920 RBL0_27 RWL_25 a_16083_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4921 VDD a_802_2446# a_709_2446# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4922 a_7963_5978# a_7762_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4923 a_3323_4898# a_3122_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4924 WBL_12 WWL_12 a_7182_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4925 WBL_3 WWL_20 a_1962_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4926 a_14343_5438# a_14142_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4927 VDD a_18202_1096# a_18109_1096# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4928 WBL_16 WWL_8 a_9502_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4929 a_10082_1906# a_9989_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4930 WBL_1 WWL_1 a_802_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4931 a_14722_6766# a_14629_6766# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4932 a_8922_1366# a_8829_1366# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4933 a_10082_5686# a_9989_5686# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4934 a_222_3256# a_129_3256# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4935 GND a_10082_7846# a_9989_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4936 a_7033_5978# RWL_9 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4937 GND a_222_5416# a_129_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4938 GND a_1382_556# a_1289_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4939 a_3702_2986# a_3609_2986# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4940 GND a_8249_3526# a_8193_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4941 VDD a_1382_7846# a_1289_7846# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4942 GND a_3029_1366# a_2973_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4943 a_10863_3818# a_10662_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4944 a_1813_7598# RWL_3 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4945 GND a_17042_826# a_16949_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4946 GND a_5442_1906# a_5349_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4947 a_13993_309# RWL_30 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4948 a_12833_8138# RWL_1 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4949 a_8829_4336# WWL_15 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4950 RBL0_28 RWL_2 a_16663_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4951 RBL0_20 RWL_6 a_12023_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4952 VDD a_5442_5686# a_5349_5686# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4953 GND a_4769_1906# a_4713_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4954 a_4189_3256# WWL_19 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4955 WBL_21 WWL_16 a_12402_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4956 RBL0_8 RWL_31 a_5063_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4957 RBL0_5 RWL_20 a_3323_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4958 a_7762_7036# a_7669_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4959 RBL0_9 RWL_16 a_5643_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4960 a_16313_39# RWL_31 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4961 GND a_14142_2446# a_14049_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4962 a_18109_5956# WWL_9 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4963 a_3553_1118# RWL_27 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4964 a_12253_4898# RWL_13 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4965 a_17529_4876# WWL_13 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4966 VDD a_14142_6226# a_14049_6226# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4967 GND a_13469_2446# a_13413_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4968 a_5873_2198# RWL_23 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4969 a_14722_826# a_14629_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4970 GND a_8249_287# a_8193_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4971 a_6223_5708# a_6022_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4972 GND a_3609_7576# a_3553_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4973 VDD a_15882_6766# a_15789_6766# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4974 a_1962_16# a_1869_16# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4975 a_5643_4628# a_5442_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4976 RBL0_27 RWL_26 a_16083_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4977 VDD a_802_2176# a_709_2176# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4978 VDD a_10662_4606# a_10569_4606# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4980 WBL_12 WWL_13 a_7182_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4981 a_14343_5168# a_14142_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4982 RBL0_30 RWL_24 a_17823_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4983 a_14722_2716# a_14629_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4984 a_15302_3796# a_15209_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4985 a_10082_1636# a_9989_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4986 a_15302_7576# a_15209_7576# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4987 a_8922_1096# a_8829_1096# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4988 WBL_15 WWL_25 a_8922_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4989 a_14722_6496# a_14629_6496# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4990 a_10082_5416# a_9989_5416# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4991 a_222_2986# a_129_2986# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4992 GND a_10082_7576# a_9989_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4993 GND a_222_5146# a_129_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4994 a_4713_8408# RWL_0 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4995 RBL0_5 RWL_9 a_3323_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4996 WBL_6 WWL_19 a_3702_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4997 GND a_8249_3256# a_8193_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4998 a_10863_3548# a_10662_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4999 GND a_17042_556# a_16949_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5000 GND a_5442_1636# a_5349_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5001 a_709_7036# WWL_5 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5002 a_9409_5146# WWL_12 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5003 a_8829_4066# WWL_16 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5004 RBL0_28 a_13963_7576# a_16663_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5005 VDD a_5442_5416# a_5349_5416# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5006 GND a_14049_826# a_13993_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5007 a_4189_2986# WWL_20 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5008 GND a_9989_3796# a_9933_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5009 GND a_4769_1636# a_4713_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5010 a_15153_5708# RWL_10 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5011 a_17473_6788# RWL_6 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5012 GND a_11149_1096# a_11093_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5013 GND a_14142_2176# a_14049_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5014 a_8773_3008# RWL_20 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5015 a_10662_7846# a_10569_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5016 VDD a_1962_3796# a_1869_3796# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5017 GND a_13469_2176# a_13413_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5018 WBL_8 WWL_6 a_4862_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5019 a_9502_826# a_9409_826# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5020 GND a_6509_8386# a_6453_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5021 a_14722_556# a_14629_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5022 GND a_15882_2716# a_15789_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5023 VDD a_15882_6496# a_15789_6496# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5024 a_6223_5438# a_6022_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5025 GND a_1962_16# a_1869_16# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5026 a_5643_4358# a_5442_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5027 a_9123_309# a_8922_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5028 VDD a_802_1906# a_709_1906# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5029 VDD a_10662_4336# a_10569_4336# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5030 a_6602_6766# a_6509_6766# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5031 a_1382_4606# a_1289_4606# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5032 GND a_1382_6766# a_1289_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5033 RBL0_30 RWL_25 a_17823_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5034 a_15302_3526# a_15209_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5035 a_7963_39# a_7762_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5036 a_10082_1366# a_9989_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5037 a_14722_2446# a_14629_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5038 a_15302_7306# a_15209_7306# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5039 GND a_12402_7306# a_12309_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5040 WBL_25 WWL_6 a_14722_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5041 a_14722_6226# a_14629_6226# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5042 WBL_15 WWL_26 a_8922_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5043 WBL_0 WWL_19 a_222_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5044 WBL_17 WWL_10 a_10082_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5045 RBL0_1 RWL_14 a_1003_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5046 GND a_11729_7306# a_11673_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5047 a_4713_8138# RWL_1 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5048 RBL0_14 RWL_2 a_8543_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5049 WBL_6 WWL_20 a_3702_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5050 a_10863_3278# a_10662_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5051 a_1233_2738# RWL_21 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5052 WBL_23 WWL_30 a_13562_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5053 a_8773_5978# RWL_9 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5054 VDD a_3122_4066# a_3029_4066# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5055 GND a_5442_1366# a_5349_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5056 a_9409_4876# WWL_13 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5057 GND a_14049_556# a_13993_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5058 GND a_9989_3526# a_9933_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5059 GND a_4769_1366# a_4713_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5060 a_4189_826# WWL_28 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5061 GND a_17042_2986# a_16949_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5062 a_15153_5438# RWL_11 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5063 RBL0_19 RWL_10 a_11443_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5064 GND a_16369_2986# a_16313_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5065 RBL0_18 RWL_14 a_10863_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5066 a_10662_7576# a_10569_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5067 a_7182_287# a_7089_287# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5068 VDD a_1962_3526# a_1869_3526# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5069 WBL_8 WWL_7 a_4862_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5070 GND a_6509_8116# a_6453_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5071 a_11673_3818# RWL_17 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5072 VDD a_13562_5146# a_13469_5146# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5073 GND a_15882_2446# a_15789_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5074 a_13993_4898# RWL_13 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5075 VDD a_15882_6226# a_15789_6226# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5076 a_6223_5168# a_6022_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5077 a_6602_2716# a_6509_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5078 a_5643_4088# a_5442_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5079 a_6602_6496# a_6509_6496# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5080 GND a_3702_6496# a_3609_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5081 a_73_7868# RWL_2 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5082 a_1382_4336# a_1289_4336# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5083 a_2449_7846# WWL_2 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5084 a_12982_5956# a_12889_5956# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5085 RBL0_30 RWL_26 a_17823_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5086 a_15302_3256# a_15209_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5087 a_14722_2176# a_14629_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5088 a_15302_7036# a_15209_7036# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5089 GND a_12402_7036# a_12309_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5090 a_7089_6766# WWL_6 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5091 WBL_26 WWL_3 a_15302_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5092 WBL_25 WWL_7 a_14722_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5093 RBL0_10 RWL_7 a_6223_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5094 WBL_15 WWL_27 a_8922_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5095 WBL_0 WWL_20 a_222_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5096 a_3122_7306# a_3029_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5097 WBL_17 WWL_11 a_10082_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5098 RBL0_1 RWL_15 a_1003_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5099 GND a_11729_7036# a_11673_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5100 RBL0_14 a_4683_7576# a_8543_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5101 a_17042_3796# a_16949_3796# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5102 GND a_17042_5956# a_16949_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5103 a_6453_4628# RWL_14 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5104 VDD a_8342_5956# a_8249_5956# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5105 GND a_16369_5956# a_16313_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5106 a_12982_826# a_12889_826# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5107 a_1233_2468# RWL_22 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5108 WBL_23 WWL_31 a_13562_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5109 GND a_9989_3256# a_9933_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5110 a_16949_6766# WWL_6 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5111 a_12309_5686# WWL_10 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5112 a_15153_5168# RWL_12 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5114 a_13562_8386# a_13469_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5115 a_11729_4606# WWL_14 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5116 RBL0_19 RWL_11 a_11443_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5117 RBL0_18 RWL_15 a_10863_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5118 a_7182_17# a_7089_17# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5119 WBL_8 WWL_8 a_4862_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5120 GND a_11729_17# a_11673_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5121 a_16893_5708# RWL_10 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5122 GND a_13562_1096# a_13469_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5123 a_11673_3548# RWL_18 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5124 VDD a_13562_4876# a_13469_4876# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5125 GND a_12889_1096# a_12833_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5126 GND a_15882_2176# a_15789_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5127 a_4282_5146# a_4189_5146# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5128 WBL_14 WWL_29 a_8342_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5129 a_6602_2446# a_6509_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5130 GND a_8922_8386# a_8829_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5131 GND a_4282_7306# a_4189_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5132 a_5643_39# a_5442_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5133 WBL_11 WWL_6 a_6602_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5134 a_6602_6226# a_6509_6226# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5135 GND a_3702_6226# a_3609_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5136 a_73_7598# RWL_3 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5137 WBL_2 WWL_14 a_1382_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5138 VDD a_17622_2716# a_17529_2716# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5139 a_17622_2986# a_17529_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5140 a_18202_7846# a_18109_7846# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5141 a_5929_287# WWL_30 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5142 a_7089_6496# WWL_7 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5143 WBL_26 WWL_4 a_15302_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5144 WBL_25 WWL_8 a_14722_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5145 RBL0_10 RWL_8 a_6223_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5146 a_3122_7036# a_3029_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5147 a_16663_309# a_16462_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5148 RBL0_1 RWL_16 a_1003_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5149 a_17042_3526# a_16949_3526# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5150 GND a_14049_4606# a_13993_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5151 a_6453_4358# RWL_15 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5152 a_1233_2198# RWL_23 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5153 a_18403_2738# a_18202_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5154 RBL0_4 RWL_14 a_2743_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5155 VDD a_11242_6766# a_11149_6766# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5156 a_8543_7868# a_8342_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5157 a_16949_6496# WWL_7 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5158 a_2973_2738# RWL_21 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5159 a_13562_8116# a_13469_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5160 a_12309_5416# WWL_11 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5161 VDD a_17042_287# a_16949_287# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5162 VDD a_4862_4066# a_4769_4066# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5163 RBL0_19 RWL_12 a_11443_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5164 RBL0_18 RWL_16 a_10863_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5165 RBL0_22 RWL_24 a_13183_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5166 a_16893_5438# RWL_11 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5167 a_17622_5956# a_17529_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5168 a_11729_826# WWL_28 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5169 a_11673_3278# RWL_19 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5170 a_12982_4876# a_12889_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5171 a_4282_1096# a_4189_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5172 a_4282_4876# a_4189_4876# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5173 GND a_129_7306# a_73_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5174 a_6602_2176# a_6509_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5175 GND a_8922_8116# a_8829_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5176 GND a_4282_7036# a_4189_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5177 a_11443_5708# a_11242_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5178 VDD a_15302_1366# a_15209_1366# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5179 WBL_11 WWL_7 a_6602_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5180 a_14722_287# a_14629_287# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5181 a_13763_6788# a_13562_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5182 GND a_6022_3796# a_5929_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5183 a_8342_2716# a_8249_2716# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5184 VDD a_6022_7576# a_5929_7576# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5185 WBL_30 WWL_5 a_17622_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5186 WBL_22 WWL_9 a_12982_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5187 GND a_5349_3796# a_5293_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5188 GND a_8342_4876# a_8249_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5189 a_5929_17# WWL_31 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5190 a_7089_6226# WWL_8 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5191 GND a_7669_4876# a_7613_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5192 a_9703_1928# a_9502_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5193 a_1003_3818# a_802_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5194 WBL_29 WWL_17 a_17042_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5195 RBL0_13 RWL_21 a_7963_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5196 a_4133_3008# RWL_20 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5197 GND a_14049_4336# a_13993_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5198 a_6453_4088# RWL_16 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5199 a_3609_4606# WWL_14 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5200 a_4862_7306# a_4769_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5201 a_18403_2468# a_18202_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5202 RBL0_4 RWL_15 a_2743_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5203 GND a_11242_2716# a_11149_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5204 a_13562_1636# a_13469_1636# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5205 a_14629_5146# WWL_12 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5206 VDD a_11242_6496# a_11149_6496# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5207 WBL_20 WWL_29 a_11822_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5208 a_1962_6766# a_1869_6766# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5209 GND a_10569_2716# a_10513_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5210 a_8543_7598# a_8342_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5211 a_16949_6226# WWL_8 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5212 a_2973_2468# RWL_22 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5213 VDD a_17042_17# a_16949_17# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5214 RBL0_31 RWL_17 a_18403_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5215 GND a_709_826# a_653_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5216 RBL0_22 RWL_25 a_13183_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5217 a_18202_6766# a_18109_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5218 a_16893_5168# RWL_12 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5219 VDD a_8922_1636# a_8829_1636# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5220 a_9502_2986# a_9409_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5221 WBL_7 WWL_12 a_4282_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5222 GND a_129_7036# a_73_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5223 a_11443_5438# a_11242_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5224 VDD a_15302_1096# a_15209_1096# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5225 WBL_11 WWL_8 a_6602_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5226 a_11822_6766# a_11729_6766# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5227 a_14722_17# a_14629_17# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5228 a_6022_1366# a_5929_1366# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5229 GND a_6022_3526# a_5929_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5230 a_4133_5978# RWL_9 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5231 WBL_31 WWL_2 a_18202_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5232 VDD a_6022_7306# a_5929_7306# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5233 GND a_5349_3526# a_5293_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5234 a_9703_1658# a_9502_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5235 a_1003_3548# a_802_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5236 GND a_2542_1906# a_2449_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5237 a_129_4606# WWL_14 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5238 VDD a_2542_5686# a_2449_5686# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5239 RBL0_13 RWL_22 a_7963_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5240 a_1289_3256# WWL_19 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5241 WBL_29 WWL_18 a_17042_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5242 a_5929_4336# WWL_15 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5243 RBL0_23 RWL_2 a_13763_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5244 GND a_1869_1906# a_1813_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5245 a_16083_1118# a_15882_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5246 GND a_14049_4066# a_13993_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5247 a_4862_7036# a_4769_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5248 a_16462_2446# a_16369_2446# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5249 a_18403_2198# a_18202_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5250 RBL0_4 RWL_16 a_2743_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5251 GND a_16462_4606# a_16369_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5252 GND a_11242_2446# a_11149_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5253 VDD a_16462_8386# a_16369_8386# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5254 a_15209_5956# WWL_9 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5255 a_1962_2716# a_1869_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5256 a_14629_4876# WWL_13 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5257 VDD a_11242_6226# a_11149_6226# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5258 GND a_15789_4606# a_15733_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5259 a_1962_6496# a_1869_6496# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5260 a_9502_5956# a_9409_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5261 GND a_10569_2446# a_10513_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5262 a_802_7846# a_709_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5263 a_2973_2198# RWL_23 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5264 a_2542_826# a_2449_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5265 RBL0_30 RWL_28 a_17823_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5266 a_3323_5708# a_3122_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5267 VDD a_7182_1366# a_7089_1366# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5268 VDD a_12982_6766# a_12889_6766# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5269 GND a_709_556# a_653_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5270 RBL0_31 RWL_18 a_18403_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5271 a_2743_4628# a_2542_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5272 RBL0_22 RWL_26 a_13183_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5273 GND a_8922_826# a_8829_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5274 WBL_16 WWL_5 a_9502_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5275 a_4133_848# RWL_28 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5276 WBL_7 WWL_13 a_4282_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5277 a_16663_7328# a_16462_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5278 a_11443_5168# a_11242_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5279 RBL0_25 RWL_24 a_14923_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5280 a_11822_2716# a_11729_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5281 a_12402_3796# a_12309_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5282 a_12402_7576# a_12309_7576# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5283 a_11822_6496# a_11729_6496# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5284 a_6022_1096# a_5929_1096# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5285 WBL_10 WWL_25 a_6022_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5286 a_9353_7868# RWL_2 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5287 GND a_6022_3256# a_5929_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5288 a_1813_8408# RWL_0 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5289 WBL_14 WWL_21 a_8342_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5290 VDD a_6022_7036# a_5929_7036# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5291 a_15882_287# a_15789_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5292 GND a_5349_3256# a_5293_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5293 RBL0_3 RWL_28 a_2163_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5294 a_9703_1388# a_9502_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5295 VDD a_3702_556# a_3609_556# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5296 a_1003_3278# a_802_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5297 GND a_7762_3796# a_7669_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5298 WBL_6 WWL_28 a_3702_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5299 GND a_2542_1636# a_2449_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5300 VDD a_7762_7576# a_7669_7576# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5301 a_6509_5146# WWL_12 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5302 RBL0_13 RWL_23 a_7963_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5303 a_5929_4066# WWL_16 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5304 RBL0_23 a_4683_7576# a_13763_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5305 VDD a_2542_5416# a_2449_5416# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5306 a_1289_2986# WWL_20 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5307 GND a_1869_1636# a_1813_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5308 a_12253_5708# RWL_10 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5309 a_17473_309# RWL_30 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5310 a_16462_2176# a_16369_2176# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5311 GND a_16462_4336# a_16369_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5312 a_14573_6788# RWL_6 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5313 GND a_11242_2176# a_11149_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5314 RBL0_16 RWL_21 a_9703_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5315 a_5873_3008# RWL_20 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5316 a_7182_4606# a_7089_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5317 VDD a_16462_8116# a_16369_8116# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5318 a_1962_2446# a_1869_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5319 GND a_15789_4336# a_15733_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5320 a_7182_8386# a_7089_8386# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5321 GND a_10569_2176# a_10513_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5322 a_802_7576# a_709_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5323 WBL_3 WWL_6 a_1962_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5324 a_1962_6226# a_1869_6226# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5325 GND a_3609_8386# a_3553_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5326 a_2542_556# a_2449_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5327 RBL0_26 RWL_30 a_15503_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5328 GND a_12982_2716# a_12889_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5329 a_7963_6518# a_7762_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5330 a_3323_5438# a_3122_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5331 RBL0_30 RWL_29 a_17823_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5332 VDD a_12982_6496# a_12889_6496# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5333 VDD a_7182_1096# a_7089_1096# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5334 RBL0_31 RWL_19 a_18403_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5335 a_2743_4358# a_2542_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5336 a_3702_6766# a_3609_6766# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5337 GND a_6602_287# a_6509_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5338 GND a_8922_556# a_8829_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5339 a_4133_578# RWL_29 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5340 a_16663_7058# a_16462_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5341 GND a_5929_826# a_5873_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5342 RBL0_25 RWL_25 a_14923_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5343 a_11822_2446# a_11729_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5344 a_12402_3526# a_12309_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5345 GND a_10082_8386# a_9989_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5346 a_7033_6518# RWL_7 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5347 a_12402_7306# a_12309_7306# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5348 a_11822_6226# a_11729_6226# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5349 WBL_10 WWL_26 a_6022_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5350 a_9353_7598# a_4683_7576# RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5351 a_1813_8138# RWL_1 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5352 RBL0_9 RWL_2 a_5643_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5353 RBL0_3 RWL_29 a_2163_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5354 a_7762_1366# a_7669_1366# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5355 RBL0_28 RWL_0 a_16663_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5356 RBL0_20 RWL_4 a_12023_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5357 VDD a_3702_286# a_3609_286# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5358 a_5873_5978# RWL_9 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5359 GND a_7762_3526# a_7669_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5360 GND a_2542_1366# a_2449_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5361 VDD a_7762_7306# a_7669_7306# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5362 a_6509_4876# WWL_13 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5363 GND a_1869_1366# a_1813_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5364 a_8249_1636# WWL_25 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5365 GND a_14142_2986# a_14049_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5366 a_12253_5438# RWL_11 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5367 a_16462_1906# a_16369_1906# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5368 WBL_28 WWL_22 a_16462_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5369 GND a_13469_2986# a_13413_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5370 GND a_16462_4066# a_16369_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5371 GND a_12402_826# a_12309_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5372 RBL0_16 RWL_22 a_9703_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5373 a_7182_4336# a_7089_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5374 a_17823_1118# a_17622_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5375 a_1962_2176# a_1869_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5376 GND a_15789_4066# a_15733_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5377 a_7182_8116# a_7089_8116# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5378 WBL_3 WWL_7 a_1962_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5379 GND a_3609_8116# a_3553_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5380 GND a_1869_16# a_1813_38# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5381 VDD a_18202_4606# a_18109_4606# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5382 VDD a_10662_5146# a_10569_5146# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5383 a_222_6766# a_129_6766# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5384 GND a_12982_2446# a_12889_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5385 a_7963_6248# a_7762_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5386 VDD a_12982_6226# a_12889_6226# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5387 a_3323_5168# a_3122_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5388 a_3702_2716# a_3609_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5389 a_2743_4088# a_2542_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5390 a_3702_6496# a_3609_6496# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5391 a_5063_1928# a_4862_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5392 GND a_3029_4876# a_2973_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5393 a_10082_5956# a_9989_5956# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5394 GND a_5929_556# a_5873_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5395 RBL0_25 RWL_26 a_14923_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5396 a_12402_3256# a_12309_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5397 GND a_10082_8116# a_9989_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5398 a_7033_6248# RWL_8 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5399 a_11822_2176# a_11729_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5400 a_12402_7036# a_12309_7036# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5401 a_4189_6766# WWL_6 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5402 WBL_21 WWL_3 a_12402_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5403 RBL0_5 RWL_7 a_3323_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5404 WBL_10 WWL_27 a_6022_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5405 a_6803_848# a_6602_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5406 RBL0_9 a_4683_7576# a_5643_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5407 a_14142_3796# a_14049_3796# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5408 GND a_14142_5956# a_14049_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5409 a_3553_4628# RWL_14 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5410 a_17529_8386# WWL_0 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5411 a_7762_1096# a_7669_1096# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5412 WBL_13 WWL_25 a_7762_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5413 RBL0_28 RWL_1 a_16663_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5414 RBL0_20 RWL_5 a_12023_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5415 VDD a_5442_5956# a_5349_5956# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5416 GND a_13469_5956# a_13413_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5417 VDD a_3702_16# a_3609_16# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5418 GND a_7762_3256# a_7669_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5419 VDD a_7762_7036# a_7669_7036# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5420 WBL_29 WWL_30 a_17042_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5421 GND a_802_1906# a_709_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5422 a_17473_7328# RWL_4 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5423 a_8249_1366# WWL_26 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5424 VDD a_9502_3796# a_9409_3796# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5425 VDD a_802_5686# a_709_5686# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5426 a_12253_5168# RWL_12 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5427 WBL_28 WWL_23 a_16462_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5428 RBL0_27 RWL_13 a_16083_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5429 a_10662_8386# a_10569_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5430 RBL0_12 RWL_27 a_7383_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5431 VDD a_7182_826# a_7089_826# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5432 GND a_12402_556# a_12309_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5433 a_6602_17# a_6509_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5434 RBL0_16 RWL_23 a_9703_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5435 a_7182_4066# a_7089_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5436 WBL_12 WWL_0 a_7182_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5437 WBL_3 WWL_8 a_1962_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5438 a_13993_5708# RWL_10 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5439 GND a_10662_1096# a_10569_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5440 a_222_2716# a_129_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5441 VDD a_18202_4336# a_18109_4336# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5442 a_8922_4606# a_8829_4606# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5443 VDD a_10662_4876# a_10569_4876# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5444 a_222_6496# a_129_6496# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5445 GND a_12982_2176# a_12889_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5446 a_1382_5146# a_1289_5146# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5447 a_3702_2446# a_3609_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5448 GND a_1382_7306# a_1289_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5449 WBL_6 WWL_6 a_3702_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5450 a_3702_6226# a_3609_6226# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5451 a_802_826# a_709_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5452 GND a_8249_6766# a_8193_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5453 a_5063_1658# a_4862_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5454 a_4862_826# a_4769_826# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5455 VDD a_10082_1636# a_9989_1636# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5456 VDD a_14722_2716# a_14629_2716# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5457 a_14722_2986# a_14629_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5458 a_15302_7846# a_15209_7846# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5459 a_8829_7576# WWL_3 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5460 RBL0_14 RWL_0 a_8543_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5461 a_4189_6496# WWL_7 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5462 WBL_21 WWL_4 a_12402_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5463 RBL0_5 RWL_8 a_3323_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5464 a_6803_578# a_6602_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5465 a_17042_17# a_16949_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5466 a_14142_3526# a_14049_3526# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5467 a_8773_6518# RWL_7 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5468 GND a_11149_4606# a_11093_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5469 a_17529_8116# WWL_1 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5470 WBL_13 WWL_26 a_7762_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5471 a_3553_4358# RWL_15 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5472 a_15503_2738# a_15302_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5473 RBL0_0 RWL_28 a_423_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5474 WBL_29 WWL_31 a_17042_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5475 GND a_802_1636# a_709_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5476 a_5643_7868# a_5442_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5477 a_17473_7058# RWL_5 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5478 VDD a_802_5416# a_709_5416# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5479 a_8249_1096# WWL_27 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5480 WBL_28 WWL_24 a_16462_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5481 VDD a_9502_3526# a_9409_3526# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5482 a_10662_8116# a_10569_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5483 VDD a_1962_4066# a_1869_4066# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5484 WBL_8 WWL_5 a_4862_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5485 a_18403_39# a_18202_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5486 WBL_12 WWL_1 a_7182_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5488 RBL0_17 RWL_24 a_10283_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5489 GND a_15882_2986# a_15789_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5490 a_13993_5438# RWL_11 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5491 a_9989_1636# WWL_25 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5492 a_14722_5956# a_14629_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5493 a_222_2446# a_129_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5494 a_10082_4876# a_9989_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5495 a_1382_1096# a_1289_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5496 WBL_0 WWL_6 a_222_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5497 a_222_6226# a_129_6226# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5498 a_8922_4336# a_8829_4336# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5499 a_73_8408# RWL_0 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5500 a_1382_4876# a_1289_4876# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5501 a_10283_848# a_10082_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5502 a_3702_2176# a_3609_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5503 GND a_1382_7036# a_1289_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5504 a_802_556# a_709_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5505 VDD a_12402_1366# a_12309_1366# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5506 WBL_6 WWL_7 a_3702_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5507 a_5063_1388# a_4862_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5508 a_10863_6788# a_10662_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5509 GND a_3122_3796# a_3029_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5510 WBL_26 WWL_29 a_15302_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5511 a_5442_2716# a_5349_2716# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5512 VDD a_3122_7576# a_3029_7576# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5513 WBL_25 WWL_5 a_14722_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5514 WBL_17 WWL_9 a_10082_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5515 GND a_2449_3796# a_2393_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5516 GND a_5442_4876# a_5349_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5517 a_9409_8386# WWL_0 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5518 RBL0_14 RWL_1 a_8543_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5519 a_8829_7306# WWL_4 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5520 a_4189_6226# WWL_8 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5521 a_6803_1928# a_6602_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5522 GND a_4769_4876# a_4713_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5523 GND a_17042_6496# a_16949_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5524 VDD a_8922_287# a_8829_287# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5525 WBL_24 WWL_17 a_14142_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5526 GND a_16369_6496# a_16313_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5527 a_12889_287# WWL_30 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5528 RBL0_8 RWL_21 a_5063_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5529 a_1233_3008# RWL_20 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5530 GND a_11149_4336# a_11093_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5531 a_8773_6248# RWL_8 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5532 WBL_13 WWL_27 a_7762_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5533 a_3553_4088# RWL_16 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5534 a_15503_2468# a_15302_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5535 a_15882_3796# a_15789_3796# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5536 RBL0_0 RWL_29 a_423_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5537 a_10662_1636# a_10569_1636# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5538 GND a_15882_5956# a_15789_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5539 a_11729_5146# WWL_12 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5540 GND a_802_1366# a_709_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5541 a_5643_7598# a_5442_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5542 GND a_1869_286# a_1813_308# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5543 a_12982_5686# a_12889_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5544 RBL0_26 RWL_17 a_15503_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5545 RBL0_17 RWL_25 a_10283_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5546 a_15302_6766# a_15209_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5547 a_13993_5168# RWL_12 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5548 a_9989_1366# WWL_26 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5549 a_222_2176# a_129_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5550 a_6602_2986# a_6509_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5551 RBL0_30 RWL_13 a_17823_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5552 WBL_15 WWL_14 a_8922_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5553 a_73_8138# RWL_1 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5554 WBL_0 WWL_7 a_222_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5555 RBL0_1 RWL_2 a_1003_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5556 WBL_2 WWL_12 a_1382_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5557 a_10283_578# a_10082_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5558 a_15733_1928# RWL_24 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5559 VDD a_14722_826# a_14629_826# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5560 VDD a_17622_3256# a_17529_3256# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5561 VDD a_12402_1096# a_12309_1096# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5562 WBL_6 WWL_8 a_3702_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5563 a_3122_1366# a_3029_1366# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5564 GND a_8342_5686# a_8249_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5565 GND a_3122_3526# a_3029_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5566 a_7089_7036# WWL_5 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5567 a_1233_5978# RWL_9 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5568 WBL_26 WWL_2 a_15302_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5569 VDD a_3122_7306# a_3029_7306# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5570 GND a_7669_5686# a_7613_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5571 GND a_2449_3526# a_2393_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5572 a_9409_8116# WWL_1 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5573 GND a_9989_6766# a_9933_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5574 a_17042_4066# a_16949_4066# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5575 a_6803_1658# a_6602_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5576 WBL_20 WWL_22 a_11822_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5577 GND a_17042_6226# a_16949_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5578 VDD a_8922_17# a_8829_17# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5579 GND a_16369_6226# a_16313_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5580 a_12889_17# WWL_31 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5581 RBL0_8 RWL_22 a_5063_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5582 WBL_24 WWL_18 a_14142_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5583 RBL0_18 RWL_2 a_10863_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5584 a_13183_1118# a_12982_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5585 GND a_11149_4066# a_11093_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5586 a_13562_2446# a_13469_2446# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5587 a_7613_848# RWL_28 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5588 a_15503_2198# a_15302_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5589 a_16083_39# a_15882_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5590 GND a_13562_4606# a_13469_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5591 a_8543_8408# a_8342_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5592 a_15882_3526# a_15789_3526# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5593 a_16949_7036# WWL_5 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5594 VDD a_13562_8386# a_13469_8386# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5595 a_12309_5956# WWL_9 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5596 GND a_12889_4606# a_12833_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5597 a_11729_4876# WWL_13 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5598 a_6602_5956# a_6509_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5599 RBL0_9 RWL_28 a_5643_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5600 a_16369_3796# WWL_17 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5601 a_17622_6496# a_17529_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5602 a_12982_5416# a_12889_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5603 VDD a_4282_1366# a_4189_1366# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5604 VDD a_8922_2446# a_8829_2446# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5605 RBL0_26 RWL_18 a_15503_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5606 RBL0_17 RWL_26 a_10283_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5607 a_7669_556# WWL_29 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5608 a_9989_1096# WWL_27 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5609 WBL_11 WWL_5 a_6602_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5610 WBL_0 WWL_8 a_222_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5611 a_16313_2738# RWL_21 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5612 RBL0_1 RWL_3 a_1003_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5613 VDD a_12402_287# a_12309_287# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5614 a_15733_1658# RWL_25 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5615 WBL_2 WWL_13 a_1382_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5616 a_13763_7328# a_13562_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5617 VDD a_17622_2986# a_17529_2986# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5618 a_8342_3256# a_8249_3256# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5619 GND a_7762_17# a_7669_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5620 a_3122_1096# a_3029_1096# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5621 WBL_5 WWL_25 a_3122_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5622 GND a_8342_5416# a_8249_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5623 a_6453_7868# RWL_2 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5624 GND a_3122_3256# a_3029_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5625 WBL_9 WWL_21 a_5442_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5626 VDD a_3122_7036# a_3029_7036# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5627 GND a_7669_5416# a_7613_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5628 GND a_2449_3256# a_2393_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5629 WBL_29 WWL_15 a_17042_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5630 a_6803_1388# a_6602_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5631 WBL_20 WWL_23 a_11822_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5632 GND a_4862_3796# a_4769_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5633 VDD a_4862_7576# a_4769_7576# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5634 a_3609_5146# WWL_12 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5635 RBL0_8 RWL_23 a_5063_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5636 RBL0_18 a_4683_7576# a_10863_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5637 a_18403_3008# a_18202_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5638 a_5293_309# RWL_30 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5639 a_13562_2176# a_13469_2176# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5640 a_7613_578# RWL_29 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5641 GND a_18109_2716# a_18053_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5642 a_11673_6788# RWL_6 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5643 GND a_13562_4336# a_13469_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5644 a_8543_8138# a_8342_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5645 RBL0_11 RWL_21 a_6803_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5646 a_2973_3008# RWL_20 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5647 a_4282_4606# a_4189_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5648 VDD a_13562_8116# a_13469_8116# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5649 a_4282_8386# a_4189_8386# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5650 GND a_12889_4336# a_12833_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5651 GND a_18202_17# a_18109_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5652 a_14049_2446# WWL_22 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5653 a_16462_556# a_16369_556# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5654 a_7613_1928# RWL_24 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5655 a_18202_7306# a_18109_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5656 RBL0_9 RWL_29 a_5643_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5657 a_16369_3526# WWL_18 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5658 a_17622_6226# a_17529_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5659 VDD a_8922_2176# a_8829_2176# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5660 a_12982_5146# a_12889_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5661 VDD a_4282_1096# a_4189_1096# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5662 RBL0_26 RWL_19 a_15503_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5663 a_6022_826# a_5929_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5664 a_16313_2468# RWL_22 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5665 VDD a_12402_17# a_12309_17# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5666 a_15733_1388# RWL_26 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5667 a_13763_7058# a_13562_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5668 a_4133_6518# RWL_7 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5669 a_8342_2986# a_8249_2986# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5670 VDD a_6022_7846# a_5929_7846# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5671 WBL_5 WWL_26 a_3122_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5672 GND a_14049_7846# a_13993_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5673 GND a_8342_5146# a_8249_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5674 a_6453_7598# a_4683_7576# RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5675 GND a_15882_826# a_15789_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5676 RBL0_4 RWL_2 a_2743_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5677 a_18403_5978# a_18202_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5678 GND a_7669_5146# a_7613_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5679 a_11093_848# RWL_28 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5680 a_129_5146# WWL_12 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5681 a_4862_1366# a_4769_1366# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5682 GND a_9409_1906# a_9353_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5683 RBL0_13 RWL_20 a_7963_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5684 GND a_709_3796# a_653_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5685 WBL_29 WWL_16 a_17042_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5686 RBL0_23 RWL_0 a_13763_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5687 WBL_20 WWL_24 a_11822_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5688 GND a_4862_3526# a_4769_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5689 a_2973_5978# RWL_9 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5690 VDD a_4862_7306# a_4769_7306# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5691 a_3609_4876# WWL_13 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5692 WBL_12 WWL_28 a_7182_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5693 VDD a_10662_556# a_10569_556# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5694 a_5349_1636# WWL_25 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5695 GND a_11242_2986# a_11149_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5696 a_13562_1906# a_13469_1906# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5697 GND a_18109_2446# a_18053_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5698 WBL_23 WWL_22 a_13562_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5699 a_11149_556# WWL_29 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5700 a_9502_6496# a_9409_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5701 a_7669_2716# WWL_21 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5702 GND a_10569_2986# a_10513_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5703 GND a_13562_4066# a_13469_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5704 a_802_8386# a_709_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5705 a_4282_4336# a_4189_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5706 RBL0_11 RWL_22 a_6803_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5707 a_14923_1118# a_14722_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5709 GND a_12889_4066# a_12833_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5710 a_4282_8116# a_4189_8116# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5711 a_14049_2176# WWL_23 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5712 VDD a_15302_4606# a_15209_4606# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5713 a_7613_1658# RWL_25 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5714 a_18202_7036# a_18109_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5715 VDD a_8922_1906# a_8829_1906# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5716 a_6022_556# a_5929_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5717 GND a_5442_17# a_5349_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5718 a_2163_1928# a_1962_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5719 a_16313_2198# RWL_23 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5720 a_9353_8408# RWL_0 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5721 a_4133_6248# RWL_8 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5722 RBL0_13 RWL_9 a_7963_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5723 WBL_14 WWL_19 a_8342_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5724 a_1289_6766# WWL_6 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5725 GND a_14049_7576# a_13993_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5726 GND a_13562_287# a_13469_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5727 WBL_5 WWL_27 a_3122_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5728 a_16083_4628# a_15882_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5729 GND a_15882_556# a_15789_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5730 GND a_9409_826# a_9353_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5731 RBL0_4 RWL_3 a_2743_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5732 a_11093_578# RWL_29 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5733 GND a_12889_826# a_12833_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5734 a_11242_3796# a_11149_3796# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5735 GND a_11242_5956# a_11149_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5736 a_14629_8386# WWL_0 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5737 a_4862_1096# a_4769_1096# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5738 GND a_9409_1636# a_9353_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5739 a_129_4876# WWL_13 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5740 RBL0_23 RWL_1 a_13763_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5741 VDD a_2542_5956# a_2449_5956# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5742 GND a_10569_5956# a_10513_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5743 GND a_709_3526# a_653_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5744 GND a_4862_3256# a_4769_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5745 VDD a_4862_7036# a_4769_7036# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5746 a_14573_7328# RWL_4 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5747 WBL_8 WWL_30 a_4862_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5748 a_5349_1366# WWL_26 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5749 VDD a_6602_3796# a_6509_3796# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5750 GND a_18109_2176# a_18053_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5751 WBL_23 WWL_23 a_13562_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5752 a_1962_2986# a_1869_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5753 RBL0_22 RWL_13 a_13183_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5754 RBL0_7 RWL_27 a_4483_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5755 a_9502_6226# a_9409_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5756 a_802_8116# a_709_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5757 a_73_308# RWL_30 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5758 RBL0_11 RWL_23 a_6803_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5759 a_4282_4066# a_4189_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5760 WBL_7 WWL_0 a_4282_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5761 RBL0_0 RWL_24 a_423_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5762 a_14049_1906# WWL_24 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5763 VDD a_15302_4336# a_15209_4336# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5764 a_7613_1388# RWL_26 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5765 a_6022_4606# a_5929_4606# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5766 a_12833_309# RWL_30 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5767 GND a_6022_6766# a_5929_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5768 GND a_3029_5686# a_2973_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5769 GND a_5349_6766# a_5293_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5770 a_7383_3818# a_7182_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5771 a_2163_1658# a_1962_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5772 a_15789_2446# WWL_22 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5773 VDD a_11822_2716# a_11729_2716# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5774 a_11822_2986# a_11729_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5775 a_9703_4898# a_9502_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5776 a_12402_7846# a_12309_7846# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5777 a_1003_6788# a_802_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5778 RBL0_18 RWL_30 a_10863_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5779 a_9353_8138# RWL_1 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5780 a_5929_7576# WWL_3 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5781 RBL0_9 RWL_0 a_5643_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5782 a_1289_6496# WWL_7 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5783 WBL_14 WWL_20 a_8342_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5784 a_16462_1906# a_16369_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5785 a_16083_4358# a_15882_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5786 GND a_9409_556# a_9353_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5788 a_16462_5686# a_16369_5686# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5789 GND a_10569_287# a_10513_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5790 GND a_12889_556# a_12833_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5791 a_11242_3526# a_11149_3526# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5792 GND a_16462_7846# a_16369_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5793 a_5873_6518# RWL_7 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5794 a_14629_8116# WWL_1 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5795 VDD a_7762_7846# a_7669_7846# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5796 GND a_15789_7846# a_15733_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5797 a_1962_5956# a_1869_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5799 GND a_9409_1366# a_9353_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5800 GND a_709_3256# a_653_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5801 a_12603_2738# a_12402_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5802 RBL0_27 RWL_10 a_16083_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5803 GND a_129_286# a_73_308# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5804 WBL_8 WWL_31 a_4862_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5805 a_802_1636# a_709_1636# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5806 a_2743_7868# a_2542_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5807 a_14573_7058# RWL_5 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5808 RBL0_31 RWL_6 a_18403_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5809 a_5349_1096# WWL_27 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5810 VDD a_6602_3526# a_6509_3526# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5811 VDD a_7182_4606# a_7089_4606# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5812 WBL_23 WWL_24 a_13562_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5813 RBL0_16 RWL_20 a_9703_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5814 WBL_3 WWL_5 a_1962_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5815 VDD a_18202_5146# a_18109_5146# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5816 WBL_7 WWL_1 a_4282_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5817 a_9933_1118# RWL_27 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5818 GND a_12982_2986# a_12889_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5819 RBL0_0 RWL_25 a_423_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5820 a_11822_5956# a_11729_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5821 a_6022_4336# a_5929_4336# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5822 WBL_25 WWL_28 a_14722_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5823 GND a_3029_5416# a_2973_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5824 VDD a_10082_2446# a_9989_2446# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5825 a_7383_3548# a_7182_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5826 a_2163_1388# a_1962_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5827 a_15789_2176# WWL_23 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5828 a_2542_2716# a_2449_2716# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5829 GND a_2542_4876# a_2449_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5830 a_6509_8386# WWL_0 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5831 RBL0_9 RWL_1 a_5643_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5832 a_5929_7306# WWL_4 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5833 a_1289_6226# WWL_8 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5834 a_8342_826# a_8249_826# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5835 a_3903_1928# a_3702_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5836 GND a_1869_4876# a_1813_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5837 a_16462_1636# a_16369_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5838 a_16083_4088# a_15882_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5839 GND a_14142_6496# a_14049_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5840 a_16462_5416# a_16369_5416# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5841 WBL_19 WWL_17 a_11242_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5842 GND a_16462_7576# a_16369_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5843 GND a_13469_6496# a_13413_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5844 RBL0_3 RWL_21 a_2163_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5845 a_7182_7846# a_7089_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5846 a_5873_6248# RWL_8 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5847 RBL0_16 RWL_9 a_9703_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5848 GND a_15789_7576# a_15733_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5849 a_17823_4628# a_17622_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5850 a_1962_286# a_1869_286# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5851 a_12603_2468# a_12402_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5852 RBL0_27 RWL_11 a_16083_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5853 GND a_12982_5956# a_12889_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5854 a_2743_7598# a_2542_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5855 VDD a_7182_4336# a_7089_4336# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5856 GND a_18202_1096# a_18109_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5857 a_10082_5686# a_9989_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5858 RBL0_21 RWL_17 a_12603_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5859 VDD a_18202_4876# a_18109_4876# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5860 a_8922_5146# a_8829_5146# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5861 GND a_17529_1096# a_17473_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5862 a_12402_6766# a_12309_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5863 RBL0_25 RWL_13 a_14923_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5864 RBL0_0 RWL_26 a_423_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5865 a_3702_2986# a_3609_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5866 WBL_10 WWL_14 a_6022_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5867 GND a_8249_7306# a_8193_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5868 a_12833_1928# RWL_24 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5869 GND a_3029_5146# a_2973_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5870 VDD a_2542_826# a_2449_826# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5871 VDD a_10082_2176# a_9989_2176# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5872 VDD a_14722_3256# a_14629_3256# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5873 a_3029_826# WWL_28 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5874 a_7383_3278# a_7182_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5875 a_15789_1906# WWL_24 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5876 GND a_5442_5686# a_5349_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5877 a_7762_4606# a_7669_4606# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5878 a_4189_7036# WWL_5 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5879 WBL_21 WWL_2 a_12402_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5880 GND a_7762_6766# a_7669_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5881 GND a_4769_5686# a_4713_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5882 GND a_9989_17# a_9933_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5883 a_6022_287# a_5929_287# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5884 a_6509_8116# WWL_1 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5885 a_14142_4066# a_14049_4066# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5886 a_16462_1366# a_16369_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5887 a_3903_1658# a_3702_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5888 GND a_14142_6226# a_14049_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5889 WBL_28 WWL_10 a_16462_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5890 a_3029_2716# WWL_21 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5891 WBL_19 WWL_18 a_11242_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5892 RBL0_12 RWL_14 a_7383_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5893 GND a_13469_6226# a_13413_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5894 RBL0_3 RWL_22 a_2163_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5895 a_7182_7576# a_7089_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5896 a_10283_1118# a_10082_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5897 VDD a_15882_287# a_15789_287# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5898 a_10662_2446# a_10569_2446# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5899 a_17823_4358# a_17622_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5900 a_12603_2198# a_12402_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5901 a_16369_287# WWL_30 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5902 a_8193_3818# RWL_17 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5903 GND a_10662_4606# a_10569_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5904 a_5643_8408# a_5442_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5905 VDD a_10662_8386# a_10569_8386# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5906 VDD a_802_5956# a_709_5956# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5907 RBL0_27 RWL_12 a_16083_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5908 VDD a_9502_4066# a_9409_4066# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5909 a_3702_5956# a_3609_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5910 RBL0_30 RWL_10 a_17823_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5911 a_8922_1096# a_8829_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5912 VDD a_222_2716# a_129_2716# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5913 a_13469_3796# WWL_17 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5914 a_14722_6496# a_14629_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5915 a_10082_5416# a_9989_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5916 VDD a_1382_1366# a_1289_1366# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5917 a_222_2986# a_129_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5918 RBL0_21 RWL_18 a_12603_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5919 a_8922_4876# a_8829_4876# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5920 WBL_6 WWL_5 a_3702_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5921 GND a_8249_7036# a_8193_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5922 a_13413_2738# RWL_21 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5923 a_12833_1658# RWL_25 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5924 a_10863_7328# a_10662_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5925 VDD a_14722_2986# a_14629_2986# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5926 VDD a_10082_1906# a_9989_1906# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5927 a_5442_3256# a_5349_3256# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5928 GND a_5442_5416# a_5349_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5929 a_3553_7868# RWL_2 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5930 a_7762_4336# a_7669_4336# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5931 a_8829_7846# WWL_2 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5932 VDD a_18202_826# a_18109_826# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5933 WBL_4 WWL_21 a_2542_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5934 GND a_4769_5416# a_4713_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5935 a_6022_17# a_5929_17# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5936 WBL_24 WWL_15 a_14142_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5937 a_3903_1388# a_3702_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5938 GND a_1962_3796# a_1869_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5939 a_8249_4606# WWL_14 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5940 VDD a_1962_7576# a_1869_7576# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5941 WBL_28 WWL_11 a_16462_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5942 a_9502_826# a_9409_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5943 RBL0_12 RWL_15 a_7383_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5944 RBL0_3 RWL_23 a_2163_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5945 WBL_18 WWL_29 a_10662_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5946 a_15503_3008# a_15302_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5947 a_10662_2176# a_10569_2176# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5948 a_17823_4088# a_17622_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5949 GND a_15882_6496# a_15789_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5950 VDD a_15882_17# a_15789_17# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5951 GND a_15209_2716# a_15153_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5952 a_16369_17# WWL_31 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5953 a_8193_3548# RWL_18 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5954 GND a_10662_4336# a_10569_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5955 a_222_5956# a_129_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5956 a_5643_8138# a_5442_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5957 RBL0_6 RWL_21 a_3903_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5958 a_1382_4606# a_1289_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5959 VDD a_10662_8116# a_10569_8116# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5960 a_1382_8386# a_1289_8386# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5961 a_11149_2446# WWL_22 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5962 a_4282_556# a_4189_556# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5963 a_4713_1928# RWL_24 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5964 a_15302_7306# a_15209_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5965 RBL0_30 RWL_11 a_17823_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5966 a_13469_3526# WWL_18 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5967 a_5063_4898# a_4862_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5968 a_14722_6226# a_14629_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5969 a_10082_5146# a_9989_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5970 VDD a_1382_1096# a_1289_1096# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5971 RBL0_21 RWL_19 a_12603_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5972 WBL_15 WWL_12 a_8922_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5973 RBL0_1 RWL_0 a_1003_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5974 WBL_0 WWL_5 a_222_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5975 RBL0_15 RWL_28 a_9123_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5976 GND a_7669_17# a_7613_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5977 a_13413_2468# RWL_22 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5978 a_12833_1388# RWL_26 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5979 a_10863_7058# a_10662_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5980 a_1233_6518# RWL_7 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5981 a_5442_2986# a_5349_2986# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5982 VDD a_3122_7846# a_3029_7846# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5983 GND a_11149_7846# a_11093_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5984 GND a_5442_5146# a_5349_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5985 a_3553_7598# RWL_3 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5986 WBL_13 WWL_14 a_7762_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5987 GND a_9989_7306# a_9933_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5988 a_15503_5978# a_15302_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5989 GND a_4769_5146# a_4713_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5990 RBL0_18 RWL_0 a_10863_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5991 GND a_6509_1906# a_6453_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5992 RBL0_8 RWL_20 a_5063_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5993 WBL_24 WWL_16 a_14142_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5994 GND a_802_4876# a_709_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5995 a_7182_287# a_7089_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5996 GND a_1962_3526# a_1869_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5997 a_9502_556# a_9409_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5998 RBL0_12 RWL_16 a_7383_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5999 VDD a_1962_7306# a_1869_7306# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6000 a_15882_4066# a_15789_4066# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6001 a_2449_1636# WWL_25 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6002 a_10662_1906# a_10569_1906# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6003 GND a_15209_2446# a_15153_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6004 WBL_18 WWL_22 a_10662_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6005 GND a_15882_6226# a_15789_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6006 GND a_18109_17# a_18053_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6007 a_8193_3278# RWL_19 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6008 a_6602_6496# a_6509_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6009 a_4769_2716# WWL_21 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6010 GND a_10662_4066# a_10569_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6011 RBL0_6 RWL_22 a_3903_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6012 a_1382_4336# a_1289_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6013 a_12023_1118# a_11822_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6014 a_1382_8116# a_1289_8116# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6015 VDD a_17622_6766# a_17529_6766# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6016 a_16369_4336# WWL_15 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6017 a_11149_2176# WWL_23 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6018 VDD a_12402_4606# a_12309_4606# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6019 a_4282_286# a_4189_286# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6020 a_4713_1658# RWL_25 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6021 a_2973_848# RWL_28 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6022 a_15302_7036# a_15209_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6023 RBL0_30 RWL_12 a_17823_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6024 WBL_15 WWL_13 a_8922_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6025 RBL0_1 RWL_1 a_1003_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6026 a_11093_1118# RWL_27 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6027 a_17042_3796# a_16949_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6028 RBL0_15 RWL_29 a_9123_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6029 a_17042_7576# a_16949_7576# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6030 a_13413_2198# RWL_23 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6031 a_12982_826# a_12889_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6032 a_6453_8408# RWL_0 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6033 a_1233_6248# RWL_8 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6034 RBL0_8 RWL_9 a_5063_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6035 WBL_9 WWL_19 a_5442_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6036 GND a_11149_7576# a_11093_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6037 a_13183_4628# a_12982_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6038 GND a_9989_7036# a_9933_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6039 a_11729_8386# WWL_0 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6040 GND a_7089_2716# a_7033_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6041 GND a_6509_1636# a_6453_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6042 RBL0_18 RWL_1 a_10863_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6043 GND a_1962_3256# a_1869_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6044 VDD a_1962_7036# a_1869_7036# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6045 a_11673_7328# RWL_4 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6046 a_2449_1366# WWL_26 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6047 VDD a_3702_3796# a_3609_3796# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6048 RBL0_2 RWL_27 a_1583_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6049 GND a_15209_2176# a_15153_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6050 WBL_18 WWL_23 a_10662_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6051 RBL0_17 RWL_13 a_10283_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6052 a_9989_4606# WWL_14 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6053 a_6602_6226# a_6509_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6054 RBL0_6 RWL_23 a_3903_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6055 a_1382_4066# a_1289_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6056 VDD a_14142_556# a_14049_556# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6057 GND a_17622_2716# a_17529_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6058 WBL_2 WWL_0 a_1382_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6059 VDD a_17622_6496# a_17529_6496# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6060 a_16369_4066# WWL_16 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6061 GND a_16949_2716# a_16893_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6062 a_8342_6766# a_8249_6766# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6063 a_11149_1906# WWL_24 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6064 VDD a_12402_4336# a_12309_4336# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6065 GND a_5349_17# a_5293_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6066 a_4282_16# a_4189_16# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6067 a_4713_1388# RWL_26 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6068 a_3122_4606# a_3029_4606# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6069 GND a_3122_6766# a_3029_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6070 a_2973_578# RWL_29 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6071 GND a_2449_6766# a_2393_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6072 a_16313_3008# RWL_20 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6073 a_17042_3526# a_16949_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6074 a_4483_3818# a_4282_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6075 a_12889_2446# WWL_22 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6076 a_17042_7306# a_16949_7306# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6077 a_6803_4898# a_6602_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6078 WBL_20 WWL_10 a_11822_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6079 GND a_14049_8386# a_13993_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6080 a_11822_556# a_11729_556# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6081 a_6453_8138# RWL_1 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6082 a_12982_556# a_12889_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6083 RBL0_4 RWL_0 a_2743_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6084 a_18403_6518# a_18202_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6085 WBL_9 WWL_20 a_5442_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6086 a_13562_1906# a_13469_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6087 a_13183_4358# a_12982_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6088 a_16893_39# RWL_31 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6089 a_13562_5686# a_13469_5686# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6090 RBL0_28 RWL_28 a_16663_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6091 GND a_13562_7846# a_13469_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6092 GND a_17042_287# a_16949_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6093 a_2973_6518# RWL_7 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6094 a_11729_8116# WWL_1 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6095 VDD a_4862_7846# a_4769_7846# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6096 GND a_12889_7846# a_12833_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6097 GND a_6509_1366# a_6453_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6098 GND a_7089_2446# a_7033_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6099 GND a_16369_826# a_16313_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6100 RBL0_22 RWL_10 a_13183_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6101 GND a_8922_1906# a_8829_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6102 GND a_18109_2986# a_18053_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6103 VDD a_8922_5686# a_8829_5686# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6104 a_7669_3256# WWL_19 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6105 a_11673_7058# RWL_5 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6106 RBL0_26 RWL_6 a_15503_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6107 a_2449_1096# WWL_27 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6108 VDD a_3702_3526# a_3609_3526# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6109 VDD a_4282_4606# a_4189_4606# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6110 WBL_18 WWL_24 a_10662_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6111 RBL0_11 RWL_20 a_6803_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6112 a_18202_1366# a_18109_1366# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6113 VDD a_15302_5146# a_15209_5146# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6114 a_14722_287# a_14629_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6115 GND a_17622_2446# a_17529_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6116 WBL_2 WWL_1 a_1382_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6117 a_16313_5978# RWL_9 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6118 a_15733_4898# RWL_13 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6119 a_8342_2716# a_8249_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6120 VDD a_17622_6226# a_17529_6226# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6121 a_8342_6496# a_8249_6496# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6122 GND a_16949_2446# a_16893_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6123 WBL_4 WWL_28 a_2542_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6124 a_3122_4336# a_3029_4336# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6125 a_9703_5708# a_9502_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6126 a_17042_3256# a_16949_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6127 a_4483_3548# a_4282_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6128 a_12889_2176# WWL_23 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6129 WBL_29 WWL_3 a_17042_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6130 a_17042_7036# a_16949_7036# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6131 RBL0_13 RWL_7 a_7963_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6132 WBL_20 WWL_11 a_11822_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6133 GND a_14049_8116# a_13993_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6134 a_3609_8386# WWL_0 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6135 RBL0_4 RWL_1 a_2743_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6136 a_18403_6248# a_18202_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6137 a_13562_1636# a_13469_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6138 a_13183_4088# a_12982_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6139 GND a_11242_6496# a_11149_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6140 GND a_18109_5956# a_18053_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6141 a_13562_5416# a_13469_5416# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6142 RBL0_28 RWL_29 a_16663_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6143 GND a_13562_7576# a_13469_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6144 GND a_10569_6496# a_10513_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6145 a_2973_6248# RWL_8 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6146 a_4282_7846# a_4189_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6147 RBL0_11 RWL_9 a_6803_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6148 GND a_12889_7576# a_12833_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6149 GND a_14049_287# a_13993_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6150 GND a_7089_2176# a_7033_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6151 a_423_1118# a_222_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6152 a_14923_4628# a_14722_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6153 GND a_16369_556# a_16313_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6154 a_6509_826# WWL_28 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6155 a_802_2446# a_709_2446# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6156 a_14049_5686# WWL_10 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6157 RBL0_22 RWL_11 a_13183_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6158 GND a_8922_1636# a_8829_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6159 VDD a_8922_5416# a_8829_5416# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6160 a_7669_2986# WWL_20 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6161 VDD a_4282_4336# a_4189_4336# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6162 GND a_15302_1096# a_15209_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6163 a_9502_287# a_9409_287# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6164 a_18202_1096# a_18109_1096# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6165 WBL_31 WWL_25 a_18202_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6166 VDD a_15302_4876# a_15209_4876# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6167 a_6022_5146# a_5929_5146# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6168 GND a_14629_1096# a_14573_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6169 GND a_17622_2176# a_17529_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6170 a_8342_2446# a_8249_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6171 GND a_6022_7306# a_5929_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6172 a_8342_6226# a_8249_6226# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6173 GND a_16949_2176# a_16893_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6174 WBL_14 WWL_6 a_8342_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6175 WBL_5 WWL_14 a_3122_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6176 GND a_5349_7306# a_5293_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6177 VDD a_11822_3256# a_11729_3256# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6178 a_9703_5438# a_9502_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6179 a_1003_7328# a_802_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6180 a_4483_3278# a_4282_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6181 a_12889_1906# WWL_24 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6182 GND a_2542_5686# a_2449_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6183 a_14573_39# RWL_31 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6184 a_129_8386# WWL_0 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6185 WBL_29 WWL_4 a_17042_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6186 a_4862_4606# a_4769_4606# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6187 a_1289_7036# WWL_5 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6188 RBL0_13 RWL_8 a_7963_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6189 GND a_4862_6766# a_4769_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6190 GND a_1869_5686# a_1813_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6191 a_3609_8116# WWL_1 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6192 a_11242_4066# a_11149_4066# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6193 GND a_16462_8386# a_16369_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6194 a_13562_1366# a_13469_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6195 GND a_11242_6226# a_11149_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6196 WBL_23 WWL_10 a_13562_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6197 GND a_15789_8386# a_15733_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6198 a_1962_6496# a_1869_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6199 RBL0_7 RWL_14 a_4483_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6200 GND a_10569_6226# a_10513_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6201 a_15302_826# a_15209_826# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6202 a_4282_7576# a_4189_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6203 a_14923_4358# a_14722_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6204 a_5293_3818# RWL_17 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6205 a_802_2176# a_709_2176# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6206 a_2743_8408# a_2542_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6207 RBL0_31 RWL_4 a_18403_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6208 a_14049_5416# WWL_11 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6209 VDD a_7182_5146# a_7089_5146# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6210 VDD a_6602_4066# a_6509_4066# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6211 RBL0_22 RWL_12 a_13183_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6212 GND a_8922_1366# a_8829_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6213 a_7613_4898# RWL_13 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6214 a_5643_848# a_5442_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6215 a_9502_17# a_9409_17# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6216 WBL_31 WWL_26 a_18202_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6217 RBL0_25 RWL_10 a_14923_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6218 a_6022_1096# a_5929_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6219 a_10569_3796# WWL_17 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6220 a_11822_6496# a_11729_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6221 a_6022_4876# a_5929_4876# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6222 a_8342_2176# a_8249_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6223 GND a_6022_7036# a_5929_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6224 WBL_14 WWL_7 a_8342_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6225 a_16083_7868# a_15882_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6226 GND a_5349_7036# a_5293_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6227 a_10513_2738# RWL_21 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6228 VDD a_11822_2986# a_11729_2986# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6229 a_9703_5168# a_9502_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6230 a_1003_7058# a_802_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6231 a_2542_3256# a_2449_3256# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6232 GND a_2542_5416# a_2449_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6233 a_129_8116# WWL_1 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6234 a_5929_7846# WWL_2 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6235 VDD a_6022_826# a_5929_826# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6236 a_4862_4336# a_4769_4336# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6237 GND a_9409_4876# a_9353_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6238 GND a_709_6766# a_653_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6239 GND a_1869_5416# a_1813_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6240 a_16462_5956# a_16369_5956# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6241 WBL_19 WWL_15 a_11242_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6242 GND a_16462_8116# a_16369_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6243 a_7182_8386# a_7089_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6244 RBL0_16 RWL_7 a_9703_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6245 WBL_23 WWL_11 a_13562_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6246 a_5349_4606# WWL_14 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6247 GND a_15789_8116# a_15733_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6248 a_1962_6226# a_1869_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6249 RBL0_7 RWL_15 a_4483_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6250 a_12982_287# a_12889_287# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6251 a_12603_3008# a_12402_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6252 a_14923_4088# a_14722_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6253 GND a_12982_6496# a_12889_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6254 GND a_7182_1096# a_7089_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6255 GND a_12309_2716# a_12253_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6256 a_9933_4628# RWL_14 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6257 a_802_1906# a_709_1906# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6258 a_5293_3548# RWL_18 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6259 a_2743_8138# a_2542_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6260 RBL0_31 RWL_5 a_18403_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6261 WBL_1 WWL_22 a_802_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6262 VDD a_7182_4876# a_7089_4876# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6263 a_5643_578# a_5442_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6264 a_15789_5686# WWL_10 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6265 WBL_31 WWL_27 a_18202_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6266 a_1813_1928# RWL_24 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6267 a_12402_7306# a_12309_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6268 RBL0_25 RWL_11 a_14923_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6269 a_10569_3526# WWL_18 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6270 a_2163_4898# a_1962_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6271 a_11822_6226# a_11729_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6272 WBL_10 WWL_12 a_6022_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6273 a_12253_39# RWL_31 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6274 WBL_14 WWL_8 a_8342_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6275 a_16083_7598# a_15882_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6276 a_10513_2468# RWL_22 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6277 GND a_3702_286# a_3609_286# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6278 a_7762_5146# a_7669_5146# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6279 VDD a_802_556# a_709_556# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6280 a_2542_2986# a_2449_2986# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6281 GND a_7762_7306# a_7669_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6282 WBL_1 WWL_28 a_802_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6283 GND a_2542_5146# a_2449_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6284 a_12603_5978# a_12402_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6285 GND a_1869_5146# a_1813_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6286 VDD a_16462_1636# a_16369_1636# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6287 a_3029_3256# WWL_19 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6288 WBL_19 WWL_16 a_11242_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6289 GND a_3609_1906# a_3553_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6290 RBL0_3 RWL_20 a_2163_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6291 a_7182_8116# a_7089_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6292 RBL0_16 RWL_8 a_9703_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6293 RBL0_7 RWL_16 a_4483_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6294 a_12982_17# a_12889_17# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6295 GND a_18202_4606# a_18109_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6296 VDD a_18202_8386# a_18109_8386# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6297 GND a_17529_4606# a_17473_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6298 GND a_12982_6226# a_12889_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6299 GND a_12309_2446# a_12253_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6300 a_9933_4358# RWL_15 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6301 a_5293_3278# RWL_19 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6302 a_3702_6496# a_3609_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6303 WBL_24 WWL_29 a_14142_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6304 WBL_1 WWL_23 a_802_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6305 a_1869_2716# WWL_21 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6306 RBL0_0 RWL_13 a_423_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6307 GND a_10082_1906# a_9989_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6308 a_5063_5708# a_4862_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6309 VDD a_14722_6766# a_14629_6766# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6310 VDD a_222_3256# a_129_3256# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6311 a_13469_4336# WWL_15 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6312 VDD a_10082_5686# a_9989_5686# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6313 a_7383_6788# a_7182_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6314 a_15789_5416# WWL_11 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6315 a_1813_1658# RWL_25 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6316 a_12402_7036# a_12309_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6317 RBL0_25 RWL_12 a_14923_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6318 a_11729_287# WWL_30 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6319 WBL_10 WWL_13 a_6022_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6320 RBL0_28 RWL_24 a_16663_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6321 a_14142_3796# a_14049_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6322 a_14142_7576# a_14049_7576# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6323 a_10513_2198# RWL_23 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6324 a_16462_4876# a_16369_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6325 a_7762_1096# a_7669_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6326 a_3553_8408# RWL_0 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6327 a_7762_4876# a_7669_4876# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6328 RBL0_3 RWL_9 a_2163_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6329 VDD a_802_286# a_709_286# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6330 WBL_4 WWL_19 a_2542_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6331 GND a_7762_7036# a_7669_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6332 a_10283_4628# a_10082_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6333 a_17823_7868# a_17622_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6334 a_18109_556# WWL_29 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6335 GND a_9502_3796# a_9409_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6336 GND a_802_5686# a_709_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6337 a_7182_1636# a_7089_1636# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6338 VDD a_9502_7576# a_9409_7576# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6339 a_8249_5146# WWL_12 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6340 GND a_7182_826# a_7089_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6341 WBL_28 WWL_9 a_16462_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6342 GND a_4189_2716# a_4133_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6343 a_3029_2986# WWL_20 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6344 GND a_8829_3796# a_8773_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6345 GND a_3609_1636# a_3553_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6346 GND a_18202_4336# a_18109_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6347 a_8922_4606# a_8829_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6348 VDD a_18202_8116# a_18109_8116# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6349 a_222_6496# a_129_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6350 WBL_27 WWL_21 a_15882_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6351 GND a_17529_4336# a_17473_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6352 a_8922_8386# a_8829_8386# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6353 GND a_12309_2176# a_12253_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6354 a_9933_4088# RWL_16 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6355 a_3702_6226# a_3609_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6356 WBL_1 WWL_24 a_802_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6357 a_4862_826# a_4769_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6358 GND a_14722_2716# a_14629_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6359 GND a_10082_1636# a_9989_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6360 VDD a_14722_6496# a_14629_6496# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6361 a_5063_5438# a_4862_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6362 VDD a_222_2986# a_129_2986# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6363 a_13469_4066# WWL_16 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6364 VDD a_10082_5416# a_9989_5416# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6365 a_5442_6766# a_5349_6766# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6366 a_1813_1388# RWL_26 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6367 a_11729_17# WWL_31 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6368 a_13413_3008# RWL_20 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6369 RBL0_28 RWL_25 a_16663_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6370 RBL0_29 RWL_21 a_17243_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6371 a_14142_3526# a_14049_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6372 a_1583_3818# a_1382_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6373 a_6453_848# RWL_28 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6374 a_14142_7306# a_14049_7306# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6375 a_3903_4898# a_3702_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6376 GND a_11149_8386# a_11093_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6377 a_3553_8138# RWL_1 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6378 RBL0_12 RWL_2 a_7383_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6379 WBL_13 WWL_12 a_7762_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6380 VDD a_802_16# a_709_16# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6381 a_15503_6518# a_15302_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6382 WBL_4 WWL_20 a_2542_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6383 a_10662_1906# a_10569_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6384 a_10283_4358# a_10082_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6385 a_17823_7598# a_17622_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6386 a_10662_5686# a_10569_5686# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6387 RBL0_7 RWL_28 a_4483_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6388 GND a_802_5416# a_709_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6389 GND a_9502_3526# a_9409_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6390 GND a_10662_7846# a_10569_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6391 a_1583_308# a_1382_286# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6392 VDD a_9502_7306# a_9409_7306# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6393 GND a_7182_556# a_7089_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6394 a_8249_4876# WWL_13 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6395 VDD a_1962_7846# a_1869_7846# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6396 GND a_4189_2446# a_4133_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6397 GND a_8829_3526# a_8773_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6398 GND a_3609_1366# a_3553_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6399 GND a_4189_826# a_4133_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6400 RBL0_17 RWL_10 a_10283_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6401 GND a_15209_2986# a_15153_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6402 GND a_18202_4066# a_18109_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6403 a_222_6226# a_129_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6404 a_4769_3256# WWL_19 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6405 a_8922_4336# a_8829_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6406 RBL0_21 RWL_6 a_12603_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6407 RBL0_6 RWL_20 a_3903_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6408 GND a_17529_4066# a_17473_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6409 VDD a_1382_4606# a_1289_4606# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6410 a_8922_8116# a_8829_8116# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6411 a_15302_1366# a_15209_1366# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6412 VDD a_12402_5146# a_12309_5146# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6413 a_13413_5978# RWL_9 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6414 a_4862_556# a_4769_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6415 GND a_14722_2446# a_14629_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6416 GND a_10082_1366# a_9989_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6417 RBL0_14 RWL_24 a_8543_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6418 a_12833_4898# RWL_13 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6419 VDD a_14722_6226# a_14629_6226# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6420 a_5063_5168# a_4862_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6421 RBL0_30 RWL_30 a_17823_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6422 a_5442_2716# a_5349_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6423 a_5442_6496# a_5349_6496# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6424 RBL0_31 RWL_31 a_18403_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6425 GND a_8922_287# a_8829_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6426 a_6803_5708# a_6602_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6427 a_18109_2716# WWL_21 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6428 RBL0_28 RWL_26 a_16663_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6429 RBL0_29 RWL_22 a_17243_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6430 a_14142_3256# a_14049_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6431 a_1583_3548# a_1382_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6432 a_6453_578# RWL_29 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6433 a_14142_7036# a_14049_7036# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6434 WBL_24 WWL_3 a_14142_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6435 RBL0_8 RWL_7 a_5063_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6436 GND a_11149_8116# a_11093_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6437 RBL0_12 a_4683_7576# a_7383_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6438 WBL_13 WWL_13 a_7762_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6439 a_15503_6248# a_15302_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6440 a_15882_3796# a_15789_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6441 a_10662_1636# a_10569_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6442 a_10283_4088# a_10082_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6443 a_15882_7576# a_15789_7576# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6444 GND a_15209_5956# a_15153_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6445 a_10662_5416# a_10569_5416# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6446 RBL0_7 RWL_29 a_4483_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6447 a_8193_6788# RWL_6 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6448 GND a_9502_3256# a_9409_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6449 GND a_10662_7576# a_10569_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6450 GND a_802_5146# a_709_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6451 a_1382_7846# a_1289_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6452 VDD a_9502_7036# a_9409_7036# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6453 RBL0_6 RWL_9 a_3903_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6454 GND a_8829_3256# a_8773_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6455 GND a_4189_2176# a_4133_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6456 a_12023_4628# a_11822_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6457 GND a_4189_556# a_4133_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6458 a_11149_5686# WWL_10 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6459 a_73_1928# RWL_24 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6460 RBL0_17 RWL_11 a_10283_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6461 a_9989_5146# WWL_12 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6462 a_4769_2986# WWL_20 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6463 a_8922_4066# a_8829_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6464 VDD a_1382_4336# a_1289_4336# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6465 WBL_15 WWL_0 a_8922_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6466 GND a_14722_826# a_14629_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6467 a_15733_5708# RWL_10 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6468 GND a_12402_1096# a_12309_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6469 a_11093_4628# RWL_14 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6470 a_15302_1096# a_15209_1096# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6471 WBL_26 WWL_25 a_15302_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6472 VDD a_12402_4876# a_12309_4876# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6473 GND a_11729_1096# a_11673_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6474 GND a_14722_2176# a_14629_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6475 a_3122_5146# a_3029_5146# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6476 a_709_3796# WWL_17 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6477 RBL0_14 RWL_25 a_8543_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6478 a_5442_2446# a_5349_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6479 GND a_3122_7306# a_3029_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6480 a_5442_6226# a_5349_6226# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6481 WBL_9 WWL_6 a_5442_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6482 GND a_2449_7306# a_2393_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6483 VDD a_17042_3796# a_16949_3796# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6484 a_17042_7846# a_16949_7846# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6485 a_6803_5438# a_6602_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6486 WBL_10 WWL_28 a_6022_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6487 RBL0_29 RWL_23 a_17243_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6488 a_1583_3278# a_1382_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6489 GND a_5929_287# a_5873_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6490 WBL_24 WWL_4 a_14142_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6491 RBL0_8 RWL_8 a_5063_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6492 RBL0_9 RWL_31 a_5643_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6493 GND a_1962_6766# a_1869_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6494 a_15882_3526# a_15789_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6495 GND a_13562_8386# a_13469_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6496 a_10662_1366# a_10569_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6497 a_15882_7306# a_15789_7306# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6498 WBL_18 WWL_10 a_10662_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6499 GND a_7089_2986# a_7033_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6500 GND a_12889_8386# a_12833_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6501 a_17243_2738# a_17042_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6502 RBL0_2 RWL_14 a_1583_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6503 a_1382_7576# a_1289_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6504 a_12023_4358# a_11822_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6505 a_2393_3818# RWL_17 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6506 a_16369_7576# WWL_3 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6507 a_73_1658# RWL_25 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6508 RBL0_26 RWL_4 a_15503_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6509 a_11149_5416# WWL_11 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6510 VDD a_4282_5146# a_4189_5146# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6511 VDD a_3702_4066# a_3609_4066# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6512 RBL0_17 RWL_12 a_10283_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6513 a_4713_4898# RWL_13 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6514 a_9989_4876# WWL_13 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6515 GND a_12402_287# a_12309_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6516 WBL_15 WWL_1 a_8922_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6517 GND a_14722_556# a_14629_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6518 RBL0_27 RWL_31 a_16083_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6519 GND a_17622_2986# a_17529_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6520 a_16313_6518# RWL_7 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6521 a_15733_5438# RWL_11 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6522 WBL_26 WWL_26 a_15302_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6523 a_11093_4358# RWL_15 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6524 a_3122_1096# a_3029_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6525 GND a_11729_826# a_11673_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6526 GND a_16949_2986# a_16893_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6527 a_709_3526# WWL_18 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6528 a_3122_4876# a_3029_4876# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6529 RBL0_14 RWL_26 a_8543_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6530 a_5442_2176# a_5349_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6531 GND a_3122_7036# a_3029_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6532 a_2393_38# RWL_31 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6533 WBL_9 WWL_7 a_5442_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6534 a_13183_7868# a_12982_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6535 GND a_2449_7036# a_2393_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6536 VDD a_17042_3526# a_16949_3526# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6537 a_6803_5168# a_6602_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6538 WBL_20 WWL_9 a_11822_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6539 GND a_7089_5956# a_7033_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6540 GND a_6509_4876# a_6453_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6541 a_8543_1928# a_8342_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6542 a_6803_309# a_6602_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6543 GND a_18109_6496# a_18053_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6544 a_13562_5956# a_13469_5956# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6545 a_15882_3256# a_15789_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6546 GND a_13562_8116# a_13469_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6547 a_7669_6766# WWL_6 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6548 a_15882_7036# a_15789_7036# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6549 a_4282_8386# a_4189_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6550 RBL0_11 RWL_7 a_6803_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6551 WBL_18 WWL_11 a_10662_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6552 a_2449_4606# WWL_14 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6553 GND a_12889_8116# a_12833_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6554 a_17243_2468# a_17042_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6555 RBL0_2 RWL_15 a_1583_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6556 a_17622_3796# a_17529_3796# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6557 a_12982_2716# a_12889_2716# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6558 GND a_17622_5956# a_17529_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6559 a_7613_5708# RWL_10 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6560 a_12023_4088# a_11822_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6561 GND a_4282_1096# a_4189_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6562 a_16369_7306# WWL_4 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6563 VDD a_8922_5956# a_8829_5956# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6564 a_73_1388# RWL_26 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6565 a_2393_3548# RWL_18 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6566 RBL0_26 RWL_5 a_15503_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6567 GND a_16949_5956# a_16893_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6568 VDD a_4282_4876# a_4189_4876# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6569 a_2393_308# RWL_30 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6570 VDD a_7182_287# a_7089_287# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6571 a_16313_6248# RWL_8 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6572 a_15733_5168# RWL_12 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6574 a_17042_6766# a_16949_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6575 a_12889_5686# WWL_10 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6576 WBL_26 WWL_27 a_15302_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6577 VDD a_8342_2716# a_8249_2716# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6578 a_8342_2986# a_8249_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6579 a_11093_4088# RWL_16 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6580 GND a_11729_556# a_11673_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6581 a_1869_826# WWL_28 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6582 WBL_5 WWL_12 a_3122_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6583 a_12603_848# a_12402_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6584 WBL_9 WWL_8 a_5442_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6585 a_17622_17# a_17529_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6586 a_13183_7598# a_12982_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6587 a_4862_287# a_4769_287# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6588 WBL_29 WWL_2 a_17042_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6589 GND a_9409_5686# a_9353_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6590 a_4862_5146# a_4769_5146# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6591 GND a_4862_7306# a_4769_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6592 a_9123_2738# a_8922_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6593 a_8543_1658# a_8342_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6594 a_423_4628# a_222_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6595 VDD a_13562_1636# a_13469_1636# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6596 GND a_18109_6226# a_18053_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6597 a_7669_6496# WWL_7 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6598 a_4282_8116# a_4189_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6599 RBL0_11 RWL_8 a_6803_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6600 a_17243_2198# a_17042_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6601 RBL0_2 RWL_16 a_1583_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6602 GND a_15302_4606# a_15209_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6603 a_18202_4606# a_18109_4606# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6604 a_17622_3526# a_17529_3526# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6605 VDD a_15302_8386# a_15209_8386# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6606 a_14049_5956# WWL_9 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6607 GND a_129_1096# a_73_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6608 GND a_14629_4606# a_14573_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6609 a_8342_5956# a_8249_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6610 a_7613_5438# RWL_11 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6611 WBL_3 WWL_29 a_1962_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6612 a_2393_3278# RWL_19 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6613 VDD a_7182_17# a_7089_17# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6614 a_2163_5708# a_1962_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6615 VDD a_11822_6766# a_11729_6766# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6616 VDD a_6022_1366# a_5929_1366# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6617 a_10569_4336# WWL_15 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6618 a_10662_826# a_10569_826# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6619 a_4483_6788# a_4282_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6620 a_12889_5416# WWL_11 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6621 WBL_14 WWL_5 a_8342_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6622 a_18053_2738# RWL_21 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6623 WBL_5 WWL_13 a_3122_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6624 a_16083_8408# a_15882_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6625 a_10283_309# a_10082_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6626 RBL0_23 RWL_24 a_13763_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6627 a_11242_3796# a_11149_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6628 a_12603_578# a_12402_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6629 a_11242_7576# a_11149_7576# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6630 a_17529_826# WWL_28 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6631 a_13562_4876# a_13469_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6632 a_4862_1096# a_4769_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6633 a_4862_17# a_4769_17# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6634 GND a_9409_5416# a_9353_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6635 a_4862_4876# a_4769_4876# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6636 GND a_709_7306# a_653_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6637 GND a_4862_7036# a_4769_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6638 VDD a_16462_2446# a_16369_2446# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6639 a_4862_17# a_4769_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6640 a_14923_7868# a_14722_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6641 a_8543_1388# a_8342_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6642 a_802_1906# a_709_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6643 a_9123_2468# a_8922_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6644 a_423_4358# a_222_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6645 GND a_6602_3796# a_6509_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6646 a_802_5686# a_709_5686# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6647 a_9502_3796# a_9409_3796# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6648 a_4282_1636# a_4189_1636# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6649 VDD a_6602_7576# a_6509_7576# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6650 WBL_23 WWL_9 a_13562_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6651 a_5349_5146# WWL_12 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6652 GND a_5929_3796# a_5873_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6653 GND a_1289_2716# a_1233_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6654 GND a_8922_4876# a_8829_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6655 a_7669_6226# WWL_8 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6656 GND a_15302_4336# a_15209_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6657 a_18202_4336# a_18109_4336# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6658 RBL0_15 RWL_17 a_9123_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6659 WBL_30 WWL_17 a_17622_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6660 a_6022_4606# a_5929_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6661 VDD a_15302_8116# a_15209_8116# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6662 RBL0_0 RWL_10 a_423_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6663 WBL_22 WWL_21 a_12982_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6664 GND a_14629_4336# a_14573_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6665 a_6022_8386# a_5929_8386# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6666 a_7613_5168# RWL_12 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6667 WBL_3 WWL_30 a_1962_286# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6668 a_9353_1928# RWL_24 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6669 GND a_11822_2716# a_11729_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6670 a_653_3818# RWL_17 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6671 a_2163_5438# a_1962_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6672 VDD a_11822_6496# a_11729_6496# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6673 VDD a_6022_1096# a_5929_1096# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6674 a_10569_4066# WWL_16 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6675 a_2542_6766# a_2449_6766# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6676 a_9989_556# WWL_29 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6677 a_18053_2468# RWL_22 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6678 a_16083_8138# a_15882_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6679 a_16462_5686# a_16369_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6680 RBL0_24 RWL_21 a_14343_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6681 a_10513_3008# RWL_20 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6682 VDD a_14722_287# a_14629_287# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6683 RBL0_23 RWL_25 a_13763_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6684 a_11242_3526# a_11149_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6685 a_11242_7306# a_11149_7306# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6686 RBL0_7 RWL_2 a_4483_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6687 GND a_709_7036# a_653_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6688 GND a_9409_5146# a_9353_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6689 a_12603_6518# a_12402_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6690 VDD a_16462_2176# a_16369_2176# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6691 a_16663_39# a_16462_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6692 a_7182_2446# a_7089_2446# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6693 a_14923_7598# a_14722_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6694 a_802_1636# a_709_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6695 a_9123_2198# a_8922_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6696 a_423_4088# a_222_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6697 GND a_7182_4606# a_7089_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6698 GND a_6602_3526# a_6509_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6699 a_9502_3526# a_9409_3526# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6700 VDD a_7182_8386# a_7089_8386# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6701 a_802_5416# a_709_5416# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6702 VDD a_6602_7306# a_6509_7306# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6703 a_5349_4876# WWL_13 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6704 GND a_1289_2446# a_1233_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6705 GND a_5929_3526# a_5873_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6706 a_7613_309# RWL_30 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6707 GND a_12309_2986# a_12253_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6708 GND a_15302_4066# a_15209_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6709 RBL0_15 RWL_18 a_9123_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6710 WBL_30 WWL_18 a_17622_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6711 WBL_31 WWL_14 a_18202_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6712 RBL0_0 RWL_11 a_423_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6713 a_1869_3256# WWL_19 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6714 a_6022_4336# a_5929_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6715 GND a_14629_4066# a_14573_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6716 a_6022_8116# a_5929_8116# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6717 a_16663_1118# a_16462_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6718 WBL_3 WWL_31 a_1962_16# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6719 a_12402_1366# a_12309_1366# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6720 a_9353_1658# RWL_25 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6721 a_10513_5978# RWL_9 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6722 GND a_11822_2446# a_11729_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6723 a_653_3548# RWL_18 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6724 a_7383_7328# a_7182_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6725 a_15789_5956# WWL_9 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6726 RBL0_9 RWL_30 a_5643_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6727 RBL0_9 RWL_24 a_5643_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6728 VDD a_11822_6226# a_11729_6226# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6729 a_2163_5168# a_1962_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6730 a_2542_2716# a_2449_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6731 a_2542_6496# a_2449_6496# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6732 a_8342_826# a_8249_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6733 a_18053_2198# RWL_23 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6734 a_15209_2716# WWL_21 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6735 a_3903_5708# a_3702_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6736 a_16462_5416# a_16369_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6737 VDD a_7762_1366# a_7669_1366# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6738 RBL0_23 RWL_26 a_13763_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6739 RBL0_24 RWL_22 a_14343_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6740 a_11242_3256# a_11149_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6741 VDD a_14722_17# a_14629_17# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6742 a_11242_7036# a_11149_7036# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6743 a_3029_6766# WWL_6 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6744 WBL_19 WWL_3 a_11242_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6745 RBL0_3 RWL_7 a_2163_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6746 RBL0_7 RWL_3 a_4483_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6747 a_17823_8408# a_17622_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6748 a_12603_6248# a_12402_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6749 VDD a_16462_1906# a_16369_1906# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6750 a_13413_848# RWL_28 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6751 a_3122_556# a_3029_556# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6752 a_7182_2176# a_7089_2176# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6753 a_9933_7868# RWL_2 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6754 GND a_12309_5956# a_12253_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6755 a_802_1366# a_709_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6756 GND a_7182_4336# a_7089_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6757 a_5293_6788# RWL_6 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6758 GND a_6602_3256# a_6509_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6759 WBL_16 WWL_17 a_9502_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6760 VDD a_7182_8116# a_7089_8116# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6761 WBL_1 WWL_10 a_802_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6762 VDD a_6602_7036# a_6509_7036# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6763 GND a_5929_3256# a_5873_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6764 RBL0_13 RWL_28 a_7963_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6765 GND a_1289_2176# a_1233_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6766 VDD a_222_6766# a_129_6766# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6767 RBL0_19 RWL_28 a_11443_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6768 VDD a_9502_556# a_9409_556# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6769 WBL_27 WWL_19 a_15882_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6770 WBL_16 WWL_28 a_9502_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6771 VDD a_12982_556# a_12889_556# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6772 RBL0_15 RWL_19 a_9123_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6773 RBL0_0 RWL_12 a_423_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6774 a_13469_556# WWL_29 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6775 a_1869_2986# WWL_20 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6776 a_6022_4066# a_5929_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6777 WBL_10 WWL_0 a_6022_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6778 GND a_2542_826# a_2449_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6779 a_12833_5708# RWL_10 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6781 a_12402_1096# a_12309_1096# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6782 WBL_21 WWL_25 a_12402_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6783 VDD a_10082_5956# a_9989_5956# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6784 a_9353_1388# RWL_26 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6785 GND a_11822_2176# a_11729_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6786 a_653_3278# RWL_19 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6787 a_7383_7058# a_7182_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6788 a_7762_4606# a_7669_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6789 RBL0_9 RWL_25 a_5643_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6790 a_2542_2446# a_2449_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6791 a_7762_8386# a_7669_8386# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6792 WBL_4 WWL_6 a_2542_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6793 a_2542_6226# a_2449_6226# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6794 a_6022_287# a_5929_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6795 a_8342_556# a_8249_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6796 a_17529_2446# WWL_22 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6797 VDD a_14142_3796# a_14049_3796# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6798 RBL0_20 RWL_27 a_12023_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6799 a_14142_7846# a_14049_7846# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6800 a_3903_5438# a_3702_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6801 a_16462_5146# a_16369_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6802 VDD a_7762_1096# a_7669_1096# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6803 RBL0_24 RWL_23 a_14343_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6804 a_14343_39# a_14142_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6805 RBL0_12 RWL_0 a_7383_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6806 a_3029_6496# WWL_7 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6807 WBL_19 WWL_4 a_11242_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6808 RBL0_3 RWL_8 a_2163_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6809 GND a_15882_287# a_15789_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6810 a_17823_8138# a_17622_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6811 a_11093_309# RWL_30 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6812 GND a_18202_7846# a_18109_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6813 a_13413_578# RWL_29 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6814 GND a_10662_8386# a_10569_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6815 a_7182_1906# a_7089_1906# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6816 WBL_12 WWL_22 a_7182_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6817 VDD a_9502_7846# a_9409_7846# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6818 GND a_17529_7846# a_17473_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6819 a_3122_286# a_3029_286# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6820 GND a_4189_2986# a_4133_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6821 GND a_7182_4066# a_7089_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6822 a_9933_7598# a_4683_7576# RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6823 a_14343_2738# a_14142_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6824 WBL_1 WWL_11 a_802_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6825 WBL_16 WWL_18 a_9502_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6826 GND a_222_2716# a_129_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6827 RBL0_13 RWL_29 a_7963_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6828 a_13469_7576# WWL_3 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6829 VDD a_222_6496# a_129_6496# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6830 RBL0_19 RWL_29 a_11443_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6831 WBL_12 WWL_30 a_7182_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6832 WBL_27 WWL_20 a_15882_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6833 RBL0_21 RWL_4 a_12603_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6834 VDD a_1382_5146# a_1289_5146# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6835 a_1813_4898# RWL_13 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6836 WBL_10 WWL_1 a_6022_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6837 a_13413_6518# RWL_7 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6838 GND a_2542_556# a_2449_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6839 GND a_14722_2986# a_14629_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6840 a_12833_5438# RWL_11 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6841 a_8829_1636# WWL_25 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6842 a_129_826# WWL_28 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6843 WBL_21 WWL_26 a_12402_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6844 a_7762_4336# a_7669_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6845 GND a_18202_826# a_18109_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6846 RBL0_9 RWL_26 a_5643_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6847 a_2542_2176# a_2449_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6848 a_7762_8116# a_7669_8116# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6849 WBL_4 WWL_7 a_2542_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6850 a_18109_3256# WWL_19 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6851 a_10283_7868# a_10082_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6852 a_17529_2176# WWL_23 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6853 RBL0_29 RWL_20 a_17243_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6854 VDD a_14142_3526# a_14049_3526# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6855 a_3903_5168# a_3702_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6856 a_8249_8386# WWL_0 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6857 RBL0_12 RWL_1 a_7383_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6858 a_3029_6226# WWL_8 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6859 GND a_4189_5956# a_4133_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6860 a_17473_1118# RWL_27 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6861 GND a_3609_4876# a_3553_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6862 a_5643_1928# a_5442_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6863 WBL_22 WWL_28 a_12982_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6864 GND a_9409_287# a_9353_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6865 GND a_18202_7576# a_18109_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6866 GND a_15209_6496# a_15153_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6867 a_10662_5956# a_10569_5956# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6868 GND a_12889_287# a_12833_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6869 a_8193_7328# RWL_4 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6870 GND a_10662_8116# a_10569_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6871 a_8922_7846# a_8829_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6872 a_4769_6766# WWL_6 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6873 a_1382_8386# a_1289_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6874 GND a_17529_7576# a_17473_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6875 a_3122_16# a_3029_16# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6876 WBL_12 WWL_23 a_7182_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6877 RBL0_6 RWL_7 a_3903_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6878 a_14343_2468# a_14142_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6880 a_14722_3796# a_14629_3796# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6881 a_10082_2716# a_9989_2716# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6882 GND a_14722_5956# a_14629_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6883 a_4713_5708# RWL_10 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6884 GND a_222_2446# a_129_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6885 GND a_10082_4876# a_9989_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6886 GND a_1382_1096# a_1289_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6887 a_13469_7306# WWL_4 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6888 VDD a_222_6226# a_129_6226# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6889 RBL0_21 RWL_5 a_12603_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6890 WBL_12 WWL_31 a_7182_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6891 VDD a_1382_4876# a_1289_4876# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6892 a_9409_2446# WWL_22 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6893 a_14142_6766# a_14049_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6894 a_13413_6248# RWL_8 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6895 RBL0_29 RWL_9 a_17243_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6896 a_12833_5168# RWL_12 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6897 a_8829_1366# WWL_26 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6898 VDD a_5442_2716# a_5349_2716# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6899 a_709_4336# WWL_15 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6900 WBL_21 WWL_27 a_12402_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6901 a_5442_2986# a_5349_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6902 RBL0_28 RWL_13 a_16663_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6903 a_7762_4066# a_7669_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6904 GND a_18202_556# a_18109_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6905 WBL_13 WWL_0 a_7762_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6906 WBL_4 WWL_8 a_2542_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6907 GND a_15209_826# a_15153_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6908 a_17529_1906# WWL_24 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6909 a_18109_2986# WWL_20 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6910 a_10283_7598# a_10082_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6911 WBL_24 WWL_2 a_14142_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6912 GND a_9502_6766# a_9409_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6913 GND a_6509_5686# a_6453_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6914 a_8249_8116# WWL_1 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6915 GND a_1962_7306# a_1869_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6916 GND a_8829_6766# a_8773_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6917 a_6223_2738# a_6022_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6918 a_5643_1658# a_5442_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6919 VDD a_15882_3796# a_15789_3796# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6920 VDD a_10662_1636# a_10569_1636# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6921 a_15882_7846# a_15789_7846# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6922 GND a_15209_6226# a_15153_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6923 a_8193_7058# RWL_5 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6924 a_8922_7576# a_8829_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6925 a_4769_6496# WWL_7 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6926 WBL_12 WWL_24 a_7182_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6927 a_1382_8116# a_1289_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6928 RBL0_6 RWL_8 a_3903_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6929 a_14343_2198# a_14142_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6930 GND a_12402_4606# a_12309_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6931 a_14722_3526# a_14629_3526# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6932 a_15302_4606# a_15209_4606# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6933 a_4282_286# a_4189_286# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6934 VDD a_12402_8386# a_12309_8386# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6935 a_11149_5956# WWL_9 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6936 RBL0_1 RWL_24 a_1003_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6937 a_4713_5438# RWL_11 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6938 GND a_222_2176# a_129_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6939 GND a_11729_4606# a_11673_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6940 a_5442_5956# a_5349_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6941 VDD a_3122_1366# a_3029_1366# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6942 a_1583_6788# a_1382_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6943 a_8829_1096# WWL_27 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6944 a_9409_2176# WWL_23 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6945 a_709_4066# WWL_16 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6946 WBL_9 WWL_5 a_5442_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6947 WBL_25 WWL_30 a_14722_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6948 a_15153_2738# RWL_21 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6949 a_13183_8408# a_12982_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6950 VDD a_17042_4066# a_16949_4066# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6951 WBL_13 WWL_1 a_7762_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6952 RBL0_18 RWL_24 a_10863_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6953 VDD a_4862_826# a_4769_826# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6954 GND a_15209_556# a_15153_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6955 a_5349_826# WWL_28 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6956 a_10662_4876# a_10569_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6957 WBL_8 WWL_17 a_4862_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6958 GND a_7089_6496# a_7033_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6959 GND a_6509_5416# a_6453_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6960 a_16083_848# a_15882_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6961 GND a_1962_7036# a_1869_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6962 VDD a_13562_2446# a_13469_2446# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6963 a_8342_287# a_8249_287# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6964 a_6223_2468# a_6022_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6965 a_12023_7868# a_11822_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6966 a_5643_1388# a_5442_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6967 VDD a_15882_3526# a_15789_3526# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6968 GND a_3702_3796# a_3609_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6969 a_6602_3796# a_6509_3796# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6970 VDD a_3702_7576# a_3609_7576# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6971 a_2449_5146# WWL_12 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6972 a_1382_1636# a_1289_1636# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6973 WBL_18 WWL_9 a_10662_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6974 a_17243_3008# a_17042_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6975 a_9989_8386# WWL_0 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6976 a_4769_6226# WWL_8 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6977 a_12982_3256# a_12889_3256# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6978 GND a_17622_6496# a_17529_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6979 a_11093_7868# RWL_2 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6980 GND a_12402_4336# a_12309_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6981 a_15302_4336# a_15209_4336# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6982 a_16369_7846# WWL_2 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6983 WBL_17 WWL_21 a_10082_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6984 RBL0_10 RWL_17 a_6223_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6985 WBL_25 WWL_17 a_14722_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6986 a_3122_4606# a_3029_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6987 VDD a_12402_8116# a_12309_8116# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6988 GND a_16949_6496# a_16893_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6989 RBL0_1 RWL_25 a_1003_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6990 a_3122_8386# a_3029_8386# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6991 GND a_11729_4336# a_11673_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6992 a_4713_5168# RWL_12 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6993 RBL0_14 RWL_13 a_8543_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6994 a_6453_1928# RWL_24 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6995 a_17042_7306# a_16949_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6996 VDD a_8342_3256# a_8249_3256# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6997 VDD a_3122_1096# a_3029_1096# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6998 a_9409_1906# WWL_24 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6999 a_14142_826# a_14049_826# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7000 a_15153_2468# RWL_22 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7001 WBL_25 WWL_31 a_14722_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7002 a_13183_8138# a_12982_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7003 a_13562_5686# a_13469_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7004 RBL0_19 RWL_21 a_11443_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7005 RBL0_18 RWL_25 a_10863_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7006 a_15882_6766# a_15789_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7007 WBL_8 WWL_18 a_4862_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7008 RBL0_2 RWL_2 a_1583_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7009 GND a_7089_6226# a_7033_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7010 a_17243_5978# a_17042_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7011 GND a_6509_5146# a_6453_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7012 a_16083_578# a_15882_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7013 VDD a_13562_2176# a_13469_2176# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7014 a_8342_17# a_8249_17# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7015 a_4282_2446# a_4189_2446# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7016 a_12023_7598# a_11822_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7017 GND a_8922_5686# a_8829_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7018 a_6223_2198# a_6022_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7019 GND a_3702_3526# a_3609_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7020 GND a_4282_4606# a_4189_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7021 a_6602_3526# a_6509_3526# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7022 a_73_4898# RWL_13 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7023 VDD a_4282_8386# a_4189_8386# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7024 a_7669_7036# WWL_5 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7025 VDD a_3702_7306# a_3609_7306# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7026 a_2449_4876# WWL_13 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7027 a_9989_8116# WWL_1 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7028 a_18202_5146# a_18109_5146# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7029 a_17622_4066# a_17529_4066# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7030 a_12982_2986# a_12889_2986# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7031 GND a_17622_6226# a_17529_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7032 a_11093_7598# a_4683_7576# RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7033 a_8342_6496# a_8249_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7034 a_7089_3796# WWL_17 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7035 GND a_12402_4066# a_12309_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7036 RBL0_10 RWL_18 a_6223_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7037 WBL_25 WWL_18 a_14722_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7038 a_3122_4336# a_3029_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7039 WBL_26 WWL_14 a_15302_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7040 GND a_16949_6226# a_16893_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7041 RBL0_1 RWL_26 a_1003_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7042 a_13763_1118# a_13562_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7043 GND a_11729_4066# a_11673_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7044 a_3122_8116# a_3029_8116# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7045 a_3122_16# a_3029_16# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7046 GND a_14049_1906# a_13993_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7047 a_6453_1658# RWL_25 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7048 a_4483_7328# a_4282_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7049 a_17042_7036# a_16949_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7050 a_12889_5956# WWL_9 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7051 a_6602_556# a_6509_556# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7052 RBL0_4 RWL_24 a_2743_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7053 VDD a_8342_2986# a_8249_2986# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7054 a_15153_2198# RWL_23 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7055 a_12309_2716# WWL_21 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7056 a_16949_3796# WWL_17 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7057 a_13562_5416# a_13469_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7058 VDD a_4862_1366# a_4769_1366# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7059 RBL0_18 RWL_26 a_10863_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7060 RBL0_19 RWL_22 a_11443_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7061 a_4483_38# a_4282_16# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7062 RBL0_2 RWL_3 a_1583_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7063 VDD a_18202_287# a_18109_287# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7064 a_16893_2738# RWL_21 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7065 a_9123_3008# a_8922_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7066 a_14923_8408# a_14722_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7067 VDD a_13562_1906# a_13469_1906# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7068 a_4282_2176# a_4189_2176# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7069 GND a_129_4606# a_73_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7070 GND a_8922_5416# a_8829_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7071 a_222_16# a_129_16# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7072 GND a_4282_4336# a_4189_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7073 a_2393_6788# RWL_6 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7074 GND a_3702_3256# a_3609_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7075 WBL_11 WWL_17 a_6602_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7076 VDD a_4282_8116# a_4189_8116# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7077 VDD a_3702_7036# a_3609_7036# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7078 a_9502_287# a_9409_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7079 a_18202_1096# a_18109_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7080 a_18202_4876# a_18109_4876# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7081 WBL_30 WWL_15 a_17622_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7082 WBL_22 WWL_19 a_12982_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7083 a_7089_3526# WWL_18 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7084 a_8342_6226# a_8249_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7085 a_1289_556# WWL_29 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7086 RBL0_10 RWL_19 a_6223_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7087 a_3122_4066# a_3029_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7088 WBL_5 WWL_0 a_3122_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7089 GND a_14049_1636# a_13993_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7090 a_6453_1388# RWL_26 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7091 a_4483_7058# a_4282_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7092 a_15302_17# a_15209_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7093 RBL0_4 RWL_25 a_2743_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7094 a_4862_4606# a_4769_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7095 a_4862_8386# a_4769_8386# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7096 a_18053_3008# RWL_20 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7097 a_14629_2446# WWL_22 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7098 VDD a_11242_3796# a_11149_3796# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7099 RBL0_15 RWL_30 a_9123_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7100 a_423_7868# a_222_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7101 a_9123_5978# a_8922_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7102 a_8543_4898# a_8342_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7103 a_11242_7846# a_11149_7846# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7104 a_16949_3526# WWL_18 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7105 a_13562_5146# a_13469_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7106 VDD a_4862_1096# a_4769_1096# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7107 RBL0_19 RWL_23 a_11443_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7108 RBL0_7 RWL_0 a_4483_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7109 a_15302_826# a_15209_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7110 a_8193_39# RWL_31 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7111 VDD a_18202_17# a_18109_17# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7112 a_16893_2468# RWL_22 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7113 a_14923_8138# a_14722_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7114 GND a_15302_7846# a_15209_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7115 a_9502_4066# a_9409_4066# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7116 a_802_5956# a_709_5956# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7117 a_4282_1906# a_4189_1906# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7118 WBL_7 WWL_22 a_4282_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7119 VDD a_6602_7846# a_6509_7846# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7120 GND a_14629_7846# a_14573_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7121 GND a_129_4336# a_73_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7122 GND a_8922_5146# a_8829_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7123 GND a_1289_2986# a_1233_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7124 GND a_4282_4066# a_4189_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7125 a_11443_2738# a_11242_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7126 WBL_11 WWL_18 a_6602_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7127 a_10082_556# a_9989_556# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7128 a_10569_7576# WWL_3 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7129 WBL_31 WWL_12 a_18202_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7130 WBL_30 WWL_16 a_17622_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7131 VDD a_6022_4606# a_5929_4606# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7132 WBL_22 WWL_20 a_12982_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7133 a_1289_286# WWL_30 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7134 WBL_5 WWL_1 a_3122_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7135 a_18053_5978# RWL_9 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7136 a_10513_6518# RWL_7 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7137 GND a_11822_2986# a_11729_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7138 VDD a_16462_556# a_16369_556# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7139 a_5929_1636# WWL_25 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7140 GND a_14049_1366# a_13993_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7141 GND a_6022_826# a_5929_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7142 a_4862_4336# a_4769_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7143 RBL0_4 RWL_26 a_2743_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7144 a_4862_8116# a_4769_8116# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7145 a_2163_38# a_1962_16# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7146 GND a_16462_1906# a_16369_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7147 VDD a_16462_5686# a_16369_5686# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7148 a_15209_3256# WWL_19 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7149 GND a_15789_1906# a_15733_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7150 a_14629_2176# WWL_23 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7151 VDD a_11242_3526# a_11149_3526# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7152 RBL0_24 RWL_20 a_14343_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7153 a_423_7598# a_222_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7154 a_1962_3796# a_1869_3796# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7155 a_5349_8386# WWL_0 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7156 a_12982_287# a_12889_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7157 RBL0_7 RWL_1 a_4483_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7158 GND a_1289_5956# a_1233_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7159 a_14573_1118# RWL_27 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7160 a_15302_556# a_15209_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7161 a_2743_1928# a_2542_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7162 a_16893_2198# RWL_23 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7163 a_9933_8408# RWL_0 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7164 GND a_15302_7576# a_15209_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7165 GND a_12309_6496# a_12253_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7166 a_5293_7328# RWL_4 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7167 WBL_16 WWL_15 a_9502_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7168 a_6022_7846# a_5929_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7169 a_1869_6766# WWL_6 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7170 GND a_14629_7576# a_14573_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7171 WBL_7 WWL_23 a_4282_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7172 GND a_129_4066# a_73_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7173 a_16663_4628# a_16462_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7174 a_11443_2468# a_11242_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7175 a_11822_3796# a_11729_3796# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7176 GND a_11822_5956# a_11729_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7177 a_1813_5708# RWL_10 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7178 GND a_5929_17# a_5873_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7179 VDD a_6022_4336# a_5929_4336# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7180 WBL_31 WWL_13 a_18202_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7181 a_10569_7306# WWL_4 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7182 a_12982_17# a_12889_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7183 a_1289_16# WWL_31 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7184 a_6509_2446# WWL_22 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7185 a_11242_6766# a_11149_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7186 a_10513_6248# RWL_8 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7187 RBL0_24 RWL_9 a_14343_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7188 a_5929_1366# WWL_26 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7189 VDD a_2542_2716# a_2449_2716# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7190 RBL0_23 RWL_13 a_13763_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7191 a_2542_2986# a_2449_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7192 GND a_6022_556# a_5929_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7193 a_4862_4066# a_4769_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7194 GND a_16462_1636# a_16369_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7195 GND a_3029_826# a_2973_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7196 a_7182_1906# a_7089_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7197 VDD a_16462_5416# a_16369_5416# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7198 GND a_15789_1636# a_15733_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7199 a_14629_1906# WWL_24 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7200 a_15209_2986# WWL_20 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7201 a_7182_5686# a_7089_5686# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7202 a_1962_3526# a_1869_3526# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7203 GND a_7182_7846# a_7089_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7204 a_3029_7036# WWL_5 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7205 a_802_4876# a_709_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7206 WBL_19 WWL_2 a_11242_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7207 GND a_6602_6766# a_6509_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7208 GND a_3609_5686# a_3553_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7209 a_5349_8116# WWL_1 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7210 GND a_5929_6766# a_5873_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7211 a_7963_3818# a_7762_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7212 a_3323_2738# a_3122_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7213 GND a_18202_8386# a_18109_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7214 a_2743_1658# a_2542_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7215 VDD a_12982_3796# a_12889_3796# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7216 WBL_27 WWL_6 a_15882_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7217 GND a_17529_8386# a_17473_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7218 GND a_12309_6226# a_12253_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7219 RBL0_28 RWL_30 a_16663_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7220 a_9933_8138# RWL_1 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7221 a_5293_7058# RWL_5 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7222 a_6022_7576# a_5929_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7223 RBL0_15 RWL_6 a_9123_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7224 a_1869_6496# WWL_7 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7225 WBL_1 WWL_9 a_802_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7226 WBL_16 WWL_16 a_9502_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7227 WBL_7 WWL_24 a_4282_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7228 a_16663_4358# a_16462_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7229 a_11443_2198# a_11242_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7230 GND a_10082_5686# a_9989_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7231 GND a_16369_287# a_16313_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7232 a_7033_3818# RWL_17 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7233 a_11822_3526# a_11729_3526# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7234 a_12402_4606# a_12309_4606# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7235 a_653_6788# RWL_6 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7236 a_9353_4898# RWL_13 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7237 a_1813_5438# RWL_11 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7238 a_2542_5956# a_2449_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7239 RBL0_28 RWL_10 a_16663_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7240 RBL0_20 RWL_14 a_12023_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7241 a_6509_2176# WWL_23 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7242 VDD a_7762_4606# a_7669_4606# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7243 a_5929_1096# WWL_27 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7244 GND a_802_286# a_709_286# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7245 WBL_4 WWL_5 a_2542_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7246 a_12253_2738# RWL_21 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7247 a_10283_8408# a_10082_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7248 VDD a_14142_4066# a_14049_4066# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7249 GND a_3029_556# a_2973_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7250 GND a_16462_1366# a_16369_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7251 a_7182_1636# a_7089_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7252 a_7182_5416# a_7089_5416# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7253 GND a_15789_1366# a_15733_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7254 WBL_3 WWL_17 a_1962_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7255 GND a_7182_7576# a_7089_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7256 GND a_4189_6496# a_4133_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7257 GND a_3609_5416# a_3553_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7258 VDD a_10662_2446# a_10569_2446# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7259 GND a_16462_17# a_16369_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7260 a_3323_2468# a_3122_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7261 a_7963_3548# a_7762_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7262 GND a_18202_8116# a_18109_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7263 a_2743_1388# a_2542_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7264 VDD a_12982_3526# a_12889_3526# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7265 a_8922_8386# a_8829_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7266 WBL_27 WWL_7 a_15882_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7267 a_3702_3796# a_3609_3796# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7268 GND a_17529_8116# a_17473_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7269 a_14343_3008# a_14142_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7270 a_1869_6226# WWL_8 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7271 a_10082_3256# a_9989_3256# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7272 a_16663_4088# a_16462_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7273 GND a_14722_6496# a_14629_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7274 GND a_10082_5416# a_9989_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7275 GND a_222_2986# a_129_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7276 a_7033_3548# RWL_18 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7277 a_12402_4336# a_12309_4336# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7278 a_13469_7846# WWL_2 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7279 GND a_8249_1096# a_8193_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7280 a_6509_287# WWL_30 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7281 RBL0_5 RWL_17 a_3323_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7282 a_7762_7846# a_7669_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7283 a_1813_5168# RWL_12 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7284 RBL0_9 RWL_13 a_5643_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7285 a_18109_6766# WWL_6 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7286 a_17529_5686# WWL_10 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7287 a_3553_1928# RWL_24 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7288 a_14142_7306# a_14049_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7289 RBL0_29 RWL_7 a_17243_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7290 VDD a_5442_3256# a_5349_3256# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7291 RBL0_28 RWL_11 a_16663_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7292 a_7963_848# a_7762_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7293 RBL0_20 RWL_15 a_12023_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7294 a_6509_1906# WWL_24 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7295 VDD a_7762_4336# a_7669_4336# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7296 a_17473_4628# RWL_14 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7297 a_1962_826# a_1869_826# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7298 a_12253_2468# RWL_22 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7299 a_10283_8138# a_10082_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7300 a_10662_5686# a_10569_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7301 a_7182_1366# a_7089_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7302 GND a_9502_7306# a_9409_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7303 WBL_12 WWL_10 a_7182_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7304 GND a_8829_7306# a_8773_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7305 WBL_3 WWL_18 a_1962_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7306 GND a_4189_6226# a_4133_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7307 a_14343_5978# a_14142_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7308 GND a_3609_5146# a_3553_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7309 VDD a_18202_1636# a_18109_1636# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7310 VDD a_8342_826# a_8249_826# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7311 VDD a_10662_2176# a_10569_2176# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7312 a_222_3796# a_129_3796# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7313 a_12309_826# WWL_28 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7314 a_1382_2446# a_1289_2446# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7315 a_7963_3278# a_7762_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7316 GND a_222_5956# a_129_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7317 a_3323_2198# a_3122_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7318 GND a_1382_4606# a_1289_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7319 a_8922_8116# a_8829_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7320 a_4769_7036# WWL_5 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7321 WBL_27 WWL_8 a_15882_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7322 a_3702_3526# a_3609_3526# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7323 VDD a_1382_8386# a_1289_8386# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7324 a_15302_5146# a_15209_5146# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7325 a_15302_287# a_15209_287# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7326 a_14722_4066# a_14629_4066# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7327 a_10082_2986# a_9989_2986# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7328 GND a_14722_6226# a_14629_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7329 GND a_10082_5146# a_9989_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7330 a_7033_3278# RWL_19 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7331 a_5442_6496# a_5349_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7332 RBL0_14 RWL_10 a_8543_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7333 a_4189_3796# WWL_17 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7334 WBL_21 WWL_14 a_12402_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7335 a_6509_17# WWL_31 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7336 RBL0_5 RWL_18 a_3323_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7337 a_7762_7576# a_7669_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7338 a_10863_1118# a_10662_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7339 GND a_11149_1906# a_11093_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7340 a_8773_3818# RWL_17 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7341 a_18109_6496# WWL_7 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7342 a_17529_5416# WWL_11 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7343 a_5643_309# a_5442_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7344 a_3553_1658# RWL_25 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7345 a_1583_7328# a_1382_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7346 RBL0_29 RWL_8 a_17243_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7347 a_14142_7036# a_14049_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7348 RBL0_28 RWL_12 a_16663_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7349 a_7963_578# a_7762_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7350 VDD a_5442_2986# a_5349_2986# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7351 RBL0_20 RWL_16 a_12023_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7352 a_17473_4358# RWL_15 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7353 a_12253_2198# RWL_23 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7354 VDD a_802_2716# a_709_2716# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7355 a_10662_5416# a_10569_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7356 VDD a_1962_1366# a_1869_1366# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7357 GND a_14142_17# a_14049_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7358 WBL_8 WWL_15 a_4862_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7359 GND a_9502_7036# a_9409_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7360 WBL_12 WWL_11 a_7182_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7361 a_1233_308# RWL_30 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7362 GND a_8829_7036# a_8773_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7363 VDD a_6022_287# a_5929_287# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7364 a_13993_2738# RWL_21 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7365 a_6223_3008# a_6022_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7366 a_12023_8408# a_11822_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7367 VDD a_15882_4066# a_15789_4066# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7368 a_8922_1636# a_8829_1636# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7369 VDD a_10662_1906# a_10569_1906# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7370 a_73_5708# RWL_10 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7371 a_222_3526# a_129_3526# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7372 a_1382_2176# a_1289_2176# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7373 GND a_1382_4336# a_1289_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7374 WBL_6 WWL_17 a_3702_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7375 VDD a_1382_8116# a_1289_8116# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7376 a_15302_1096# a_15209_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7377 a_11443_848# a_11242_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7378 a_11093_8408# RWL_0 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7379 a_15302_17# a_15209_17# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7380 a_15302_4876# a_15209_4876# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7381 WBL_17 WWL_19 a_10082_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7382 WBL_25 WWL_15 a_14722_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7383 a_709_7576# WWL_3 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7384 a_9409_5686# WWL_10 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7385 a_8829_4606# WWL_14 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7386 a_5442_6226# a_5349_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7387 RBL0_14 RWL_11 a_8543_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7388 a_4189_3526# WWL_18 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7389 RBL0_5 RWL_19 a_3323_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7390 a_12833_39# RWL_31 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7391 WBL_28 WWL_29 a_16462_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7392 GND a_17042_3796# a_16949_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7393 VDD a_17042_7576# a_16949_7576# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7394 GND a_16369_3796# a_16313_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7395 GND a_11149_1636# a_11093_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7396 a_8773_3548# RWL_18 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7397 a_18109_6226# WWL_8 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7398 a_3553_1388# RWL_26 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7399 a_1583_7058# a_1382_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7400 GND a_9989_1096# a_9933_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7401 a_15153_3008# RWL_20 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7402 a_11729_2446# WWL_22 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7403 a_6223_5978# a_6022_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7404 a_17473_4088# RWL_16 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7405 a_5643_4898# a_5442_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7406 a_15882_7306# a_15789_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7407 a_10662_5146# a_10569_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7408 VDD a_1962_1096# a_1869_1096# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7409 WBL_8 WWL_16 a_4862_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7410 RBL0_2 RWL_0 a_1583_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7411 a_17243_6518# a_17042_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7412 a_12982_6766# a_12889_6766# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7413 VDD a_6022_17# a_5929_17# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7414 a_13993_2468# RWL_22 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7415 a_12023_8138# a_11822_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7416 GND a_12402_7846# a_12309_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7417 a_73_5438# RWL_11 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7418 WBL_0 WWL_17 a_222_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7419 a_6602_4066# a_6509_4066# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7420 a_1382_1906# a_1289_1906# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7421 WBL_2 WWL_22 a_1382_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7422 VDD a_3702_7846# a_3609_7846# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7423 GND a_11729_7846# a_11673_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7424 GND a_1382_4066# a_1289_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7425 WBL_6 WWL_18 a_3702_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7426 a_11093_8138# RWL_1 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7427 VDD a_8342_6766# a_8249_6766# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7428 WBL_26 WWL_12 a_15302_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7429 a_11443_578# a_11242_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7430 a_7089_4336# WWL_15 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7431 WBL_25 WWL_16 a_14722_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7432 VDD a_3122_4606# a_3029_4606# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7433 WBL_17 WWL_20 a_10082_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7434 a_709_7306# WWL_4 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7435 a_9409_5416# WWL_11 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7436 RBL0_14 RWL_12 a_8543_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7437 a_17042_1366# a_16949_1366# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7438 GND a_17042_3526# a_16949_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7439 a_15153_5978# RWL_9 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7440 VDD a_17042_7306# a_16949_7306# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7441 VDD a_4282_556# a_4189_556# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7442 GND a_16369_3526# a_16313_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7443 GND a_11149_1366# a_11093_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7444 a_8773_3278# RWL_19 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7445 GND a_13562_1906# a_13469_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7446 a_8543_5708# a_8342_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7447 VDD a_13562_5686# a_13469_5686# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7448 a_12309_3256# WWL_19 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7449 a_16949_4336# WWL_15 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7450 GND a_12889_1906# a_12833_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7451 a_11729_2176# WWL_23 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7452 RBL0_19 RWL_20 a_11443_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7453 a_15882_7036# a_15789_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7454 a_8773_848# RWL_28 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7455 a_2449_8386# WWL_0 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7456 RBL0_2 RWL_1 a_1583_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7457 a_17243_6248# a_17042_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7458 a_17622_3796# a_17529_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7459 a_11673_1118# RWL_27 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7460 a_12982_2716# a_12889_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7461 a_17622_7576# a_17529_7576# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7462 a_12982_6496# a_12889_6496# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7463 a_13993_2198# RWL_23 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7464 GND a_12402_7576# a_12309_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7465 a_2393_7328# RWL_4 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7466 RBL0_11 RWL_28 a_6803_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7467 WBL_0 WWL_18 a_222_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7468 WBL_11 WWL_15 a_6602_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7469 a_3122_7846# a_3029_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7470 a_73_5168# RWL_12 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7471 WBL_2 WWL_23 a_1382_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7472 RBL0_1 RWL_13 a_1003_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7473 GND a_11729_7576# a_11673_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7474 a_3903_308# a_3702_286# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7475 GND a_7182_287# a_7089_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7476 a_13763_4628# a_13562_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7477 a_8829_556# WWL_29 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7478 GND a_8342_2716# a_8249_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7479 VDD a_8342_6496# a_8249_6496# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7480 a_7089_4066# WWL_16 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7481 GND a_7669_2716# a_7613_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7482 VDD a_3122_4336# a_3029_4336# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7483 WBL_26 WWL_13 a_15302_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7484 a_17042_1096# a_16949_1096# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7485 WBL_29 WWL_25 a_17042_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7486 GND a_17042_3256# a_16949_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7487 VDD a_17042_7036# a_16949_7036# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7488 a_4862_287# a_4769_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7489 a_3609_2446# WWL_22 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7490 RBL0_19 RWL_9 a_11443_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7491 VDD a_4282_286# a_4189_286# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7492 GND a_16369_3256# a_16313_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7493 RBL0_18 RWL_13 a_10863_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7494 GND a_13562_1636# a_13469_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7495 a_423_8408# a_222_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7496 a_9123_6518# a_8922_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7497 a_8543_5438# a_8342_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7498 VDD a_13562_5416# a_13469_5416# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7499 a_4282_1906# a_4189_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7500 a_12309_2986# WWL_20 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7501 a_16949_4066# WWL_16 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7502 GND a_12889_1636# a_12833_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7503 a_11729_1906# WWL_24 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7504 a_4282_5686# a_4189_5686# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7505 a_6453_309# RWL_30 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7506 GND a_4282_7846# a_4189_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7507 a_8773_578# RWL_29 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7508 GND a_3702_6766# a_3609_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7509 a_2449_8116# WWL_1 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7510 a_16893_3008# RWL_20 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7511 a_18202_4606# a_18109_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7512 a_12982_2446# a_12889_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7513 a_17622_3526# a_17529_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7514 a_18202_8386# a_18109_8386# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7515 GND a_15302_8386# a_15209_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7516 a_17622_7306# a_17529_7306# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7517 a_12982_6226# a_12889_6226# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7518 WBL_22 WWL_6 a_12982_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7519 GND a_14629_8386# a_14573_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7520 a_17622_556# a_17529_556# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7521 a_2393_7058# RWL_5 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7522 RBL0_10 RWL_6 a_6223_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7523 RBL0_11 RWL_29 a_6803_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7524 a_3122_7576# a_3029_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7525 WBL_11 WWL_16 a_6602_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7526 WBL_2 WWL_24 a_1382_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7527 a_13763_4358# a_13562_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7528 a_4133_3818# RWL_17 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7529 a_10662_826# a_10569_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7530 VDD a_6022_5146# a_5929_5146# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7531 GND a_8342_2446# a_8249_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7532 a_6453_4898# RWL_13 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7533 VDD a_8342_6226# a_8249_6226# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7534 GND a_7669_2446# a_7613_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7535 a_18053_6518# RWL_7 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7536 WBL_29 WWL_26 a_17042_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7537 a_129_2446# WWL_22 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7538 RBL0_23 RWL_10 a_13763_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7539 a_12253_848# RWL_28 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7540 a_3609_2176# WWL_23 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7541 VDD a_4862_4606# a_4769_4606# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7542 VDD a_4282_16# a_4189_16# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7543 VDD a_11242_4066# a_11149_4066# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7544 a_16893_5978# RWL_9 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7545 GND a_13562_1366# a_13469_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7546 a_423_8138# a_222_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7547 a_9123_6248# a_8922_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7548 a_802_5686# a_709_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7549 a_8543_5168# a_8342_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7550 a_9502_3796# a_9409_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7551 RBL0_17 RWL_28 a_10283_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7552 a_4282_1636# a_4189_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7553 a_9502_7576# a_9409_7576# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7554 a_4282_5416# a_4189_5416# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7555 GND a_12889_1366# a_12833_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7556 GND a_129_7846# a_73_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7557 WBL_14 WWL_28 a_8342_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7558 VDD a_11822_556# a_11729_556# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7559 GND a_4282_7576# a_4189_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7560 GND a_1289_6496# a_1233_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7561 a_18202_4336# a_18109_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7563 a_12982_2176# a_12889_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7564 a_17622_3256# a_17529_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7565 GND a_15302_8116# a_15209_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7566 a_18202_8116# a_18109_8116# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7567 WBL_30 WWL_3 a_17622_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7568 a_17622_7036# a_17529_7036# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7569 a_6022_8386# a_5929_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7570 WBL_22 WWL_7 a_12982_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7571 GND a_14629_8116# a_14573_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7572 a_11443_3008# a_11242_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7573 a_13763_4088# a_13562_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7574 GND a_11822_6496# a_11729_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7575 a_9353_5708# RWL_10 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7576 GND a_6022_1096# a_5929_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7577 a_10662_556# a_10569_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7578 a_4133_3548# RWL_18 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7579 GND a_14049_4876# a_13993_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7580 VDD a_6022_4876# a_5929_4876# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7581 a_10569_7846# WWL_2 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7582 GND a_5349_1096# a_5293_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7583 a_16083_1928# a_15882_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7584 GND a_8342_2176# a_8249_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7585 a_4862_7846# a_4769_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7586 GND a_7669_2176# a_7613_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7587 RBL0_4 RWL_13 a_2743_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7588 a_1003_1118# a_802_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7589 a_18053_6248# RWL_8 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7590 GND a_14722_287# a_14629_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7591 a_15209_6766# WWL_6 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7592 a_14629_5686# WWL_10 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7593 a_129_2176# WWL_23 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7594 a_11242_7306# a_11149_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7595 RBL0_24 RWL_7 a_14343_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7596 RBL0_23 RWL_11 a_13763_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7597 WBL_29 WWL_27 a_17042_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7598 VDD a_2542_3256# a_2449_3256# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7599 a_12253_578# RWL_29 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7600 a_3609_1906# WWL_24 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7601 VDD a_4862_4336# a_4769_4336# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7602 a_8922_17# a_8829_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7603 a_14573_4628# RWL_14 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7604 VDD a_16462_5956# a_16369_5956# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7605 a_9502_3526# a_9409_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7606 a_1962_4066# a_1869_4066# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7607 GND a_7182_8386# a_7089_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7608 a_802_5416# a_709_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7609 a_4282_1366# a_4189_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7610 a_9502_7306# a_9409_7306# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7611 GND a_6602_7306# a_6509_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7612 RBL0_17 RWL_29 a_10283_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7613 WBL_10 WWL_30 a_6022_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7614 GND a_4282_16# a_4189_16# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7615 WBL_7 WWL_10 a_4282_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7616 GND a_129_7576# a_73_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7617 GND a_5929_7306# a_5873_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7618 GND a_16369_17# a_16313_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7619 GND a_1289_6226# a_1233_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7620 a_11443_5978# a_11242_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7621 RBL0_31 RWL_27 a_18403_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7622 VDD a_15302_1636# a_15209_1636# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7623 a_18202_4066# a_18109_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7624 WBL_31 WWL_0 a_18202_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7625 RBL0_15 RWL_4 a_9123_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7626 a_6022_8116# a_5929_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7627 WBL_30 WWL_4 a_17622_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7628 a_1869_7036# WWL_5 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7629 WBL_22 WWL_8 a_12982_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7630 RBL0_28 RWL_31 a_16663_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7631 a_12402_5146# a_12309_5146# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7632 a_11822_4066# a_11729_4066# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7633 a_653_7328# RWL_4 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7634 GND a_11822_6226# a_11729_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7635 a_9353_5438# RWL_11 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7636 a_4133_3278# RWL_19 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7637 a_1289_3796# WWL_17 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7638 a_2542_6496# a_2449_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7639 RBL0_9 RWL_10 a_5643_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7640 a_16083_1658# a_15882_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7641 a_4862_7576# a_4769_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7642 a_2973_38# RWL_31 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7643 a_5873_3818# RWL_17 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7644 a_15209_6496# WWL_7 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7645 a_14629_5416# WWL_11 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7646 VDD a_7762_5146# a_7669_5146# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7647 a_11242_7036# a_11149_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7648 RBL0_24 RWL_8 a_14343_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7649 WBL_20 WWL_28 a_11822_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7650 a_129_1906# WWL_24 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7651 VDD a_2542_2986# a_2449_2986# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7652 RBL0_23 RWL_12 a_13763_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7653 GND a_11729_287# a_11673_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7654 RBL0_4 RWL_30 a_2743_308# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7655 a_14573_4358# RWL_15 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7656 a_14923_848# a_14722_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7657 a_7182_5956# a_7089_5956# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7658 a_9502_3256# a_9409_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7659 a_802_5146# a_709_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7660 WBL_3 WWL_15 a_1962_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7661 GND a_7182_8116# a_7089_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7662 GND a_6602_7036# a_6509_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7663 VDD a_18202_2446# a_18109_2446# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7664 WBL_16 WWL_3 a_9502_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7665 a_9502_7036# a_9409_7036# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7666 WBL_10 WWL_31 a_6022_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7667 WBL_7 WWL_11 a_4282_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7668 a_16663_7868# a_16462_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7669 GND a_5929_7036# a_5873_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7670 a_3323_3008# a_3122_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7671 VDD a_12982_4066# a_12889_4066# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7672 a_6022_1636# a_5929_1636# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7673 WBL_27 WWL_5 a_15882_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7674 GND a_3029_2716# a_2973_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7675 WBL_31 WWL_1 a_18202_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7676 RBL0_15 RWL_5 a_9123_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7677 a_12402_1096# a_12309_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7678 a_12402_4876# a_12309_4876# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7679 a_9353_5168# RWL_12 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7680 a_7762_8386# a_7669_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7681 a_653_7058# RWL_5 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7682 a_6509_5686# WWL_10 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7683 a_5929_4606# WWL_14 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7684 a_2542_6226# a_2449_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7685 RBL0_9 RWL_11 a_5643_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7686 a_1289_3526# WWL_18 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7687 a_16083_1388# a_15882_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7688 WBL_7 WWL_29 a_4282_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7689 GND a_14142_3796# a_14049_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7690 a_16462_2716# a_16369_2716# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7691 VDD a_14142_7576# a_14049_7576# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7692 GND a_7762_1096# a_7669_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7693 GND a_13469_3796# a_13413_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7694 GND a_16462_4876# a_16369_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7695 a_5873_3548# RWL_18 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7696 a_15209_6226# WWL_8 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7697 a_17823_1928# a_17622_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7698 GND a_15789_4876# a_15733_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7699 VDD a_7762_4876# a_7669_4876# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7700 a_12253_3008# RWL_20 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7701 RBL0_27 RWL_21 a_16083_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7702 a_3323_5978# a_3122_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7703 GND a_14049_17# a_13993_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7704 a_12603_309# a_12402_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7705 a_14923_578# a_14722_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7706 VDD a_7182_1636# a_7089_1636# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7707 a_14573_4088# RWL_16 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7708 a_2743_4898# a_2542_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7709 a_3122_286# a_3029_286# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7710 a_222_556# a_129_556# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7711 WBL_3 WWL_16 a_1962_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7712 a_14343_6518# a_14142_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7713 VDD a_18202_2176# a_18109_2176# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7714 WBL_16 WWL_4 a_9502_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7715 a_8922_2446# a_8829_2446# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7716 a_16663_7598# a_16462_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7717 a_10082_6766# a_9989_6766# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7718 GND a_222_6496# a_129_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7719 a_3702_4066# a_3609_4066# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7720 GND a_8249_4606# a_8193_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7721 GND a_3029_2446# a_2973_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7722 RBL0_20 RWL_2 a_12023_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7723 VDD a_5442_6766# a_5349_6766# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7724 WBL_21 WWL_12 a_12402_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7725 VDD a_3702_826# a_3609_826# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7726 a_4189_4336# WWL_15 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7727 a_7762_8116# a_7669_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7728 a_6509_5416# WWL_11 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7729 RBL0_9 RWL_12 a_5643_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7730 a_14142_1366# a_14049_1366# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7731 WBL_7 WWL_30 a_4282_286# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7732 GND a_14142_3526# a_14049_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7733 a_18109_7036# WWL_5 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7734 a_17529_5956# WWL_9 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7735 a_12253_5978# RWL_9 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7736 RBL0_12 RWL_24 a_7383_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7737 VDD a_14142_7306# a_14049_7306# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7738 GND a_13469_3526# a_13413_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7739 a_10662_287# a_10569_287# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7740 a_5873_3278# RWL_19 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7741 a_7182_4876# a_7089_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7742 a_17823_1658# a_17622_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7743 GND a_10662_1906# a_10569_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7744 a_5643_5708# a_5442_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7745 VDD a_9502_1366# a_9409_1366# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7746 VDD a_10662_5686# a_10569_5686# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7747 RBL0_27 RWL_22 a_16083_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7748 VDD a_802_3256# a_709_3256# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7749 a_7963_6788# a_7762_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7750 a_222_286# a_129_286# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7751 a_17529_287# WWL_30 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7752 WBL_12 WWL_9 a_7182_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7753 a_14343_6248# a_14142_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7754 a_14722_3796# a_14629_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7755 VDD a_18202_1906# a_18109_1906# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7756 a_10082_2716# a_9989_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7757 a_8922_2176# a_8829_2176# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7758 a_14722_7576# a_14629_7576# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7759 a_10082_6496# a_9989_6496# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7760 a_222_4066# a_129_4066# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7761 a_7033_6788# RWL_6 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7762 GND a_222_6226# a_129_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7763 WBL_6 WWL_15 a_3702_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7764 GND a_8249_4336# a_8193_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7765 GND a_3029_2176# a_2973_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7766 a_10863_4628# a_10662_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7767 GND a_5442_2716# a_5349_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7768 a_8829_5146# WWL_12 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7769 a_7762_1636# a_7669_1636# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7770 RBL0_20 a_4683_7576# a_12023_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7771 VDD a_5442_6496# a_5349_6496# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7772 a_4189_4066# WWL_16 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7773 GND a_4769_2716# a_4713_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7774 WBL_21 WWL_13 a_12402_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7775 a_14142_1096# a_14049_1096# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7776 WBL_24 WWL_25 a_14142_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7777 a_17473_7868# RWL_2 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7778 WBL_7 WWL_31 a_4282_16# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7779 GND a_14142_3256# a_14049_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7780 WBL_28 WWL_21 a_16462_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7781 VDD a_14142_7036# a_14049_7036# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7782 RBL0_12 RWL_25 a_7383_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7783 GND a_13469_3256# a_13413_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7784 a_10662_17# a_10569_17# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7785 a_17823_1388# a_17622_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7786 GND a_15882_3796# a_15789_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7787 GND a_10662_1636# a_10569_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7788 VDD a_15882_7576# a_15789_7576# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7789 a_6223_6518# a_6022_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7790 a_5643_5438# a_5442_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7791 VDD a_9502_1096# a_9409_1096# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7792 VDD a_10662_5416# a_10569_5416# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7793 a_1382_1906# a_1289_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7794 RBL0_27 RWL_23 a_16083_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7795 VDD a_802_2986# a_709_2986# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7796 a_1382_5686# a_1289_5686# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7797 GND a_1382_7846# a_1289_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7798 a_17529_17# WWL_31 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7799 a_222_16# a_129_16# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7800 RBL0_30 RWL_21 a_17823_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7801 a_13993_3008# RWL_20 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7802 a_15302_4606# a_15209_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7803 a_10082_2446# a_9989_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7804 a_14722_3526# a_14629_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7805 a_15302_8386# a_15209_8386# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7806 GND a_12402_8386# a_12309_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7807 a_8922_1906# a_8829_1906# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7808 a_14722_7306# a_14629_7306# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7809 a_10082_6226# a_9989_6226# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7810 WBL_15 WWL_22 a_8922_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7811 WBL_0 WWL_15 a_222_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7812 WBL_17 WWL_6 a_10082_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7813 RBL0_1 RWL_10 a_1003_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7814 GND a_11729_8386# a_11673_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7815 a_5442_556# a_5349_556# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7816 RBL0_5 RWL_6 a_3323_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7817 WBL_6 WWL_16 a_3702_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7818 GND a_8249_4066# a_8193_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7819 a_10863_4358# a_10662_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7820 a_1233_3818# RWL_17 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7821 VDD a_3122_5146# a_3029_5146# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7822 GND a_5442_2446# a_5349_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7823 a_709_7846# WWL_2 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7824 a_9409_5956# WWL_9 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7825 a_3553_4898# RWL_13 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7826 a_8829_4876# WWL_13 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7827 VDD a_5442_6226# a_5349_6226# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7828 GND a_9989_4606# a_9933_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7829 GND a_4769_2446# a_4713_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7830 a_15789_556# WWL_29 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7831 a_15153_6518# RWL_7 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7832 VDD a_17042_7846# a_16949_7846# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7833 GND a_4862_826# a_4769_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7834 WBL_24 WWL_26 a_14142_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7835 RBL0_18 RWL_10 a_10863_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7836 a_17473_7598# a_13963_7576# RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7837 RBL0_12 RWL_26 a_7383_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7838 VDD a_1962_4606# a_1869_4606# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7839 WBL_8 WWL_3 a_4862_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7840 a_15882_1366# a_15789_1366# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7841 a_8342_287# a_8249_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7842 GND a_15882_3526# a_15789_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7843 a_13993_5978# RWL_9 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7844 GND a_10662_1366# a_10569_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7845 VDD a_15882_7306# a_15789_7306# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7846 a_6223_6248# a_6022_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7847 a_5643_5168# a_5442_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7848 a_6602_3796# a_6509_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7849 a_1382_1636# a_1289_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7850 a_6602_7576# a_6509_7576# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7851 a_1382_5416# a_1289_5416# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7852 GND a_1382_7576# a_1289_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7853 a_16369_1636# WWL_25 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7854 RBL0_30 RWL_22 a_17823_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7855 a_15302_4336# a_15209_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7856 a_10082_2176# a_9989_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7857 a_14722_3256# a_14629_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7858 a_15302_8116# a_15209_8116# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7859 GND a_12402_8116# a_12309_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7860 a_13413_309# RWL_30 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7861 WBL_25 WWL_3 a_14722_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7862 a_14722_7036# a_14629_7036# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7863 WBL_15 WWL_23 a_8922_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7864 WBL_0 WWL_16 a_222_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7865 a_3122_8386# a_3029_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7866 WBL_17 WWL_7 a_10082_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7867 RBL0_1 RWL_11 a_1003_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7868 GND a_11729_8116# a_11673_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7869 a_6453_5708# RWL_10 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7870 a_10513_39# RWL_31 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7871 a_10863_4088# a_10662_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7872 GND a_3122_1096# a_3029_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7873 RBL0_13 RWL_30 a_7963_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7874 a_1233_3548# RWL_18 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7875 RBL0_19 RWL_30 a_11443_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7876 GND a_11149_4876# a_11093_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7877 VDD a_3122_4876# a_3029_4876# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7878 a_8773_6788# RWL_6 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7879 GND a_2449_1096# a_2393_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7880 a_13183_1928# a_12982_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7881 GND a_5442_2176# a_5349_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7882 WBL_16 WWL_30 a_9502_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7883 GND a_9989_4336# a_9933_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7884 a_14142_826# a_14049_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7885 GND a_4769_2176# a_4713_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7886 a_12309_6766# WWL_6 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7887 a_15153_6248# RWL_8 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7888 a_11729_5686# WWL_10 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7889 GND a_4862_556# a_4769_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7890 WBL_24 WWL_27 a_14142_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7891 RBL0_19 RWL_7 a_11443_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7892 RBL0_18 RWL_11 a_10863_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7893 GND a_1869_826# a_1813_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7894 VDD a_1962_4336# a_1869_4336# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7895 WBL_8 WWL_4 a_4862_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7896 a_15882_1096# a_15789_1096# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7897 a_11673_4628# RWL_14 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7898 VDD a_13562_5956# a_13469_5956# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7899 GND a_15882_3256# a_15789_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7900 a_6602_3526# a_6509_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7901 GND a_4282_8386# a_4189_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7902 VDD a_15882_7036# a_15789_7036# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7903 a_1382_1366# a_1289_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7904 a_6602_7306# a_6509_7306# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7905 GND a_3702_7306# a_3609_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7906 WBL_2 WWL_10 a_1382_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7907 a_16369_1366# WWL_26 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7908 VDD a_17622_3796# a_17529_3796# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7909 RBL0_26 RWL_27 a_15503_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7910 VDD a_12402_1636# a_12309_1636# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7911 a_12982_2986# a_12889_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7912 a_17622_7846# a_17529_7846# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7913 a_15302_4066# a_15209_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7914 VDD a_15302_556# a_15209_556# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7915 RBL0_30 RWL_23 a_17823_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7916 a_7089_7576# WWL_3 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7917 WBL_26 WWL_28 a_15302_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7918 WBL_26 WWL_0 a_15302_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7919 WBL_25 WWL_4 a_14722_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7920 RBL0_10 RWL_4 a_6223_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7921 WBL_15 WWL_24 a_8922_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7922 a_3122_8116# a_3029_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7923 WBL_17 WWL_8 a_10082_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7924 RBL0_1 RWL_12 a_1003_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7925 a_17042_4606# a_16949_4606# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7926 GND a_17042_6766# a_16949_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7927 GND a_14049_5686# a_13993_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7929 GND a_8342_2986# a_8249_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7930 a_6453_5438# RWL_11 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7931 GND a_16369_6766# a_16313_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7932 a_1233_3278# RWL_19 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7933 RBL0_4 RWL_10 a_2743_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7934 GND a_7669_2986# a_7613_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7935 a_18403_3818# a_18202_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7936 a_13183_1658# a_12982_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7937 WBL_16 WWL_31 a_9502_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7938 GND a_9989_4066# a_9933_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7939 a_14142_556# a_14049_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7940 a_16949_7576# WWL_3 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7941 a_2973_3818# RWL_17 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7942 a_12309_6496# WWL_7 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7943 a_11729_5416# WWL_11 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7944 VDD a_4862_5146# a_4769_5146# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7945 RBL0_19 RWL_8 a_11443_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7946 RBL0_18 RWL_12 a_10863_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7948 GND a_1869_556# a_1813_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7949 GND a_18202_287# a_18109_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7950 a_16893_6518# RWL_7 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7951 a_12982_5956# a_12889_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7952 a_11673_4358# RWL_15 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7953 GND a_17529_826# a_17473_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7954 GND a_4189_16# a_4133_38# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7955 a_4282_5956# a_4189_5956# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7956 GND a_129_8386# a_73_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7957 a_6602_3256# a_6509_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7958 GND a_4282_8116# a_4189_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7959 a_6602_7036# a_6509_7036# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7960 GND a_3702_7036# a_3609_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7961 VDD a_15302_2446# a_15209_2446# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7962 WBL_11 WWL_3 a_6602_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7963 WBL_2 WWL_11 a_1382_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7964 a_13763_7868# a_13562_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7965 a_16369_1096# WWL_27 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7966 VDD a_17622_3526# a_17529_3526# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7967 a_8342_3796# a_8249_3796# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7968 RBL0_7 RWL_31 a_4483_38# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7969 a_3122_1636# a_3029_1636# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7970 WBL_22 WWL_5 a_12982_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7971 GND a_8342_5956# a_8249_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7972 WBL_22 WWL_30 a_12982_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7973 a_7089_7306# WWL_4 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7974 WBL_26 WWL_1 a_15302_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7975 GND a_7669_5956# a_7613_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7976 RBL0_10 RWL_5 a_6223_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7977 a_17042_4336# a_16949_4336# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7978 RBL0_13 RWL_17 a_7963_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7979 GND a_14049_5416# a_13993_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7980 WBL_20 WWL_21 a_11822_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7981 a_3609_5686# WWL_10 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7982 a_6453_5168# RWL_12 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7983 a_4862_8386# a_4769_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7984 RBL0_4 RWL_11 a_2743_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7985 a_18403_3548# a_18202_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7986 a_13183_1388# a_12982_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7987 GND a_11242_3796# a_11149_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7988 a_13562_2716# a_13469_2716# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7989 VDD a_11242_7576# a_11149_7576# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7990 GND a_4862_1096# a_4769_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7991 GND a_10569_3796# a_10513_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7992 GND a_13562_4876# a_13469_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7993 a_16949_7306# WWL_4 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7994 a_2973_3548# RWL_18 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7995 a_12309_6226# WWL_8 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7996 VDD a_4862_4876# a_4769_4876# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7997 a_14923_1928# a_14722_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7998 GND a_12889_4876# a_12833_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7999 RBL0_22 RWL_21 a_13183_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8000 a_18202_7846# a_18109_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8001 a_16893_6248# RWL_8 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8002 a_17622_6766# a_17529_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8003 GND a_15209_287# a_15153_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8004 VDD a_8922_2716# a_8829_2716# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8005 a_11673_4088# RWL_16 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8006 VDD a_4282_1636# a_4189_1636# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8007 a_9502_7846# a_9409_7846# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8008 GND a_17529_556# a_17473_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8009 a_7669_826# WWL_28 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8010 GND a_129_8116# a_73_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8011 a_11443_6518# a_11242_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8012 VDD a_15302_2176# a_15209_2176# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8013 WBL_11 WWL_4 a_6602_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8014 a_18403_848# a_18202_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8015 a_6022_2446# a_5929_2446# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8016 a_13763_7598# a_13562_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8017 GND a_6022_4606# a_5929_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8018 a_8342_3526# a_8249_3526# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8019 VDD a_6022_8386# a_5929_8386# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8020 WBL_30 WWL_2 a_17622_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8021 GND a_5349_4606# a_5293_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8022 WBL_22 WWL_31 a_12982_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8023 a_9703_2738# a_9502_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8024 a_1003_4628# a_802_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8025 a_129_5686# WWL_10 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8026 VDD a_2542_6766# a_2449_6766# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8028 RBL0_13 RWL_18 a_7963_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8029 a_1289_4336# WWL_15 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8030 WBL_29 WWL_14 a_17042_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8031 GND a_14049_5146# a_13993_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8032 a_4862_8116# a_4769_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8033 a_3609_5416# WWL_11 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8034 RBL0_4 RWL_12 a_2743_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8035 a_11242_1366# a_11149_1366# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8036 a_18403_3278# a_18202_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8037 GND a_16462_5686# a_16369_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8038 GND a_11242_3526# a_11149_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8039 a_15209_7036# WWL_5 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8040 a_14629_5956# WWL_9 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8041 RBL0_7 RWL_24 a_4483_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8042 a_1962_3796# a_1869_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8043 VDD a_11242_7306# a_11149_7306# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8044 GND a_15789_5686# a_15733_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8045 GND a_709_1096# a_653_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8046 a_1962_7576# a_1869_7576# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8047 GND a_10569_3526# a_10513_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8048 a_2973_3278# RWL_19 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8049 a_4282_4876# a_4189_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8050 a_14923_1658# a_14722_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8051 VDD a_7182_2446# a_7089_2446# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8052 a_14049_2716# WWL_21 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8053 a_2743_5708# a_2542_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8054 VDD a_6602_1366# a_6509_1366# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8055 RBL0_31 RWL_14 a_18403_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8056 a_16462_826# a_16369_826# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8057 RBL0_22 RWL_22 a_13183_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8058 a_18202_7576# a_18109_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8059 VDD a_4862_287# a_4769_287# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8060 a_5349_287# WWL_30 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8061 RBL0_3 RWL_31 a_2163_38# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8062 WBL_7 WWL_9 a_4282_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8063 a_16663_8408# a_16462_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8064 a_11443_6248# a_11242_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8065 a_16083_309# a_15882_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8066 VDD a_15302_1906# a_15209_1906# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8067 a_11822_3796# a_11729_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8068 a_18403_578# a_18202_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8069 a_11822_7576# a_11729_7576# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8070 a_6022_2176# a_5929_2176# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8071 GND a_6022_4336# a_5929_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8072 a_4133_6788# RWL_6 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8073 WBL_14 WWL_17 a_8342_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8074 VDD a_6022_8116# a_5929_8116# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8075 GND a_5349_4336# a_5293_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8076 a_9703_2468# a_9502_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8077 a_1003_4358# a_802_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8078 GND a_2542_2716# a_2449_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8079 a_4862_1636# a_4769_1636# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8080 a_129_5416# WWL_11 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8081 a_5929_5146# WWL_12 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8082 RBL0_13 RWL_19 a_7963_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8083 VDD a_2542_6496# a_2449_6496# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8084 a_1289_4066# WWL_16 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8085 GND a_1869_2716# a_1813_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8086 a_16462_3256# a_16369_3256# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8087 a_11242_1096# a_11149_1096# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8088 WBL_19 WWL_25 a_11242_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8089 a_14573_7868# RWL_2 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8090 GND a_16462_5416# a_16369_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8091 a_7182_5686# a_7089_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8092 GND a_11242_3256# a_11149_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8093 RBL0_16 RWL_17 a_9703_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8094 VDD a_10662_826# a_10569_826# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8095 WBL_23 WWL_21 a_13562_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8096 a_1962_3526# a_1869_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8097 VDD a_11242_7036# a_11149_7036# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8098 GND a_15789_5416# a_15733_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8099 a_11149_826# WWL_28 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8100 RBL0_7 RWL_25 a_4483_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8101 a_9502_6766# a_9409_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8102 GND a_10569_3256# a_10513_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8103 a_1962_7306# a_1869_7306# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8104 a_73_848# RWL_28 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8105 a_14923_1388# a_14722_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8106 a_9933_1928# RWL_24 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8107 GND a_12982_3796# a_12889_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8108 a_3323_6518# a_3122_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8109 VDD a_12982_7576# a_12889_7576# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8110 a_2743_5438# a_2542_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8111 a_14142_287# a_14049_287# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8112 VDD a_6602_1096# a_6509_1096# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8113 VDD a_7182_2176# a_7089_2176# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8114 RBL0_31 RWL_15 a_18403_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8115 RBL0_22 RWL_23 a_13183_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8116 VDD a_4862_17# a_4769_17# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8117 a_5349_17# WWL_31 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8118 WBL_16 WWL_2 a_9502_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8119 a_16663_8138# a_16462_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8120 RBL0_25 RWL_21 a_14923_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8121 a_11822_3526# a_11729_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8122 a_12402_4606# a_12309_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8123 a_12402_8386# a_12309_8386# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8124 a_6022_1906# a_5929_1906# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8125 a_11822_7306# a_11729_7306# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8126 RBL0_24 RWL_31 a_14343_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8127 WBL_10 WWL_22 a_6022_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8128 GND a_3029_2986# a_2973_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8129 GND a_6022_4066# a_5929_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8130 WBL_14 WWL_18 a_8342_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8131 a_16083_4898# a_15882_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8132 a_7383_1118# a_7182_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8133 GND a_5349_4066# a_5293_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8134 a_7762_2446# a_7669_2446# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8135 a_9703_2198# a_9502_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8136 RBL0_20 RWL_0 a_12023_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8137 a_1003_4088# a_802_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8138 GND a_7762_4606# a_7669_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8139 GND a_2542_2446# a_2449_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8140 VDD a_7762_8386# a_7669_8386# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8141 a_6509_5956# WWL_9 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8142 a_5929_4876# WWL_13 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8143 VDD a_2542_6226# a_2449_6226# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8144 GND a_1869_2446# a_1813_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8145 a_3609_556# WWL_29 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8146 a_12253_6518# RWL_7 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8147 a_16462_2986# a_16369_2986# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8148 VDD a_14142_7846# a_14049_7846# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8149 GND a_129_826# a_73_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8150 WBL_19 WWL_26 a_11242_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8151 GND a_16462_5146# a_16369_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8152 a_14573_7598# a_13963_7576# RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8153 a_7182_5416# a_7089_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8154 RBL0_16 RWL_18 a_9703_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8155 GND a_15789_5146# a_15733_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8156 RBL0_7 RWL_26 a_4483_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8157 a_1962_3256# a_1869_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8158 GND a_18202_1906# a_18109_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8159 WBL_3 WWL_3 a_1962_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8160 a_1962_7036# a_1869_7036# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8161 a_73_578# RWL_29 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8162 VDD a_18202_5686# a_18109_5686# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8163 GND a_17529_1906# a_17473_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8164 RBL0_27 RWL_20 a_16083_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8165 a_9933_1658# RWL_25 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8166 GND a_12982_3526# a_12889_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8167 a_7963_7328# a_7762_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8168 VDD a_12982_7306# a_12889_7306# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8169 a_3323_6248# a_3122_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8170 a_2743_5168# a_2542_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8171 a_14142_17# a_14049_17# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8172 VDD a_7182_1906# a_7089_1906# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8173 a_3702_3796# a_3609_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8174 RBL0_31 RWL_16 a_18403_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8175 a_3702_7576# a_3609_7576# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8176 GND a_3029_5956# a_2973_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8177 a_13469_1636# WWL_25 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8178 a_15789_2716# WWL_21 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8179 RBL0_25 RWL_22 a_14923_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8180 a_12402_4336# a_12309_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8181 a_7033_7328# RWL_4 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8182 a_11822_3256# a_11729_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8183 a_12402_8116# a_12309_8116# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8184 a_11822_7036# a_11729_7036# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8185 WBL_10 WWL_23 a_6022_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8186 a_3553_5708# RWL_10 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8187 a_7762_2176# a_7669_2176# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8188 a_8922_556# a_8829_556# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8189 RBL0_20 RWL_1 a_12023_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8190 a_12402_556# a_12309_556# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8191 a_15882_17# a_15789_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8192 GND a_7762_4336# a_7669_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8193 a_5873_6788# RWL_6 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8194 a_10283_1928# a_10082_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8195 GND a_2542_2176# a_2449_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8196 VDD a_7762_8116# a_7669_8116# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8197 a_1962_826# a_1869_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8198 GND a_1869_2176# a_1813_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8199 a_3609_286# WWL_30 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8200 a_17473_8408# RWL_0 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8201 a_8249_2446# WWL_22 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8202 VDD a_802_6766# a_709_6766# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8203 a_12253_6248# RWL_8 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8204 RBL0_27 RWL_9 a_16083_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8205 RBL0_29 RWL_28 a_17243_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8206 WBL_28 WWL_19 a_16462_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8207 WBL_19 WWL_27 a_11242_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8208 GND a_129_556# a_73_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8209 a_7182_5146# a_7089_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8210 RBL0_16 RWL_19 a_9703_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8211 GND a_18202_1636# a_18109_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8212 WBL_3 WWL_4 a_1962_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8213 GND a_8342_826# a_8249_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8214 a_8773_39# RWL_31 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8215 a_8922_1906# a_8829_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8216 VDD a_18202_5416# a_18109_5416# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8217 a_222_3796# a_129_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8218 VDD a_10662_5956# a_10569_5956# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8219 a_8922_5686# a_8829_5686# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8220 GND a_17529_1636# a_17473_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8221 a_222_7576# a_129_7576# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8222 a_9933_1388# RWL_26 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8223 GND a_12982_3256# a_12889_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8224 a_7963_7058# a_7762_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8225 a_3702_3526# a_3609_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8226 GND a_1382_8386# a_1289_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8227 VDD a_12982_7036# a_12889_7036# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8228 a_3702_7306# a_3609_7306# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8229 GND a_8249_7846# a_8193_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8230 RBL0_20 RWL_31 a_12023_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8231 a_5063_2738# a_4862_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8232 a_15302_287# a_15209_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8233 a_13469_1366# WWL_26 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8234 VDD a_10082_2716# a_9989_2716# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8235 VDD a_14722_3796# a_14629_3796# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8236 RBL0_21 RWL_27 a_12603_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8237 a_10082_2986# a_9989_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8238 a_14722_7846# a_14629_7846# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8239 VDD a_3122_556# a_3029_556# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8240 RBL0_25 RWL_23 a_14923_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8241 a_12402_4066# a_12309_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8242 a_7033_7058# RWL_5 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8243 a_4189_7576# WWL_3 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8244 WBL_21 WWL_0 a_12402_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8245 RBL0_5 RWL_4 a_3323_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8246 WBL_10 WWL_24 a_6022_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8247 a_14142_4606# a_14049_4606# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8248 GND a_14142_6766# a_14049_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8249 GND a_11149_5686# a_11093_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8250 GND a_5442_2986# a_5349_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8251 a_3553_5438# RWL_11 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8252 a_7762_1906# a_7669_1906# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8253 WBL_13 WWL_22 a_7762_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8254 GND a_13469_6766# a_13413_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8255 GND a_4769_2986# a_4713_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8256 a_15503_3818# a_15302_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8257 GND a_7762_4066# a_7669_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8258 a_10283_1658# a_10082_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8259 a_2743_38# a_2542_16# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8260 a_17823_4898# a_17622_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8261 a_1962_556# a_1869_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8262 a_3609_16# WWL_31 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8263 GND a_802_2716# a_709_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8264 a_17473_8138# RWL_1 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8265 VDD a_802_6496# a_709_6496# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8266 RBL0_29 RWL_29 a_17243_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8267 a_8249_2176# WWL_23 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8268 WBL_28 WWL_20 a_16462_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8269 VDD a_9502_4606# a_9409_4606# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8270 VDD a_1962_5146# a_1869_5146# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8271 a_2743_308# a_2542_286# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8272 GND a_6022_287# a_5929_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8273 GND a_8342_556# a_8249_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8274 GND a_18202_1366# a_18109_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8275 a_13993_6518# RWL_7 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8276 a_8193_1118# RWL_27 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8277 a_8922_1636# a_8829_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8278 VDD a_15882_7846# a_15789_7846# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8279 a_10082_5956# a_9989_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8280 a_222_3526# a_129_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8281 GND a_5349_826# a_5293_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8282 GND a_17529_1366# a_17473_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8283 a_222_7306# a_129_7306# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8284 a_8922_5416# a_8829_5416# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8285 a_1382_5956# a_1289_5956# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8286 a_3702_3256# a_3609_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8287 GND a_1382_8116# a_1289_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8288 a_3702_7036# a_3609_7036# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8289 VDD a_12402_2446# a_12309_2446# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8290 WBL_6 WWL_3 a_3702_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8291 GND a_8249_7576# a_8193_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8292 a_5063_2468# a_4862_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8293 a_10863_7868# a_10662_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8294 a_13469_1096# WWL_27 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8295 RBL0_30 RWL_20 a_17823_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8296 VDD a_14722_3526# a_14629_3526# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8297 a_5442_3796# a_5349_3796# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8298 WBL_17 WWL_5 a_10082_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8299 GND a_5442_5956# a_5349_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8300 VDD a_3122_286# a_3029_286# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8301 a_8829_8386# WWL_0 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8302 a_4189_7306# WWL_4 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8303 WBL_21 WWL_1 a_12402_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8304 GND a_4769_5956# a_4713_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8305 RBL0_5 RWL_5 a_3323_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8306 a_13562_17# a_13469_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8307 a_14142_4336# a_14049_4336# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8308 RBL0_8 RWL_17 a_5063_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8309 GND a_11149_5416# a_11093_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8310 a_8773_7328# RWL_4 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8311 a_3553_5168# RWL_12 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8312 WBL_13 WWL_23 a_7762_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8313 RBL0_12 RWL_13 a_7383_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8314 a_15503_3548# a_15302_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8316 a_10283_1388# a_10082_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8317 a_10662_2716# a_10569_2716# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8318 a_6453_39# RWL_31 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8319 GND a_802_2446# a_709_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8320 GND a_10662_4876# a_10569_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8321 GND a_1962_1096# a_1869_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8322 VDD a_802_6226# a_709_6226# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8323 a_8249_1906# WWL_24 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8324 VDD a_9502_4336# a_9409_4336# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8325 a_14923_39# a_14722_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8326 VDD a_1962_4876# a_1869_4876# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8327 a_12023_1928# a_11822_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8328 WBL_8 WWL_2 a_4862_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8329 RBL0_17 RWL_21 a_10283_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8330 a_15302_7846# a_15209_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8331 a_13993_6248# RWL_8 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8332 RBL0_30 RWL_9 a_17823_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8333 a_9989_2446# WWL_22 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8334 a_14722_6766# a_14629_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8335 a_8922_1366# a_8829_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8336 VDD a_1382_1636# a_1289_1636# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8337 a_222_3256# a_129_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8338 GND a_5349_556# a_5293_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8339 a_6602_7846# a_6509_7846# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8340 a_222_7036# a_129_7036# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8341 WBL_15 WWL_10 a_8922_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8342 WBL_0 WWL_3 a_222_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8343 a_11093_1928# RWL_24 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8344 a_6223_848# a_6022_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8345 VDD a_12402_2176# a_12309_2176# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8346 WBL_6 WWL_4 a_3702_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8347 a_3122_2446# a_3029_2446# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8348 a_10863_7598# a_10662_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8349 a_5063_2198# a_4862_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8350 GND a_3122_4606# a_3029_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8351 a_5442_3526# a_5349_3526# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8352 VDD a_3122_8386# a_3029_8386# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8353 WBL_25 WWL_2 a_14722_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8354 GND a_2449_4606# a_2393_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8355 VDD a_3122_16# a_3029_16# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8356 a_8829_8116# WWL_1 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8357 GND a_9989_7846# a_9933_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8358 a_17042_5146# a_16949_5146# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8359 a_6803_2738# a_6602_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8360 GND a_17042_7306# a_16949_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8361 GND a_16369_7306# a_16313_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8362 RBL0_8 RWL_18 a_5063_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8363 WBL_24 WWL_14 a_14142_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8364 GND a_11149_5146# a_11093_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8365 a_8773_7058# RWL_5 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8366 WBL_13 WWL_24 a_7762_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8367 a_15503_3278# a_15302_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8368 GND a_13562_5686# a_13469_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8369 WBL_18 WWL_28 a_10662_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8370 a_15882_4606# a_15789_4606# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8371 a_12309_7036# WWL_5 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8372 a_11729_5956# WWL_9 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8373 GND a_12889_5686# a_12833_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8374 RBL0_2 RWL_24 a_1583_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8375 GND a_15882_6766# a_15789_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8376 GND a_802_2176# a_709_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8377 a_1382_4876# a_1289_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8378 a_12023_1658# a_11822_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8379 a_12982_6496# a_12889_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8380 VDD a_4282_2446# a_4189_2446# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8381 a_11149_2716# WWL_21 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8382 RBL0_26 RWL_14 a_15503_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8383 VDD a_3702_1366# a_3609_1366# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8384 a_4282_826# a_4189_826# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8385 RBL0_17 RWL_22 a_10283_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8386 a_9989_2176# WWL_23 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8387 a_15302_7576# a_15209_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8388 WBL_15 WWL_11 a_8922_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8389 WBL_0 WWL_4 a_222_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8390 a_16313_3818# RWL_17 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8391 WBL_2 WWL_9 a_1382_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8392 a_11093_1658# RWL_25 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8393 a_15733_2738# RWL_21 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8394 a_13763_8408# a_13562_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8395 VDD a_17622_4066# a_17529_4066# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8396 VDD a_12402_1906# a_12309_1906# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8397 a_6223_578# a_6022_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8398 a_11242_17# a_11149_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8399 a_3122_2176# a_3029_2176# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8400 GND a_8342_6496# a_8249_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8401 GND a_3122_4336# a_3029_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8402 a_7089_7846# WWL_2 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8403 a_1233_6788# RWL_6 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8404 WBL_9 WWL_17 a_5442_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8405 VDD a_3122_8116# a_3029_8116# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8406 GND a_7669_6496# a_7613_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8407 GND a_2449_4336# a_2393_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8408 a_17042_1096# a_16949_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8409 GND a_9989_7576# a_9933_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8410 a_17042_4876# a_16949_4876# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8411 a_6803_2468# a_6602_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8412 GND a_17042_7036# a_16949_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8413 WBL_20 WWL_19 a_11822_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8414 GND a_4282_286# a_4189_286# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8415 RBL0_8 RWL_19 a_5063_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8416 GND a_16369_7036# a_16313_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8417 a_12603_39# a_12402_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8418 a_13562_3256# a_13469_3256# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8419 GND a_18109_3796# a_18053_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8420 a_11673_7868# RWL_2 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8421 GND a_13562_5416# a_13469_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8422 a_16949_7846# WWL_2 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8423 a_4282_5686# a_4189_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8424 RBL0_11 RWL_17 a_6803_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8425 a_15882_4336# a_15789_4336# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8426 RBL0_2 RWL_25 a_1583_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8427 WBL_18 WWL_21 a_10662_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8428 GND a_12889_5416# a_12833_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8429 a_7963_309# a_7762_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8430 a_6602_6766# a_6509_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8431 a_12023_1388# a_11822_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8432 a_18202_8386# a_18109_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8433 a_16369_4606# WWL_14 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8434 a_17622_7306# a_17529_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8435 VDD a_8922_3256# a_8829_3256# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8436 a_12982_6226# a_12889_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8437 VDD a_3702_1096# a_3609_1096# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8438 VDD a_4282_2176# a_4189_2176# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8439 RBL0_26 RWL_15 a_15503_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8440 RBL0_17 RWL_23 a_10283_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8441 a_9989_1906# WWL_24 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8442 WBL_11 WWL_2 a_6602_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8443 a_1003_308# a_802_286# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8444 a_16313_3548# RWL_18 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8445 a_15733_2468# RWL_22 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8446 a_13763_8138# a_13562_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8447 a_3553_308# RWL_30 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8448 a_11093_1388# RWL_26 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8449 VDD a_8342_287# a_8249_287# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8450 a_8342_4066# a_8249_4066# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8451 a_3122_1906# a_3029_1906# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8452 WBL_5 WWL_22 a_3122_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8453 GND a_8342_6226# a_8249_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8454 a_12309_287# WWL_30 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8455 GND a_3122_4066# a_3029_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8456 GND a_7669_6226# a_7613_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8457 WBL_9 WWL_18 a_5442_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8458 a_13183_4898# a_12982_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8459 a_4483_1118# a_4282_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8460 GND a_2449_4066# a_2393_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8461 RBL0_2 RWL_30 a_1583_308# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8462 a_4862_2446# a_4769_2446# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8463 WBL_29 WWL_12 a_17042_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8464 a_6803_2198# a_6602_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8465 a_13763_848# a_13562_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8466 WBL_20 WWL_20 a_11822_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8467 GND a_4862_4606# a_4769_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8468 VDD a_4862_8386# a_4769_8386# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8469 a_3609_5956# WWL_9 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8470 a_423_1928# a_222_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8471 GND a_1289_286# a_1233_308# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8472 a_13562_2986# a_13469_2986# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8473 GND a_18109_3526# a_18053_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8474 VDD a_11242_7846# a_11149_7846# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8475 GND a_13562_5146# a_13469_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8476 a_7669_3796# WWL_17 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8477 a_11673_7598# a_4683_7576# RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8478 a_4282_5416# a_4189_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8479 GND a_14722_17# a_14629_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8480 RBL0_11 RWL_18 a_6803_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8481 GND a_12889_5146# a_12833_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8482 RBL0_2 RWL_26 a_1583_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8483 GND a_15302_1906# a_15209_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8484 VDD a_15302_5686# a_15209_5686# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8485 a_14049_3256# WWL_19 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8486 VDD a_14142_826# a_14049_826# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8487 GND a_14629_1906# a_14573_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8488 a_7613_2738# RWL_21 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8489 RBL0_22 RWL_20 a_13183_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8490 a_18202_8116# a_18109_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8491 a_17622_7036# a_17529_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8492 VDD a_8922_2986# a_8829_2986# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8493 VDD a_4282_1906# a_4189_1906# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8494 RBL0_26 RWL_16 a_15503_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8495 a_10569_1636# WWL_25 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8496 WBL_5 WWL_29 a_3122_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8497 a_15733_2198# RWL_23 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8498 a_16313_3278# RWL_19 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8499 a_12889_2716# WWL_21 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8500 a_4133_7328# RWL_4 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8501 VDD a_8342_17# a_8249_17# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8502 WBL_14 WWL_15 a_8342_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8503 a_16083_5708# a_15882_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8504 a_11822_826# a_11729_826# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8505 WBL_5 WWL_23 a_3122_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8506 a_12309_17# WWL_31 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8507 a_18403_6788# a_18202_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8508 a_9703_3008# a_9502_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8509 a_10283_39# a_10082_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8510 a_4862_2176# a_4769_2176# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8511 a_129_5956# WWL_9 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8512 a_11443_309# a_11242_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8513 GND a_9409_2716# a_9353_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8514 WBL_29 WWL_13 a_17042_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8515 a_13763_578# a_13562_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8516 GND a_709_4606# a_653_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8517 a_2973_6788# RWL_6 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8518 GND a_4862_4336# a_4769_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8519 VDD a_4862_8116# a_4769_8116# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8520 a_423_1658# a_222_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8521 a_14573_8408# RWL_0 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8522 a_5349_2446# WWL_22 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8523 RBL0_22 RWL_9 a_13183_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8524 GND a_18109_3256# a_18053_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8525 WBL_23 WWL_19 a_13562_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8526 a_9502_7306# a_9409_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8527 a_7669_3526# WWL_18 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8528 a_1962_7846# a_1869_7846# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8529 a_4282_5146# a_4189_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8530 a_7089_556# WWL_29 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8531 RBL0_11 RWL_19 a_6803_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8532 GND a_15302_1636# a_15209_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8533 a_18202_1636# a_18109_1636# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8534 a_6022_1906# a_5929_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8535 VDD a_15302_5416# a_15209_5416# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8536 a_14049_2986# WWL_20 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8537 a_6022_5686# a_5929_5686# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8538 GND a_14629_1636# a_14573_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8539 a_7613_2468# RWL_22 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8540 GND a_6022_7846# a_5929_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8541 GND a_5349_7846# a_5293_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8542 a_2163_2738# a_1962_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8543 a_10569_1366# WWL_26 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8544 VDD a_11822_3796# a_11729_3796# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8545 a_9703_5978# a_9502_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8546 a_1003_7868# a_802_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8547 WBL_5 WWL_30 a_3122_286# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8548 a_11822_7846# a_11729_7846# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8549 a_4133_7058# RWL_5 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8550 a_1289_7576# WWL_3 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8551 RBL0_13 RWL_6 a_7963_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8552 WBL_14 WWL_16 a_8342_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8553 a_16083_5438# a_15882_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8554 WBL_5 WWL_24 a_3122_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8555 a_3702_16# a_3609_16# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8556 a_16462_6766# a_16369_6766# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8557 a_11242_4606# a_11149_4606# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8558 GND a_11242_6766# a_11149_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8559 GND a_2542_2986# a_2449_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8560 a_4862_1906# a_4769_1906# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8561 GND a_9409_2446# a_9353_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8562 GND a_10569_6766# a_10513_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8563 GND a_709_4336# a_653_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8564 GND a_1869_2986# a_1813_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8565 a_12603_3818# a_12402_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8566 GND a_4862_4066# a_4769_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8567 GND a_12402_17# a_12309_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8568 a_423_1388# a_222_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8569 a_14923_4898# a_14722_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8570 GND a_7182_1906# a_7089_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8571 a_802_2716# a_709_2716# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8572 a_14573_8138# RWL_1 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8573 RBL0_31 RWL_2 a_18403_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8574 VDD a_7182_5686# a_7089_5686# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8575 a_5349_2176# WWL_23 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8576 VDD a_6602_4606# a_6509_4606# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8577 WBL_23 WWL_20 a_13562_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8578 a_9502_7036# a_9409_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8579 a_5293_1118# RWL_27 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8580 GND a_15302_1366# a_15209_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8581 a_6022_1636# a_5929_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8582 RBL0_0 RWL_21 a_423_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8583 VDD a_12982_7846# a_12889_7846# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8584 a_6022_5416# a_5929_5416# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8585 GND a_14629_1366# a_14573_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8586 a_7613_2198# RWL_23 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8587 a_802_16# a_709_16# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8588 GND a_6022_7576# a_5929_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8589 GND a_3029_6496# a_2973_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8590 a_8773_309# RWL_30 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8591 GND a_5349_7576# a_5293_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8592 a_7383_4628# a_7182_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8593 a_2163_2468# a_1962_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8594 a_15789_3256# WWL_19 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8595 a_10569_1096# WWL_27 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8596 RBL0_25 RWL_20 a_14923_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8597 VDD a_11822_3526# a_11729_3526# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8598 a_1003_7598# a_802_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8599 WBL_5 WWL_31 a_3122_16# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8600 a_2542_3796# a_2449_3796# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8601 GND a_2542_5956# a_2449_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8602 a_5929_8386# WWL_0 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8603 a_1289_7306# WWL_4 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8604 RBL0_11 RWL_30 a_6803_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8605 GND a_1869_5956# a_1813_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8606 a_16083_5168# a_15882_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8607 a_16462_2716# a_16369_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8608 a_16462_6496# a_16369_6496# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8609 a_11242_4336# a_11149_4336# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8610 VDD a_10082_556# a_9989_556# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8611 RBL0_3 RWL_17 a_2163_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8612 a_5873_7328# RWL_4 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8613 a_1962_6766# a_1869_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8614 GND a_9409_2176# a_9353_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8615 RBL0_7 RWL_13 a_4483_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8616 a_17823_5708# a_17622_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8617 GND a_709_4066# a_653_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8618 a_12603_3548# a_12402_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8619 RBL0_27 RWL_7 a_16083_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8620 GND a_7182_1636# a_7089_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8621 RBL0_31 a_13963_7576# a_18403_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8622 VDD a_7182_5416# a_7089_5416# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8623 a_14573_848# RWL_28 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8624 a_5349_1906# WWL_24 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8625 VDD a_6602_4336# a_6509_4336# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8626 WBL_3 WWL_2 a_1962_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8627 VDD a_18202_5956# a_18109_5956# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8628 a_12402_7846# a_12309_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8629 RBL0_25 RWL_9 a_14923_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8630 a_6022_1366# a_5929_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8631 a_11822_6766# a_11729_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8632 RBL0_0 RWL_22 a_423_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8633 a_3702_7846# a_3609_7846# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8634 WBL_10 WWL_10 a_6022_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8635 RBL0_21 RWL_28 a_12603_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8636 GND a_8249_8386# a_8193_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8637 GND a_3029_6226# a_2973_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8638 VDD a_10082_3256# a_9989_3256# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8639 a_14629_556# WWL_29 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8640 a_7762_1906# a_7669_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8641 a_7383_4358# a_7182_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8642 a_1382_16# a_1289_16# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8643 a_15789_2986# WWL_20 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8644 GND a_3702_826# a_3609_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8645 a_2163_2198# a_1962_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8646 a_7762_5686# a_7669_5686# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8647 a_2542_3526# a_2449_3526# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8648 GND a_7762_7846# a_7669_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8649 RBL0_13 RWL_31 a_7963_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8650 a_5929_8116# WWL_1 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8651 a_14142_5146# a_14049_5146# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8652 a_16462_2446# a_16369_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8653 a_3903_2738# a_3702_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8654 GND a_14142_7306# a_14049_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8655 WBL_28 WWL_6 a_16462_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8656 a_16462_6226# a_16369_6226# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8657 RBL0_12 RWL_10 a_7383_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8658 a_10662_287# a_10569_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8659 a_3029_3796# WWL_17 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8660 WBL_19 WWL_14 a_11242_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8661 GND a_13469_7306# a_13413_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8662 RBL0_3 RWL_18 a_2163_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8663 a_5873_7058# RWL_5 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8664 RBL0_16 RWL_6 a_9703_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8665 a_17823_5438# a_17622_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8666 a_12603_3278# a_12402_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8667 GND a_10662_5686# a_10569_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8668 RBL0_27 RWL_8 a_16083_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8669 VDD a_9502_5146# a_9409_5146# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8670 GND a_12982_6766# a_12889_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8671 GND a_7182_1366# a_7089_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8672 a_9933_4898# RWL_13 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8673 a_222_286# a_129_286# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8674 a_12253_309# RWL_30 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8675 WBL_1 WWL_21 a_802_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8676 a_14573_578# RWL_29 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8677 VDD a_222_3796# a_129_3796# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8678 a_10082_6496# a_9989_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8679 VDD a_1382_2446# a_1289_2446# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8680 RBL0_21 RWL_14 a_12603_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8681 a_8922_5956# a_8829_5956# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8682 a_222_7846# a_129_7846# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8683 a_12402_7576# a_12309_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8684 RBL0_0 RWL_23 a_423_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8685 RBL0_17 RWL_30 a_10283_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8686 WBL_10 WWL_11 a_6022_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8687 GND a_8249_8116# a_8193_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8688 RBL0_21 RWL_29 a_12603_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8689 WBL_14 WWL_30 a_8342_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8690 a_13413_3818# RWL_17 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8691 a_12833_2738# RWL_21 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8692 a_5063_3008# a_4862_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8693 a_10863_8408# a_10662_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8694 VDD a_14722_4066# a_14629_4066# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8695 VDD a_10082_2986# a_9989_2986# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8696 a_7762_1636# a_7669_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8697 a_7383_4088# a_7182_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8698 GND a_5442_6496# a_5349_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8699 a_7762_5416# a_7669_5416# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8700 GND a_3702_556# a_3609_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8701 a_4189_7846# WWL_2 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8702 VDD a_802_826# a_709_826# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8703 WBL_4 WWL_17 a_2542_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8704 GND a_7762_7576# a_7669_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8705 GND a_4769_6496# a_4713_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8706 a_14142_1096# a_14049_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8707 a_14142_4876# a_14049_4876# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8708 a_16462_2176# a_16369_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8709 a_3903_2468# a_3702_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8710 GND a_14142_7036# a_14049_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8711 a_8249_5686# WWL_10 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8712 WBL_28 WWL_7 a_16462_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8713 RBL0_12 RWL_11 a_7383_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8714 a_3029_3526# WWL_18 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8715 GND a_13469_7036# a_13413_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8716 RBL0_3 RWL_19 a_2163_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8717 a_10662_3256# a_10569_3256# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8718 a_17823_5168# a_17622_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8719 GND a_9502_1096# a_9409_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8720 GND a_15209_3796# a_15153_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8721 GND a_18202_4876# a_18109_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8722 GND a_10662_5416# a_10569_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8723 GND a_802_2986# a_709_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8724 a_8193_4628# RWL_14 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8725 a_1382_5686# a_1289_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8726 RBL0_6 RWL_17 a_3903_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8727 GND a_17529_4876# a_17473_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8728 VDD a_9502_4876# a_9409_4876# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8729 GND a_8829_1096# a_8773_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8730 a_3702_6766# a_3609_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8731 WBL_24 WWL_28 a_14142_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8732 GND a_16949_17# a_16893_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8733 a_15302_8386# a_15209_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8734 RBL0_30 RWL_7 a_17823_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8735 a_5063_5978# a_4862_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8736 VDD a_222_3526# a_129_3526# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8737 a_13469_4606# WWL_14 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8738 a_14722_7306# a_14629_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8739 a_10082_6226# a_9989_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8740 VDD a_1382_2176# a_1289_2176# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8742 RBL0_21 RWL_15 a_12603_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8743 WBL_6 WWL_2 a_3702_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8744 WBL_14 WWL_31 a_8342_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8745 a_709_1636# WWL_25 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8746 a_13413_3548# RWL_18 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8747 a_12833_2468# RWL_22 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8748 a_10863_8138# a_10662_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8749 a_5442_4066# a_5349_4066# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8750 a_7762_1366# a_7669_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8751 GND a_5442_6226# a_5349_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8752 WBL_13 WWL_10 a_7762_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8753 GND a_9989_8386# a_9933_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8755 GND a_4769_6226# a_4713_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8756 WBL_4 WWL_18 a_2542_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8757 a_10283_4898# a_10082_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8758 a_1583_1118# a_1382_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8759 a_18109_826# WWL_28 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8760 GND a_802_5956# a_709_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8761 WBL_24 WWL_12 a_14142_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8762 a_3903_2198# a_3702_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8763 a_1583_848# a_1382_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8764 GND a_1962_4606# a_1869_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8765 a_8249_5416# WWL_11 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8766 WBL_28 WWL_8 a_16462_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8767 RBL0_12 RWL_12 a_7383_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8768 VDD a_1962_8386# a_1869_8386# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8769 a_15882_5146# a_15789_5146# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8770 WBL_11 WWL_29 a_6602_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8771 a_10662_2986# a_10569_2986# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8772 GND a_15209_3526# a_15153_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8773 GND a_15882_7306# a_15789_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8774 a_8193_4358# RWL_15 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8775 a_222_6766# a_129_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8776 GND a_10662_5146# a_10569_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8777 a_4769_3796# WWL_17 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8778 a_8922_4876# a_8829_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8779 a_1382_5416# a_1289_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8780 RBL0_6 RWL_18 a_3903_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8781 WBL_20 WWL_30 a_11822_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8782 GND a_12402_1906# a_12309_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8783 VDD a_12402_5686# a_12309_5686# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8784 a_11149_3256# WWL_19 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8785 GND a_11729_1906# a_11673_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8786 a_4713_2738# RWL_21 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8787 RBL0_17 RWL_20 a_10283_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8788 a_15302_8116# a_15209_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8789 a_14722_7036# a_14629_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8790 RBL0_30 RWL_8 a_17823_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8791 a_14923_309# a_14722_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8792 VDD a_1382_1906# a_1289_1906# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8793 RBL0_21 RWL_16 a_12603_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8794 WBL_15 WWL_9 a_8922_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8795 WBL_0 WWL_2 a_222_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8796 a_709_1366# WWL_26 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8797 a_12833_2198# RWL_23 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8798 a_13413_3278# RWL_19 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8799 a_1233_7328# RWL_4 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8800 WBL_9 WWL_15 a_5442_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8801 a_13183_5708# a_12982_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8802 VDD a_17042_1366# a_16949_1366# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8803 GND a_9989_8116# a_9933_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8804 WBL_13 WWL_11 a_7762_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8805 a_15503_6788# a_15302_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8806 a_6803_3008# a_6602_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8807 GND a_7089_3796# a_7033_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8808 GND a_6509_2716# a_6453_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8809 WBL_24 WWL_13 a_14142_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8810 a_1583_578# a_1382_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8811 GND a_1962_4336# a_1869_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8812 VDD a_1962_8116# a_1869_8116# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8813 GND a_2542_16# a_2449_16# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8814 a_15882_1096# a_15789_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8815 a_11673_8408# RWL_0 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8816 a_17243_848# a_17042_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8817 GND a_14629_17# a_14573_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8818 a_2449_2446# WWL_22 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8819 a_15882_4876# a_15789_4876# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8820 RBL0_17 RWL_9 a_10283_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8821 GND a_15209_3256# a_15153_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8822 WBL_18 WWL_19 a_10662_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8823 GND a_15882_7036# a_15789_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8824 a_9989_5686# WWL_10 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8825 a_8193_4088# RWL_16 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8826 a_6602_7306# a_6509_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8827 a_4769_3526# WWL_18 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8828 a_1382_5146# a_1289_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8829 RBL0_6 RWL_19 a_3903_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8830 WBL_20 WWL_31 a_11822_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8831 GND a_17622_3796# a_17529_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8832 a_8543_39# a_8342_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8833 GND a_12402_1636# a_12309_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8834 VDD a_17622_7576# a_17529_7576# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8835 a_16369_5146# WWL_12 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8836 a_15302_1636# a_15209_1636# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8837 a_3122_1906# a_3029_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8838 GND a_16949_3796# a_16893_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8839 VDD a_12402_5416# a_12309_5416# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8840 GND a_11729_1636# a_11673_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8841 a_11149_2986# WWL_20 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8842 a_3122_5686# a_3029_5686# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8843 a_4713_2468# RWL_22 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8844 GND a_3122_7846# a_3029_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8845 GND a_2449_7846# a_2393_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8846 a_15733_3008# RWL_20 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8847 a_17042_4606# a_16949_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8848 a_17042_8386# a_16949_8386# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8849 a_6803_5978# a_6602_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8850 WBL_20 WWL_6 a_11822_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8851 a_709_1096# WWL_27 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8852 a_1233_7058# RWL_5 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8853 RBL0_8 RWL_6 a_5063_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8854 WBL_9 WWL_16 a_5442_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8855 a_13183_5438# a_12982_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8856 VDD a_17042_1096# a_16949_1096# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8857 a_13562_6766# a_13469_6766# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8858 WBL_17 WWL_29 a_10082_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8859 GND a_7089_3526# a_7033_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8860 GND a_6509_2446# a_6453_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8861 GND a_1962_4066# a_1869_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8862 GND a_4282_1906# a_4189_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8863 a_12023_4898# a_11822_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8864 VDD a_8922_6766# a_8829_6766# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8865 a_17243_578# a_17042_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8866 a_7669_4336# WWL_15 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8867 a_11673_8138# RWL_1 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8868 RBL0_26 RWL_2 a_15503_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8869 VDD a_4282_5686# a_4189_5686# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8870 a_2449_2176# WWL_23 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8871 VDD a_3702_4606# a_3609_4606# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8872 WBL_18 WWL_20 a_10662_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8873 a_9989_5416# WWL_11 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8874 a_6602_7036# a_6509_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8875 a_17622_1366# a_17529_1366# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8876 a_18202_2446# a_18109_2446# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8877 GND a_17622_3526# a_17529_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8878 a_15733_5978# RWL_9 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8879 GND a_12402_1366# a_12309_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8880 a_2393_1118# RWL_27 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8881 a_8342_3796# a_8249_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8882 a_11093_4898# RWL_13 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8883 VDD a_17622_7306# a_17529_7306# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8884 a_3122_1636# a_3029_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8885 GND a_16949_3526# a_16893_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8886 a_16369_4876# WWL_13 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8887 a_8342_7576# a_8249_7576# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8888 a_3122_5416# a_3029_5416# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8889 GND a_11729_1366# a_11673_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8890 a_4713_2198# RWL_23 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8891 GND a_3122_7576# a_3029_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8892 GND a_2449_7576# a_2393_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8893 a_17042_4336# a_16949_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8894 a_4483_4628# a_4282_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8895 a_12889_3256# WWL_19 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8896 a_17042_8116# a_16949_8116# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8897 WBL_20 WWL_7 a_11822_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8898 a_18403_7328# a_18202_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8899 a_7762_556# a_7669_556# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8900 a_13183_5168# a_12982_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8901 a_13562_2716# a_13469_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8902 a_13562_6496# a_13469_6496# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8903 a_2973_7328# RWL_4 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8904 GND a_12309_17# a_12253_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8905 a_14923_5708# a_14722_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8906 GND a_6509_2176# a_6453_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8907 GND a_7089_3256# a_7033_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8908 RBL0_2 RWL_13 a_1583_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8909 a_14049_6766# WWL_6 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8910 RBL0_22 RWL_7 a_13183_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8911 GND a_129_1906# a_73_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8912 GND a_8922_2716# a_8829_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8913 GND a_4282_1636# a_4189_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8914 VDD a_8922_6496# a_8829_6496# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8915 a_7669_4066# WWL_16 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8916 RBL0_26 a_13963_7576# a_15503_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8917 VDD a_4282_5416# a_4189_5416# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8918 a_2393_848# RWL_28 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8919 a_2449_1906# WWL_24 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8920 VDD a_3702_4336# a_3609_4336# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8921 a_17622_1096# a_17529_1096# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8922 a_18202_2176# a_18109_2176# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8923 WBL_30 WWL_25 a_17622_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8924 VDD a_15302_5956# a_15209_5956# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8925 a_16313_6788# RWL_6 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8926 a_7613_3008# RWL_20 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8927 GND a_17622_3256# a_17529_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8928 a_8342_3526# a_8249_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8929 GND a_6022_8386# a_5929_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8930 VDD a_17622_7036# a_17529_7036# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8931 a_3122_1366# a_3029_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8932 a_8342_7306# a_8249_7306# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8933 GND a_16949_3256# a_16893_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8934 WBL_5 WWL_10 a_3122_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8935 GND a_5349_8386# a_5293_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8936 VDD a_1962_556# a_1869_556# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8937 a_9703_6518# a_9502_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8938 a_2449_556# WWL_29 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8939 a_1003_8408# a_802_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8940 a_4862_1906# a_4769_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8941 a_4483_4358# a_4282_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8942 a_12889_2986# WWL_20 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8943 a_17042_4066# a_16949_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8944 WBL_29 WWL_0 a_17042_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8945 a_4862_5686# a_4769_5686# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8946 RBL0_13 RWL_4 a_7963_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8947 WBL_20 WWL_8 a_11822_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8948 GND a_4862_7846# a_4769_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8949 a_18403_7058# a_18202_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8950 a_11242_5146# a_11149_5146# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8951 a_13562_2446# a_13469_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8952 GND a_11242_7306# a_11149_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8953 WBL_23 WWL_6 a_13562_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8954 a_13562_6226# a_13469_6226# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8955 GND a_18109_6766# a_18053_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8956 RBL0_7 RWL_10 a_4483_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8957 GND a_9409_2986# a_9353_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8958 GND a_10569_7306# a_10513_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8959 a_2973_7058# RWL_5 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8960 RBL0_11 RWL_6 a_6803_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8961 a_14923_5438# a_14722_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8962 a_16462_826# a_16369_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8963 a_9502_1366# a_9409_1366# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8964 a_802_3256# a_709_3256# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8965 RBL0_31 RWL_0 a_18403_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8966 a_14049_6496# WWL_7 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8967 VDD a_6602_5146# a_6509_5146# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8968 RBL0_22 RWL_8 a_13183_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8969 GND a_129_1636# a_73_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8970 GND a_8922_2446# a_8829_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8971 a_7613_5978# RWL_9 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8972 GND a_4862_287# a_4769_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8973 GND a_4282_1366# a_4189_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8974 VDD a_8922_6226# a_8829_6226# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8975 a_2393_578# RWL_29 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8976 a_18202_1906# a_18109_1906# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8977 WBL_31 WWL_22 a_18202_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8978 WBL_30 WWL_26 a_17622_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8979 a_6022_5956# a_5929_5956# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8980 a_18053_848# RWL_28 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8981 a_8342_3256# a_8249_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8982 GND a_6022_8116# a_5929_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8983 WBL_14 WWL_3 a_8342_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8984 a_8342_7036# a_8249_7036# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8985 a_11242_556# a_11149_556# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8986 WBL_5 WWL_11 a_3122_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8987 GND a_5349_8116# a_5293_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8988 a_10513_3818# RWL_17 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8989 a_2163_3008# a_1962_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8990 VDD a_1962_286# a_1869_286# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8991 VDD a_11822_4066# a_11729_4066# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8992 a_9703_6248# a_9502_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8993 a_2449_286# WWL_30 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8994 a_1003_8138# a_802_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8995 RBL0_27 RWL_28 a_16083_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8996 a_4862_1636# a_4769_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8997 a_4483_4088# a_4282_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8998 GND a_2542_6496# a_2449_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8999 WBL_29 WWL_1 a_17042_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9000 GND a_9409_5956# a_9353_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9001 a_4862_5416# a_4769_5416# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9002 a_1289_7846# WWL_2 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9003 GND a_709_7846# a_653_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9004 RBL0_13 RWL_5 a_7963_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9005 VDD a_17622_556# a_17529_556# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9006 GND a_4862_7576# a_4769_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9007 GND a_1869_6496# a_1813_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9008 a_11242_1096# a_11149_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9009 a_423_4898# a_222_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9010 a_11242_4876# a_11149_4876# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9011 GND a_10662_826# a_10569_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9012 a_13562_2176# a_13469_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9013 GND a_11242_7036# a_11149_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9014 WBL_23 WWL_7 a_13562_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9015 a_5349_5686# WWL_10 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9017 a_1962_7306# a_1869_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9018 RBL0_7 RWL_11 a_4483_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9019 GND a_10569_7036# a_10513_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9020 a_14923_5168# a_14722_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9021 a_9933_5708# RWL_10 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9022 GND a_6602_1096# a_6509_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9023 a_14142_287# a_14049_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9024 GND a_12309_3796# a_12253_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9025 GND a_15302_4876# a_15209_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9026 a_16462_556# a_16369_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9027 a_9502_1096# a_9409_1096# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9028 WBL_16 WWL_25 a_9502_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9029 a_802_2986# a_709_2986# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9030 a_5293_4628# RWL_14 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9031 RBL0_31 RWL_1 a_18403_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9032 a_14049_6226# WWL_8 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9033 VDD a_7182_5956# a_7089_5956# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9034 GND a_129_1366# a_73_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9035 a_16663_1928# a_16462_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9036 GND a_14629_4876# a_14573_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9037 VDD a_6602_4876# a_6509_4876# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9038 GND a_5929_1096# a_5873_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9039 GND a_8922_2176# a_8829_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9040 WBL_3 WWL_28 a_1962_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9042 a_15789_6766# WWL_6 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9043 WBL_31 WWL_23 a_18202_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9044 a_12402_8386# a_12309_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9045 RBL0_25 RWL_7 a_14923_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9046 a_2163_5978# a_1962_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9047 WBL_30 WWL_27 a_17622_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9048 RBL0_15 RWL_27 a_9123_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9049 VDD a_6022_1636# a_5929_1636# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9050 a_10569_4606# WWL_14 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9051 a_11822_7306# a_11729_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9052 RBL0_0 RWL_20 a_423_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9053 a_18053_578# RWL_29 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9054 WBL_14 WWL_4 a_8342_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9055 a_653_1118# RWL_27 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9056 a_10513_3548# RWL_18 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9057 VDD a_1962_16# a_1869_16# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9058 a_2449_16# WWL_31 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9059 a_2542_4066# a_2449_4066# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9060 GND a_7762_8386# a_7669_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9061 RBL0_27 RWL_29 a_16083_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9062 a_4862_1366# a_4769_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9063 GND a_2542_6226# a_2449_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9064 GND a_709_7576# a_653_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9065 WBL_26 WWL_30 a_15302_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9066 GND a_1869_6226# a_1813_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9067 VDD a_16462_2716# a_16369_2716# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9068 a_16462_2986# a_16369_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9069 WBL_19 WWL_12 a_11242_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9070 GND a_10082_17# a_9989_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9071 a_3029_4336# WWL_15 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9072 GND a_10662_556# a_10569_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9073 RBL0_16 RWL_4 a_9703_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9074 a_5349_5416# WWL_11 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9075 a_1962_7036# a_1869_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9076 WBL_23 WWL_8 a_13562_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9077 RBL0_7 RWL_12 a_4483_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9078 GND a_18202_5686# a_18109_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9079 GND a_17529_5686# a_17473_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9080 GND a_12982_7306# a_12889_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9081 a_9933_5438# RWL_11 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9082 GND a_12309_3526# a_12253_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9083 WBL_16 WWL_26 a_9502_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9084 a_5293_4358# RWL_15 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9085 RBL0_0 RWL_9 a_423_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9086 WBL_1 WWL_19 a_802_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9087 a_1869_3796# WWL_17 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9088 a_6022_4876# a_5929_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9089 a_16663_1658# a_16462_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9090 VDD a_10082_6766# a_9989_6766# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9091 a_7383_7868# a_7182_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9092 a_15789_6496# WWL_7 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9093 a_1813_2738# RWL_21 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9094 a_12402_8116# a_12309_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9095 WBL_31 WWL_24 a_18202_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9096 a_11822_7036# a_11729_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9097 RBL0_25 RWL_8 a_14923_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9098 GND a_17529_287# a_17473_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9099 WBL_10 WWL_9 a_6022_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9100 a_9989_826# WWL_28 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9101 RBL0_20 RWL_24 a_12023_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9102 a_16462_5956# a_16369_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9103 a_10513_3278# RWL_19 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9104 a_7762_5956# a_7669_5956# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9105 WBL_4 WWL_15 a_2542_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9106 GND a_7762_8116# a_7669_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9107 a_10283_5708# a_10082_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9108 VDD a_14142_1366# a_14049_1366# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9109 WBL_26 WWL_31 a_15302_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9110 a_12603_6788# a_12402_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9111 a_709_556# WWL_29 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9112 a_3903_3008# a_3702_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9113 a_7182_2716# a_7089_2716# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9114 WBL_28 WWL_5 a_16462_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9115 GND a_4189_3796# a_4133_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9116 a_3029_4066# WWL_16 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9117 GND a_7182_4876# a_7089_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9118 GND a_3609_2716# a_3553_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9119 WBL_19 WWL_13 a_11242_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9121 RBL0_16 RWL_5 a_9703_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9122 a_9502_17# a_9409_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9123 GND a_18202_5416# a_18109_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9124 a_8922_5686# a_8829_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9125 a_5063_848# a_4862_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9126 WBL_27 WWL_17 a_15882_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9127 GND a_17529_5416# a_17473_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9128 GND a_12309_3256# a_12253_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9129 GND a_12982_7036# a_12889_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9130 a_9933_5168# RWL_12 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9131 WBL_16 WWL_27 a_9502_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9132 a_5293_4088# RWL_16 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9133 a_3702_7306# a_3609_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9134 WBL_1 WWL_20 a_802_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9135 a_1869_3526# WWL_18 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9136 a_16663_1388# a_16462_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9137 GND a_14722_3796# a_14629_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9138 GND a_10082_2716# a_9989_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9139 VDD a_14722_7576# a_14629_7576# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9140 a_5063_6518# a_4862_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9141 a_13469_5146# WWL_12 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9142 a_12402_1636# a_12309_1636# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9143 VDD a_222_4066# a_129_4066# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9144 VDD a_10082_6496# a_9989_6496# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9145 a_7383_7598# a_7182_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9146 a_15789_6226# WWL_8 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9147 a_1813_2468# RWL_22 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9148 a_7669_287# WWL_30 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9149 RBL0_28 RWL_21 a_16663_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9150 a_12833_3008# RWL_20 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9151 RBL0_29 RWL_17 a_17243_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9152 a_14142_4606# a_14049_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9153 RBL0_20 RWL_25 a_12023_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9154 a_14142_8386# a_14049_8386# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9155 a_18403_309# a_18202_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9156 a_3903_5978# a_3702_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9157 VDD a_7762_1636# a_7669_1636# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9158 RBL0_3 RWL_6 a_2163_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9159 a_17473_1928# RWL_24 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9160 WBL_4 WWL_16 a_2542_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9161 a_10283_5438# a_10082_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9162 VDD a_14142_1096# a_14049_1096# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9163 a_10662_6766# a_10569_6766# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9164 GND a_802_6496# a_709_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9165 a_709_286# WWL_30 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9166 GND a_9502_4606# a_9409_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9167 VDD a_9502_8386# a_9409_8386# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9168 a_8249_5956# WWL_9 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9169 a_3122_826# a_3029_826# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9170 GND a_2449_16# a_2393_38# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9171 GND a_4189_3526# a_4133_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9172 GND a_8829_4606# a_8773_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9173 GND a_3609_2446# a_3553_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9174 GND a_1382_1906# a_1289_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9175 GND a_18202_5146# a_18109_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9176 a_222_7306# a_129_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9177 a_8922_5416# a_8829_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9178 a_5063_578# a_4862_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9179 WBL_27 WWL_18 a_15882_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9180 a_4769_4336# WWL_15 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9181 RBL0_21 RWL_2 a_12603_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9182 VDD a_1382_5686# a_1289_5686# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9183 VDD a_9502_826# a_9409_826# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9184 GND a_17529_5146# a_17473_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9185 VDD a_12982_826# a_12889_826# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9186 a_3702_7036# a_3609_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9187 a_13469_826# WWL_28 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9188 a_15302_2446# a_15209_2446# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9189 a_14722_1366# a_14629_1366# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9190 GND a_14722_3526# a_14629_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9191 a_12833_5978# RWL_9 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9192 GND a_10082_2446# a_9989_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9193 VDD a_14722_7306# a_14629_7306# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9194 a_5063_6248# a_4862_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9195 a_5442_3796# a_5349_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9196 a_13469_4876# WWL_13 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9197 VDD a_10082_6226# a_9989_6226# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9198 a_5442_7576# a_5349_7576# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9199 a_16462_287# a_16369_287# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9200 GND a_3122_286# a_3029_286# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9201 a_1813_2198# RWL_23 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9202 a_7762_4876# a_7669_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9203 VDD a_222_556# a_129_556# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9204 a_18109_3796# WWL_17 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9205 a_7669_17# WWL_31 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9206 a_17529_2716# WWL_21 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9207 RBL0_28 RWL_22 a_16663_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9208 RBL0_29 RWL_18 a_17243_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9209 a_14142_4336# a_14049_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9210 a_1583_4628# a_1382_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9211 RBL0_20 RWL_26 a_12023_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9212 a_14142_8116# a_14049_8116# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9213 WBL_13 WWL_9 a_7762_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9214 a_17473_1658# RWL_25 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9215 a_15503_7328# a_15302_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9216 a_10283_5168# a_10082_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9217 a_10662_2716# a_10569_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9218 WBL_8 WWL_25 a_4862_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9219 a_10662_6496# a_10569_6496# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9220 a_7182_17# a_7089_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9221 a_8193_7868# RWL_2 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9222 GND a_802_6226# a_709_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9223 a_709_16# WWL_31 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9224 GND a_9502_4336# a_9409_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9225 VDD a_9502_8116# a_9409_8116# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9226 WBL_12 WWL_21 a_7182_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9227 GND a_8829_4336# a_8773_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9228 a_12023_5708# a_11822_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9229 GND a_3609_2176# a_3553_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9230 GND a_4189_3256# a_4133_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9231 VDD a_15882_1366# a_15789_1366# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9232 a_11149_6766# WWL_6 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9233 RBL0_17 RWL_7 a_10283_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9234 GND a_1382_1636# a_1289_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9235 a_222_7036# a_129_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9236 a_8922_5146# a_8829_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9237 a_4769_4066# WWL_16 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9238 RBL0_21 a_4683_7576# a_12603_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9239 VDD a_1382_5416# a_1289_5416# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9240 VDD a_10662_287# a_10569_287# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9241 a_11149_287# WWL_30 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9242 a_11093_5708# RWL_10 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9243 a_14722_1096# a_14629_1096# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9244 WBL_25 WWL_25 a_14722_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9245 a_15302_2176# a_15209_2176# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9246 VDD a_12402_5956# a_12309_5956# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9247 GND a_14722_3256# a_14629_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9248 a_13413_6788# RWL_6 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9249 GND a_10082_2176# a_9989_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9250 a_4713_3008# RWL_20 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9251 RBL0_14 RWL_21 a_8543_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9252 a_5442_3526# a_5349_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9253 GND a_3122_8386# a_3029_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9254 VDD a_14722_7036# a_14629_7036# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9255 RBL0_25 RWL_31 a_14923_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9256 a_5442_7306# a_5349_7306# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9257 a_16462_17# a_16369_17# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9258 GND a_2449_8386# a_2393_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9259 VDD a_222_286# a_129_286# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9260 a_6803_6518# a_6602_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9261 a_18109_3526# WWL_18 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9262 RBL0_29 RWL_19 a_17243_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9263 a_14142_4066# a_14049_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9264 a_1583_4358# a_1382_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9265 WBL_30 WWL_29 a_17622_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9266 RBL0_28 RWL_23 a_16663_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9267 WBL_24 WWL_0 a_14142_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9268 RBL0_8 RWL_4 a_5063_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9269 GND a_1962_7846# a_1869_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9270 a_17473_1388# RWL_26 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9271 a_15503_7058# a_15302_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9272 a_15882_4606# a_15789_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9273 a_10662_2446# a_10569_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9274 a_15882_8386# a_15789_8386# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9275 WBL_18 WWL_6 a_10662_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9276 GND a_15209_6766# a_15153_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9277 a_10662_6226# a_10569_6226# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9278 WBL_8 WWL_26 a_4862_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9279 a_8193_7598# a_4683_7576# RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9280 RBL0_2 RWL_10 a_1583_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9281 GND a_6509_2986# a_6453_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9282 a_17243_3818# a_17042_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9283 GND a_9502_4066# a_9409_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9284 RBL0_6 RWL_6 a_3903_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9285 GND a_8829_4066# a_8773_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9286 a_12023_5438# a_11822_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9287 VDD a_15882_1096# a_15789_1096# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9288 a_6602_1366# a_6509_1366# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9289 a_4282_826# a_4189_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9290 a_73_2738# RWL_21 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9291 RBL0_26 RWL_0 a_15503_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9292 a_11149_6496# WWL_7 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9293 VDD a_3702_5146# a_3609_5146# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9294 RBL0_17 RWL_8 a_10283_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9295 a_4713_5978# RWL_9 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9296 a_9989_5956# WWL_9 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9297 GND a_1382_1366# a_1289_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9298 VDD a_10662_17# a_10569_17# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9299 a_11149_17# WWL_31 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9300 a_15733_6518# RWL_7 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9301 a_7089_1636# WWL_25 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9302 a_11093_5438# RWL_11 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9303 a_15302_1906# a_15209_1906# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9304 WBL_26 WWL_22 a_15302_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9305 VDD a_17622_7846# a_17529_7846# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9306 WBL_25 WWL_26 a_14722_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9307 a_3122_5956# a_3029_5956# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9308 a_9409_2716# WWL_21 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9309 a_709_4606# WWL_14 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9310 RBL0_14 RWL_22 a_8543_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9311 a_5442_3256# a_5349_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9312 GND a_3122_8116# a_3029_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9313 WBL_9 WWL_3 a_5442_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9314 a_5442_7036# a_5349_7036# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9315 VDD a_222_16# a_129_16# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9316 GND a_2449_8116# a_2393_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9317 VDD a_17042_4606# a_16949_4606# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9318 a_6803_6248# a_6602_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9319 WBL_20 WWL_5 a_11822_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9320 a_1583_4088# a_1382_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9321 WBL_24 WWL_1 a_14142_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9322 GND a_6509_5956# a_6453_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9323 VDD a_5442_556# a_5349_556# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9324 RBL0_8 RWL_5 a_5063_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9325 a_16949_1636# WWL_25 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9326 GND a_1962_7576# a_1869_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9327 a_15882_4336# a_15789_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9328 a_10662_2176# a_10569_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9329 a_15882_8116# a_15789_8116# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9330 WBL_18 WWL_7 a_10662_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9331 a_2449_5686# WWL_10 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9332 WBL_8 WWL_27 a_4862_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9333 RBL0_2 RWL_11 a_1583_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9334 a_17243_3548# a_17042_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9335 a_9933_848# RWL_28 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9336 a_12982_3796# a_12889_3796# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9337 a_12023_5168# a_11822_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9338 GND a_3702_1096# a_3609_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9339 a_2393_4628# RWL_14 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9340 GND a_12402_4876# a_12309_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9341 a_16369_8386# WWL_0 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9342 a_4282_556# a_4189_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9343 a_6223_39# a_6022_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9344 a_6602_1096# a_6509_1096# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9345 WBL_11 WWL_25 a_6602_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9346 a_73_2468# RWL_22 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9347 RBL0_26 RWL_1 a_15503_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9348 a_11149_6226# WWL_8 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9349 VDD a_4282_5956# a_4189_5956# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9350 RBL0_29 RWL_30 a_17243_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9351 a_13763_1928# a_13562_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9352 GND a_11729_4876# a_11673_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9353 VDD a_3702_4876# a_3609_4876# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9354 RBL0_21 RWL_31 a_12603_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9355 a_17042_7846# a_16949_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9356 a_16313_7328# RWL_4 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9357 a_15733_6248# RWL_8 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9358 GND a_8342_287# a_8249_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9359 a_12889_6766# WWL_6 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9360 a_11093_5168# RWL_12 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9361 a_7089_1366# WWL_26 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9362 WBL_26 WWL_23 a_15302_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9363 VDD a_8342_3796# a_8249_3796# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9364 RBL0_10 RWL_27 a_6223_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9365 WBL_25 WWL_27 a_14722_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9366 VDD a_3122_1636# a_3029_1636# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9367 a_8342_7846# a_8249_7846# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9368 GND a_7669_826# a_7613_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9369 RBL0_14 RWL_23 a_8543_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9370 WBL_9 WWL_4 a_5442_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9371 VDD a_17042_4336# a_16949_4336# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9372 GND a_4862_8386# a_4769_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9373 GND a_7089_6766# a_7033_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9374 a_9123_3818# a_8922_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9375 a_423_5708# a_222_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9376 a_8543_2738# a_8342_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9377 a_16949_1366# WWL_26 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9378 VDD a_13562_2716# a_13469_2716# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9379 a_13562_2986# a_13469_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9380 GND a_18109_7306# a_18053_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9381 a_15882_4066# a_15789_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9382 a_7669_7576# WWL_3 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9383 RBL0_11 RWL_4 a_6803_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9384 a_2449_5416# WWL_11 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9385 WBL_18 WWL_8 a_10662_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9386 RBL0_2 RWL_12 a_1583_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9387 a_18202_1906# a_18109_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9388 a_17243_3278# a_17042_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9389 GND a_15302_5686# a_15209_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9390 a_18202_5686# a_18109_5686# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9391 GND a_14142_826# a_14049_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9392 a_17622_4606# a_17529_4606# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9393 a_9933_578# RWL_29 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9394 a_12982_3526# a_12889_3526# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9395 a_14049_7036# WWL_5 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9396 GND a_17622_6766# a_17529_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9397 GND a_14629_5686# a_14573_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9398 GND a_8922_2986# a_8829_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9399 a_7613_6518# RWL_7 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9400 a_16369_8116# WWL_1 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9401 WBL_11 WWL_26 a_6602_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9402 a_73_2198# RWL_23 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9403 a_2393_4358# RWL_15 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9404 a_3122_4876# a_3029_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9405 GND a_16949_6766# a_16893_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9406 a_13763_1658# a_13562_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9407 GND a_8342_17# a_8249_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9408 VDD a_6022_2446# a_5929_2446# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9409 a_4483_7868# a_4282_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9410 a_16313_7058# RWL_5 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9411 a_653_308# RWL_30 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9412 a_17042_7576# a_16949_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9413 a_12889_6496# WWL_7 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9414 a_7089_1096# WWL_27 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9415 VDD a_8342_3526# a_8249_3526# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9416 WBL_26 WWL_24 a_15302_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9417 GND a_5349_287# a_5293_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9418 a_11822_826# a_11729_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9419 a_18053_3818# RWL_17 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9420 WBL_5 WWL_9 a_3122_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9421 GND a_7669_556# a_7613_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9422 a_13562_5956# a_13469_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9423 GND a_9409_6496# a_9353_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9424 a_4862_5956# a_4769_5956# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9425 GND a_709_8386# a_653_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9426 GND a_4862_8116# a_4769_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9427 VDD a_11242_1366# a_11149_1366# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9428 a_9123_3548# a_8922_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9429 a_423_5438# a_222_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9430 a_8543_2468# a_8342_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9431 a_16949_1096# WWL_27 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9432 a_802_6766# a_709_6766# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9433 a_4282_2716# a_4189_2716# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9434 WBL_23 WWL_5 a_13562_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9435 GND a_18109_7036# a_18053_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9436 GND a_8922_5956# a_8829_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9437 GND a_1289_3796# a_1233_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9438 GND a_4282_4876# a_4189_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9439 a_7669_7306# WWL_4 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9440 RBL0_11 RWL_5 a_6803_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9441 a_18202_1636# a_18109_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9442 a_18202_5416# a_18109_5416# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9443 GND a_15302_5416# a_15209_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9444 a_6022_5686# a_5929_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9445 GND a_14142_556# a_14049_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9446 RBL0_17 RWL_31 a_10283_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9447 a_17622_4336# a_17529_4336# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9448 WBL_22 WWL_17 a_12982_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9449 GND a_14629_5416# a_14573_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9450 GND a_11149_826# a_11093_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9451 a_7613_6248# RWL_8 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9452 a_8342_6766# a_8249_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9453 WBL_11 WWL_27 a_6602_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9454 a_2393_4088# RWL_16 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9455 a_13763_1388# a_13562_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9456 GND a_11822_3796# a_11729_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9457 a_2163_6518# a_1962_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9458 VDD a_11822_7576# a_11729_7576# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9459 a_10569_5146# WWL_12 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9460 VDD a_6022_2176# a_5929_2176# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9461 WBL_0 WWL_29 a_222_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9462 a_4483_7598# a_4282_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9463 a_12889_6226# WWL_8 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9464 a_6602_826# a_6509_826# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9465 WBL_14 WWL_2 a_8342_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9466 a_11822_556# a_11729_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9467 a_18053_3548# RWL_18 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9468 RBL0_24 RWL_17 a_14343_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9469 RBL0_23 RWL_21 a_13763_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9470 a_11242_4606# a_11149_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9471 a_11242_8386# a_11149_8386# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9472 a_6223_309# a_6022_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9473 VDD a_4862_1636# a_4769_1636# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9474 GND a_709_8116# a_653_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9475 GND a_9409_6226# a_9353_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9476 a_14573_1928# RWL_24 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9477 VDD a_16462_3256# a_16369_3256# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9478 VDD a_11242_1096# a_11149_1096# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9479 a_423_5168# a_222_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9480 a_1962_1366# a_1869_1366# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9481 a_8543_2198# a_8342_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9482 a_802_2716# a_709_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9483 a_9123_3278# a_8922_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9484 GND a_7182_5686# a_7089_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9485 GND a_6602_4606# a_6509_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9486 a_9502_4606# a_9409_4606# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9487 a_802_6496# a_709_6496# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9488 VDD a_6602_8386# a_6509_8386# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9489 a_5349_5956# WWL_9 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9490 GND a_129_4876# a_73_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9491 GND a_1289_3526# a_1233_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9492 GND a_5929_4606# a_5873_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9493 a_18202_1366# a_18109_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9494 GND a_15302_5146# a_15209_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9495 WBL_18 WWL_30 a_10662_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9496 WBL_31 WWL_10 a_18202_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9497 GND a_6022_17# a_5929_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9498 RBL0_15 RWL_14 a_9123_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9499 WBL_30 WWL_14 a_17622_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9500 RBL0_0 RWL_7 a_423_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9501 a_6022_5416# a_5929_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9502 WBL_22 WWL_18 a_12982_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9503 a_1869_4336# WWL_15 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9504 GND a_14629_5146# a_14573_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9505 GND a_11149_556# a_11093_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9506 a_1289_826# WWL_28 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9507 a_12402_2446# a_12309_2446# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9508 a_11822_1366# a_11729_1366# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9509 a_9353_2738# RWL_21 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9510 GND a_11822_3526# a_11729_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9511 a_653_4628# RWL_14 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9512 a_7383_8408# a_7182_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9513 a_15789_7036# WWL_5 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9514 a_11822_17# a_11729_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9515 VDD a_11822_7306# a_11729_7306# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9516 a_2163_6248# a_1962_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9517 VDD a_6022_1906# a_5929_1906# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9518 a_2542_3796# a_2449_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9519 a_10569_4876# WWL_13 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9520 WBL_0 WWL_30 a_222_286# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9521 a_2542_7576# a_2449_7576# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9522 a_4862_4876# a_4769_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9523 a_18053_3278# RWL_19 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9524 a_15209_3796# WWL_17 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9525 a_16462_6496# a_16369_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9526 VDD a_7762_2446# a_7669_2446# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9527 a_14629_2716# WWL_21 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9528 RBL0_23 RWL_22 a_13763_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9529 RBL0_24 RWL_18 a_14343_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9530 a_11242_4336# a_11149_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9531 a_11242_8116# a_11149_8116# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9532 a_14573_1658# RWL_25 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9533 a_12603_7328# a_12402_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9534 VDD a_16462_2986# a_16369_2986# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9535 a_7182_3256# a_7089_3256# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9536 a_1962_1096# a_1869_1096# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9537 WBL_3 WWL_25 a_1962_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9538 GND a_7182_5416# a_7089_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9539 RBL0_6 RWL_30 a_3903_308# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9540 a_802_2446# a_709_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9541 a_5293_7868# RWL_2 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9542 GND a_6602_4336# a_6509_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9543 a_9502_4336# a_9409_4336# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9544 WBL_1 WWL_6 a_802_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9545 a_802_6226# a_709_6226# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9546 VDD a_6602_8116# a_6509_8116# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9547 WBL_7 WWL_21 a_4282_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9548 GND a_1289_3256# a_1233_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9549 GND a_5929_4336# a_5873_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9550 VDD a_12982_1366# a_12889_1366# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9551 WBL_27 WWL_15 a_15882_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9552 a_10082_826# a_9989_826# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9553 WBL_18 WWL_31 a_10662_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9554 WBL_31 WWL_11 a_18202_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9555 RBL0_15 RWL_15 a_9123_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9556 RBL0_0 RWL_8 a_423_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9557 a_6022_5146# a_5929_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9558 a_1869_4066# WWL_16 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9559 a_11822_1096# a_11729_1096# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9560 a_12402_2176# a_12309_2176# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9561 a_9353_2468# RWL_22 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9562 GND a_11822_3256# a_11729_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9563 a_653_4358# RWL_15 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9564 a_7383_8138# a_7182_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9565 a_10513_6788# RWL_6 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9566 a_7762_5686# a_7669_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9567 VDD a_16462_826# a_16369_826# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9568 RBL0_9 RWL_21 a_5643_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9569 a_1813_3008# RWL_20 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9570 a_2542_3526# a_2449_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9571 VDD a_11822_7036# a_11729_7036# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9572 WBL_0 WWL_31 a_222_16# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9573 a_2542_7306# a_2449_7306# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9574 a_3903_6518# a_3702_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9575 a_16462_6226# a_16369_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9576 VDD a_7762_2176# a_7669_2176# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9577 a_15209_3526# WWL_18 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9578 WBL_9 WWL_29 a_5442_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9579 RBL0_24 RWL_19 a_14343_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9580 a_11242_4066# a_11149_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9581 RBL0_23 RWL_23 a_13763_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9582 a_3029_7576# WWL_3 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9583 WBL_19 WWL_0 a_11242_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9584 RBL0_3 RWL_4 a_2163_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9585 a_14573_1388# RWL_26 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9586 a_12603_7058# a_12402_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9587 a_7182_2986# a_7089_2986# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9588 GND a_12309_6766# a_12253_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9589 GND a_7182_5146# a_7089_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9590 WBL_3 WWL_26 a_1962_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9591 a_802_2176# a_709_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9592 a_5293_7598# a_4683_7576# RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9593 GND a_3609_2986# a_3553_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9594 a_14343_3818# a_14142_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9595 GND a_6602_4066# a_6509_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9596 WBL_1 WWL_7 a_802_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9597 a_13763_309# a_13562_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9598 WBL_16 WWL_14 a_9502_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9599 GND a_5929_4066# a_5873_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9600 a_16663_4898# a_16462_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9601 a_7963_1118# a_7762_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9602 GND a_222_3796# a_129_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9603 VDD a_12982_1096# a_12889_1096# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9604 a_3702_1366# a_3609_1366# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9605 VDD a_222_7576# a_129_7576# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9606 GND a_8249_1906# a_8193_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9607 WBL_27 WWL_16 a_15882_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9608 RBL0_21 RWL_0 a_12603_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9609 a_1813_5978# RWL_9 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9610 RBL0_15 RWL_16 a_9123_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9611 RBL0_4 RWL_31 a_2743_38# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9612 a_9409_556# WWL_29 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9613 a_12833_6518# RWL_7 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9614 a_7033_1118# RWL_27 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9615 a_4189_1636# WWL_25 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9616 GND a_10082_2986# a_9989_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9617 VDD a_14722_7846# a_14629_7846# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9618 a_12402_1906# a_12309_1906# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9619 WBL_21 WWL_22 a_12402_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9620 VDD a_14142_287# a_14049_287# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9621 a_9353_2198# RWL_23 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9622 a_6509_2716# WWL_21 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9623 a_653_4088# RWL_16 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9624 a_7762_5416# a_7669_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9625 GND a_802_826# a_709_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9626 RBL0_9 RWL_22 a_5643_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9627 a_2542_3256# a_2449_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9628 a_2542_7036# a_2449_7036# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9629 WBL_4 WWL_3 a_2542_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9630 a_18109_4336# WWL_15 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9631 a_17529_3256# WWL_19 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9632 RBL0_28 RWL_20 a_16663_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9633 VDD a_14142_4606# a_14049_4606# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9634 a_10863_39# a_10662_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9635 a_3903_6248# a_3702_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9636 VDD a_7762_1906# a_7669_1906# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9637 a_3029_7306# WWL_4 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9638 WBL_19 WWL_1 a_11242_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9639 GND a_3609_5956# a_3553_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9640 RBL0_3 RWL_5 a_2163_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9641 a_11822_287# a_11729_287# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9642 a_8193_8408# RWL_0 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9643 WBL_12 WWL_19 a_7182_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9644 WBL_3 WWL_27 a_1962_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9645 a_14343_3548# a_14142_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9646 WBL_1 WWL_8 a_802_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9647 a_222_1366# a_129_1366# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9648 a_10082_3796# a_9989_3796# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9649 GND a_10082_5956# a_9989_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9650 GND a_222_3526# a_129_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9651 a_13469_8386# WWL_0 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9652 VDD a_222_7306# a_129_7306# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9653 a_3702_1096# a_3609_1096# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9654 GND a_8249_1636# a_8193_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9655 WBL_6 WWL_25 a_3702_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9656 RBL0_21 RWL_1 a_12603_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9657 VDD a_1382_5956# a_1289_5956# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9658 a_18202_556# a_18109_556# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9659 a_10863_1928# a_10662_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9660 a_14142_7846# a_14049_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9661 a_13413_7328# RWL_4 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9662 a_12833_6248# RWL_8 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9663 a_4189_1366# WWL_26 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9664 a_8829_2446# WWL_22 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9665 VDD a_5442_3796# a_5349_3796# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9666 RBL0_28 RWL_9 a_16663_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9667 WBL_21 WWL_23 a_12402_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9668 RBL0_20 RWL_13 a_12023_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9669 RBL0_5 RWL_27 a_3323_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9670 a_5442_7846# a_5349_7846# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9671 VDD a_14142_17# a_14049_17# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9672 a_7762_5146# a_7669_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9673 GND a_802_556# a_709_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9674 RBL0_9 RWL_23 a_5643_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9675 WBL_4 WWL_4 a_2542_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9676 a_17529_2986# WWL_20 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9677 a_18109_4066# WWL_16 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9678 VDD a_14142_4336# a_14049_4336# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9679 GND a_9502_7846# a_9409_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9680 GND a_1962_8386# a_1869_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9681 GND a_8829_7846# a_8773_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9682 GND a_4189_6766# a_4133_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9683 a_6223_3818# a_6022_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9684 a_5643_2738# a_5442_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9685 a_11822_17# a_11729_17# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9686 VDD a_10662_2716# a_10569_2716# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9687 a_10662_2986# a_10569_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9688 GND a_15209_7306# a_15153_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9689 a_8193_8138# RWL_1 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9690 a_4769_7576# WWL_3 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9691 WBL_12 WWL_20 a_7182_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9692 RBL0_6 RWL_4 a_3903_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9693 a_15302_1906# a_15209_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9694 a_14343_3278# a_14142_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9695 GND a_12402_5686# a_12309_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9696 a_15302_5686# a_15209_5686# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9697 a_14722_4606# a_14629_4606# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9698 a_222_1096# a_129_1096# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9699 WBL_0 WWL_25 a_222_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9700 a_10082_3526# a_9989_3526# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9701 a_11149_7036# WWL_5 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9703 GND a_14722_6766# a_14629_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9704 a_4713_6518# RWL_7 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9705 GND a_11729_5686# a_11673_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9706 GND a_222_3256# a_129_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9707 a_13469_8116# WWL_1 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9708 VDD a_222_7036# a_129_7036# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9709 GND a_8249_1366# a_8193_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9710 WBL_6 WWL_26 a_3702_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9711 a_10863_1658# a_10662_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9712 a_16893_848# RWL_28 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9713 VDD a_3122_2446# a_3029_2446# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9714 a_9409_3256# WWL_19 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9715 a_1583_7868# a_1382_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9716 a_13413_7058# RWL_5 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9717 RBL0_29 RWL_6 a_17243_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9718 a_709_5146# WWL_12 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9719 GND a_9989_1906# a_9933_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9720 a_8829_2176# WWL_23 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9721 a_14142_7576# a_14049_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9722 a_4189_1096# WWL_27 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9723 WBL_21 WWL_24 a_12402_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9724 RBL0_14 RWL_20 a_8543_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9725 VDD a_5442_3526# a_5349_3526# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9726 a_15153_3818# RWL_17 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9727 VDD a_17042_5146# a_16949_5146# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9728 RBL0_25 RWL_28 a_14923_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9729 a_17473_4898# RWL_13 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9730 a_8773_1118# RWL_27 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9731 a_10662_5956# a_10569_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9732 a_16949_556# WWL_29 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9733 GND a_9502_7576# a_9409_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9734 GND a_6509_6496# a_6453_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9735 GND a_1962_8116# a_1869_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9736 a_1233_848# RWL_28 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9737 GND a_8829_7576# a_8773_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9738 a_6223_3548# a_6022_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9739 a_5643_2468# a_5442_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9740 VDD a_15882_4606# a_15789_4606# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9741 a_1382_2716# a_1289_2716# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9742 WBL_18 WWL_5 a_10662_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9743 GND a_15209_7036# a_15153_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9744 GND a_1382_4876# a_1289_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9745 a_4769_7306# WWL_4 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9746 RBL0_6 RWL_5 a_3903_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9747 a_15302_1636# a_15209_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9748 a_15302_5416# a_15209_5416# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9749 GND a_12402_5416# a_12309_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9750 a_3122_5686# a_3029_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9751 WBL_0 WWL_26 a_222_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9752 a_73_3008# RWL_20 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9753 WBL_17 WWL_17 a_10082_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9754 a_14722_4336# a_14629_4336# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9755 RBL0_1 RWL_21 a_1003_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9756 GND a_11729_5416# a_11673_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9757 a_5442_6766# a_5349_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9758 a_4713_6248# RWL_8 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9759 RBL0_14 RWL_9 a_8543_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9760 GND a_8249_17# a_8193_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9761 WBL_6 WWL_27 a_3702_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9762 a_14573_309# RWL_30 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9763 a_16893_578# RWL_29 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9764 a_10863_1388# a_10662_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9765 a_17042_8386# a_16949_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9766 VDD a_3122_2176# a_3029_2176# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9767 a_8829_1906# WWL_24 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9768 a_9409_2986# WWL_20 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9769 a_709_4876# WWL_13 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9770 a_1583_7598# a_1382_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9771 GND a_9989_1636# a_9933_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9772 WBL_9 WWL_2 a_5442_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9773 GND a_17042_1096# a_16949_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9774 a_15153_3548# RWL_18 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9775 RBL0_21 RWL_30 a_12603_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9776 RBL0_25 RWL_29 a_14923_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9777 RBL0_19 RWL_17 a_11443_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9778 VDD a_17042_4876# a_16949_4876# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9779 GND a_16369_1096# a_16313_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9780 RBL0_18 RWL_21 a_10863_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9781 a_15882_7846# a_15789_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9782 VDD a_1962_1636# a_1869_1636# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9783 WBL_8 WWL_14 a_4862_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9784 GND a_7089_7306# a_7033_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9785 GND a_6509_6226# a_6453_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9786 a_11673_1928# RWL_24 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9787 a_1233_578# RWL_29 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9788 VDD a_13562_3256# a_13469_3256# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9789 a_5643_2198# a_5442_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9790 a_6223_3278# a_6022_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9791 VDD a_15882_4336# a_15789_4336# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9792 GND a_4282_5686# a_4189_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9793 GND a_3702_4606# a_3609_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9794 a_73_5978# RWL_9 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9795 a_6602_4606# a_6509_4606# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9796 VDD a_3702_8386# a_3609_8386# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9797 a_2449_5956# WWL_9 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9798 a_17622_5146# a_17529_5146# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9799 a_12982_4066# a_12889_4066# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9800 a_15302_1366# a_15209_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9801 GND a_17622_7306# a_17529_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9802 WBL_26 WWL_10 a_15302_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9803 GND a_12402_5146# a_12309_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9804 a_3122_5416# a_3029_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9805 WBL_0 WWL_27 a_222_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9806 RBL0_10 RWL_14 a_6223_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9807 WBL_25 WWL_14 a_14722_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9808 GND a_16949_7306# a_16893_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9809 RBL0_1 RWL_22 a_1003_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9810 WBL_17 WWL_18 a_10082_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9811 GND a_11729_5146# a_11673_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9812 WBL_28 WWL_28 a_16462_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9813 a_6453_2738# RWL_21 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9814 a_4483_8408# a_4282_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9815 a_17042_8116# a_16949_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9816 a_12889_7036# WWL_5 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9817 VDD a_8342_4066# a_8249_4066# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9818 VDD a_3122_1906# a_3029_1906# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9820 GND a_9989_1366# a_9933_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9821 a_15153_3278# RWL_19 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9822 a_12309_3796# WWL_17 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9823 a_13562_6496# a_13469_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9824 VDD a_4862_2446# a_4769_2446# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9825 a_11729_2716# WWL_21 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9826 RBL0_18 RWL_22 a_10863_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9827 RBL0_19 RWL_18 a_11443_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9828 a_15882_7576# a_15789_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9829 GND a_7089_7036# a_7033_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9830 a_17243_6788# a_17042_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9831 a_16893_3818# RWL_17 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9832 a_11673_1658# RWL_25 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9833 a_8543_3008# a_8342_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9835 VDD a_13562_2986# a_13469_2986# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9836 a_4282_3256# a_4189_3256# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9837 GND a_129_5686# a_73_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9838 GND a_8922_6496# a_8829_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9839 GND a_4282_5416# a_4189_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9840 a_2393_7868# RWL_2 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9841 GND a_3702_4336# a_3609_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9842 a_6602_4336# a_6509_4336# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9843 a_7669_7846# WWL_2 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9844 WBL_2 WWL_21 a_1382_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9845 VDD a_3702_8116# a_3609_8116# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9846 a_3903_848# a_3702_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9847 a_17622_1096# a_17529_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9848 a_18202_5956# a_18109_5956# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9849 WBL_22 WWL_15 a_12982_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9850 a_17622_4876# a_17529_4876# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9851 GND a_17622_7036# a_17529_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9852 a_8342_7306# a_8249_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9853 a_7089_4606# WWL_14 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9854 WBL_26 WWL_11 a_15302_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9855 RBL0_10 RWL_15 a_6223_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9856 GND a_16949_7036# a_16893_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9857 a_3122_5146# a_3029_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9858 RBL0_1 RWL_23 a_1003_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9859 a_17042_1636# a_16949_1636# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9860 WBL_24 WWL_30 a_14142_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9861 GND a_14049_2716# a_13993_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9862 a_6453_2468# RWL_22 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9863 a_4483_8138# a_4282_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9864 a_4862_5686# a_4769_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9865 VDD a_4282_826# a_4189_826# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9866 RBL0_4 RWL_21 a_2743_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9867 a_17473_39# RWL_31 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9868 a_8543_5978# a_8342_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9869 a_12309_3526# WWL_18 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9870 a_16949_4606# WWL_14 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9871 a_13562_6226# a_13469_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9872 VDD a_4862_2176# a_4769_2176# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9873 RBL0_18 RWL_23 a_10863_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9874 RBL0_19 RWL_19 a_11443_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9875 a_16893_3548# RWL_18 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9876 a_11673_1388# RWL_26 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9877 a_9502_5146# a_9409_5146# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9878 a_4282_2986# a_4189_2986# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9879 GND a_129_5416# a_73_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9880 GND a_8922_6226# a_8829_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9881 GND a_4282_5146# a_4189_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9882 a_18109_287# WWL_30 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9883 a_2393_7598# RWL_3 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9884 a_11443_3818# a_11242_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9885 GND a_3702_4066# a_3609_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9886 WBL_11 WWL_14 a_6602_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9887 a_3903_578# a_3702_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9888 a_13763_4898# a_13562_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9889 a_8829_826# WWL_28 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9890 GND a_6022_1906# a_5929_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9891 VDD a_6022_5686# a_5929_5686# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9892 WBL_30 WWL_12 a_17622_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9893 GND a_5349_1906# a_5293_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9894 WBL_22 WWL_16 a_12982_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9895 a_8342_7036# a_8249_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9896 RBL0_10 RWL_16 a_6223_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9897 a_1003_1928# a_802_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9898 a_4133_1118# RWL_27 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9899 GND a_1962_286# a_1869_286# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9900 WBL_24 WWL_31 a_14142_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9901 a_1289_1636# WWL_25 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9902 VDD a_11822_7846# a_11729_7846# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9903 GND a_14049_2446# a_13993_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9904 a_6453_2198# RWL_23 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9905 a_3609_2716# WWL_21 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9906 a_4862_5416# a_4769_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9907 RBL0_4 RWL_22 a_2743_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9909 VDD a_16462_6766# a_16369_6766# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9910 a_15209_4336# WWL_15 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9911 a_14629_3256# WWL_19 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9912 VDD a_11242_4606# a_11149_4606# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9913 RBL0_23 RWL_20 a_13763_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9914 a_9123_6788# a_8922_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9915 VDD a_4862_1906# a_4769_1906# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9916 a_4713_39# RWL_31 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9917 RBL0_31 RWL_24 a_18403_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9918 WBL_15 WWL_29 a_8922_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9919 a_16893_3278# RWL_19 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9920 a_18202_4876# a_18109_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9921 a_9502_1096# a_9409_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9922 a_802_2986# a_709_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9923 WBL_21 WWL_29 a_12402_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9924 a_5293_8408# RWL_0 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9925 a_9502_4876# a_9409_4876# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9926 GND a_129_5146# a_73_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9927 WBL_7 WWL_19 a_4282_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9928 a_16663_5708# a_16462_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9929 a_17622_826# a_17529_826# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9930 a_18109_17# WWL_31 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9931 a_11443_3548# a_11242_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9932 GND a_6022_1636# a_5929_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9933 WBL_31 WWL_9 a_18202_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9934 VDD a_6022_5416# a_5929_5416# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9935 a_17243_309# a_17042_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9936 WBL_30 WWL_13 a_17622_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9937 a_10569_8386# WWL_0 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9938 GND a_5349_1636# a_5293_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9939 a_1003_1658# a_802_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9940 a_18053_6788# RWL_6 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9941 a_15153_39# RWL_31 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9942 a_129_2716# WWL_21 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9943 a_9353_3008# RWL_20 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9944 a_11242_7846# a_11149_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9945 a_10513_7328# RWL_4 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9946 RBL0_23 RWL_9 a_13763_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9947 a_1289_1366# WWL_26 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9948 a_5929_2446# WWL_22 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9949 VDD a_2542_3796# a_2449_3796# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9950 GND a_14049_2176# a_13993_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9951 a_2542_7846# a_2449_7846# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9952 a_4862_5146# a_4769_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9953 RBL0_4 RWL_23 a_2743_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9954 GND a_16462_2716# a_16369_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9955 VDD a_16462_6496# a_16369_6496# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9956 GND a_15789_2716# a_15733_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9957 a_14629_2986# WWL_20 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9958 a_15209_4066# WWL_16 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9959 a_7182_6766# a_7089_6766# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9960 VDD a_11242_4336# a_11149_4336# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9961 a_1962_4606# a_1869_4606# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9962 a_802_5956# a_709_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9963 GND a_6602_7846# a_6509_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9964 GND a_5929_7846# a_5873_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9965 VDD a_11822_826# a_11729_826# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9966 GND a_1289_6766# a_1233_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9967 RBL0_31 RWL_25 a_18403_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9968 a_3323_3818# a_3122_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9969 a_2743_2738# a_2542_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9970 GND a_12309_7306# a_12253_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9971 a_5293_8138# RWL_1 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9972 RBL0_15 RWL_2 a_9123_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9973 a_1869_7576# WWL_3 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9974 WBL_1 WWL_5 a_802_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9975 WBL_16 WWL_12 a_9502_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9976 WBL_7 WWL_20 a_4282_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9977 a_16663_5438# a_16462_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9978 a_12402_1906# a_12309_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9979 a_11443_3278# a_11242_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9980 a_12402_5686# a_12309_5686# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9981 a_11822_4606# a_11729_4606# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9982 a_653_7868# RWL_2 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9983 a_9353_5978# RWL_9 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9984 GND a_6022_1366# a_5929_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9985 GND a_11822_6766# a_11729_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9986 a_1813_6518# RWL_7 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9987 a_10569_8116# WWL_1 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9988 GND a_5349_1366# a_5293_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9989 a_4713_848# RWL_28 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9990 a_1003_1388# a_802_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9991 RBL0_20 RWL_10 a_12023_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9992 GND a_7762_1906# a_7669_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9993 VDD a_7762_5686# a_7669_5686# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9994 a_6509_3256# WWL_19 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9995 a_11242_7576# a_11149_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9996 a_10513_7058# RWL_5 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9997 RBL0_24 RWL_6 a_14343_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9998 a_5929_2176# WWL_23 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9999 a_1289_1096# WWL_27 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10000 RBL0_9 RWL_20 a_5643_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10001 VDD a_2542_3526# a_2449_3526# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10002 a_12253_3818# RWL_17 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10003 VDD a_14142_5146# a_14049_5146# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10004 RBL0_4 RWL_28 a_2743_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10005 GND a_16462_2446# a_16369_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10006 a_14573_4898# RWL_13 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10007 a_5873_1118# RWL_27 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10008 a_7182_2716# a_7089_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10009 VDD a_16462_6226# a_16369_6226# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10010 a_7182_6496# a_7089_6496# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10011 a_4769_556# WWL_29 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10012 GND a_15789_2446# a_15733_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10013 a_3029_7846# WWL_2 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10014 a_1962_4336# a_1869_4336# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10015 GND a_6602_7576# a_6509_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10016 GND a_3609_6496# a_3553_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10017 GND a_5929_7576# a_5873_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10018 a_3323_3548# a_3122_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10019 a_7963_4628# a_7762_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10020 RBL0_31 RWL_26 a_18403_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10021 a_2743_2468# a_2542_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10022 VDD a_12982_4606# a_12889_4606# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10023 WBL_27 WWL_3 a_15882_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10024 GND a_12309_7036# a_12253_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10025 RBL0_15 a_4683_7576# a_9123_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10026 WBL_16 WWL_13 a_9502_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10027 a_1869_7306# WWL_4 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10028 a_16663_5168# a_16462_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10029 a_12402_1636# a_12309_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10030 GND a_10082_6496# a_9989_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10031 a_7033_4628# RWL_14 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10032 a_12402_5416# a_12309_5416# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10033 VDD a_222_7846# a_129_7846# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10034 a_11822_4336# a_11729_4336# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10035 a_653_7598# RWL_3 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10036 a_2542_6766# a_2449_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10037 a_1813_6248# RWL_8 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10038 RBL0_9 RWL_9 a_5643_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10039 a_17529_6766# WWL_6 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10040 a_4713_578# RWL_29 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10041 a_14142_8386# a_14049_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10042 RBL0_28 RWL_7 a_16663_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10043 RBL0_20 RWL_11 a_12023_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10044 GND a_7762_1636# a_7669_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10045 VDD a_7762_5416# a_7669_5416# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10046 a_5929_1906# WWL_24 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10047 a_6509_2986# WWL_20 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10048 a_17473_5708# RWL_10 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10049 WBL_4 WWL_2 a_2542_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10050 GND a_14142_1096# a_14049_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10051 a_12253_3548# RWL_18 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10052 a_13562_556# a_13469_556# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10053 RBL0_4 RWL_29 a_2743_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10054 VDD a_14142_4876# a_14049_4876# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10055 GND a_13469_1096# a_13413_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10056 GND a_16462_2176# a_16369_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10057 a_7182_2446# a_7089_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10058 GND a_9502_8386# a_9409_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10059 a_3122_826# a_3029_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10060 GND a_15789_2176# a_15733_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10061 WBL_12 WWL_6 a_7182_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10062 a_7182_6226# a_7089_6226# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10063 GND a_8829_8386# a_8773_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10064 RBL0_31 RWL_28 a_18403_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10065 WBL_3 WWL_14 a_1962_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10066 GND a_4189_7306# a_4133_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10067 GND a_3609_6226# a_3553_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10068 VDD a_18202_2716# a_18109_2716# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10069 GND a_12982_17# a_12889_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10070 VDD a_10662_3256# a_10569_3256# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10071 a_3323_3278# a_3122_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10072 a_7963_4358# a_7762_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10073 a_2743_2198# a_2542_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10074 VDD a_12982_4336# a_12889_4336# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10075 GND a_1382_5686# a_1289_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10076 GND a_9502_826# a_9409_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10077 WBL_27 WWL_4 a_15882_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10078 a_3702_4606# a_3609_4606# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10079 GND a_12982_826# a_12889_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10080 a_14722_5146# a_14629_5146# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10081 a_10082_4066# a_9989_4066# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10082 a_12402_1366# a_12309_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10083 GND a_14722_7306# a_14629_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10084 GND a_10082_6226# a_9989_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10085 a_7033_4358# RWL_15 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10086 WBL_21 WWL_10 a_12402_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10087 a_16462_287# a_16369_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10088 RBL0_5 RWL_14 a_3323_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10089 WBL_7 WWL_28 a_4282_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10090 a_18109_7576# WWL_3 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10091 a_17529_6496# WWL_7 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10092 a_3553_2738# RWL_21 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10093 a_1583_8408# a_1382_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10094 RBL0_29 RWL_4 a_17243_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10095 a_14142_8116# a_14049_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10096 RBL0_28 RWL_8 a_16663_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10097 RBL0_20 RWL_12 a_12023_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10098 VDD a_5442_4066# a_5349_4066# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10099 GND a_7762_1366# a_7669_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10100 a_18053_309# RWL_30 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10101 a_17473_5438# RWL_11 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10102 a_12253_3278# RWL_19 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10103 VDD a_802_3796# a_709_3796# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10104 a_10662_6496# a_10569_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10105 VDD a_1962_2446# a_1869_2446# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10106 GND a_9502_8116# a_9409_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10107 a_3122_556# a_3029_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10108 a_7182_2176# a_7089_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10109 a_222_826# a_129_826# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10110 RBL0_27 RWL_30 a_16083_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10111 WBL_12 WWL_7 a_7182_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10112 GND a_8829_8116# a_8773_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10113 RBL0_31 RWL_29 a_18403_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10114 GND a_4189_7036# a_4133_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10115 a_14343_6788# a_14142_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10116 a_13993_3818# RWL_17 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10117 VDD a_15882_5146# a_15789_5146# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10118 a_5643_3008# a_5442_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10119 a_8922_2716# a_8829_2716# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10120 VDD a_10662_2986# a_10569_2986# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10121 a_222_4606# a_129_4606# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10122 a_1382_3256# a_1289_3256# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10123 a_7963_4088# a_7762_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10124 GND a_222_6766# a_129_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10125 GND a_1382_5416# a_1289_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10126 GND a_9502_556# a_9409_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10127 GND a_10662_287# a_10569_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10128 a_3702_4336# a_3609_4336# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10129 a_4769_7846# WWL_2 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10130 GND a_12982_556# a_12889_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10131 GND a_8249_4876# a_8193_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10132 GND a_6509_826# a_6453_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10133 a_14722_1096# a_14629_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10134 a_15302_5956# a_15209_5956# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10135 WBL_17 WWL_15 a_10082_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10136 a_14722_4876# a_14629_4876# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10137 GND a_14722_7036# a_14629_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10138 a_9409_6766# WWL_6 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10139 a_8829_5686# WWL_10 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10140 a_7033_4088# RWL_16 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10141 a_5442_7306# a_5349_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10142 RBL0_14 RWL_7 a_8543_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10143 a_4189_4606# WWL_14 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10144 WBL_21 WWL_11 a_12402_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10145 RBL0_5 RWL_15 a_3323_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10146 GND a_222_286# a_129_286# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10147 a_14142_1636# a_14049_1636# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10148 GND a_11149_2716# a_11093_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10149 a_8773_4628# RWL_14 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10150 a_18109_7306# WWL_4 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10151 a_3553_2468# RWL_22 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10152 RBL0_29 RWL_5 a_17243_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10153 a_17529_6226# WWL_8 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10154 a_1583_8138# a_1382_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10155 RBL0_14 RWL_31 a_8543_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10156 a_5643_5978# a_5442_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10157 VDD a_9502_1636# a_9409_1636# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10158 a_17473_5168# RWL_12 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10159 a_15882_8386# a_15789_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10160 VDD a_802_3526# a_709_3526# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10161 a_10662_6226# a_10569_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10162 GND a_10662_17# a_10569_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10163 VDD a_1962_2176# a_1869_2176# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10164 WBL_8 WWL_12 a_4862_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10165 WBL_12 WWL_8 a_7182_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10166 GND a_15882_1096# a_15789_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10167 a_13993_3548# RWL_18 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10168 VDD a_15882_4876# a_15789_4876# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10169 a_73_6518# RWL_7 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10170 a_6602_5146# a_6509_5146# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10171 a_222_4336# a_129_4336# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10172 a_1382_2986# a_1289_2986# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10173 GND a_1382_5146# a_1289_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10174 WBL_6 WWL_14 a_3702_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10175 GND a_6509_556# a_6453_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10177 a_10863_4898# a_10662_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10178 GND a_3122_1906# a_3029_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10179 VDD a_3122_5686# a_3029_5686# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10180 WBL_25 WWL_12 a_14722_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10181 a_7383_848# a_7182_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10182 GND a_2449_1906# a_2393_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10183 RBL0_1 RWL_20 a_1003_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10184 WBL_17 WWL_16 a_10082_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10185 a_709_8386# WWL_0 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10186 a_9409_6496# WWL_7 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10187 a_8829_5416# WWL_11 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10188 RBL0_14 RWL_8 a_8543_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10189 a_5442_7036# a_5349_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10190 a_17042_2446# a_16949_2446# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10191 RBL0_5 RWL_16 a_3323_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10192 GND a_17042_4606# a_16949_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10193 VDD a_17042_8386# a_16949_8386# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10194 a_1233_1118# RWL_27 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10195 GND a_16369_4606# a_16313_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10196 GND a_11149_2446# a_11093_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10197 a_8773_4358# RWL_15 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10198 a_3553_2198# RWL_23 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10199 VDD a_13562_6766# a_13469_6766# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10200 a_12309_4336# WWL_15 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10201 a_11729_3256# WWL_19 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10202 a_9989_287# WWL_30 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10203 RBL0_18 RWL_20 a_10863_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10204 a_6223_6788# a_6022_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10205 a_15882_8116# a_15789_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10206 VDD a_1962_1906# a_1869_1906# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10207 WBL_8 WWL_13 a_4862_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10208 a_17243_7328# a_17042_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10209 RBL0_26 RWL_24 a_15503_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10210 a_12982_3796# a_12889_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10211 a_12982_7576# a_12889_7576# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10212 a_13993_3278# RWL_19 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10213 a_15302_4876# a_15209_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10214 a_6602_1096# a_6509_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10215 a_2393_8408# RWL_0 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10216 WBL_15 WWL_21 a_8922_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10217 WBL_0 WWL_14 a_222_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10218 a_6602_4876# a_6509_4876# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10219 a_73_6248# RWL_8 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10220 RBL0_1 RWL_9 a_1003_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10221 WBL_2 WWL_19 a_1382_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10222 a_5442_826# a_5349_826# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10223 a_13763_5708# a_13562_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10224 VDD a_17622_1366# a_17529_1366# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10225 GND a_8342_3796# a_8249_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10226 GND a_3122_1636# a_3029_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10227 VDD a_8342_7576# a_8249_7576# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10228 a_7089_5146# WWL_12 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10229 WBL_26 WWL_9 a_15302_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10230 VDD a_3122_5416# a_3029_5416# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10231 a_5063_309# a_4862_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10232 GND a_7669_3796# a_7613_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10233 WBL_25 WWL_13 a_14722_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10234 a_7383_578# a_7182_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10235 GND a_2449_1636# a_2393_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10236 a_9409_6226# WWL_8 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10237 a_709_8116# WWL_1 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10238 GND a_9989_4876# a_9933_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10239 a_17042_2176# a_16949_2176# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10240 a_15789_826# WWL_28 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10241 GND a_17042_4336# a_16949_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10242 a_15153_6788# RWL_6 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10243 a_6453_3008# RWL_20 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10244 VDD a_17042_8116# a_16949_8116# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10245 RBL0_10 RWL_31 a_6223_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10246 RBL0_18 RWL_9 a_10863_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10247 GND a_16369_4336# a_16313_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10248 GND a_11149_2176# a_11093_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10249 a_8773_4088# RWL_16 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10250 GND a_13562_2716# a_13469_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10251 a_8543_6518# a_8342_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10252 a_15882_1636# a_15789_1636# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10253 VDD a_13562_6496# a_13469_6496# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10254 a_16949_5146# WWL_12 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10255 a_12309_4066# WWL_16 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10256 GND a_12889_2716# a_12833_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10257 a_11729_2986# WWL_20 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10258 a_4282_6766# a_4189_6766# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10259 a_9989_17# WWL_31 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10260 GND a_3702_7846# a_3609_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10261 a_18202_5686# a_18109_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10262 a_17243_7058# a_17042_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10263 RBL0_26 RWL_25 a_15503_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10264 a_12982_3526# a_12889_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10265 a_17622_4606# a_17529_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10266 a_17622_8386# a_17529_8386# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10267 a_12982_7306# a_12889_7306# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10268 a_2393_8138# RWL_1 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10269 RBL0_10 RWL_2 a_6223_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10270 WBL_11 WWL_12 a_6602_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10271 WBL_2 WWL_20 a_1382_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10272 a_13763_5438# a_13562_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10273 VDD a_17622_1096# a_17529_1096# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10274 WBL_27 WWL_29 a_15882_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10275 a_8342_1366# a_8249_1366# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10276 GND a_8342_3526# a_8249_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10277 a_6453_5978# RWL_9 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10278 GND a_3122_1366# a_3029_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10279 VDD a_8342_7306# a_8249_7306# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10280 a_7089_4876# WWL_13 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10281 GND a_7669_3526# a_7613_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10282 VDD a_9502_287# a_9409_287# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10283 GND a_2449_1366# a_2393_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10284 VDD a_12982_287# a_12889_287# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10285 a_13469_287# WWL_30 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10286 a_17042_1906# a_16949_1906# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10287 WBL_29 WWL_22 a_17042_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10288 GND a_4862_1906# a_4769_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10289 GND a_14049_2986# a_13993_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10290 GND a_17042_4066# a_16949_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10291 VDD a_4862_5686# a_4769_5686# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10292 a_3609_3256# WWL_19 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10293 RBL0_19 RWL_6 a_11443_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10294 GND a_16369_4066# a_16313_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10295 a_18403_1118# a_18202_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10296 RBL0_4 RWL_20 a_2743_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10297 VDD a_11242_5146# a_11149_5146# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10298 GND a_13562_2446# a_13469_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10299 a_9123_7328# a_8922_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10300 a_8543_6248# a_8342_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10301 a_11673_4898# RWL_13 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10302 a_2973_1118# RWL_27 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10303 GND a_2449_286# a_2393_308# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10304 a_4282_2716# a_4189_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10305 a_16949_4876# WWL_13 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10306 VDD a_13562_6226# a_13469_6226# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10307 a_7762_17# a_7669_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10308 a_4282_6496# a_4189_6496# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10309 GND a_12889_2446# a_12833_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10310 GND a_3702_7576# a_3609_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10311 a_18202_5416# a_18109_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10312 a_12982_3256# a_12889_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10313 a_17622_4336# a_17529_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10314 RBL0_26 RWL_26 a_15503_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10315 a_17622_8116# a_17529_8116# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10316 WBL_22 WWL_3 a_12982_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10317 a_12982_7036# a_12889_7036# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10318 VDD a_15302_826# a_15209_826# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10319 RBL0_10 a_4683_7576# a_6223_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10320 WBL_11 WWL_13 a_6602_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10321 a_13763_5168# a_13562_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10322 a_8342_1096# a_8249_1096# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10323 WBL_14 WWL_25 a_8342_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10324 a_4133_4628# RWL_14 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10325 VDD a_6022_5956# a_5929_5956# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10326 GND a_14049_5956# a_13993_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10327 a_6602_826# a_6509_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10328 GND a_8342_3256# a_8249_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10329 VDD a_8342_7036# a_8249_7036# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10330 RBL0_4 RWL_9 a_2743_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10331 GND a_7669_3256# a_7613_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10332 VDD a_9502_17# a_9409_17# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10333 a_18053_7328# RWL_4 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10334 VDD a_12982_17# a_12889_17# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10335 a_14629_6766# WWL_6 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10336 a_129_3256# WWL_19 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10337 a_11242_8386# a_11149_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10338 RBL0_23 RWL_7 a_13763_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10339 RBL0_13 RWL_27 a_7963_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10340 a_13469_17# WWL_31 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10341 GND a_709_1906# a_653_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10342 WBL_29 WWL_23 a_17042_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10343 GND a_4862_1636# a_4769_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10344 VDD a_4862_5416# a_4769_5416# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10345 a_3609_2986# WWL_20 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10346 a_8193_848# RWL_28 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10347 a_14573_5708# RWL_10 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10348 GND a_11242_1096# a_11149_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10349 a_1382_556# a_1289_556# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10350 a_16893_6788# RWL_6 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10351 VDD a_11242_4876# a_11149_4876# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10352 a_9123_7058# a_8922_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10353 a_1962_5146# a_1869_5146# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10354 GND a_10569_1096# a_10513_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10355 GND a_13562_2176# a_13469_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10356 a_9502_4606# a_9409_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10357 a_802_6496# a_709_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10358 a_4282_2446# a_4189_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10359 a_9502_8386# a_9409_8386# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10360 GND a_6602_8386# a_6509_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10361 a_4282_6226# a_4189_6226# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10362 GND a_12889_2176# a_12833_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10363 WBL_7 WWL_6 a_4282_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10364 RBL0_10 RWL_28 a_6223_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10365 GND a_5929_8386# a_5873_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10366 GND a_1289_7306# a_1233_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10367 a_3323_308# a_3122_286# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10368 VDD a_15302_2716# a_15209_2716# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10369 VDD a_7762_556# a_7669_556# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10370 a_8249_556# WWL_29 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10371 a_18202_5146# a_18109_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10372 a_17622_4066# a_17529_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10373 RBL0_15 RWL_0 a_9123_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10374 WBL_30 WWL_0 a_17622_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10375 WBL_22 WWL_4 a_12982_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10376 a_11822_5146# a_11729_5146# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10377 a_653_8408# RWL_0 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10378 GND a_11822_7306# a_11729_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10379 a_9353_6518# RWL_7 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10380 WBL_14 WWL_26 a_8342_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10381 a_4133_4358# RWL_15 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10382 a_16083_2738# a_15882_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10383 a_6602_556# a_6509_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10384 a_18053_7058# RWL_5 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10385 a_15209_7576# WWL_3 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10386 a_14629_6496# WWL_7 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10387 a_11242_8116# a_11149_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10388 RBL0_24 RWL_4 a_14343_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10389 GND a_709_1636# a_653_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10390 WBL_29 WWL_24 a_17042_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10391 a_129_2986# WWL_20 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10392 VDD a_2542_4066# a_2449_4066# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10393 RBL0_23 RWL_8 a_13763_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10394 GND a_4862_1366# a_4769_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10395 a_5442_17# a_5349_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10396 a_8193_578# RWL_29 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10397 GND a_9989_826# a_9933_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10398 GND a_16462_2986# a_16369_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10399 a_14573_5438# RWL_11 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10400 a_1382_286# a_1289_286# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10401 a_1962_1096# a_1869_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10402 GND a_15789_2986# a_15733_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10403 a_9502_4336# a_9409_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10404 a_1962_4876# a_1869_4876# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10405 a_802_6226# a_709_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10406 a_4282_2176# a_4189_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10407 GND a_6602_8116# a_6509_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10408 a_9502_8116# a_9409_8116# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10409 a_17042_556# a_16949_556# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10410 GND a_12889_17# a_12833_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10411 WBL_7 WWL_7 a_4282_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10412 RBL0_10 RWL_29 a_6223_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10413 GND a_5929_8116# a_5873_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10414 GND a_1289_7036# a_1233_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10415 a_11443_6788# a_11242_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10416 VDD a_12982_5146# a_12889_5146# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10417 a_2743_3008# a_2542_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10418 a_6022_2716# a_5929_2716# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10419 a_10082_826# a_9989_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10420 a_6803_39# a_6602_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10421 GND a_3029_3796# a_2973_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10422 GND a_6022_4876# a_5929_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10423 WBL_30 WWL_1 a_17622_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10424 RBL0_15 RWL_1 a_9123_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10425 GND a_5349_4876# a_5293_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10426 a_1869_7846# WWL_2 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10427 a_7383_1928# a_7182_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10428 a_11822_1096# a_11729_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10429 a_12402_5956# a_12309_5956# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10430 a_9933_309# RWL_30 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10431 a_1003_4898# a_802_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10432 a_11822_4876# a_11729_4876# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10433 GND a_16462_826# a_16369_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10434 a_9353_6248# RWL_8 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10435 a_653_8138# RWL_1 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10436 GND a_11822_7036# a_11729_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10437 a_6509_6766# WWL_6 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10438 a_5929_5686# WWL_10 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10439 a_4133_4088# RWL_16 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10440 a_2542_7306# a_2449_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10441 RBL0_9 RWL_7 a_5643_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10442 WBL_14 WWL_27 a_8342_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10443 a_1289_4606# WWL_14 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10444 a_16083_2468# a_15882_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10445 a_16462_3796# a_16369_3796# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10446 a_11242_1636# a_11149_1636# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10447 GND a_16462_5956# a_16369_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10448 a_5873_4628# RWL_14 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10449 a_15209_7306# WWL_4 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10450 RBL0_24 RWL_5 a_14343_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10451 a_14629_6226# WWL_8 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10452 VDD a_7762_5956# a_7669_5956# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10453 GND a_15789_5956# a_15733_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10454 GND a_709_1366# a_653_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10455 a_17243_39# a_17042_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10456 VDD a_11242_556# a_11149_556# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10457 GND a_7669_287# a_7613_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10458 RBL0_27 RWL_17 a_16083_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10459 GND a_9989_556# a_9933_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10460 a_2743_5978# a_2542_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10461 a_14573_5168# RWL_12 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10462 RBL0_16 RWL_27 a_9703_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10463 a_1382_16# a_1289_16# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10464 VDD a_6602_1636# a_6509_1636# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10465 VDD a_7182_2716# a_7089_2716# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10466 a_7182_2986# a_7089_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10467 RBL0_31 RWL_13 a_18403_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10469 WBL_3 WWL_12 a_1962_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10470 a_9502_4066# a_9409_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10471 VDD a_18202_3256# a_18109_3256# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10472 WBL_16 WWL_0 a_9502_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10473 WBL_7 WWL_8 a_4282_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10474 GND a_12982_1096# a_12889_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10475 a_15733_848# RWL_28 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10476 VDD a_12982_4876# a_12889_4876# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10477 WBL_27 WWL_2 a_15882_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10478 GND a_8249_5686# a_8193_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10479 a_3702_5146# a_3609_5146# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10480 a_10082_556# a_9989_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10481 GND a_3029_3526# a_2973_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10482 a_7383_1658# a_7182_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10483 GND a_8922_17# a_8829_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10484 RBL0_23 RWL_28 a_13763_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10485 GND a_14142_287# a_14049_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10486 GND a_16462_556# a_16369_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10487 a_6509_6496# WWL_7 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10488 a_5929_5416# WWL_11 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10489 RBL0_9 RWL_8 a_5643_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10490 GND a_13469_826# a_13413_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10491 a_14142_2446# a_14049_2446# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10492 a_2542_7036# a_2449_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10493 a_16083_2198# a_15882_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10494 GND a_14142_4606# a_14049_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10495 a_17529_7036# WWL_5 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10496 a_16462_3526# a_16369_3526# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10497 VDD a_14142_8386# a_14049_8386# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10498 GND a_13469_4606# a_13413_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10499 a_7182_5956# a_7089_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10500 a_5873_4358# RWL_15 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10501 a_17823_2738# a_17622_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10502 a_11822_287# a_11729_287# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10503 VDD a_9502_2446# a_9409_2446# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10504 VDD a_10662_6766# a_10569_6766# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10505 GND a_10569_17# a_10513_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10506 RBL0_27 RWL_18 a_16083_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10507 a_7963_7868# a_7762_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10508 a_3323_6788# a_3122_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10509 WBL_12 WWL_5 a_7182_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10510 WBL_3 WWL_13 a_1962_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10511 a_14343_7328# a_14142_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10512 WBL_16 WWL_1 a_9502_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10513 RBL0_21 RWL_24 a_12603_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10514 VDD a_18202_2986# a_18109_2986# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10515 a_10082_3796# a_9989_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10516 a_8922_3256# a_8829_3256# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10517 a_10082_7576# a_9989_7576# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10518 a_222_5146# a_129_5146# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10519 RBL0_18 RWL_31 a_10863_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10520 a_15733_578# RWL_29 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10521 a_12402_4876# a_12309_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10522 a_7033_7868# RWL_2 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10523 GND a_222_7306# a_129_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10524 a_3702_1096# a_3609_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10525 GND a_8249_5416# a_8193_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10526 WBL_10 WWL_21 a_6022_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10527 a_3702_4876# a_3609_4876# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10528 a_10863_5708# a_10662_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10529 GND a_3029_3256# a_2973_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10530 VDD a_14722_1366# a_14629_1366# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10531 a_7383_1388# a_7182_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10532 RBL0_23 RWL_29 a_13763_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10533 GND a_5442_3796# a_5349_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10534 a_7762_2716# a_7669_2716# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10535 VDD a_5442_7576# a_5349_7576# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10536 a_4189_5146# WWL_12 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10537 WBL_21 WWL_9 a_12402_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10538 GND a_4769_3796# a_4713_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10539 GND a_7762_4876# a_7669_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10540 a_6509_6226# WWL_8 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10542 GND a_11149_287# a_11093_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10543 GND a_13469_556# a_13413_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10544 a_14142_2176# a_14049_2176# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10545 a_3609_826# WWL_28 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10546 GND a_14142_4336# a_14049_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10547 a_18109_7846# WWL_2 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10548 a_12253_6788# RWL_6 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10549 a_3553_3008# RWL_20 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10550 WBL_28 WWL_17 a_16462_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10551 VDD a_14142_8116# a_14049_8116# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10552 RBL0_12 RWL_21 a_7383_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10553 GND a_13469_4336# a_13413_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10554 a_5873_4088# RWL_16 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10555 a_6602_287# a_6509_287# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10556 a_17823_2468# a_17622_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10557 a_8193_1928# RWL_24 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10558 GND a_10662_2716# a_10569_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10559 a_5643_6518# a_5442_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10560 VDD a_9502_2176# a_9409_2176# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10561 VDD a_10662_6496# a_10569_6496# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10562 RBL0_27 RWL_19 a_16083_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10563 VDD a_802_4066# a_709_4066# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10564 a_7963_7598# a_7762_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10565 a_1382_6766# a_1289_6766# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10566 a_15302_5686# a_15209_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10567 RBL0_30 RWL_17 a_17823_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10568 a_14722_4606# a_14629_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10569 a_14343_7058# a_14142_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10570 a_222_1096# a_129_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10571 RBL0_21 RWL_25 a_12603_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10572 a_10082_3526# a_9989_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10573 a_8922_2986# a_8829_2986# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10574 a_14722_8386# a_14629_8386# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10575 a_10082_7306# a_9989_7306# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10576 a_222_4876# a_129_4876# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10577 GND a_6602_17# a_6509_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10578 a_7033_7598# a_4683_7576# RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10579 GND a_222_7036# a_129_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10580 RBL0_5 RWL_2 a_3323_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10581 WBL_6 WWL_12 a_3702_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10582 GND a_8249_5146# a_8193_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10583 a_10863_5438# a_10662_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10584 VDD a_14722_1096# a_14629_1096# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10585 a_5442_1366# a_5349_1366# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10586 GND a_5442_3526# a_5349_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10587 a_9409_7036# WWL_5 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10588 a_8829_5956# WWL_9 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10589 a_3553_5978# RWL_9 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10590 a_8922_826# a_8829_826# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10591 VDD a_5442_7306# a_5349_7306# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10592 GND a_9989_5686# a_9933_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10593 a_4189_4876# WWL_13 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10594 a_12402_826# a_12309_826# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10595 GND a_4769_3526# a_4713_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10596 a_14142_1906# a_14049_1906# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10597 WBL_24 WWL_22 a_14142_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10598 GND a_1962_1906# a_1869_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10599 GND a_11149_2986# a_11093_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10600 GND a_14142_4066# a_14049_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10601 a_8249_2716# WWL_21 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10602 WBL_28 WWL_18 a_16462_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10603 VDD a_1962_5686# a_1869_5686# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10604 RBL0_12 RWL_22 a_7383_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10605 GND a_13469_4066# a_13413_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10606 a_15503_1118# a_15302_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10607 a_15882_2446# a_15789_2446# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10608 a_2743_848# a_2542_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10609 a_6602_17# a_6509_17# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10610 a_17823_2198# a_17622_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10611 GND a_15882_4606# a_15789_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10612 a_8193_1658# RWL_25 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10613 GND a_10662_2446# a_10569_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10614 VDD a_15882_8386# a_15789_8386# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10615 a_6223_7328# a_6022_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10616 a_5643_6248# a_5442_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10617 VDD a_9502_1906# a_9409_1906# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10618 a_1382_2716# a_1289_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10619 VDD a_10662_6226# a_10569_6226# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10620 a_1382_6496# a_1289_6496# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10621 WBL_13 WWL_29 a_7762_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10622 a_15302_5416# a_15209_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10623 RBL0_30 RWL_18 a_17823_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10624 RBL0_21 RWL_26 a_12603_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10625 a_10082_3256# a_9989_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10626 a_14722_4336# a_14629_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10627 a_14722_8116# a_14629_8116# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10628 WBL_0 WWL_12 a_222_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10629 WBL_15 WWL_19 a_8922_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10630 WBL_17 WWL_3 a_10082_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10631 a_10082_7036# a_9989_7036# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10632 RBL0_1 RWL_7 a_1003_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10633 VDD a_3122_826# a_3029_826# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10634 RBL0_5 RWL_3 a_3323_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10635 WBL_6 WWL_13 a_3702_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10636 a_10863_5168# a_10662_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10637 a_5442_1096# a_5349_1096# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10638 WBL_9 WWL_25 a_5442_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10639 a_1233_4628# RWL_14 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10640 VDD a_3122_5956# a_3029_5956# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10641 GND a_11149_5956# a_11093_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10642 a_8773_7868# RWL_2 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10643 GND a_5442_3256# a_5349_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10644 WBL_13 WWL_21 a_7762_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10645 VDD a_5442_7036# a_5349_7036# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10646 GND a_9989_5416# a_9933_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10647 a_10082_287# a_9989_287# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10648 GND a_4769_3256# a_4713_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10649 a_15153_7328# RWL_4 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10650 a_11729_6766# WWL_6 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10651 WBL_24 WWL_23 a_14142_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10652 RBL0_18 RWL_7 a_10863_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10653 RBL0_8 RWL_27 a_5063_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10654 GND a_1962_1636# a_1869_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10655 VDD a_1962_5416# a_1869_5416# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10656 RBL0_12 RWL_23 a_7383_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10657 VDD a_16462_287# a_16369_287# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10658 WBL_8 WWL_0 a_4862_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10659 a_11673_5708# RWL_10 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10660 a_15882_2176# a_15789_2176# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10661 a_2743_578# a_2542_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10662 GND a_15882_4336# a_15789_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10663 a_13993_6788# RWL_6 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10664 a_8193_1388# RWL_26 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10665 a_6223_7058# a_6022_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10666 GND a_10662_2176# a_10569_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10667 a_6602_4606# a_6509_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10668 VDD a_15882_8116# a_15789_8116# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10669 a_1382_2446# a_1289_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10670 a_6602_8386# a_6509_8386# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10671 GND a_3702_8386# a_3609_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10672 a_1382_6226# a_1289_6226# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10673 WBL_2 WWL_6 a_1382_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10674 a_16369_2446# WWL_22 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10675 VDD a_12402_2716# a_12309_2716# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10676 a_12982_7846# a_12889_7846# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10677 a_15302_5146# a_15209_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10678 RBL0_30 RWL_19 a_17823_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10679 a_14722_4066# a_14629_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10680 WBL_25 WWL_0 a_14722_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10681 RBL0_10 RWL_0 a_6223_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10682 WBL_15 WWL_20 a_8922_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10683 WBL_17 WWL_4 a_10082_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10684 WBL_0 WWL_13 a_222_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10685 RBL0_1 RWL_8 a_1003_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10686 a_17042_1906# a_16949_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10687 a_17042_5686# a_16949_5686# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10688 GND a_17042_7846# a_16949_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10689 a_6453_6518# RWL_7 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10690 VDD a_8342_7846# a_8249_7846# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10691 GND a_16369_7846# a_16313_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10692 WBL_9 WWL_26 a_5442_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10693 a_1233_4358# RWL_15 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10694 a_8773_7598# a_4683_7576# RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10695 a_13183_2738# a_12982_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10696 GND a_9989_5146# a_9933_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10697 a_10082_17# a_9989_17# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10698 a_15153_7058# RWL_5 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10699 a_12309_7576# WWL_3 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10700 a_11729_6496# WWL_7 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10701 RBL0_19 RWL_4 a_11443_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10702 WBL_24 WWL_24 a_14142_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10703 RBL0_18 RWL_8 a_10863_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10704 WBL_19 WWL_29 a_11242_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10705 GND a_1962_1366# a_1869_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10706 VDD a_16462_17# a_16369_17# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10707 WBL_8 WWL_1 a_4862_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10708 GND a_13562_2986# a_13469_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10709 a_11673_5438# RWL_11 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10710 a_7669_1636# WWL_25 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10711 a_15882_1906# a_15789_1906# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10712 a_9989_2716# WWL_21 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10713 GND a_12889_2986# a_12833_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10714 GND a_15882_4066# a_15789_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10715 a_6602_4336# a_6509_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10716 a_1382_2176# a_1289_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10717 a_6602_8116# a_6509_8116# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10718 GND a_3702_8116# a_3609_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10719 WBL_2 WWL_7 a_1382_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10720 a_16369_2176# WWL_23 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10721 VDD a_17622_4606# a_17529_4606# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10722 a_3122_2716# a_3029_2716# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10723 GND a_3122_4876# a_3029_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10724 a_7089_8386# WWL_0 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10725 WBL_25 WWL_1 a_14722_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10726 RBL0_10 RWL_1 a_6223_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10727 a_16313_1118# RWL_27 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10728 GND a_2449_4876# a_2393_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10729 a_17042_1636# a_16949_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10730 a_4483_1928# a_4282_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10731 a_17042_5416# a_16949_5416# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10732 a_15209_556# WWL_29 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10733 GND a_17042_7576# a_16949_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10734 GND a_14049_6496# a_13993_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10735 WBL_20 WWL_17 a_11822_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10736 GND a_4282_826# a_4189_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10737 a_3609_6766# WWL_6 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10738 a_6453_6248# RWL_8 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10739 WBL_9 WWL_27 a_5442_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10740 a_1233_4088# RWL_16 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10741 GND a_16369_7576# a_16313_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10742 RBL0_4 RWL_7 a_2743_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10743 a_18403_4628# a_18202_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10744 a_13183_2468# a_12982_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10745 a_18202_17# a_18109_17# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10746 a_13562_3796# a_13469_3796# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10747 GND a_13562_5956# a_13469_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10748 a_16949_8386# WWL_0 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10749 a_2973_4628# RWL_14 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10750 a_12309_7306# WWL_4 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10751 a_11729_6226# WWL_8 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10752 VDD a_4862_5956# a_4769_5956# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10753 RBL0_19 RWL_5 a_11443_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10754 GND a_12889_5956# a_12833_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10755 GND a_18109_1096# a_18053_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10756 RBL0_22 RWL_17 a_13183_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10757 a_16893_7328# RWL_4 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10758 a_17622_7846# a_17529_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10759 a_11673_5168# RWL_12 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10760 a_7669_1366# WWL_26 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10761 VDD a_8922_3796# a_8829_3796# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10762 a_12982_6766# a_12889_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10763 RBL0_11 RWL_27 a_6803_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10764 VDD a_3702_1636# a_3609_1636# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10765 VDD a_4282_2716# a_4189_2716# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10766 a_4282_2986# a_4189_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10767 RBL0_26 RWL_13 a_15503_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10768 a_6602_4066# a_6509_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10769 VDD a_15302_3256# a_15209_3256# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10770 WBL_11 WWL_0 a_6602_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10771 a_1003_848# a_802_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10772 WBL_2 WWL_8 a_1382_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10773 a_3553_848# RWL_28 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10774 a_16369_1906# WWL_24 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10775 VDD a_17622_4336# a_17529_4336# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10776 GND a_6022_5686# a_5929_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10777 a_8342_4606# a_8249_4606# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10778 WBL_22 WWL_2 a_12982_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10779 GND a_8342_6766# a_8249_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10780 GND a_5349_5686# a_5293_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10781 a_7089_8116# WWL_1 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10782 GND a_7669_6766# a_7613_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10783 a_1003_5708# a_802_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10784 a_9703_3818# a_9502_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10785 a_17042_1366# a_16949_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10786 a_4483_1658# a_4282_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10787 a_129_6766# WWL_6 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10788 RBL0_2 RWL_28 a_1583_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10789 WBL_29 WWL_10 a_17042_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10790 RBL0_13 RWL_14 a_7963_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10791 WBL_20 WWL_18 a_11822_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10792 GND a_14049_6226# a_13993_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10793 GND a_4282_556# a_4189_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10794 a_3609_6496# WWL_7 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10795 RBL0_4 RWL_8 a_2743_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10796 GND a_1289_826# a_1233_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10797 a_11242_2446# a_11149_2446# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10798 a_18403_4358# a_18202_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10799 a_13183_2198# a_12982_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10800 GND a_11242_4606# a_11149_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10801 a_14629_7036# WWL_5 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10802 a_16893_309# RWL_30 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10803 a_13562_3526# a_13469_3526# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10804 VDD a_11242_8386# a_11149_8386# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10805 GND a_10569_4606# a_10513_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10806 a_4282_5956# a_4189_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10807 a_2973_4358# RWL_15 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10808 a_16949_8116# WWL_1 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10809 a_14923_2738# a_14722_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10810 a_14049_3796# WWL_17 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10811 RBL0_31 RWL_10 a_18403_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10812 VDD a_6602_2446# a_6509_2446# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10813 RBL0_22 RWL_18 a_13183_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10814 a_16893_7058# RWL_5 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10815 RBL0_25 RWL_30 a_14923_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10816 a_17622_7576# a_17529_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10817 a_7669_1096# WWL_27 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10818 VDD a_8922_3526# a_8829_3526# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10819 a_17622_826# a_17529_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10820 WBL_7 WWL_5 a_4282_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10821 a_11443_7328# a_11242_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10822 VDD a_15302_2986# a_15209_2986# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10823 WBL_11 WWL_1 a_6602_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10824 a_1003_578# a_802_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10825 a_6022_3256# a_5929_3256# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10826 a_3553_578# RWL_29 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10827 GND a_6022_5416# a_5929_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10829 a_4133_7868# RWL_2 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10830 a_8342_4336# a_8249_4336# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10831 GND a_5349_5416# a_5293_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10832 WBL_5 WWL_21 a_3122_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10833 GND a_8829_17# a_8773_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10834 VDD a_11822_1366# a_11729_1366# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10835 a_9703_3548# a_9502_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10836 a_1003_5438# a_802_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10837 a_4483_1388# a_4282_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10838 GND a_2542_3796# a_2449_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10839 RBL0_2 RWL_29 a_1583_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10840 a_4862_2716# a_4769_2716# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10841 a_129_6496# WWL_7 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10842 WBL_29 WWL_11 a_17042_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10843 RBL0_13 RWL_15 a_7963_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10844 VDD a_2542_7576# a_2449_7576# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10845 a_1289_5146# WWL_12 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10846 a_16083_3008# a_15882_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10847 GND a_1869_3796# a_1813_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10848 GND a_4862_4876# a_4769_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10850 a_3609_6226# WWL_8 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10851 GND a_1289_556# a_1233_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10852 a_18403_4088# a_18202_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10853 a_11242_2176# a_11149_2176# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10854 GND a_16462_6496# a_16369_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10855 GND a_11242_4336# a_11149_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10856 a_15209_7846# WWL_2 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10857 WBL_23 WWL_17 a_13562_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10858 a_1962_4606# a_1869_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10859 VDD a_11242_8116# a_11149_8116# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10860 GND a_15789_6496# a_15733_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10861 RBL0_7 RWL_21 a_4483_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10862 a_9502_7846# a_9409_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10863 GND a_10569_4336# a_10513_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10864 a_1962_8386# a_1869_8386# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10865 a_2973_4088# RWL_16 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10866 GND a_11822_826# a_11729_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10867 a_14923_2468# a_14722_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10868 a_5293_1928# RWL_24 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10869 a_2743_6518# a_2542_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10870 RBL0_31 RWL_11 a_18403_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10871 VDD a_6602_2176# a_6509_2176# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10872 VDD a_7182_3256# a_7089_3256# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10873 a_14049_3526# WWL_18 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10874 RBL0_22 RWL_19 a_13183_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10875 a_17622_556# a_17529_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10876 a_11443_7058# a_11242_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10877 a_12402_5686# a_12309_5686# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10878 RBL0_25 RWL_17 a_14923_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10879 a_11822_4606# a_11729_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10880 WBL_5 WWL_28 a_3122_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10881 a_6022_2986# a_5929_2986# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10882 a_11822_8386# a_11729_8386# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10883 GND a_6022_5146# a_5929_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10884 a_4133_7598# RWL_3 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10885 WBL_14 WWL_14 a_8342_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10886 a_16083_5978# a_15882_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10887 GND a_5349_5146# a_5293_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10888 VDD a_11822_1096# a_11729_1096# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10889 a_2542_1366# a_2449_1366# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10890 a_9703_3278# a_9502_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10891 GND a_7762_5686# a_7669_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10892 a_1003_5168# a_802_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10893 GND a_2542_3526# a_2449_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10894 a_6509_7036# WWL_5 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10895 a_129_6226# WWL_8 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10896 a_5929_5956# WWL_9 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10897 VDD a_2542_7306# a_2449_7306# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10898 RBL0_13 RWL_16 a_7963_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10899 GND a_709_4876# a_653_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10900 a_1289_4876# WWL_13 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10901 GND a_1869_3526# a_1813_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10902 a_3029_1636# WWL_25 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10903 a_16462_4066# a_16369_4066# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10904 a_11242_1906# a_11149_1906# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10905 WBL_19 WWL_22 a_11242_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10906 GND a_16462_6226# a_16369_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10907 a_7182_6496# a_7089_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10908 WBL_28 WWL_30 a_16462_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10909 a_5349_2716# WWL_21 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10910 GND a_11242_4066# a_11149_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10911 WBL_23 WWL_18 a_13562_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10912 RBL0_16 RWL_14 a_9703_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10913 GND a_15789_6226# a_15733_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10914 RBL0_7 RWL_22 a_4483_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10915 a_1962_4336# a_1869_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10916 GND a_10569_4066# a_10513_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10917 a_1962_8116# a_1869_8116# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10918 a_9502_7576# a_9409_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10919 a_12603_1118# a_12402_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10920 VDD a_18202_6766# a_18109_6766# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10921 a_7089_826# WWL_28 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10922 GND a_11822_556# a_11729_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10923 a_14923_2198# a_14722_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10924 a_5293_1658# RWL_25 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10925 a_9933_2738# RWL_21 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10926 GND a_12982_4606# a_12889_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10927 a_7963_8408# a_7762_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10928 VDD a_12982_8386# a_12889_8386# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10929 a_3323_7328# a_3122_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10930 a_2743_6248# a_2542_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10931 VDD a_6602_1906# a_6509_1906# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10932 VDD a_7182_2986# a_7089_2986# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10933 RBL0_31 RWL_12 a_18403_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10934 GND a_6509_17# a_6453_39# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10935 a_15789_3796# WWL_17 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10936 a_12402_5416# a_12309_5416# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10937 RBL0_25 RWL_18 a_14923_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10938 a_7033_8408# RWL_0 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10939 a_11822_4336# a_11729_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10940 a_11822_8116# a_11729_8116# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10941 WBL_10 WWL_19 a_6022_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10942 a_7762_3256# a_7669_3256# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10943 a_2542_1096# a_2449_1096# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10944 WBL_4 WWL_25 a_2542_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10945 GND a_7762_5416# a_7669_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10946 a_5873_7868# RWL_2 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10947 GND a_2542_3256# a_2449_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10948 VDD a_2542_7036# a_2449_7036# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10949 GND a_1869_3256# a_1813_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10950 a_12253_7328# RWL_4 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10951 a_3029_1366# WWL_26 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10952 WBL_28 WWL_15 a_16462_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10953 WBL_19 WWL_23 a_11242_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10954 RBL0_3 RWL_27 a_2163_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10955 WBL_28 WWL_31 a_16462_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10956 a_7182_6226# a_7089_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10957 RBL0_16 RWL_15 a_9703_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10958 RBL0_7 RWL_23 a_4483_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10959 a_1962_4066# a_1869_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10960 GND a_18202_2716# a_18109_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10961 a_17823_3008# a_17622_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10962 WBL_3 WWL_0 a_1962_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10963 VDD a_18202_6496# a_18109_6496# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10964 a_8922_6766# a_8829_6766# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10966 GND a_17529_2716# a_17473_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10967 a_9933_2468# RWL_22 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10968 GND a_12982_4336# a_12889_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10969 a_7963_8138# a_7762_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10970 a_5293_1388# RWL_26 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10971 a_3323_7058# a_3122_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10972 a_3702_4606# a_3609_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10973 VDD a_12982_8116# a_12889_8116# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10974 a_3702_8386# a_3609_8386# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10975 GND a_3029_6766# a_2973_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10976 a_5063_3818# a_4862_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10977 VDD a_222_1366# a_129_1366# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10978 a_13469_2446# WWL_22 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10979 VDD a_10082_3796# a_9989_3796# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10980 a_7383_4898# a_7182_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10981 a_10082_7846# a_9989_7846# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10982 a_15789_3526# WWL_18 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10983 a_12402_5146# a_12309_5146# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10984 RBL0_25 RWL_19 a_14923_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10985 a_7033_8138# RWL_1 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10986 a_11822_4066# a_11729_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10987 RBL0_5 RWL_0 a_3323_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10988 WBL_10 WWL_20 a_6022_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10989 a_14142_1906# a_14049_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10990 a_14142_5686# a_14049_5686# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10991 GND a_14142_7846# a_14049_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10992 a_3553_6518# RWL_7 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10993 a_8829_287# WWL_30 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10994 a_7762_2986# a_7669_2986# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10995 VDD a_5442_7846# a_5349_7846# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10996 GND a_13469_7846# a_13413_7868# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10997 VDD a_10082_826# a_9989_826# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10998 WBL_4 WWL_26 a_2542_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10999 GND a_7762_5146# a_7669_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11000 a_5873_7598# a_4683_7576# RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11001 a_10283_2738# a_10082_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11002 a_17823_5978# a_17622_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11003 GND a_9502_1906# a_9409_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11004 GND a_802_3796# a_709_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11005 VDD a_802_7576# a_709_7576# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11006 a_12253_7058# RWL_5 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11007 RBL0_27 RWL_6 a_16083_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11008 VDD a_9502_5686# a_9409_5686# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11009 GND a_8829_1906# a_8773_1928# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11010 a_8249_3256# WWL_19 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11011 WBL_28 WWL_16 a_16462_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11012 a_3029_1096# WWL_27 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11013 RBL0_12 RWL_20 a_7383_3008# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11014 WBL_19 WWL_24 a_11242_1906# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11015 a_222_826# a_129_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11016 RBL0_16 RWL_16 a_9703_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11017 GND a_17042_17# a_16949_17# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11018 GND a_18202_2446# a_18109_2446# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11019 WBL_3 WWL_1 a_1962_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11020 a_8922_2716# a_8829_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11021 GND a_10662_2986# a_10569_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11022 VDD a_18202_6226# a_18109_6226# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11023 a_4769_1636# WWL_25 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11024 a_222_4606# a_129_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11025 GND a_17529_2446# a_17473_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11026 a_222_8386# a_129_8386# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11027 a_8922_6496# a_8829_6496# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11028 a_9933_2198# RWL_23 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11029 GND a_12982_4066# a_12889_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11030 a_3702_4336# a_3609_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11031 a_3702_8116# a_3609_8116# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11032 a_5063_3548# a_4862_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11033 VDD a_222_1096# a_129_1096# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11034 a_13469_2176# WWL_23 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11035 VDD a_14722_4606# a_14629_4606# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11036 VDD a_10082_3526# a_9989_3526# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11037 a_14629_826# WWL_28 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11038 a_4189_8386# WWL_0 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11039 RBL0_5 RWL_1 a_3323_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11040 a_13413_1118# RWL_27 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11041 a_14142_1636# a_14049_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11042 a_1583_1928# a_1382_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11043 a_17622_287# a_17529_287# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11044 a_14142_5416# a_14049_5416# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11045 a_15733_39# RWL_31 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11046 GND a_14142_7576# a_14049_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11047 GND a_11149_6496# a_11093_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11048 a_8773_8408# RWL_0 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11049 a_3553_6248# RWL_8 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11050 RBL0_12 RWL_9 a_7383_5978# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11051 a_8829_17# WWL_31 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11052 WBL_13 WWL_19 a_7762_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11053 GND a_13469_7576# a_13413_7598# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11054 WBL_4 WWL_27 a_2542_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11055 a_15503_4628# a_15302_4606# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11056 a_10283_2468# a_10082_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11057 a_10662_3796# a_10569_3796# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11058 GND a_10662_5956# a_10569_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11059 GND a_9502_1636# a_9409_1636# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11060 GND a_802_3526# a_709_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11061 VDD a_802_7306# a_709_7306# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11062 VDD a_9502_5416# a_9409_5416# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11063 a_8249_2986# WWL_20 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11064 VDD a_1962_5956# a_1869_5956# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11065 GND a_8829_1636# a_8773_1658# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11066 a_222_556# a_129_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11067 RBL0_17 RWL_17 a_10283_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11068 GND a_15209_1096# a_15153_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11069 GND a_18202_2176# a_18109_2176# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11070 a_13993_7328# RWL_4 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11071 a_8922_2446# a_8829_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11072 a_14722_7846# a_14629_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11073 a_10082_6766# a_9989_6766# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11074 a_4769_1366# WWL_26 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11075 VDD a_1382_2716# a_1289_2716# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11076 a_222_4336# a_129_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11077 RBL0_6 RWL_27 a_3903_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11078 GND a_17529_2176# a_17473_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11079 a_1382_2986# a_1289_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11080 RBL0_21 RWL_13 a_12603_4898# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11081 a_222_8116# a_129_8116# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11082 WBL_15 WWL_6 a_8922_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11083 a_8922_6226# a_8829_6226# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11084 a_3702_4066# a_3609_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11085 VDD a_12402_3256# a_12309_3256# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11086 WBL_6 WWL_0 a_3702_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11087 VDD a_11822_287# a_11729_287# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11088 a_13469_1906# WWL_24 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11089 a_5063_3278# a_4862_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11090 VDD a_14722_4336# a_14629_4336# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11091 GND a_3122_5686# a_3029_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11092 a_5442_4606# a_5349_4606# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11093 WBL_17 WWL_2 a_10082_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11094 GND a_5442_6766# a_5349_6766# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11095 GND a_2449_5686# a_2393_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11096 a_4189_8116# WWL_1 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11097 GND a_4769_6766# a_4713_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11098 a_6803_3818# a_6602_3796# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11099 GND a_17042_8386# a_16949_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11100 a_14142_1366# a_14049_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11101 a_1583_1658# a_1382_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11102 a_17622_17# a_17529_17# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11103 GND a_16369_8386# a_16313_8408# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11104 WBL_24 WWL_10 a_14142_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11105 RBL0_8 RWL_14 a_5063_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11106 GND a_11149_6226# a_11093_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11107 a_8773_8138# RWL_1 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11108 WBL_13 WWL_20 a_7762_2986# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11109 a_15882_1906# a_15789_1906# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11110 a_15503_4358# a_15302_4336# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11111 a_10283_2198# a_10082_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11112 a_15882_5686# a_15789_5686# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11113 a_4713_309# RWL_30 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11114 a_10662_3526# a_10569_3526# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11115 a_11729_7036# WWL_5 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11116 GND a_15882_7846# a_15789_7846# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11117 GND a_9502_1366# a_9409_1366# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11118 GND a_802_3256# a_709_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11119 a_8193_4898# RWL_13 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11120 a_1382_5956# a_1289_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11121 VDD a_802_7036# a_709_7036# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11122 GND a_8829_1366# a_8773_1388# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11123 a_12023_2738# a_11822_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11124 RBL0_26 RWL_10 a_15503_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11125 a_11149_3796# WWL_17 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11126 VDD a_3702_2446# a_3609_2446# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11127 a_15882_556# a_15789_556# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11128 RBL0_17 RWL_18 a_10283_3548# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11129 a_13993_7058# RWL_5 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11130 a_9989_3256# WWL_19 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11131 a_14722_7576# a_14629_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11132 RBL0_30 RWL_6 a_17823_6788# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11133 a_4769_1096# WWL_27 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11134 a_8922_2176# a_8829_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11135 a_222_4066# a_129_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11136 WBL_15 WWL_7 a_8922_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11137 WBL_0 WWL_0 a_222_8386# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11138 a_5442_826# a_5349_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11139 WBL_2 WWL_5 a_1382_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11140 a_11093_2738# RWL_21 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11141 a_15733_3818# RWL_17 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11142 VDD a_17622_5146# a_17529_5146# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11143 VDD a_12402_2986# a_12309_2986# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11144 WBL_6 WWL_1 a_3702_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11145 VDD a_11822_17# a_11729_17# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11146 a_3122_3256# a_3029_3256# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11147 GND a_3122_5416# a_3029_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11148 a_1233_7868# RWL_2 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11149 a_5442_4336# a_5349_4336# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11150 GND a_2449_5416# a_2393_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11151 a_7033_848# RWL_28 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11152 a_17042_5956# a_16949_5956# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11153 a_10513_848# RWL_28 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11154 a_6803_3548# a_6602_3526# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11155 GND a_17042_8116# a_16949_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11156 a_1583_1388# a_1382_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11157 WBL_20 WWL_15 a_11822_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11158 WBL_24 WWL_11 a_14142_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11159 RBL0_8 RWL_15 a_5063_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11160 GND a_16369_8116# a_16313_8138# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11161 a_13183_3008# a_12982_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11162 GND a_1962_4876# a_1869_4876# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11163 RBL0_8 RWL_28 a_5063_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11164 a_15882_1636# a_15789_1636# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11165 a_15503_4088# a_15302_4066# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11166 a_2163_308# a_1962_286# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11167 GND a_13562_6496# a_13469_6496# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11168 VDD a_6602_556# a_6509_556# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11169 a_15882_5416# a_15789_5416# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11170 WBL_11 WWL_28 a_6602_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11171 a_12309_7846# WWL_2 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11172 GND a_7089_1096# a_7033_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11173 RBL0_2 RWL_21 a_1583_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11174 WBL_18 WWL_17 a_10662_3796# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11175 GND a_15882_7576# a_15789_7576# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11176 GND a_12889_6496# a_12833_6518# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11177 a_10569_556# WWL_29 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11178 a_6602_7846# a_6509_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11179 a_12023_2468# a_11822_2446# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11181 a_16369_5686# WWL_10 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11182 a_2393_1928# RWL_24 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11183 a_17622_8386# a_17529_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11184 a_12982_7306# a_12889_7306# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11185 RBL0_26 RWL_11 a_15503_5438# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11186 VDD a_3702_2176# a_3609_2176# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11187 VDD a_4282_3256# a_4189_3256# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11188 a_11149_3526# WWL_18 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11189 RBL0_17 RWL_19 a_10283_3278# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11190 a_9989_2986# WWL_20 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11191 WBL_15 WWL_8 a_8922_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11192 WBL_0 WWL_1 a_222_8116# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11193 GND a_17622_1096# a_17529_1096# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11194 a_5442_556# a_5349_556# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11195 a_16313_4628# RWL_14 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11196 RBL0_31 RWL_30 a_18403_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11197 a_15733_3548# RWL_18 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11198 a_11093_2468# RWL_22 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11199 VDD a_17622_4876# a_17529_4876# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11200 GND a_16949_1096# a_16893_1118# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11201 a_8342_5146# a_8249_5146# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11202 a_3122_2986# a_3029_2986# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11203 GND a_8342_7306# a_8249_7306# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11204 GND a_3122_5146# a_3029_5146# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11205 a_1233_7598# RWL_3 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11206 GND a_9502_287# a_9409_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11207 GND a_7669_7306# a_7613_7328# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11208 WBL_9 WWL_14 a_5442_4606# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11209 a_13183_5978# a_12982_5956# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11210 GND a_2449_5146# a_2393_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11211 GND a_12982_287# a_12889_287# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11212 VDD a_17042_1636# a_16949_1636# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11213 a_7033_578# RWL_29 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11214 GND a_8829_826# a_8773_848# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11215 a_10513_578# RWL_29 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11216 a_6803_3278# a_6602_3256# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11217 GND a_4862_5686# a_4769_5686# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11218 WBL_20 WWL_16 a_11822_4066# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11219 a_3609_7036# WWL_5 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11220 RBL0_8 RWL_16 a_5063_4088# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11221 RBL0_8 RWL_29 a_5063_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11222 a_13562_4066# a_13469_4066# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11223 GND a_18109_4606# a_18053_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11224 a_15882_1366# a_15789_1366# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11225 GND a_13562_6226# a_13469_6226# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11226 a_4282_6496# a_4189_6496# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11227 a_2449_2716# WWL_21 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11228 WBL_18 WWL_18 a_10662_3526# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11229 RBL0_11 RWL_14 a_6803_4628# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11230 GND a_12889_6226# a_12833_6248# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11231 RBL0_2 RWL_22 a_1583_2468# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11232 a_6602_7576# a_6509_7576# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11233 VDD a_15302_6766# a_15209_6766# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11234 a_14049_4336# WWL_15 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11235 a_12023_2198# a_11822_2176# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11236 a_7613_3818# RWL_17 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11237 a_2393_1658# RWL_25 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11238 a_17622_8116# a_17529_8116# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11239 a_16369_5416# WWL_11 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11240 VDD a_8922_4066# a_8829_4066# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11241 a_12982_7036# a_12889_7036# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11242 RBL0_26 RWL_12 a_15503_5168# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11243 VDD a_3702_1906# a_3609_1906# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11244 VDD a_4282_2986# a_4189_2986# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11245 GND a_15302_826# a_15209_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11246 a_15733_3278# RWL_19 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11247 a_16313_4358# RWL_15 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11248 a_17042_4876# a_16949_4876# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11249 a_8342_1096# a_8249_1096# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11250 a_11093_2198# RWL_23 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11251 a_12889_3796# WWL_17 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11252 a_4133_8408# RWL_0 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11253 a_8342_4876# a_8249_4876# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11254 GND a_8342_7036# a_8249_7036# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11255 WBL_5 WWL_19 a_3122_3256# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11256 a_18403_7868# a_18202_7846# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11257 GND a_7669_7036# a_7613_7058# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11258 GND a_6509_287# a_6453_309# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11259 WBL_17 WWL_28 a_10082_826# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11260 GND a_8829_556# a_8773_578# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11261 a_4862_3256# a_4769_3256# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11262 a_129_7036# WWL_5 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11263 WBL_29 WWL_9 a_17042_5956# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11264 GND a_9409_3796# a_9353_3818# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11265 GND a_709_5686# a_653_5708# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11266 a_2973_7868# RWL_2 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11267 GND a_4862_5416# a_4769_5416# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11268 a_9703_848# a_9502_826# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11269 a_423_2738# a_222_2716# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11270 GND a_18109_4336# a_18053_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11271 WBL_23 WWL_15 a_13562_4336# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11272 a_9502_8386# a_9409_8386# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11273 a_7669_4606# WWL_14 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11274 a_4282_6226# a_4189_6226# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11275 RBL0_11 RWL_15 a_6803_4358# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11276 RBL0_2 RWL_23 a_1583_2198# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11277 GND a_15302_2716# a_15209_2716# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11278 a_14923_3008# a_14722_2986# GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11279 a_17622_1636# a_17529_1636# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11280 a_18202_2716# a_18109_2716# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11281 VDD a_15302_6496# a_15209_6496# VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11282 GND a_14629_2716# a_14573_2738# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11283 a_14049_4066# WWL_16 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11284 a_6022_6766# a_5929_6766# VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11285 a_7613_3548# RWL_18 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11286 a_2393_1388# RWL_26 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11287 GND a_15302_556# a_15209_556# GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

.ends

