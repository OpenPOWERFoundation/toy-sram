magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< nwell >>
rect 0 0 720 1214
<< pmos >>
rect 204 102 240 1112
rect 296 102 332 1112
rect 388 102 424 1112
rect 480 102 516 1112
<< pdiff >>
rect 148 1100 204 1112
rect 148 1066 159 1100
rect 193 1066 204 1100
rect 148 1032 204 1066
rect 148 998 159 1032
rect 193 998 204 1032
rect 148 964 204 998
rect 148 930 159 964
rect 193 930 204 964
rect 148 896 204 930
rect 148 862 159 896
rect 193 862 204 896
rect 148 828 204 862
rect 148 794 159 828
rect 193 794 204 828
rect 148 760 204 794
rect 148 726 159 760
rect 193 726 204 760
rect 148 692 204 726
rect 148 658 159 692
rect 193 658 204 692
rect 148 624 204 658
rect 148 590 159 624
rect 193 590 204 624
rect 148 556 204 590
rect 148 522 159 556
rect 193 522 204 556
rect 148 488 204 522
rect 148 454 159 488
rect 193 454 204 488
rect 148 420 204 454
rect 148 386 159 420
rect 193 386 204 420
rect 148 352 204 386
rect 148 318 159 352
rect 193 318 204 352
rect 148 284 204 318
rect 148 250 159 284
rect 193 250 204 284
rect 148 216 204 250
rect 148 182 159 216
rect 193 182 204 216
rect 148 148 204 182
rect 148 114 159 148
rect 193 114 204 148
rect 148 102 204 114
rect 240 1100 296 1112
rect 240 1066 251 1100
rect 285 1066 296 1100
rect 240 1032 296 1066
rect 240 998 251 1032
rect 285 998 296 1032
rect 240 964 296 998
rect 240 930 251 964
rect 285 930 296 964
rect 240 896 296 930
rect 240 862 251 896
rect 285 862 296 896
rect 240 828 296 862
rect 240 794 251 828
rect 285 794 296 828
rect 240 760 296 794
rect 240 726 251 760
rect 285 726 296 760
rect 240 692 296 726
rect 240 658 251 692
rect 285 658 296 692
rect 240 624 296 658
rect 240 590 251 624
rect 285 590 296 624
rect 240 556 296 590
rect 240 522 251 556
rect 285 522 296 556
rect 240 488 296 522
rect 240 454 251 488
rect 285 454 296 488
rect 240 420 296 454
rect 240 386 251 420
rect 285 386 296 420
rect 240 352 296 386
rect 240 318 251 352
rect 285 318 296 352
rect 240 284 296 318
rect 240 250 251 284
rect 285 250 296 284
rect 240 216 296 250
rect 240 182 251 216
rect 285 182 296 216
rect 240 148 296 182
rect 240 114 251 148
rect 285 114 296 148
rect 240 102 296 114
rect 332 1100 388 1112
rect 332 1066 343 1100
rect 377 1066 388 1100
rect 332 1032 388 1066
rect 332 998 343 1032
rect 377 998 388 1032
rect 332 964 388 998
rect 332 930 343 964
rect 377 930 388 964
rect 332 896 388 930
rect 332 862 343 896
rect 377 862 388 896
rect 332 828 388 862
rect 332 794 343 828
rect 377 794 388 828
rect 332 760 388 794
rect 332 726 343 760
rect 377 726 388 760
rect 332 692 388 726
rect 332 658 343 692
rect 377 658 388 692
rect 332 624 388 658
rect 332 590 343 624
rect 377 590 388 624
rect 332 556 388 590
rect 332 522 343 556
rect 377 522 388 556
rect 332 488 388 522
rect 332 454 343 488
rect 377 454 388 488
rect 332 420 388 454
rect 332 386 343 420
rect 377 386 388 420
rect 332 352 388 386
rect 332 318 343 352
rect 377 318 388 352
rect 332 284 388 318
rect 332 250 343 284
rect 377 250 388 284
rect 332 216 388 250
rect 332 182 343 216
rect 377 182 388 216
rect 332 148 388 182
rect 332 114 343 148
rect 377 114 388 148
rect 332 102 388 114
rect 424 1100 480 1112
rect 424 1066 435 1100
rect 469 1066 480 1100
rect 424 1032 480 1066
rect 424 998 435 1032
rect 469 998 480 1032
rect 424 964 480 998
rect 424 930 435 964
rect 469 930 480 964
rect 424 896 480 930
rect 424 862 435 896
rect 469 862 480 896
rect 424 828 480 862
rect 424 794 435 828
rect 469 794 480 828
rect 424 760 480 794
rect 424 726 435 760
rect 469 726 480 760
rect 424 692 480 726
rect 424 658 435 692
rect 469 658 480 692
rect 424 624 480 658
rect 424 590 435 624
rect 469 590 480 624
rect 424 556 480 590
rect 424 522 435 556
rect 469 522 480 556
rect 424 488 480 522
rect 424 454 435 488
rect 469 454 480 488
rect 424 420 480 454
rect 424 386 435 420
rect 469 386 480 420
rect 424 352 480 386
rect 424 318 435 352
rect 469 318 480 352
rect 424 284 480 318
rect 424 250 435 284
rect 469 250 480 284
rect 424 216 480 250
rect 424 182 435 216
rect 469 182 480 216
rect 424 148 480 182
rect 424 114 435 148
rect 469 114 480 148
rect 424 102 480 114
rect 516 1100 572 1112
rect 516 1066 527 1100
rect 561 1066 572 1100
rect 516 1032 572 1066
rect 516 998 527 1032
rect 561 998 572 1032
rect 516 964 572 998
rect 516 930 527 964
rect 561 930 572 964
rect 516 896 572 930
rect 516 862 527 896
rect 561 862 572 896
rect 516 828 572 862
rect 516 794 527 828
rect 561 794 572 828
rect 516 760 572 794
rect 516 726 527 760
rect 561 726 572 760
rect 516 692 572 726
rect 516 658 527 692
rect 561 658 572 692
rect 516 624 572 658
rect 516 590 527 624
rect 561 590 572 624
rect 516 556 572 590
rect 516 522 527 556
rect 561 522 572 556
rect 516 488 572 522
rect 516 454 527 488
rect 561 454 572 488
rect 516 420 572 454
rect 516 386 527 420
rect 561 386 572 420
rect 516 352 572 386
rect 516 318 527 352
rect 561 318 572 352
rect 516 284 572 318
rect 516 250 527 284
rect 561 250 572 284
rect 516 216 572 250
rect 516 182 527 216
rect 561 182 572 216
rect 516 148 572 182
rect 516 114 527 148
rect 561 114 572 148
rect 516 102 572 114
<< pdiffc >>
rect 159 1066 193 1100
rect 159 998 193 1032
rect 159 930 193 964
rect 159 862 193 896
rect 159 794 193 828
rect 159 726 193 760
rect 159 658 193 692
rect 159 590 193 624
rect 159 522 193 556
rect 159 454 193 488
rect 159 386 193 420
rect 159 318 193 352
rect 159 250 193 284
rect 159 182 193 216
rect 159 114 193 148
rect 251 1066 285 1100
rect 251 998 285 1032
rect 251 930 285 964
rect 251 862 285 896
rect 251 794 285 828
rect 251 726 285 760
rect 251 658 285 692
rect 251 590 285 624
rect 251 522 285 556
rect 251 454 285 488
rect 251 386 285 420
rect 251 318 285 352
rect 251 250 285 284
rect 251 182 285 216
rect 251 114 285 148
rect 343 1066 377 1100
rect 343 998 377 1032
rect 343 930 377 964
rect 343 862 377 896
rect 343 794 377 828
rect 343 726 377 760
rect 343 658 377 692
rect 343 590 377 624
rect 343 522 377 556
rect 343 454 377 488
rect 343 386 377 420
rect 343 318 377 352
rect 343 250 377 284
rect 343 182 377 216
rect 343 114 377 148
rect 435 1066 469 1100
rect 435 998 469 1032
rect 435 930 469 964
rect 435 862 469 896
rect 435 794 469 828
rect 435 726 469 760
rect 435 658 469 692
rect 435 590 469 624
rect 435 522 469 556
rect 435 454 469 488
rect 435 386 469 420
rect 435 318 469 352
rect 435 250 469 284
rect 435 182 469 216
rect 435 114 469 148
rect 527 1066 561 1100
rect 527 998 561 1032
rect 527 930 561 964
rect 527 862 561 896
rect 527 794 561 828
rect 527 726 561 760
rect 527 658 561 692
rect 527 590 561 624
rect 527 522 561 556
rect 527 454 561 488
rect 527 386 561 420
rect 527 318 561 352
rect 527 250 561 284
rect 527 182 561 216
rect 527 114 561 148
<< nsubdiff >>
rect 36 1066 94 1112
rect 36 1032 48 1066
rect 82 1032 94 1066
rect 36 998 94 1032
rect 36 964 48 998
rect 82 964 94 998
rect 36 930 94 964
rect 36 896 48 930
rect 82 896 94 930
rect 36 862 94 896
rect 36 828 48 862
rect 82 828 94 862
rect 36 794 94 828
rect 36 760 48 794
rect 82 760 94 794
rect 36 726 94 760
rect 36 692 48 726
rect 82 692 94 726
rect 36 658 94 692
rect 36 624 48 658
rect 82 624 94 658
rect 36 590 94 624
rect 36 556 48 590
rect 82 556 94 590
rect 36 522 94 556
rect 36 488 48 522
rect 82 488 94 522
rect 36 454 94 488
rect 36 420 48 454
rect 82 420 94 454
rect 36 386 94 420
rect 36 352 48 386
rect 82 352 94 386
rect 36 318 94 352
rect 36 284 48 318
rect 82 284 94 318
rect 36 250 94 284
rect 36 216 48 250
rect 82 216 94 250
rect 36 182 94 216
rect 36 148 48 182
rect 82 148 94 182
rect 36 102 94 148
rect 626 1066 684 1112
rect 626 1032 638 1066
rect 672 1032 684 1066
rect 626 998 684 1032
rect 626 964 638 998
rect 672 964 684 998
rect 626 930 684 964
rect 626 896 638 930
rect 672 896 684 930
rect 626 862 684 896
rect 626 828 638 862
rect 672 828 684 862
rect 626 794 684 828
rect 626 760 638 794
rect 672 760 684 794
rect 626 726 684 760
rect 626 692 638 726
rect 672 692 684 726
rect 626 658 684 692
rect 626 624 638 658
rect 672 624 684 658
rect 626 590 684 624
rect 626 556 638 590
rect 672 556 684 590
rect 626 522 684 556
rect 626 488 638 522
rect 672 488 684 522
rect 626 454 684 488
rect 626 420 638 454
rect 672 420 684 454
rect 626 386 684 420
rect 626 352 638 386
rect 672 352 684 386
rect 626 318 684 352
rect 626 284 638 318
rect 672 284 684 318
rect 626 250 684 284
rect 626 216 638 250
rect 672 216 684 250
rect 626 182 684 216
rect 626 148 638 182
rect 672 148 684 182
rect 626 102 684 148
<< nsubdiffcont >>
rect 48 1032 82 1066
rect 48 964 82 998
rect 48 896 82 930
rect 48 828 82 862
rect 48 760 82 794
rect 48 692 82 726
rect 48 624 82 658
rect 48 556 82 590
rect 48 488 82 522
rect 48 420 82 454
rect 48 352 82 386
rect 48 284 82 318
rect 48 216 82 250
rect 48 148 82 182
rect 638 1032 672 1066
rect 638 964 672 998
rect 638 896 672 930
rect 638 828 672 862
rect 638 760 672 794
rect 638 692 672 726
rect 638 624 672 658
rect 638 556 672 590
rect 638 488 672 522
rect 638 420 672 454
rect 638 352 672 386
rect 638 284 672 318
rect 638 216 672 250
rect 638 148 672 182
<< poly >>
rect 191 1194 529 1214
rect 191 1160 207 1194
rect 241 1160 275 1194
rect 309 1160 343 1194
rect 377 1160 411 1194
rect 445 1160 479 1194
rect 513 1160 529 1194
rect 191 1144 529 1160
rect 204 1112 240 1144
rect 296 1112 332 1144
rect 388 1112 424 1144
rect 480 1112 516 1144
rect 204 70 240 102
rect 296 70 332 102
rect 388 70 424 102
rect 480 70 516 102
rect 191 54 529 70
rect 191 20 207 54
rect 241 20 275 54
rect 309 20 343 54
rect 377 20 411 54
rect 445 20 479 54
rect 513 20 529 54
rect 191 0 529 20
<< polycont >>
rect 207 1160 241 1194
rect 275 1160 309 1194
rect 343 1160 377 1194
rect 411 1160 445 1194
rect 479 1160 513 1194
rect 207 20 241 54
rect 275 20 309 54
rect 343 20 377 54
rect 411 20 445 54
rect 479 20 513 54
<< locali >>
rect 191 1160 199 1194
rect 241 1160 271 1194
rect 309 1160 343 1194
rect 377 1160 411 1194
rect 449 1160 479 1194
rect 521 1160 529 1194
rect 159 1100 193 1116
rect 48 1020 82 1032
rect 48 948 82 964
rect 48 876 82 896
rect 48 804 82 828
rect 48 732 82 760
rect 48 660 82 692
rect 48 590 82 624
rect 48 522 82 554
rect 48 454 82 482
rect 48 386 82 410
rect 48 318 82 338
rect 48 250 82 266
rect 48 182 82 194
rect 159 1032 193 1058
rect 159 964 193 986
rect 159 896 193 914
rect 159 828 193 842
rect 159 760 193 770
rect 159 692 193 698
rect 159 624 193 626
rect 159 588 193 590
rect 159 516 193 522
rect 159 444 193 454
rect 159 372 193 386
rect 159 300 193 318
rect 159 228 193 250
rect 159 156 193 182
rect 159 98 193 114
rect 251 1100 285 1116
rect 251 1032 285 1058
rect 251 964 285 986
rect 251 896 285 914
rect 251 828 285 842
rect 251 760 285 770
rect 251 692 285 698
rect 251 624 285 626
rect 251 588 285 590
rect 251 516 285 522
rect 251 444 285 454
rect 251 372 285 386
rect 251 300 285 318
rect 251 228 285 250
rect 251 156 285 182
rect 251 98 285 114
rect 343 1100 377 1116
rect 343 1032 377 1058
rect 343 964 377 986
rect 343 896 377 914
rect 343 828 377 842
rect 343 760 377 770
rect 343 692 377 698
rect 343 624 377 626
rect 343 588 377 590
rect 343 516 377 522
rect 343 444 377 454
rect 343 372 377 386
rect 343 300 377 318
rect 343 228 377 250
rect 343 156 377 182
rect 343 98 377 114
rect 435 1100 469 1116
rect 435 1032 469 1058
rect 435 964 469 986
rect 435 896 469 914
rect 435 828 469 842
rect 435 760 469 770
rect 435 692 469 698
rect 435 624 469 626
rect 435 588 469 590
rect 435 516 469 522
rect 435 444 469 454
rect 435 372 469 386
rect 435 300 469 318
rect 435 228 469 250
rect 435 156 469 182
rect 435 98 469 114
rect 527 1100 561 1116
rect 527 1032 561 1058
rect 527 964 561 986
rect 527 896 561 914
rect 527 828 561 842
rect 527 760 561 770
rect 527 692 561 698
rect 527 624 561 626
rect 527 588 561 590
rect 527 516 561 522
rect 527 444 561 454
rect 527 372 561 386
rect 527 300 561 318
rect 527 228 561 250
rect 527 156 561 182
rect 638 1020 672 1032
rect 638 948 672 964
rect 638 876 672 896
rect 638 804 672 828
rect 638 732 672 760
rect 638 660 672 692
rect 638 590 672 624
rect 638 522 672 554
rect 638 454 672 482
rect 638 386 672 410
rect 638 318 672 338
rect 638 250 672 266
rect 638 182 672 194
rect 527 98 561 114
rect 191 20 199 54
rect 241 20 271 54
rect 309 20 343 54
rect 377 20 411 54
rect 449 20 479 54
rect 521 20 529 54
<< viali >>
rect 199 1160 207 1194
rect 207 1160 233 1194
rect 271 1160 275 1194
rect 275 1160 305 1194
rect 343 1160 377 1194
rect 415 1160 445 1194
rect 445 1160 449 1194
rect 487 1160 513 1194
rect 513 1160 521 1194
rect 48 1066 82 1092
rect 48 1058 82 1066
rect 48 998 82 1020
rect 48 986 82 998
rect 48 930 82 948
rect 48 914 82 930
rect 48 862 82 876
rect 48 842 82 862
rect 48 794 82 804
rect 48 770 82 794
rect 48 726 82 732
rect 48 698 82 726
rect 48 658 82 660
rect 48 626 82 658
rect 48 556 82 588
rect 48 554 82 556
rect 48 488 82 516
rect 48 482 82 488
rect 48 420 82 444
rect 48 410 82 420
rect 48 352 82 372
rect 48 338 82 352
rect 48 284 82 300
rect 48 266 82 284
rect 48 216 82 228
rect 48 194 82 216
rect 48 148 82 156
rect 48 122 82 148
rect 159 1066 193 1092
rect 159 1058 193 1066
rect 159 998 193 1020
rect 159 986 193 998
rect 159 930 193 948
rect 159 914 193 930
rect 159 862 193 876
rect 159 842 193 862
rect 159 794 193 804
rect 159 770 193 794
rect 159 726 193 732
rect 159 698 193 726
rect 159 658 193 660
rect 159 626 193 658
rect 159 556 193 588
rect 159 554 193 556
rect 159 488 193 516
rect 159 482 193 488
rect 159 420 193 444
rect 159 410 193 420
rect 159 352 193 372
rect 159 338 193 352
rect 159 284 193 300
rect 159 266 193 284
rect 159 216 193 228
rect 159 194 193 216
rect 159 148 193 156
rect 159 122 193 148
rect 251 1066 285 1092
rect 251 1058 285 1066
rect 251 998 285 1020
rect 251 986 285 998
rect 251 930 285 948
rect 251 914 285 930
rect 251 862 285 876
rect 251 842 285 862
rect 251 794 285 804
rect 251 770 285 794
rect 251 726 285 732
rect 251 698 285 726
rect 251 658 285 660
rect 251 626 285 658
rect 251 556 285 588
rect 251 554 285 556
rect 251 488 285 516
rect 251 482 285 488
rect 251 420 285 444
rect 251 410 285 420
rect 251 352 285 372
rect 251 338 285 352
rect 251 284 285 300
rect 251 266 285 284
rect 251 216 285 228
rect 251 194 285 216
rect 251 148 285 156
rect 251 122 285 148
rect 343 1066 377 1092
rect 343 1058 377 1066
rect 343 998 377 1020
rect 343 986 377 998
rect 343 930 377 948
rect 343 914 377 930
rect 343 862 377 876
rect 343 842 377 862
rect 343 794 377 804
rect 343 770 377 794
rect 343 726 377 732
rect 343 698 377 726
rect 343 658 377 660
rect 343 626 377 658
rect 343 556 377 588
rect 343 554 377 556
rect 343 488 377 516
rect 343 482 377 488
rect 343 420 377 444
rect 343 410 377 420
rect 343 352 377 372
rect 343 338 377 352
rect 343 284 377 300
rect 343 266 377 284
rect 343 216 377 228
rect 343 194 377 216
rect 343 148 377 156
rect 343 122 377 148
rect 435 1066 469 1092
rect 435 1058 469 1066
rect 435 998 469 1020
rect 435 986 469 998
rect 435 930 469 948
rect 435 914 469 930
rect 435 862 469 876
rect 435 842 469 862
rect 435 794 469 804
rect 435 770 469 794
rect 435 726 469 732
rect 435 698 469 726
rect 435 658 469 660
rect 435 626 469 658
rect 435 556 469 588
rect 435 554 469 556
rect 435 488 469 516
rect 435 482 469 488
rect 435 420 469 444
rect 435 410 469 420
rect 435 352 469 372
rect 435 338 469 352
rect 435 284 469 300
rect 435 266 469 284
rect 435 216 469 228
rect 435 194 469 216
rect 435 148 469 156
rect 435 122 469 148
rect 527 1066 561 1092
rect 527 1058 561 1066
rect 527 998 561 1020
rect 527 986 561 998
rect 527 930 561 948
rect 527 914 561 930
rect 527 862 561 876
rect 527 842 561 862
rect 527 794 561 804
rect 527 770 561 794
rect 527 726 561 732
rect 527 698 561 726
rect 527 658 561 660
rect 527 626 561 658
rect 527 556 561 588
rect 527 554 561 556
rect 527 488 561 516
rect 527 482 561 488
rect 527 420 561 444
rect 527 410 561 420
rect 527 352 561 372
rect 527 338 561 352
rect 527 284 561 300
rect 527 266 561 284
rect 527 216 561 228
rect 527 194 561 216
rect 527 148 561 156
rect 527 122 561 148
rect 638 1066 672 1092
rect 638 1058 672 1066
rect 638 998 672 1020
rect 638 986 672 998
rect 638 930 672 948
rect 638 914 672 930
rect 638 862 672 876
rect 638 842 672 862
rect 638 794 672 804
rect 638 770 672 794
rect 638 726 672 732
rect 638 698 672 726
rect 638 658 672 660
rect 638 626 672 658
rect 638 556 672 588
rect 638 554 672 556
rect 638 488 672 516
rect 638 482 672 488
rect 638 420 672 444
rect 638 410 672 420
rect 638 352 672 372
rect 638 338 672 352
rect 638 284 672 300
rect 638 266 672 284
rect 638 216 672 228
rect 638 194 672 216
rect 638 148 672 156
rect 638 122 672 148
rect 199 20 207 54
rect 207 20 233 54
rect 271 20 275 54
rect 275 20 305 54
rect 343 20 377 54
rect 415 20 445 54
rect 445 20 449 54
rect 487 20 513 54
rect 513 20 521 54
<< metal1 >>
rect 187 1194 533 1214
rect 187 1160 199 1194
rect 233 1160 271 1194
rect 305 1160 343 1194
rect 377 1160 415 1194
rect 449 1160 487 1194
rect 521 1160 533 1194
rect 187 1148 533 1160
rect 36 1092 94 1104
rect 36 1058 48 1092
rect 82 1058 94 1092
rect 36 1020 94 1058
rect 36 986 48 1020
rect 82 986 94 1020
rect 36 948 94 986
rect 36 914 48 948
rect 82 914 94 948
rect 36 876 94 914
rect 36 842 48 876
rect 82 842 94 876
rect 36 804 94 842
rect 36 770 48 804
rect 82 770 94 804
rect 36 732 94 770
rect 36 698 48 732
rect 82 698 94 732
rect 36 660 94 698
rect 36 626 48 660
rect 82 626 94 660
rect 36 588 94 626
rect 36 554 48 588
rect 82 554 94 588
rect 36 516 94 554
rect 36 482 48 516
rect 82 482 94 516
rect 36 444 94 482
rect 36 410 48 444
rect 82 410 94 444
rect 36 372 94 410
rect 36 338 48 372
rect 82 338 94 372
rect 36 300 94 338
rect 36 266 48 300
rect 82 266 94 300
rect 36 228 94 266
rect 36 194 48 228
rect 82 194 94 228
rect 36 156 94 194
rect 36 122 48 156
rect 82 122 94 156
rect 36 110 94 122
rect 150 1092 202 1104
rect 150 1058 159 1092
rect 193 1058 202 1092
rect 150 1020 202 1058
rect 150 986 159 1020
rect 193 986 202 1020
rect 150 948 202 986
rect 150 914 159 948
rect 193 914 202 948
rect 150 876 202 914
rect 150 842 159 876
rect 193 842 202 876
rect 150 804 202 842
rect 150 770 159 804
rect 193 770 202 804
rect 150 732 202 770
rect 150 698 159 732
rect 193 698 202 732
rect 150 660 202 698
rect 150 626 159 660
rect 193 626 202 660
rect 150 588 202 626
rect 150 554 159 588
rect 193 554 202 588
rect 150 552 202 554
rect 150 488 159 500
rect 193 488 202 500
rect 150 424 159 436
rect 193 424 202 436
rect 150 360 159 372
rect 193 360 202 372
rect 150 300 202 308
rect 150 296 159 300
rect 193 296 202 300
rect 150 232 202 244
rect 150 168 202 180
rect 150 110 202 116
rect 242 1098 294 1104
rect 242 1034 294 1046
rect 242 970 294 982
rect 242 914 251 918
rect 285 914 294 918
rect 242 906 294 914
rect 242 842 251 854
rect 285 842 294 854
rect 242 778 251 790
rect 285 778 294 790
rect 242 714 251 726
rect 285 714 294 726
rect 242 660 294 662
rect 242 626 251 660
rect 285 626 294 660
rect 242 588 294 626
rect 242 554 251 588
rect 285 554 294 588
rect 242 516 294 554
rect 242 482 251 516
rect 285 482 294 516
rect 242 444 294 482
rect 242 410 251 444
rect 285 410 294 444
rect 242 372 294 410
rect 242 338 251 372
rect 285 338 294 372
rect 242 300 294 338
rect 242 266 251 300
rect 285 266 294 300
rect 242 228 294 266
rect 242 194 251 228
rect 285 194 294 228
rect 242 156 294 194
rect 242 122 251 156
rect 285 122 294 156
rect 242 110 294 122
rect 334 1092 386 1104
rect 334 1058 343 1092
rect 377 1058 386 1092
rect 334 1020 386 1058
rect 334 986 343 1020
rect 377 986 386 1020
rect 334 948 386 986
rect 334 914 343 948
rect 377 914 386 948
rect 334 876 386 914
rect 334 842 343 876
rect 377 842 386 876
rect 334 804 386 842
rect 334 770 343 804
rect 377 770 386 804
rect 334 732 386 770
rect 334 698 343 732
rect 377 698 386 732
rect 334 660 386 698
rect 334 626 343 660
rect 377 626 386 660
rect 334 588 386 626
rect 334 554 343 588
rect 377 554 386 588
rect 334 552 386 554
rect 334 488 343 500
rect 377 488 386 500
rect 334 424 343 436
rect 377 424 386 436
rect 334 360 343 372
rect 377 360 386 372
rect 334 300 386 308
rect 334 296 343 300
rect 377 296 386 300
rect 334 232 386 244
rect 334 168 386 180
rect 334 110 386 116
rect 426 1098 478 1104
rect 426 1034 478 1046
rect 426 970 478 982
rect 426 914 435 918
rect 469 914 478 918
rect 426 906 478 914
rect 426 842 435 854
rect 469 842 478 854
rect 426 778 435 790
rect 469 778 478 790
rect 426 714 435 726
rect 469 714 478 726
rect 426 660 478 662
rect 426 626 435 660
rect 469 626 478 660
rect 426 588 478 626
rect 426 554 435 588
rect 469 554 478 588
rect 426 516 478 554
rect 426 482 435 516
rect 469 482 478 516
rect 426 444 478 482
rect 426 410 435 444
rect 469 410 478 444
rect 426 372 478 410
rect 426 338 435 372
rect 469 338 478 372
rect 426 300 478 338
rect 426 266 435 300
rect 469 266 478 300
rect 426 228 478 266
rect 426 194 435 228
rect 469 194 478 228
rect 426 156 478 194
rect 426 122 435 156
rect 469 122 478 156
rect 426 110 478 122
rect 518 1092 570 1104
rect 518 1058 527 1092
rect 561 1058 570 1092
rect 518 1020 570 1058
rect 518 986 527 1020
rect 561 986 570 1020
rect 518 948 570 986
rect 518 914 527 948
rect 561 914 570 948
rect 518 876 570 914
rect 518 842 527 876
rect 561 842 570 876
rect 518 804 570 842
rect 518 770 527 804
rect 561 770 570 804
rect 518 732 570 770
rect 518 698 527 732
rect 561 698 570 732
rect 518 660 570 698
rect 518 626 527 660
rect 561 626 570 660
rect 518 588 570 626
rect 518 554 527 588
rect 561 554 570 588
rect 518 552 570 554
rect 518 488 527 500
rect 561 488 570 500
rect 518 424 527 436
rect 561 424 570 436
rect 518 360 527 372
rect 561 360 570 372
rect 518 300 570 308
rect 518 296 527 300
rect 561 296 570 300
rect 518 232 570 244
rect 518 168 570 180
rect 518 110 570 116
rect 626 1092 684 1104
rect 626 1058 638 1092
rect 672 1058 684 1092
rect 626 1020 684 1058
rect 626 986 638 1020
rect 672 986 684 1020
rect 626 948 684 986
rect 626 914 638 948
rect 672 914 684 948
rect 626 876 684 914
rect 626 842 638 876
rect 672 842 684 876
rect 626 804 684 842
rect 626 770 638 804
rect 672 770 684 804
rect 626 732 684 770
rect 626 698 638 732
rect 672 698 684 732
rect 626 660 684 698
rect 626 626 638 660
rect 672 626 684 660
rect 626 588 684 626
rect 626 554 638 588
rect 672 554 684 588
rect 626 516 684 554
rect 626 482 638 516
rect 672 482 684 516
rect 626 444 684 482
rect 626 410 638 444
rect 672 410 684 444
rect 626 372 684 410
rect 626 338 638 372
rect 672 338 684 372
rect 626 300 684 338
rect 626 266 638 300
rect 672 266 684 300
rect 626 228 684 266
rect 626 194 638 228
rect 672 194 684 228
rect 626 156 684 194
rect 626 122 638 156
rect 672 122 684 156
rect 626 110 684 122
rect 187 54 533 66
rect 187 20 199 54
rect 233 20 271 54
rect 305 20 343 54
rect 377 20 415 54
rect 449 20 487 54
rect 521 20 533 54
rect 187 0 533 20
<< via1 >>
rect 150 516 202 552
rect 150 500 159 516
rect 159 500 193 516
rect 193 500 202 516
rect 150 482 159 488
rect 159 482 193 488
rect 193 482 202 488
rect 150 444 202 482
rect 150 436 159 444
rect 159 436 193 444
rect 193 436 202 444
rect 150 410 159 424
rect 159 410 193 424
rect 193 410 202 424
rect 150 372 202 410
rect 150 338 159 360
rect 159 338 193 360
rect 193 338 202 360
rect 150 308 202 338
rect 150 266 159 296
rect 159 266 193 296
rect 193 266 202 296
rect 150 244 202 266
rect 150 228 202 232
rect 150 194 159 228
rect 159 194 193 228
rect 193 194 202 228
rect 150 180 202 194
rect 150 156 202 168
rect 150 122 159 156
rect 159 122 193 156
rect 193 122 202 156
rect 150 116 202 122
rect 242 1092 294 1098
rect 242 1058 251 1092
rect 251 1058 285 1092
rect 285 1058 294 1092
rect 242 1046 294 1058
rect 242 1020 294 1034
rect 242 986 251 1020
rect 251 986 285 1020
rect 285 986 294 1020
rect 242 982 294 986
rect 242 948 294 970
rect 242 918 251 948
rect 251 918 285 948
rect 285 918 294 948
rect 242 876 294 906
rect 242 854 251 876
rect 251 854 285 876
rect 285 854 294 876
rect 242 804 294 842
rect 242 790 251 804
rect 251 790 285 804
rect 285 790 294 804
rect 242 770 251 778
rect 251 770 285 778
rect 285 770 294 778
rect 242 732 294 770
rect 242 726 251 732
rect 251 726 285 732
rect 285 726 294 732
rect 242 698 251 714
rect 251 698 285 714
rect 285 698 294 714
rect 242 662 294 698
rect 334 516 386 552
rect 334 500 343 516
rect 343 500 377 516
rect 377 500 386 516
rect 334 482 343 488
rect 343 482 377 488
rect 377 482 386 488
rect 334 444 386 482
rect 334 436 343 444
rect 343 436 377 444
rect 377 436 386 444
rect 334 410 343 424
rect 343 410 377 424
rect 377 410 386 424
rect 334 372 386 410
rect 334 338 343 360
rect 343 338 377 360
rect 377 338 386 360
rect 334 308 386 338
rect 334 266 343 296
rect 343 266 377 296
rect 377 266 386 296
rect 334 244 386 266
rect 334 228 386 232
rect 334 194 343 228
rect 343 194 377 228
rect 377 194 386 228
rect 334 180 386 194
rect 334 156 386 168
rect 334 122 343 156
rect 343 122 377 156
rect 377 122 386 156
rect 334 116 386 122
rect 426 1092 478 1098
rect 426 1058 435 1092
rect 435 1058 469 1092
rect 469 1058 478 1092
rect 426 1046 478 1058
rect 426 1020 478 1034
rect 426 986 435 1020
rect 435 986 469 1020
rect 469 986 478 1020
rect 426 982 478 986
rect 426 948 478 970
rect 426 918 435 948
rect 435 918 469 948
rect 469 918 478 948
rect 426 876 478 906
rect 426 854 435 876
rect 435 854 469 876
rect 469 854 478 876
rect 426 804 478 842
rect 426 790 435 804
rect 435 790 469 804
rect 469 790 478 804
rect 426 770 435 778
rect 435 770 469 778
rect 469 770 478 778
rect 426 732 478 770
rect 426 726 435 732
rect 435 726 469 732
rect 469 726 478 732
rect 426 698 435 714
rect 435 698 469 714
rect 469 698 478 714
rect 426 662 478 698
rect 518 516 570 552
rect 518 500 527 516
rect 527 500 561 516
rect 561 500 570 516
rect 518 482 527 488
rect 527 482 561 488
rect 561 482 570 488
rect 518 444 570 482
rect 518 436 527 444
rect 527 436 561 444
rect 561 436 570 444
rect 518 410 527 424
rect 527 410 561 424
rect 561 410 570 424
rect 518 372 570 410
rect 518 338 527 360
rect 527 338 561 360
rect 561 338 570 360
rect 518 308 570 338
rect 518 266 527 296
rect 527 266 561 296
rect 561 266 570 296
rect 518 244 570 266
rect 518 228 570 232
rect 518 194 527 228
rect 527 194 561 228
rect 561 194 570 228
rect 518 180 570 194
rect 518 156 570 168
rect 518 122 527 156
rect 527 122 561 156
rect 561 122 570 156
rect 518 116 570 122
<< metal2 >>
rect 10 1098 710 1104
rect 10 1046 242 1098
rect 294 1046 426 1098
rect 478 1046 710 1098
rect 10 1034 710 1046
rect 10 982 242 1034
rect 294 982 426 1034
rect 478 982 710 1034
rect 10 970 710 982
rect 10 918 242 970
rect 294 918 426 970
rect 478 918 710 970
rect 10 906 710 918
rect 10 854 242 906
rect 294 854 426 906
rect 478 854 710 906
rect 10 842 710 854
rect 10 790 242 842
rect 294 790 426 842
rect 478 790 710 842
rect 10 778 710 790
rect 10 726 242 778
rect 294 726 426 778
rect 478 726 710 778
rect 10 714 710 726
rect 10 662 242 714
rect 294 662 426 714
rect 478 662 710 714
rect 10 632 710 662
rect 10 552 710 582
rect 10 500 150 552
rect 202 500 334 552
rect 386 500 518 552
rect 570 500 710 552
rect 10 488 710 500
rect 10 436 150 488
rect 202 436 334 488
rect 386 436 518 488
rect 570 436 710 488
rect 10 424 710 436
rect 10 372 150 424
rect 202 372 334 424
rect 386 372 518 424
rect 570 372 710 424
rect 10 360 710 372
rect 10 308 150 360
rect 202 308 334 360
rect 386 308 518 360
rect 570 308 710 360
rect 10 296 710 308
rect 10 244 150 296
rect 202 244 334 296
rect 386 244 518 296
rect 570 244 710 296
rect 10 232 710 244
rect 10 180 150 232
rect 202 180 334 232
rect 386 180 518 232
rect 570 180 710 232
rect 10 168 710 180
rect 10 116 150 168
rect 202 116 334 168
rect 386 116 518 168
rect 570 116 710 168
rect 10 110 710 116
<< labels >>
flabel comment s 176 607 176 607 0 FreeSans 300 0 0 0 S
flabel comment s 176 607 176 607 0 FreeSans 300 0 0 0 S
flabel comment s 268 607 268 607 0 FreeSans 300 0 0 0 S
flabel comment s 268 607 268 607 0 FreeSans 300 0 0 0 D
flabel comment s 360 607 360 607 0 FreeSans 300 0 0 0 S
flabel comment s 360 607 360 607 0 FreeSans 300 0 0 0 S
flabel comment s 452 607 452 607 0 FreeSans 300 0 0 0 S
flabel comment s 452 607 452 607 0 FreeSans 300 0 0 0 D
flabel comment s 544 607 544 607 0 FreeSans 300 0 0 0 S
flabel metal1 s 48 610 82 621 0 FreeSans 100 0 0 0 BULK
port 1 nsew
flabel metal1 s 339 1167 397 1192 0 FreeSans 100 0 0 0 GATE
port 3 nsew
flabel metal1 s 335 24 393 49 0 FreeSans 100 0 0 0 GATE
port 3 nsew
flabel metal1 s 636 612 670 623 0 FreeSans 100 0 0 0 BULK
port 1 nsew
flabel metal2 s 56 886 71 952 0 FreeSans 100 0 0 0 DRAIN
port 2 nsew
flabel metal2 s 59 312 73 375 0 FreeSans 100 0 0 0 SOURCE
port 4 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 9582762
string GDS_START 9560732
<< end >>
