magic
tech sky130A
magscale 1 2
timestamp 1658881652
<< error_s >>
rect 15 254 28 270
rect 83 254 98 268
rect 117 256 130 270
rect 198 266 351 312
rect 180 254 372 266
rect 451 254 464 270
rect 546 254 565 270
rect 580 254 586 270
rect 595 254 608 270
rect 663 254 678 268
rect 697 256 710 270
rect 778 266 931 312
rect 760 254 952 266
rect 1031 254 1044 270
rect 1126 254 1145 270
rect 1160 254 1166 270
rect 1175 254 1188 270
rect 1243 254 1258 268
rect 1277 256 1290 270
rect 1358 266 1511 312
rect 1340 254 1532 266
rect 1611 254 1624 270
rect 1706 254 1725 270
rect 1740 254 1746 270
rect 1755 254 1768 270
rect 1823 254 1838 268
rect 1857 256 1870 270
rect 1938 266 2091 312
rect 1920 254 2112 266
rect 2191 254 2204 270
rect 2286 254 2305 270
rect 2320 254 2326 270
rect 2335 254 2348 270
rect 2403 254 2418 268
rect 2437 256 2450 270
rect 2518 266 2671 312
rect 2500 254 2692 266
rect 2771 254 2784 270
rect 2866 254 2885 270
rect 2900 254 2906 270
rect 2915 254 2928 270
rect 2983 254 2998 268
rect 3017 256 3030 270
rect 3098 266 3251 312
rect 3080 254 3272 266
rect 3351 254 3364 270
rect 3446 254 3465 270
rect 3480 254 3486 270
rect 3495 254 3508 270
rect 3563 254 3578 268
rect 3597 256 3610 270
rect 3678 266 3831 312
rect 3660 254 3852 266
rect 3931 254 3944 270
rect 4026 254 4045 270
rect 4060 254 4066 270
rect 4075 254 4088 270
rect 4143 254 4158 268
rect 4177 256 4190 270
rect 4258 266 4411 312
rect 4240 254 4432 266
rect 4511 254 4524 270
rect 4612 254 4625 270
rect 0 240 4625 254
rect 15 170 28 240
rect 73 214 102 228
rect 155 214 171 228
rect 209 218 215 226
rect 222 224 330 240
rect 73 212 171 214
rect 57 204 108 212
rect 155 204 189 212
rect 57 192 82 204
rect 89 192 108 204
rect 162 202 189 204
rect 198 204 215 218
rect 260 204 292 224
rect 337 218 343 226
rect 351 218 366 240
rect 432 234 451 237
rect 337 212 366 218
rect 381 214 397 228
rect 432 215 454 234
rect 464 228 480 229
rect 463 226 480 228
rect 464 221 480 226
rect 454 214 460 215
rect 463 214 492 221
rect 381 213 492 214
rect 381 212 498 213
rect 337 204 419 212
rect 454 209 460 212
rect 198 202 419 204
rect 162 198 234 202
rect 262 200 290 202
rect 315 198 419 202
rect 57 184 108 192
rect 155 190 287 198
rect 290 190 419 198
rect 463 204 498 212
rect 155 188 234 190
rect 315 188 419 190
rect 155 184 252 188
rect 9 136 28 170
rect 73 176 102 184
rect 73 170 90 176
rect 73 168 107 170
rect 155 168 171 184
rect 172 180 252 184
rect 300 184 419 188
rect 300 180 380 184
rect 172 174 380 180
rect 381 174 397 184
rect 445 180 460 195
rect 463 192 464 204
rect 471 192 498 204
rect 463 184 498 192
rect 463 183 492 184
rect 183 170 287 174
rect 74 164 107 168
rect 70 162 107 164
rect 70 161 137 162
rect 70 156 101 161
rect 107 156 137 161
rect 198 158 213 170
rect 70 152 137 156
rect 43 149 137 152
rect 43 142 92 149
rect 43 136 73 142
rect 92 137 97 142
rect 9 120 89 136
rect 101 128 137 149
rect 222 148 252 157
rect 275 152 293 170
rect 351 168 397 174
rect 432 170 445 180
rect 463 170 480 183
rect 432 168 480 170
rect 313 162 315 164
rect 315 157 327 162
rect 300 150 330 157
rect 300 148 331 150
rect 351 148 387 168
rect 432 167 479 168
rect 445 162 479 167
rect 198 144 387 148
rect 213 141 387 144
rect 206 138 387 141
rect 415 161 479 162
rect 9 118 28 120
rect 43 118 77 120
rect 9 102 89 118
rect 9 96 28 102
rect -1 80 28 96
rect 43 86 73 102
rect 101 80 107 128
rect 110 122 129 128
rect 144 122 174 130
rect 110 114 174 122
rect 110 98 190 114
rect 206 107 268 138
rect 284 107 346 138
rect 415 136 464 161
rect 479 136 509 152
rect 378 122 408 130
rect 415 128 525 136
rect 378 114 423 122
rect 110 96 129 98
rect 144 96 190 98
rect 110 80 190 96
rect 217 94 252 107
rect 293 104 330 107
rect 293 102 335 104
rect 222 91 252 94
rect 231 87 238 91
rect 238 86 239 87
rect 197 80 207 86
rect -7 72 34 80
rect -7 46 8 72
rect 15 46 34 72
rect 98 68 129 80
rect 144 68 247 80
rect 259 70 285 96
rect 300 91 330 102
rect 362 98 424 114
rect 362 96 408 98
rect 362 80 424 96
rect 436 80 442 128
rect 445 120 525 128
rect 445 118 464 120
rect 479 118 513 120
rect 445 102 525 118
rect 445 80 464 102
rect 479 86 509 102
rect 537 96 543 170
rect 546 96 565 240
rect 580 96 586 240
rect 595 170 608 240
rect 653 214 682 228
rect 735 214 751 228
rect 789 218 795 226
rect 802 224 910 240
rect 653 212 751 214
rect 637 204 688 212
rect 735 204 769 212
rect 637 192 662 204
rect 669 192 688 204
rect 742 202 769 204
rect 778 204 795 218
rect 840 204 872 224
rect 917 218 923 226
rect 931 218 946 240
rect 1012 234 1031 237
rect 917 212 946 218
rect 961 214 977 228
rect 1012 215 1034 234
rect 1044 228 1060 229
rect 1043 226 1060 228
rect 1044 221 1060 226
rect 1034 214 1040 215
rect 1043 214 1072 221
rect 961 213 1072 214
rect 961 212 1078 213
rect 917 204 999 212
rect 1034 209 1040 212
rect 778 202 999 204
rect 742 198 814 202
rect 842 200 870 202
rect 895 198 999 202
rect 637 184 688 192
rect 735 190 867 198
rect 870 190 999 198
rect 1043 204 1078 212
rect 735 188 814 190
rect 895 188 999 190
rect 735 184 832 188
rect 589 136 608 170
rect 653 176 682 184
rect 653 170 670 176
rect 653 168 687 170
rect 735 168 751 184
rect 752 180 832 184
rect 880 184 999 188
rect 880 180 960 184
rect 752 174 960 180
rect 961 174 977 184
rect 1025 180 1040 195
rect 1043 192 1044 204
rect 1051 192 1078 204
rect 1043 184 1078 192
rect 1043 183 1072 184
rect 763 170 867 174
rect 654 164 687 168
rect 650 162 687 164
rect 650 161 717 162
rect 650 156 681 161
rect 687 156 717 161
rect 778 158 793 170
rect 650 152 717 156
rect 623 149 717 152
rect 623 142 672 149
rect 623 136 653 142
rect 672 137 677 142
rect 589 120 669 136
rect 681 128 717 149
rect 802 148 832 157
rect 855 152 873 170
rect 931 168 977 174
rect 1012 170 1025 180
rect 1043 170 1060 183
rect 1012 168 1060 170
rect 893 162 895 164
rect 895 157 907 162
rect 880 150 910 157
rect 880 148 911 150
rect 931 148 967 168
rect 1012 167 1059 168
rect 1025 162 1059 167
rect 778 144 967 148
rect 793 141 967 144
rect 786 138 967 141
rect 995 161 1059 162
rect 589 118 608 120
rect 623 118 657 120
rect 589 102 669 118
rect 589 96 608 102
rect 305 70 408 80
rect 259 68 408 70
rect 429 68 464 80
rect 98 66 260 68
rect 110 46 129 66
rect 144 64 174 66
rect -7 38 34 46
rect -1 28 28 38
rect 116 28 129 46
rect 181 50 260 66
rect 292 66 464 68
rect 292 50 371 66
rect 378 64 408 66
rect 181 42 371 50
rect 436 46 442 66
rect 181 38 260 42
rect 262 38 290 42
rect 292 38 371 42
rect 166 28 174 38
rect 193 30 196 38
rect 197 30 215 38
rect 260 30 292 38
rect 337 30 355 38
rect 193 28 359 30
rect 378 28 389 38
rect 451 28 464 66
rect 536 80 565 96
rect 579 80 608 96
rect 623 86 653 102
rect 681 80 687 128
rect 690 122 709 128
rect 724 122 754 130
rect 690 114 754 122
rect 690 98 770 114
rect 786 107 848 138
rect 864 107 926 138
rect 995 136 1044 161
rect 1059 136 1089 152
rect 958 122 988 130
rect 995 128 1105 136
rect 958 114 1003 122
rect 690 96 709 98
rect 724 96 770 98
rect 690 80 770 96
rect 797 94 832 107
rect 873 104 910 107
rect 873 102 915 104
rect 802 91 832 94
rect 811 87 818 91
rect 818 86 819 87
rect 777 80 787 86
rect 536 72 571 80
rect 536 46 537 72
rect 544 46 571 72
rect 536 38 571 46
rect 573 72 614 80
rect 573 46 588 72
rect 595 46 614 72
rect 678 68 709 80
rect 724 68 827 80
rect 839 70 865 96
rect 880 91 910 102
rect 942 98 1004 114
rect 942 96 988 98
rect 942 80 1004 96
rect 1016 80 1022 128
rect 1025 120 1105 128
rect 1025 118 1044 120
rect 1059 118 1093 120
rect 1025 102 1105 118
rect 1025 80 1044 102
rect 1059 86 1089 102
rect 1117 96 1123 170
rect 1126 96 1145 240
rect 1160 96 1166 240
rect 1175 170 1188 240
rect 1233 214 1262 228
rect 1315 214 1331 228
rect 1369 218 1375 226
rect 1382 224 1490 240
rect 1233 212 1331 214
rect 1217 204 1268 212
rect 1315 204 1349 212
rect 1217 192 1242 204
rect 1249 192 1268 204
rect 1322 202 1349 204
rect 1358 204 1375 218
rect 1420 204 1452 224
rect 1497 218 1503 226
rect 1511 218 1526 240
rect 1592 234 1611 237
rect 1497 212 1526 218
rect 1541 214 1557 228
rect 1592 215 1614 234
rect 1624 228 1640 229
rect 1623 226 1640 228
rect 1624 221 1640 226
rect 1614 214 1620 215
rect 1623 214 1652 221
rect 1541 213 1652 214
rect 1541 212 1658 213
rect 1497 204 1579 212
rect 1614 209 1620 212
rect 1358 202 1579 204
rect 1322 198 1394 202
rect 1422 200 1450 202
rect 1475 198 1579 202
rect 1217 184 1268 192
rect 1315 190 1447 198
rect 1450 190 1579 198
rect 1623 204 1658 212
rect 1315 188 1394 190
rect 1475 188 1579 190
rect 1315 184 1412 188
rect 1169 136 1188 170
rect 1233 176 1262 184
rect 1233 170 1250 176
rect 1233 168 1267 170
rect 1315 168 1331 184
rect 1332 180 1412 184
rect 1460 184 1579 188
rect 1460 180 1540 184
rect 1332 174 1540 180
rect 1541 174 1557 184
rect 1605 180 1620 195
rect 1623 192 1624 204
rect 1631 192 1658 204
rect 1623 184 1658 192
rect 1623 183 1652 184
rect 1343 170 1447 174
rect 1234 164 1267 168
rect 1230 162 1267 164
rect 1230 161 1297 162
rect 1230 156 1261 161
rect 1267 156 1297 161
rect 1358 158 1373 170
rect 1230 152 1297 156
rect 1203 149 1297 152
rect 1203 142 1252 149
rect 1203 136 1233 142
rect 1252 137 1257 142
rect 1169 120 1249 136
rect 1261 128 1297 149
rect 1382 148 1412 157
rect 1435 152 1453 170
rect 1511 168 1557 174
rect 1592 170 1605 180
rect 1623 170 1640 183
rect 1592 168 1640 170
rect 1473 162 1475 164
rect 1475 157 1487 162
rect 1460 150 1490 157
rect 1460 148 1491 150
rect 1511 148 1547 168
rect 1592 167 1639 168
rect 1605 162 1639 167
rect 1358 144 1547 148
rect 1373 141 1547 144
rect 1366 138 1547 141
rect 1575 161 1639 162
rect 1169 118 1188 120
rect 1203 118 1237 120
rect 1169 102 1249 118
rect 1169 96 1188 102
rect 885 70 988 80
rect 839 68 988 70
rect 1009 68 1044 80
rect 678 66 840 68
rect 690 46 709 66
rect 724 64 754 66
rect 573 38 614 46
rect 536 28 565 38
rect 579 28 608 38
rect 696 28 709 46
rect 761 50 840 66
rect 872 66 1044 68
rect 872 50 951 66
rect 958 64 988 66
rect 761 42 951 50
rect 1016 46 1022 66
rect 761 38 840 42
rect 842 38 870 42
rect 872 38 951 42
rect 746 28 754 38
rect 773 30 776 38
rect 777 30 795 38
rect 840 30 872 38
rect 917 30 935 38
rect 773 28 939 30
rect 958 28 969 38
rect 1031 28 1044 66
rect 1116 80 1145 96
rect 1159 80 1188 96
rect 1203 86 1233 102
rect 1261 80 1267 128
rect 1270 122 1289 128
rect 1304 122 1334 130
rect 1270 114 1334 122
rect 1270 98 1350 114
rect 1366 107 1428 138
rect 1444 107 1506 138
rect 1575 136 1624 161
rect 1639 136 1669 152
rect 1538 122 1568 130
rect 1575 128 1685 136
rect 1538 114 1583 122
rect 1270 96 1289 98
rect 1304 96 1350 98
rect 1270 80 1350 96
rect 1377 94 1412 107
rect 1453 104 1490 107
rect 1453 102 1495 104
rect 1382 91 1412 94
rect 1391 87 1398 91
rect 1398 86 1399 87
rect 1357 80 1367 86
rect 1116 72 1151 80
rect 1116 46 1117 72
rect 1124 46 1151 72
rect 1116 38 1151 46
rect 1153 72 1194 80
rect 1153 46 1168 72
rect 1175 46 1194 72
rect 1258 68 1289 80
rect 1304 68 1407 80
rect 1419 70 1445 96
rect 1460 91 1490 102
rect 1522 98 1584 114
rect 1522 96 1568 98
rect 1522 80 1584 96
rect 1596 80 1602 128
rect 1605 120 1685 128
rect 1605 118 1624 120
rect 1639 118 1673 120
rect 1605 102 1685 118
rect 1605 80 1624 102
rect 1639 86 1669 102
rect 1697 96 1703 170
rect 1706 96 1725 240
rect 1740 96 1746 240
rect 1755 170 1768 240
rect 1813 214 1842 228
rect 1895 214 1911 228
rect 1949 218 1955 226
rect 1962 224 2070 240
rect 1813 212 1911 214
rect 1797 204 1848 212
rect 1895 204 1929 212
rect 1797 192 1822 204
rect 1829 192 1848 204
rect 1902 202 1929 204
rect 1938 204 1955 218
rect 2000 204 2032 224
rect 2077 218 2083 226
rect 2091 218 2106 240
rect 2172 234 2191 237
rect 2077 212 2106 218
rect 2121 214 2137 228
rect 2172 215 2194 234
rect 2204 228 2220 229
rect 2203 226 2220 228
rect 2204 221 2220 226
rect 2194 214 2200 215
rect 2203 214 2232 221
rect 2121 213 2232 214
rect 2121 212 2238 213
rect 2077 204 2159 212
rect 2194 209 2200 212
rect 1938 202 2159 204
rect 1902 198 1974 202
rect 2002 200 2030 202
rect 2055 198 2159 202
rect 1797 184 1848 192
rect 1895 190 2027 198
rect 2030 190 2159 198
rect 2203 204 2238 212
rect 1895 188 1974 190
rect 2055 188 2159 190
rect 1895 184 1992 188
rect 1749 136 1768 170
rect 1813 176 1842 184
rect 1813 170 1830 176
rect 1813 168 1847 170
rect 1895 168 1911 184
rect 1912 180 1992 184
rect 2040 184 2159 188
rect 2040 180 2120 184
rect 1912 174 2120 180
rect 2121 174 2137 184
rect 2185 180 2200 195
rect 2203 192 2204 204
rect 2211 192 2238 204
rect 2203 184 2238 192
rect 2203 183 2232 184
rect 1923 170 2027 174
rect 1814 164 1847 168
rect 1810 162 1847 164
rect 1810 161 1877 162
rect 1810 156 1841 161
rect 1847 156 1877 161
rect 1938 158 1953 170
rect 1810 152 1877 156
rect 1783 149 1877 152
rect 1783 142 1832 149
rect 1783 136 1813 142
rect 1832 137 1837 142
rect 1749 120 1829 136
rect 1841 128 1877 149
rect 1962 148 1992 157
rect 2015 152 2033 170
rect 2091 168 2137 174
rect 2172 170 2185 180
rect 2203 170 2220 183
rect 2172 168 2220 170
rect 2053 162 2055 164
rect 2055 157 2067 162
rect 2040 150 2070 157
rect 2040 148 2071 150
rect 2091 148 2127 168
rect 2172 167 2219 168
rect 2185 162 2219 167
rect 1938 144 2127 148
rect 1953 141 2127 144
rect 1946 138 2127 141
rect 2155 161 2219 162
rect 1749 118 1768 120
rect 1783 118 1817 120
rect 1749 102 1829 118
rect 1749 96 1768 102
rect 1465 70 1568 80
rect 1419 68 1568 70
rect 1589 68 1624 80
rect 1258 66 1420 68
rect 1270 46 1289 66
rect 1304 64 1334 66
rect 1153 38 1194 46
rect 1116 28 1145 38
rect 1159 28 1188 38
rect 1276 28 1289 46
rect 1341 50 1420 66
rect 1452 66 1624 68
rect 1452 50 1531 66
rect 1538 64 1568 66
rect 1341 42 1531 50
rect 1596 46 1602 66
rect 1341 38 1420 42
rect 1422 38 1450 42
rect 1452 38 1531 42
rect 1326 28 1334 38
rect 1353 30 1356 38
rect 1357 30 1375 38
rect 1420 30 1452 38
rect 1497 30 1515 38
rect 1353 28 1519 30
rect 1538 28 1549 38
rect 1611 28 1624 66
rect 1696 80 1725 96
rect 1739 80 1768 96
rect 1783 86 1813 102
rect 1841 80 1847 128
rect 1850 122 1869 128
rect 1884 122 1914 130
rect 1850 114 1914 122
rect 1850 98 1930 114
rect 1946 107 2008 138
rect 2024 107 2086 138
rect 2155 136 2204 161
rect 2219 136 2249 152
rect 2118 122 2148 130
rect 2155 128 2265 136
rect 2118 114 2163 122
rect 1850 96 1869 98
rect 1884 96 1930 98
rect 1850 80 1930 96
rect 1957 94 1992 107
rect 2033 104 2070 107
rect 2033 102 2075 104
rect 1962 91 1992 94
rect 1971 87 1978 91
rect 1978 86 1979 87
rect 1937 80 1947 86
rect 1696 72 1731 80
rect 1696 46 1697 72
rect 1704 46 1731 72
rect 1696 38 1731 46
rect 1733 72 1774 80
rect 1733 46 1748 72
rect 1755 46 1774 72
rect 1838 68 1869 80
rect 1884 68 1987 80
rect 1999 70 2025 96
rect 2040 91 2070 102
rect 2102 98 2164 114
rect 2102 96 2148 98
rect 2102 80 2164 96
rect 2176 80 2182 128
rect 2185 120 2265 128
rect 2185 118 2204 120
rect 2219 118 2253 120
rect 2185 102 2265 118
rect 2185 80 2204 102
rect 2219 86 2249 102
rect 2277 96 2283 170
rect 2286 96 2305 240
rect 2320 96 2326 240
rect 2335 170 2348 240
rect 2393 214 2422 228
rect 2475 214 2491 228
rect 2529 218 2535 226
rect 2542 224 2650 240
rect 2393 212 2491 214
rect 2377 204 2428 212
rect 2475 204 2509 212
rect 2377 192 2402 204
rect 2409 192 2428 204
rect 2482 202 2509 204
rect 2518 204 2535 218
rect 2580 204 2612 224
rect 2657 218 2663 226
rect 2671 218 2686 240
rect 2752 234 2771 237
rect 2657 212 2686 218
rect 2701 214 2717 228
rect 2752 215 2774 234
rect 2784 228 2800 229
rect 2783 226 2800 228
rect 2784 221 2800 226
rect 2774 214 2780 215
rect 2783 214 2812 221
rect 2701 213 2812 214
rect 2701 212 2818 213
rect 2657 204 2739 212
rect 2774 209 2780 212
rect 2518 202 2739 204
rect 2482 198 2554 202
rect 2582 200 2610 202
rect 2635 198 2739 202
rect 2377 184 2428 192
rect 2475 190 2607 198
rect 2610 190 2739 198
rect 2783 204 2818 212
rect 2475 188 2554 190
rect 2635 188 2739 190
rect 2475 184 2572 188
rect 2329 136 2348 170
rect 2393 176 2422 184
rect 2393 170 2410 176
rect 2393 168 2427 170
rect 2475 168 2491 184
rect 2492 180 2572 184
rect 2620 184 2739 188
rect 2620 180 2700 184
rect 2492 174 2700 180
rect 2701 174 2717 184
rect 2765 180 2780 195
rect 2783 192 2784 204
rect 2791 192 2818 204
rect 2783 184 2818 192
rect 2783 183 2812 184
rect 2503 170 2607 174
rect 2394 164 2427 168
rect 2390 162 2427 164
rect 2390 161 2457 162
rect 2390 156 2421 161
rect 2427 156 2457 161
rect 2518 158 2533 170
rect 2390 152 2457 156
rect 2363 149 2457 152
rect 2363 142 2412 149
rect 2363 136 2393 142
rect 2412 137 2417 142
rect 2329 120 2409 136
rect 2421 128 2457 149
rect 2542 148 2572 157
rect 2595 152 2613 170
rect 2671 168 2717 174
rect 2752 170 2765 180
rect 2783 170 2800 183
rect 2752 168 2800 170
rect 2633 162 2635 164
rect 2635 157 2647 162
rect 2620 150 2650 157
rect 2620 148 2651 150
rect 2671 148 2707 168
rect 2752 167 2799 168
rect 2765 162 2799 167
rect 2518 144 2707 148
rect 2533 141 2707 144
rect 2526 138 2707 141
rect 2735 161 2799 162
rect 2329 118 2348 120
rect 2363 118 2397 120
rect 2329 102 2409 118
rect 2329 96 2348 102
rect 2045 70 2148 80
rect 1999 68 2148 70
rect 2169 68 2204 80
rect 1838 66 2000 68
rect 1850 46 1869 66
rect 1884 64 1914 66
rect 1733 38 1774 46
rect 1696 28 1725 38
rect 1739 28 1768 38
rect 1856 28 1869 46
rect 1921 50 2000 66
rect 2032 66 2204 68
rect 2032 50 2111 66
rect 2118 64 2148 66
rect 1921 42 2111 50
rect 2176 46 2182 66
rect 1921 38 2000 42
rect 2002 38 2030 42
rect 2032 38 2111 42
rect 1906 28 1914 38
rect 1933 30 1936 38
rect 1937 30 1955 38
rect 2000 30 2032 38
rect 2077 30 2095 38
rect 1933 28 2099 30
rect 2118 28 2129 38
rect 2191 28 2204 66
rect 2276 80 2305 96
rect 2319 80 2348 96
rect 2363 86 2393 102
rect 2421 80 2427 128
rect 2430 122 2449 128
rect 2464 122 2494 130
rect 2430 114 2494 122
rect 2430 98 2510 114
rect 2526 107 2588 138
rect 2604 107 2666 138
rect 2735 136 2784 161
rect 2799 136 2829 152
rect 2698 122 2728 130
rect 2735 128 2845 136
rect 2698 114 2743 122
rect 2430 96 2449 98
rect 2464 96 2510 98
rect 2430 80 2510 96
rect 2537 94 2572 107
rect 2613 104 2650 107
rect 2613 102 2655 104
rect 2542 91 2572 94
rect 2551 87 2558 91
rect 2558 86 2559 87
rect 2517 80 2527 86
rect 2276 72 2311 80
rect 2276 46 2277 72
rect 2284 46 2311 72
rect 2276 38 2311 46
rect 2313 72 2354 80
rect 2313 46 2328 72
rect 2335 46 2354 72
rect 2418 68 2449 80
rect 2464 68 2567 80
rect 2579 70 2605 96
rect 2620 91 2650 102
rect 2682 98 2744 114
rect 2682 96 2728 98
rect 2682 80 2744 96
rect 2756 80 2762 128
rect 2765 120 2845 128
rect 2765 118 2784 120
rect 2799 118 2833 120
rect 2765 102 2845 118
rect 2765 80 2784 102
rect 2799 86 2829 102
rect 2857 96 2863 170
rect 2866 96 2885 240
rect 2900 96 2906 240
rect 2915 170 2928 240
rect 2973 214 3002 228
rect 3055 214 3071 228
rect 3109 218 3115 226
rect 3122 224 3230 240
rect 2973 212 3071 214
rect 2957 204 3008 212
rect 3055 204 3089 212
rect 2957 192 2982 204
rect 2989 192 3008 204
rect 3062 202 3089 204
rect 3098 204 3115 218
rect 3160 204 3192 224
rect 3237 218 3243 226
rect 3251 218 3266 240
rect 3332 234 3351 237
rect 3237 212 3266 218
rect 3281 214 3297 228
rect 3332 215 3354 234
rect 3364 228 3380 229
rect 3363 226 3380 228
rect 3364 221 3380 226
rect 3354 214 3360 215
rect 3363 214 3392 221
rect 3281 213 3392 214
rect 3281 212 3398 213
rect 3237 204 3319 212
rect 3354 209 3360 212
rect 3098 202 3319 204
rect 3062 198 3134 202
rect 3162 200 3190 202
rect 3215 198 3319 202
rect 2957 184 3008 192
rect 3055 190 3187 198
rect 3190 190 3319 198
rect 3363 204 3398 212
rect 3055 188 3134 190
rect 3215 188 3319 190
rect 3055 184 3152 188
rect 2909 136 2928 170
rect 2973 176 3002 184
rect 2973 170 2990 176
rect 2973 168 3007 170
rect 3055 168 3071 184
rect 3072 180 3152 184
rect 3200 184 3319 188
rect 3200 180 3280 184
rect 3072 174 3280 180
rect 3281 174 3297 184
rect 3345 180 3360 195
rect 3363 192 3364 204
rect 3371 192 3398 204
rect 3363 184 3398 192
rect 3363 183 3392 184
rect 3083 170 3187 174
rect 2974 164 3007 168
rect 2970 162 3007 164
rect 2970 161 3037 162
rect 2970 156 3001 161
rect 3007 156 3037 161
rect 3098 158 3113 170
rect 2970 152 3037 156
rect 2943 149 3037 152
rect 2943 142 2992 149
rect 2943 136 2973 142
rect 2992 137 2997 142
rect 2909 120 2989 136
rect 3001 128 3037 149
rect 3122 148 3152 157
rect 3175 152 3193 170
rect 3251 168 3297 174
rect 3332 170 3345 180
rect 3363 170 3380 183
rect 3332 168 3380 170
rect 3213 162 3215 164
rect 3215 157 3227 162
rect 3200 150 3230 157
rect 3200 148 3231 150
rect 3251 148 3287 168
rect 3332 167 3379 168
rect 3345 162 3379 167
rect 3098 144 3287 148
rect 3113 141 3287 144
rect 3106 138 3287 141
rect 3315 161 3379 162
rect 2909 118 2928 120
rect 2943 118 2977 120
rect 2909 102 2989 118
rect 2909 96 2928 102
rect 2625 70 2728 80
rect 2579 68 2728 70
rect 2749 68 2784 80
rect 2418 66 2580 68
rect 2430 46 2449 66
rect 2464 64 2494 66
rect 2313 38 2354 46
rect 2276 28 2305 38
rect 2319 28 2348 38
rect 2436 28 2449 46
rect 2501 50 2580 66
rect 2612 66 2784 68
rect 2612 50 2691 66
rect 2698 64 2728 66
rect 2501 42 2691 50
rect 2756 46 2762 66
rect 2501 38 2580 42
rect 2582 38 2610 42
rect 2612 38 2691 42
rect 2486 28 2494 38
rect 2513 30 2516 38
rect 2517 30 2535 38
rect 2580 30 2612 38
rect 2657 30 2675 38
rect 2513 28 2679 30
rect 2698 28 2709 38
rect 2771 28 2784 66
rect 2856 80 2885 96
rect 2899 80 2928 96
rect 2943 86 2973 102
rect 3001 80 3007 128
rect 3010 122 3029 128
rect 3044 122 3074 130
rect 3010 114 3074 122
rect 3010 98 3090 114
rect 3106 107 3168 138
rect 3184 107 3246 138
rect 3315 136 3364 161
rect 3379 136 3409 152
rect 3278 122 3308 130
rect 3315 128 3425 136
rect 3278 114 3323 122
rect 3010 96 3029 98
rect 3044 96 3090 98
rect 3010 80 3090 96
rect 3117 94 3152 107
rect 3193 104 3230 107
rect 3193 102 3235 104
rect 3122 91 3152 94
rect 3131 87 3138 91
rect 3138 86 3139 87
rect 3097 80 3107 86
rect 2856 72 2891 80
rect 2856 46 2857 72
rect 2864 46 2891 72
rect 2856 38 2891 46
rect 2893 72 2934 80
rect 2893 46 2908 72
rect 2915 46 2934 72
rect 2998 68 3029 80
rect 3044 68 3147 80
rect 3159 70 3185 96
rect 3200 91 3230 102
rect 3262 98 3324 114
rect 3262 96 3308 98
rect 3262 80 3324 96
rect 3336 80 3342 128
rect 3345 120 3425 128
rect 3345 118 3364 120
rect 3379 118 3413 120
rect 3345 102 3425 118
rect 3345 80 3364 102
rect 3379 86 3409 102
rect 3437 96 3443 170
rect 3446 96 3465 240
rect 3480 96 3486 240
rect 3495 170 3508 240
rect 3553 214 3582 228
rect 3635 214 3651 228
rect 3689 218 3695 226
rect 3702 224 3810 240
rect 3553 212 3651 214
rect 3537 204 3588 212
rect 3635 204 3669 212
rect 3537 192 3562 204
rect 3569 192 3588 204
rect 3642 202 3669 204
rect 3678 204 3695 218
rect 3740 204 3772 224
rect 3817 218 3823 226
rect 3831 218 3846 240
rect 3912 234 3931 237
rect 3817 212 3846 218
rect 3861 214 3877 228
rect 3912 215 3934 234
rect 3944 228 3960 229
rect 3943 226 3960 228
rect 3944 221 3960 226
rect 3934 214 3940 215
rect 3943 214 3972 221
rect 3861 213 3972 214
rect 3861 212 3978 213
rect 3817 204 3899 212
rect 3934 209 3940 212
rect 3678 202 3899 204
rect 3642 198 3714 202
rect 3742 200 3770 202
rect 3795 198 3899 202
rect 3537 184 3588 192
rect 3635 190 3767 198
rect 3770 190 3899 198
rect 3943 204 3978 212
rect 3635 188 3714 190
rect 3795 188 3899 190
rect 3635 184 3732 188
rect 3489 136 3508 170
rect 3553 176 3582 184
rect 3553 170 3570 176
rect 3553 168 3587 170
rect 3635 168 3651 184
rect 3652 180 3732 184
rect 3780 184 3899 188
rect 3780 180 3860 184
rect 3652 174 3860 180
rect 3861 174 3877 184
rect 3925 180 3940 195
rect 3943 192 3944 204
rect 3951 192 3978 204
rect 3943 184 3978 192
rect 3943 183 3972 184
rect 3663 170 3767 174
rect 3554 164 3587 168
rect 3550 162 3587 164
rect 3550 161 3617 162
rect 3550 156 3581 161
rect 3587 156 3617 161
rect 3678 158 3693 170
rect 3550 152 3617 156
rect 3523 149 3617 152
rect 3523 142 3572 149
rect 3523 136 3553 142
rect 3572 137 3577 142
rect 3489 120 3569 136
rect 3581 128 3617 149
rect 3702 148 3732 157
rect 3755 152 3773 170
rect 3831 168 3877 174
rect 3912 170 3925 180
rect 3943 170 3960 183
rect 3912 168 3960 170
rect 3793 162 3795 164
rect 3795 157 3807 162
rect 3780 150 3810 157
rect 3780 148 3811 150
rect 3831 148 3867 168
rect 3912 167 3959 168
rect 3925 162 3959 167
rect 3678 144 3867 148
rect 3693 141 3867 144
rect 3686 138 3867 141
rect 3895 161 3959 162
rect 3489 118 3508 120
rect 3523 118 3557 120
rect 3489 102 3569 118
rect 3489 96 3508 102
rect 3205 70 3308 80
rect 3159 68 3308 70
rect 3329 68 3364 80
rect 2998 66 3160 68
rect 3010 46 3029 66
rect 3044 64 3074 66
rect 2893 38 2934 46
rect 2856 28 2885 38
rect 2899 28 2928 38
rect 3016 28 3029 46
rect 3081 50 3160 66
rect 3192 66 3364 68
rect 3192 50 3271 66
rect 3278 64 3308 66
rect 3081 42 3271 50
rect 3336 46 3342 66
rect 3081 38 3160 42
rect 3162 38 3190 42
rect 3192 38 3271 42
rect 3066 28 3074 38
rect 3093 30 3096 38
rect 3097 30 3115 38
rect 3160 30 3192 38
rect 3237 30 3255 38
rect 3093 28 3259 30
rect 3278 28 3289 38
rect 3351 28 3364 66
rect 3436 80 3465 96
rect 3479 80 3508 96
rect 3523 86 3553 102
rect 3581 80 3587 128
rect 3590 122 3609 128
rect 3624 122 3654 130
rect 3590 114 3654 122
rect 3590 98 3670 114
rect 3686 107 3748 138
rect 3764 107 3826 138
rect 3895 136 3944 161
rect 3959 136 3989 152
rect 3858 122 3888 130
rect 3895 128 4005 136
rect 3858 114 3903 122
rect 3590 96 3609 98
rect 3624 96 3670 98
rect 3590 80 3670 96
rect 3697 94 3732 107
rect 3773 104 3810 107
rect 3773 102 3815 104
rect 3702 91 3732 94
rect 3711 87 3718 91
rect 3718 86 3719 87
rect 3677 80 3687 86
rect 3436 72 3471 80
rect 3436 46 3437 72
rect 3444 46 3471 72
rect 3436 38 3471 46
rect 3473 72 3514 80
rect 3473 46 3488 72
rect 3495 46 3514 72
rect 3578 68 3609 80
rect 3624 68 3727 80
rect 3739 70 3765 96
rect 3780 91 3810 102
rect 3842 98 3904 114
rect 3842 96 3888 98
rect 3842 80 3904 96
rect 3916 80 3922 128
rect 3925 120 4005 128
rect 3925 118 3944 120
rect 3959 118 3993 120
rect 3925 102 4005 118
rect 3925 80 3944 102
rect 3959 86 3989 102
rect 4017 96 4023 170
rect 4026 96 4045 240
rect 4060 96 4066 240
rect 4075 170 4088 240
rect 4133 214 4162 228
rect 4215 214 4231 228
rect 4269 218 4275 226
rect 4282 224 4390 240
rect 4133 212 4231 214
rect 4117 204 4168 212
rect 4215 204 4249 212
rect 4117 192 4142 204
rect 4149 192 4168 204
rect 4222 202 4249 204
rect 4258 204 4275 218
rect 4320 204 4352 224
rect 4397 218 4403 226
rect 4411 218 4426 240
rect 4492 234 4511 237
rect 4397 212 4426 218
rect 4441 214 4457 228
rect 4492 215 4514 234
rect 4524 228 4540 229
rect 4523 226 4540 228
rect 4524 221 4540 226
rect 4514 214 4520 215
rect 4523 214 4552 221
rect 4441 213 4552 214
rect 4441 212 4558 213
rect 4397 204 4479 212
rect 4514 209 4520 212
rect 4258 202 4479 204
rect 4222 198 4294 202
rect 4322 200 4350 202
rect 4375 198 4479 202
rect 4117 184 4168 192
rect 4215 190 4347 198
rect 4350 190 4479 198
rect 4523 204 4558 212
rect 4215 188 4294 190
rect 4375 188 4479 190
rect 4215 184 4312 188
rect 4069 136 4088 170
rect 4133 176 4162 184
rect 4133 170 4150 176
rect 4133 168 4167 170
rect 4215 168 4231 184
rect 4232 180 4312 184
rect 4360 184 4479 188
rect 4360 180 4440 184
rect 4232 174 4440 180
rect 4441 174 4457 184
rect 4505 180 4520 195
rect 4523 192 4524 204
rect 4531 192 4558 204
rect 4523 184 4558 192
rect 4523 183 4552 184
rect 4243 170 4347 174
rect 4134 164 4167 168
rect 4130 162 4167 164
rect 4130 161 4197 162
rect 4130 156 4161 161
rect 4167 156 4197 161
rect 4258 158 4273 170
rect 4130 152 4197 156
rect 4103 149 4197 152
rect 4103 142 4152 149
rect 4103 136 4133 142
rect 4152 137 4157 142
rect 4069 120 4149 136
rect 4161 128 4197 149
rect 4282 148 4312 157
rect 4335 152 4353 170
rect 4411 168 4457 174
rect 4492 170 4505 180
rect 4523 170 4540 183
rect 4492 168 4540 170
rect 4373 162 4375 164
rect 4375 157 4387 162
rect 4360 150 4390 157
rect 4360 148 4391 150
rect 4411 148 4447 168
rect 4492 167 4539 168
rect 4505 162 4539 167
rect 4258 144 4447 148
rect 4273 141 4447 144
rect 4266 138 4447 141
rect 4475 161 4539 162
rect 4069 118 4088 120
rect 4103 118 4137 120
rect 4069 102 4149 118
rect 4069 96 4088 102
rect 3785 70 3888 80
rect 3739 68 3888 70
rect 3909 68 3944 80
rect 3578 66 3740 68
rect 3590 46 3609 66
rect 3624 64 3654 66
rect 3473 38 3514 46
rect 3436 28 3465 38
rect 3479 28 3508 38
rect 3596 28 3609 46
rect 3661 50 3740 66
rect 3772 66 3944 68
rect 3772 50 3851 66
rect 3858 64 3888 66
rect 3661 42 3851 50
rect 3916 46 3922 66
rect 3661 38 3740 42
rect 3742 38 3770 42
rect 3772 38 3851 42
rect 3646 28 3654 38
rect 3673 30 3676 38
rect 3677 30 3695 38
rect 3740 30 3772 38
rect 3817 30 3835 38
rect 3673 28 3839 30
rect 3858 28 3869 38
rect 3931 28 3944 66
rect 4016 80 4045 96
rect 4059 80 4088 96
rect 4103 86 4133 102
rect 4161 80 4167 128
rect 4170 122 4189 128
rect 4204 122 4234 130
rect 4170 114 4234 122
rect 4170 98 4250 114
rect 4266 107 4328 138
rect 4344 107 4406 138
rect 4475 136 4524 161
rect 4539 136 4569 152
rect 4438 122 4468 130
rect 4475 128 4585 136
rect 4438 114 4483 122
rect 4170 96 4189 98
rect 4204 96 4250 98
rect 4170 80 4250 96
rect 4277 94 4312 107
rect 4353 104 4390 107
rect 4353 102 4395 104
rect 4282 91 4312 94
rect 4291 87 4298 91
rect 4298 86 4299 87
rect 4257 80 4267 86
rect 4016 72 4051 80
rect 4016 46 4017 72
rect 4024 46 4051 72
rect 4016 38 4051 46
rect 4053 72 4094 80
rect 4053 46 4068 72
rect 4075 46 4094 72
rect 4158 68 4189 80
rect 4204 68 4307 80
rect 4319 70 4345 96
rect 4360 91 4390 102
rect 4422 98 4484 114
rect 4422 96 4468 98
rect 4422 80 4484 96
rect 4496 80 4502 128
rect 4505 120 4585 128
rect 4505 118 4524 120
rect 4539 118 4573 120
rect 4505 102 4585 118
rect 4505 80 4524 102
rect 4539 86 4569 102
rect 4597 96 4603 170
rect 4612 96 4625 240
rect 4365 70 4468 80
rect 4319 68 4468 70
rect 4489 68 4524 80
rect 4158 66 4320 68
rect 4170 46 4189 66
rect 4204 64 4234 66
rect 4053 38 4094 46
rect 4016 28 4045 38
rect 4059 28 4088 38
rect 4176 28 4189 46
rect 4241 50 4320 66
rect 4352 66 4524 68
rect 4352 50 4431 66
rect 4438 64 4468 66
rect 4241 42 4431 50
rect 4496 46 4502 66
rect 4241 38 4320 42
rect 4322 38 4350 42
rect 4352 38 4431 42
rect 4226 28 4234 38
rect 4253 30 4256 38
rect 4257 30 4275 38
rect 4320 30 4352 38
rect 4397 30 4415 38
rect 4253 28 4419 30
rect 4438 28 4449 38
rect 4511 28 4524 66
rect 4596 80 4625 96
rect 4596 72 4631 80
rect 4596 46 4597 72
rect 4604 46 4631 72
rect 4596 38 4631 46
rect 4596 28 4625 38
rect -1 22 4625 28
rect 0 14 4625 22
rect 15 0 28 14
rect 43 -4 73 14
rect 116 0 159 14
rect 166 1 174 14
rect 207 1 345 14
rect 378 1 386 14
rect 129 -18 159 0
rect 222 -2 330 1
rect 222 -4 252 -2
rect 300 -4 330 -2
rect 393 -18 423 14
rect 451 0 464 14
rect 479 -4 509 14
rect 546 0 565 14
rect 580 0 586 14
rect 595 0 608 14
rect 623 -4 653 14
rect 696 0 739 14
rect 746 1 754 14
rect 787 1 925 14
rect 958 1 966 14
rect 709 -18 739 0
rect 802 -2 910 1
rect 802 -4 832 -2
rect 880 -4 910 -2
rect 973 -18 1003 14
rect 1031 0 1044 14
rect 1059 -4 1089 14
rect 1126 0 1145 14
rect 1160 0 1166 14
rect 1175 0 1188 14
rect 1203 -4 1233 14
rect 1276 0 1319 14
rect 1326 1 1334 14
rect 1367 1 1505 14
rect 1538 1 1546 14
rect 1289 -18 1319 0
rect 1382 -2 1490 1
rect 1382 -4 1412 -2
rect 1460 -4 1490 -2
rect 1553 -18 1583 14
rect 1611 0 1624 14
rect 1639 -4 1669 14
rect 1706 0 1725 14
rect 1740 0 1746 14
rect 1755 0 1768 14
rect 1783 -4 1813 14
rect 1856 0 1899 14
rect 1906 1 1914 14
rect 1947 1 2085 14
rect 2118 1 2126 14
rect 1869 -18 1899 0
rect 1962 -2 2070 1
rect 1962 -4 1992 -2
rect 2040 -4 2070 -2
rect 2133 -18 2163 14
rect 2191 0 2204 14
rect 2219 -4 2249 14
rect 2286 0 2305 14
rect 2320 0 2326 14
rect 2335 0 2348 14
rect 2363 -4 2393 14
rect 2436 0 2479 14
rect 2486 1 2494 14
rect 2527 1 2665 14
rect 2698 1 2706 14
rect 2449 -18 2479 0
rect 2542 -2 2650 1
rect 2542 -4 2572 -2
rect 2620 -4 2650 -2
rect 2713 -18 2743 14
rect 2771 0 2784 14
rect 2799 -4 2829 14
rect 2866 0 2885 14
rect 2900 0 2906 14
rect 2915 0 2928 14
rect 2943 -4 2973 14
rect 3016 0 3059 14
rect 3066 1 3074 14
rect 3107 1 3245 14
rect 3278 1 3286 14
rect 3029 -18 3059 0
rect 3122 -2 3230 1
rect 3122 -4 3152 -2
rect 3200 -4 3230 -2
rect 3293 -18 3323 14
rect 3351 0 3364 14
rect 3379 -4 3409 14
rect 3446 0 3465 14
rect 3480 0 3486 14
rect 3495 0 3508 14
rect 3523 -4 3553 14
rect 3596 0 3639 14
rect 3646 1 3654 14
rect 3687 1 3825 14
rect 3858 1 3866 14
rect 3609 -18 3639 0
rect 3702 -2 3810 1
rect 3702 -4 3732 -2
rect 3780 -4 3810 -2
rect 3873 -18 3903 14
rect 3931 0 3944 14
rect 3959 -4 3989 14
rect 4026 0 4045 14
rect 4060 0 4066 14
rect 4075 0 4088 14
rect 4103 -4 4133 14
rect 4176 0 4219 14
rect 4226 1 4234 14
rect 4267 1 4405 14
rect 4438 1 4446 14
rect 4189 -18 4219 0
rect 4282 -2 4390 1
rect 4282 -4 4312 -2
rect 4360 -4 4390 -2
rect 4453 -18 4483 14
rect 4511 0 4524 14
rect 4539 -4 4569 14
rect 4612 0 4625 14
<< pwell >>
rect 552 0 580 270
rect 1132 0 1160 270
rect 1712 0 1740 270
rect 2292 0 2320 270
rect 2872 0 2900 270
rect 3452 0 3480 270
rect 4032 0 4060 270
<< poly >>
rect 552 240 580 270
rect 1132 240 1160 270
rect 1712 240 1740 270
rect 2292 240 2320 270
rect 2872 240 2900 270
rect 3452 240 3480 270
rect 4032 240 4060 270
<< polycont >>
rect 623 102 653 136
rect 1059 102 1089 136
rect 1203 102 1233 136
rect 1639 102 1669 136
rect 1783 102 1813 136
rect 2219 102 2249 136
rect 2363 102 2393 136
rect 2799 102 2829 136
rect 2943 102 2973 136
rect 3379 102 3409 136
rect 3523 102 3553 136
rect 3959 102 3989 136
rect 4103 102 4133 136
rect 4539 102 4569 136
<< viali >>
rect 43 102 73 136
rect 479 102 509 136
rect 623 102 653 136
rect 1059 102 1089 136
rect 1203 102 1233 136
rect 1639 102 1669 136
rect 1783 102 1813 136
rect 2219 102 2249 136
rect 2363 102 2393 136
rect 2799 102 2829 136
rect 2943 102 2973 136
rect 3379 102 3409 136
rect 3523 102 3553 136
rect 3959 102 3989 136
rect 4103 102 4133 136
rect 4539 102 4569 136
<< metal1 >>
rect 552 226 580 240
rect 1132 226 1160 240
rect 1712 226 1740 240
rect 2292 226 2320 240
rect 2872 226 2900 240
rect 3452 226 3480 240
rect 4032 226 4060 240
rect 0 102 43 136
rect 73 102 479 136
rect 509 102 623 136
rect 653 102 1059 136
rect 1089 102 1203 136
rect 1233 102 1639 136
rect 1669 102 1783 136
rect 1813 102 2219 136
rect 2249 102 2363 136
rect 2393 102 2799 136
rect 2829 102 2943 136
rect 2973 102 3379 136
rect 3409 102 3523 136
rect 3553 102 3959 136
rect 3989 102 4103 136
rect 4133 102 4539 136
rect 552 0 580 14
rect 1132 0 1160 14
rect 1712 0 1740 14
rect 2292 0 2320 14
rect 2872 0 2900 14
rect 3452 0 3480 14
rect 4032 0 4060 14
use 10T_toy_magic  10T_toy_magic_0
timestamp 1658880696
transform 1 0 3580 0 1 19
box -100 -19 452 251
use 10T_toy_magic  10T_toy_magic_1
timestamp 1658880696
transform 1 0 4160 0 1 19
box -100 -19 452 251
use 10T_toy_magic  10T_toy_magic_2
timestamp 1658880696
transform 1 0 3000 0 1 19
box -100 -19 452 251
use 10T_toy_magic  10T_toy_magic_3
timestamp 1658880696
transform 1 0 2420 0 1 19
box -100 -19 452 251
use 10T_toy_magic  10T_toy_magic_4
timestamp 1658880696
transform 1 0 1840 0 1 19
box -100 -19 452 251
use 10T_toy_magic  10T_toy_magic_5
timestamp 1658880696
transform 1 0 1260 0 1 19
box -100 -19 452 251
use 10T_toy_magic  10T_toy_magic_6
timestamp 1658880696
transform 1 0 680 0 1 19
box -100 -19 452 251
use 10T_toy_magic  10T_toy_magic_7
timestamp 1658880696
transform 1 0 100 0 1 19
box -100 -19 452 251
<< labels >>
rlabel poly 0 240 30 270 1 WWL
port 17 ew signal input
rlabel metal1 0 102 15 136 1 RWL
port 18 ew signal input
rlabel corelocali 74 184 89 212 1 WBLb_0
port 19 ns signal input
rlabel corelocali 464 184 479 213 1 WBL_0
port 20 ns signal input
rlabel corelocali 0 38 15 80 1 RBL1_0
port 1 ns signal output
rlabel corelocali 537 38 552 80 1 RBL0_0
port 2 ns signal output
rlabel corelocali 654 184 669 212 1 WBLb_1
port 21 ns signal input
rlabel corelocali 1044 184 1059 213 1 WBL_1
port 22 ns signal input
rlabel corelocali 580 38 595 80 1 RBL1_1
port 3 ns signal output
rlabel corelocali 1117 38 1132 80 1 RBL0_1
port 4 ns signal output
rlabel corelocali 1234 184 1249 212 1 WBLb_2
port 23 ns signal input
rlabel corelocali 1624 184 1639 213 1 WBL_2
port 24 ns signal input
rlabel corelocali 1160 38 1175 80 1 RBL1_2
port 5 ns signal output
rlabel corelocali 1697 38 1712 80 1 RBL0_2
port 6 ns signal output
rlabel corelocali 1814 184 1829 212 1 WBLb_3
port 25 ns signal input
rlabel corelocali 2204 184 2219 213 1 WBL_3
port 26 ns signal input
rlabel corelocali 1740 38 1755 80 1 RBL1_3
port 7 ns signal output
rlabel corelocali 2277 38 2292 80 1 RBL0_3
port 8 ns signal output
rlabel corelocali 2394 184 2409 212 1 WBLb_4
port 27 ns signal input
rlabel corelocali 2784 184 2799 213 1 WBL_4
port 28 ns signal input
rlabel corelocali 2320 38 2335 80 1 RBL1_4
port 8 ns signal output
rlabel corelocali 2857 38 2872 80 1 RBL0_4
port 10 ns signal output
rlabel corelocali 2974 184 2989 212 1 WBLb_5
port 29 ns signal input
rlabel corelocali 3364 184 3379 213 1 WBL_5
port 30 ns signal input
rlabel corelocali 2900 38 2915 80 1 RBL1_5
port 11 ns signal output
rlabel corelocali 3437 38 3452 80 1 RBL0_5
port 12 ns signal output
rlabel corelocali 3554 184 3569 212 1 WBLb_6
port 31 ns signal input
rlabel corelocali 3944 184 3959 213 1 WBL_6
port 32 ns signal input
rlabel corelocali 3480 38 3495 80 1 RBL1_6
port 13 ns signal output
rlabel corelocali 4017 38 4032 80 1 RBL0_6
port 14 ns signal output
rlabel corelocali 4134 184 4149 212 1 WBLb_7
port 33 ns signal input
rlabel corelocali 4524 184 4539 213 1 WBL_7
port 34 ns signal input
rlabel corelocali 4060 38 4075 80 1 RBL1_7
port 15 ns signal output
rlabel corelocali 4597 38 4612 80 1 RBL0_7
port 16 ns signal output
rlabel metal1 0 226 15 240 1 VDD
port 35 ns power bidirectional abutment
rlabel metal1 0 0 15 14 1 GND
port 36 ns ground bidirectional abutment
<< end >>
