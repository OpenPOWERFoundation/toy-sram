// Global Parameters for ToySRAM Testsite

`include "defines.v"

`define GENMODE 0      // 0=NoDelay, 1=Delay

// RA LCB
`define LCBSDR_CONFIGWIDTH 16
`define LCBDDR_CONFIGWIDTH 32

