* HSPICE file created from 10T_32x32_magic.ext - technology: sky130A

.option scale=0.005u

.subckt x10T_32x32_magic RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL0_3 RBL1_4
+ RBL0_4 RBL1_5 RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10
+ RBL0_10 RBL1_11 RBL0_11 RBL1_12 RBL0_12 RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15
+ RBL0_15 WWL_0 RWL_0 WWL_1 RWL_1 WWL_2 RWL_2 WWL_3 RWL_3 WWL_4 RWL_4 WWL_5 RWL_5
+ WWL_6 RWL_6 WWL_7 RWL_7 WWL_8 RWL_8 WWL_9 RWL_9 WWL_10 RWL_10 WWL_11 RWL_11 WWL_12
+ RWL_12 WWL_13 RWL_13 WWL_14 RWL_14 WWL_15 RWL_15 WWL_16 RWL_16 WWL_17 RWL_17 WWL_18
+ RWL_18 WWL_19 RWL_19 WWL_20 RWL_20 WWL_21 RWL_21 WWL_22 RWL_22 WWL_23 RWL_23 WWL_24
+ RWL_24 WWL_25 RWL_25 WWL_26 RWL_26 WWL_27 RWL_27 WWL_28 RWL_28 WWL_29 RWL_29 WWL_30
+ RWL_30 WWL_31 RWL_31 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL0_19
+ RBL1_20 RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 RBL1_24 RBL0_24
+ RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL0_27 RBL1_28 RBL0_28 RBL1_29 RBL0_29
+ RBL1_30 RBL0_30 RBL1_31 RBL0_31 WBL_0 WBLb_0 WBL_1 WBLb_1 WBL_2 WBLb_2 WBL_3 WBLb_19
+ WBL_4 WBLb_4 WBL_5 WBLb_5 WBL_22 WBLb_6 WBL_23 WBLb_7 WBL_24 WBLb_8 WBL_25 WBLb_9
+ WBL_26 WBLb_10 WBL_11 WBLb_11 WBL_12 WBLb_12 WBL_13 WBLb_13 WBL_14 WBLb_30 WBL_15
+ WBLb_31 VDD GND
C0 RWL_11 x0/VDD 2.32fF
C1 RBL0_12 RBL1_13 2.23fF
C2 x1/VDD RWL_8 2.32fF
C3 RWL_12 x2/VDD 2.32fF
C4 x3/VDD RWL_21 2.32fF
C5 x4/VDD RWL_22 2.32fF
C6 x5/VDD RWL_14 2.32fF
C7 x6/VDD RWL_26 2.32fF
C8 x7/VDD RWL_0 2.32fF
C9 x8/VDD RWL_16 2.32fF
C10 RWL_30 x9/VDD 2.32fF
C11 RWL_17 x10/VDD 2.28fF
C12 RWL_24 RWL_23 4.09fF
C13 RWL_26 RWL_27 4.09fF
C14 RWL_24 VDD 2.79fF
C15 RBL0_4 RBL1_5 2.23fF
C16 RWL_7 RWL_8 4.09fF
C17 RWL_30 RWL_31 4.09fF
C18 RWL_9 RWL_8 4.09fF
C19 RWL_7 x11/VDD 2.28fF
C20 x12/VDD RWL_29 2.32fF
C21 x13/VDD RWL_8 2.32fF
C22 RWL_26 x14/VDD 2.32fF
C23 RWL_15 RWL_14 4.09fF
C24 RBL0_8 RBL1_9 2.23fF
C25 x15/VDD RWL_31 2.32fF
C26 x16/VDD RWL_25 2.32fF
C27 RBL0_30 RBL1_31 2.23fF
C28 RWL_7 x17/VDD 2.32fF
C29 RWL_0 x18/VDD 2.28fF
C30 x19/VDD RWL_3 2.28fF
C31 WBLb_8 RBL0_7 2.11fF
C32 RBL1_8 WBL_7 2.42fF
C33 RWL_15 x20/VDD 2.32fF
C34 RBL0_0 RBL1_1 2.23fF
C35 RBL0_20 RBL1_21 2.23fF
C36 x21/VDD RWL_31 2.32fF
C37 x22/VDD RWL_8 2.32fF
C38 RWL_7 RWL_6 4.09fF
C39 RWL_17 RWL_18 4.09fF
C40 x23/VDD RWL_31 2.28fF
C41 x24/VDD RWL_26 2.28fF
C42 RBL0_26 RBL1_27 2.23fF
C43 x25/VDD RWL_29 2.32fF
C44 x26/VDD RWL_6 2.32fF
C45 RWL_2 x27/VDD 2.32fF
C46 RBL0_16 RBL1_17 2.23fF
C47 x28/VDD RWL_22 2.32fF
C48 RWL_28 RWL_29 4.09fF
C49 RWL_13 x29/VDD 2.28fF
C50 RWL_2 x19/RWL 2.04fF
C51 x30/VDD RWL_6 2.32fF
C52 RWL_2 x31/VDD 2.32fF
C53 x32/VDD RWL_24 2.28fF
C54 x33/VDD RWL_8 2.28fF
C55 x34/VDD RWL_4 2.32fF
C56 RWL_11 x35/VDD 2.32fF
C57 RWL_23 VDD 9.89fF
C58 RBL0_11 RBL1_12 2.23fF
C59 x36/VDD RWL_26 2.32fF
C60 RWL_30 RWL_29 4.11fF
C61 RWL_9 x37/VDD 2.32fF
C62 RBL1_8 RBL0_7 10.18fF
C63 RWL_6 RWL_5 4.09fF
C64 x38/VDD RWL_12 2.32fF
C65 x39/VDD RWL_27 2.32fF
C66 RWL_4 RWL_5 4.09fF
C67 x40/VDD RWL_5 2.32fF
C68 x41/VDD RWL_11 2.32fF
C69 RBL0_3 RBL1_4 2.23fF
C70 x42/VDD RWL_7 2.32fF
C71 RWL_1 x43/VDD 2.32fF
C72 x44/VDD RWL_24 2.32fF
C73 RWL_21 VDD 2.79fF
C74 x45/VDD RWL_9 2.32fF
C75 x46/VDD RWL_27 2.32fF
C76 x47/VDD RWL_27 2.28fF
C77 RWL_4 x48/VDD 2.28fF
C78 RWL_17 x49/VDD 2.32fF
C79 RBL0_29 RBL1_30 2.23fF
C80 RWL_19 x50/VDD 2.32fF
C81 RWL_9 x51/VDD 2.32fF
C82 RWL_15 x52/VDD 2.28fF
C83 RWL_12 x53/VDD 2.32fF
C84 RWL_30 x54/VDD 2.32fF
C85 RBL0_19 RBL1_20 2.23fF
C86 RWL_0 x55/VDD 2.32fF
C87 x56/VDD RWL_13 2.32fF
C88 RWL_25 RWL_26 4.09fF
C89 RBL0_25 RBL1_26 2.23fF
C90 RWL_28 x57/VDD 2.32fF
C91 x58/VDD RWL_29 2.32fF
C92 RWL_4 x19/RWL 2.04fF
C93 RBL0_23 WBLb_24 2.11fF
C94 WBL_23 RBL1_24 2.42fF
C95 x59/VDD RWL_24 2.32fF
C96 x60/VDD RWL_14 2.28fF
C97 RWL_9 x61/VDD 2.28fF
C98 RBL0_14 RBL1_15 2.23fF
C99 x62/VDD RWL_15 2.32fF
C100 RWL_30 x63/VDD 2.28fF
C101 RWL_18 RWL_19 4.09fF
C102 x64/VDD RWL_19 2.32fF
C103 x65/VDD RWL_21 2.28fF
C104 RWL_2 x66/VDD 2.28fF
C105 RBL0_6 RBL1_7 2.23fF
C106 RWL_19 x67/VDD 2.28fF
C107 RWL_10 x68/VDD 2.32fF
C108 RWL_4 x69/VDD 2.32fF
C109 x70/VDD RWL_28 2.32fF
C110 x71/VDD RWL_22 2.28fF
C111 RBL0_10 RBL1_11 2.23fF
C112 RWL_17 x72/VDD 2.32fF
C113 RWL_10 x73/VDD 2.32fF
C114 RWL_1 RWL_2 4.09fF
C115 RWL_19 VDD 6.48fF
C116 x74/VDD RWL_16 2.28fF
C117 RWL_17 RWL_16 4.09fF
C118 RWL_4 x75/VDD 2.32fF
C119 x76/VDD RWL_1 2.32fF
C120 x77/VDD RWL_28 2.28fF
C121 x78/VDD RWL_16 2.32fF
C122 RWL_5 x79/VDD 2.32fF
C123 RBL0_2 RBL1_3 2.23fF
C124 RBL0_22 RBL1_23 2.23fF
C125 x80/VDD RWL_24 2.32fF
C126 RWL_25 x81/VDD 2.32fF
C127 RBL0_28 RBL1_29 2.23fF
C128 RWL_7 x82/VDD 2.32fF
C129 x83/VDD RWL_5 2.32fF
C130 RWL_25 RWL_24 4.09fF
C131 VDD RWL_20 9.89fF
C132 RBL0_23 RBL1_24 10.18fF
C133 x84/VDD RWL_22 2.32fF
C134 WBLb_16 RBL0_15 2.11fF
C135 RBL1_16 WBL_15 2.42fF
C136 RWL_12 x85/VDD 2.28fF
C137 x86/VDD RWL_28 2.32fF
C138 RBL0_18 RBL1_19 2.23fF
C139 x87/VDD RWL_30 2.32fF
C140 RWL_11 RWL_12 4.09fF
C141 RWL_1 RWL_0 4.23fF
C142 x88/VDD RWL_16 2.32fF
C143 RBL0_24 RBL1_25 2.23fF
C144 RWL_21 RWL_20 4.09fF
C145 RWL_10 x89/VDD 2.28fF
C146 x90/VDD RWL_10 2.32fF
C147 RWL_1 x91/VDD 2.32fF
C148 x92/VDD RWL_31 2.32fF
C149 RBL0_13 RBL1_14 2.23fF
C150 x93/VDD RWL_18 2.32fF
C151 x19/RWL x94/VDD 2.28fF
C152 x95/VDD RWL_14 2.32fF
C153 RWL_13 RWL_14 4.09fF
C154 x96/VDD RWL_29 2.28fF
C155 RWL_25 x97/VDD 2.28fF
C156 x98/VDD x94/RWL 2.28fF
C157 x99/VDD RWL_18 2.28fF
C158 RBL0_5 RBL1_6 2.23fF
C159 RWL_28 RWL_27 4.09fF
C160 GND VDD 76.06fF
C161 RWL_5 x100/VDD 2.28fF
C162 RBL0_9 RBL1_10 2.23fF
C163 x101/VDD RWL_15 2.32fF
C164 x102/VDD RWL_2 2.32fF
C165 x103/VDD RWL_27 2.32fF
C166 RWL_22 RWL_23 4.09fF
C167 x104/VDD RWL_17 2.32fF
C168 RWL_22 VDD 6.48fF
C169 RBL1_16 RBL0_15 10.18fF
C170 RWL_18 x105/VDD 2.32fF
C171 x106/VDD RWL_13 2.32fF
C172 RBL0_1 RBL1_2 2.23fF
C173 RBL0_21 RBL1_22 2.23fF
C174 x107/VDD RWL_6 2.28fF
C175 RWL_19 x108/VDD 2.32fF
C176 x109/VDD RWL_6 2.32fF
C177 RWL_11 RWL_10 4.09fF
C178 RBL0_27 RBL1_28 2.23fF
C179 RWL_21 RWL_22 4.09fF
C180 RWL_10 RWL_9 4.09fF
C181 x110/VDD RWL_18 2.32fF
C182 RWL_15 RWL_16 4.09fF
C183 x111/VDD x19/RWL 2.32fF
C184 RWL_11 x112/VDD 2.28fF
C185 x113/VDD RWL_21 2.32fF
C186 RBL0_17 RBL1_18 2.23fF
C187 RWL_21 x114/VDD 2.32fF
C188 RWL_19 RWL_20 4.09fF
C189 RWL_12 RWL_13 4.09fF
C190 x115/VDD RWL_0 2.32fF
C191 x116/VDD RWL_14 2.32fF
C192 RWL_1 x117/VDD 2.28fF
C193 x118/VDD RWL_13 2.32fF
C194 RWL_25 x119/VDD 2.32fF
X10T_1x8_magic_0 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_2 RWL_2 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x10T_1x8_magic
X10T_1x8_magic_1 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_3 RWL_3 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x10T_1x8_magic
X10T_1x8_magic_2 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_0 RWL_0 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x10T_1x8_magic
X10T_1x8_magic_3 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_1 RWL_1 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x10T_1x8_magic
X10T_1x8_magic_4 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_7 RWL_7 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x10T_1x8_magic
X10T_1x8_magic_5 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_6 RWL_6 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x10T_1x8_magic
X10T_1x8_magic_6 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_4 RWL_4 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x10T_1x8_magic
X10T_1x8_magic_7 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_5 RWL_5 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x10T_1x8_magic
X10T_1x8_magic_90 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x72/WWL RWL_17 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x72/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_8 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_14 RWL_14 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x10T_1x8_magic
X10T_1x8_magic_80 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x120/WWL RWL_23 WBLb_16
+ WBL_16 WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21
+ WBLb_22 WBL_22 WBLb_23 WBL_23 VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_91 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x105/WWL RWL_18 WBLb_16
+ WBL_16 WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21
+ WBLb_22 WBL_22 WBLb_23 WBL_23 x105/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_70 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x57/WWL RWL_28 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x57/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_81 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x121/WWL RWL_23 WBLb_24
+ WBL_24 WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29
+ WBLb_30 WBL_30 WBLb_31 WBL_31 VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_92 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x104/WWL RWL_17 WBLb_24
+ WBL_24 WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29
+ WBLb_30 WBL_30 WBLb_31 WBL_31 x104/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_9 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_15 RWL_15 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x10T_1x8_magic
X10T_1x8_magic_60 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x19/WWL x19/RWL WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x19/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_71 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x86/WWL RWL_28 WBLb_24 WBL_24
+ WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29 WBLb_30
+ WBL_30 WBLb_31 WBL_31 x86/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_82 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x84/WWL RWL_22 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x84/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_93 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x110/WWL RWL_18 WBLb_24
+ WBL_24 WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29
+ WBLb_30 WBL_30 WBLb_31 WBL_31 x110/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_61 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x102/WWL RWL_2 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x102/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_72 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x39/WWL RWL_27 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x39/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_83 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x28/WWL RWL_22 WBLb_24 WBL_24
+ WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29 WBLb_30
+ WBL_30 WBLb_31 WBL_31 x28/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_94 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x78/WWL RWL_16 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x78/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_50 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x106/WWL RWL_13 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x106/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_62 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x76/WWL RWL_1 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x76/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_120 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x111/WWL x19/RWL WBLb_16
+ WBL_16 WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21
+ WBLb_22 WBL_22 WBLb_23 WBL_23 x111/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_73 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x103/WWL RWL_27 WBLb_24
+ WBL_24 WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29
+ WBLb_30 WBL_30 WBLb_31 WBL_31 x103/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_40 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x81/WWL RWL_25 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x81/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_84 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x3/WWL RWL_21 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x3/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_95 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x88/WWL RWL_16 WBLb_24 WBL_24
+ WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29 WBLb_30
+ WBL_30 WBLb_31 WBL_31 x88/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_51 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x2/WWL RWL_12 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x2/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_63 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x115/WWL RWL_0 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x115/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_121 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x94/WWL x94/RWL WBLb_24
+ WBL_24 WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29
+ WBLb_30 WBL_30 WBLb_31 WBL_31 x94/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_74 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x14/WWL RWL_26 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x14/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_41 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x4/WWL RWL_22 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x4/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_85 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x113/WWL RWL_21 WBLb_24
+ WBL_24 WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29
+ WBLb_30 WBL_30 WBLb_31 WBL_31 x113/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_30 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_18 RWL_18 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x10T_1x8_magic
X10T_1x8_magic_96 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x20/WWL RWL_15 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x20/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_52 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x41/WWL RWL_11 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x41/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_110 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x22/WWL RWL_8 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x22/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_122 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x27/WWL RWL_2 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x27/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_64 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x21/WWL RWL_31 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x21/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_20 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_28 RWL_28 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x10T_1x8_magic
X10T_1x8_magic_75 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x36/WWL RWL_26 WBLb_24 WBL_24
+ WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29 WBLb_30
+ WBL_30 WBLb_31 WBL_31 x36/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_42 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x114/WWL RWL_21 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x114/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_86 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x122/WWL RWL_20 WBLb_16
+ WBL_16 WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21
+ WBLb_22 WBL_22 WBLb_23 WBL_23 VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_31 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_16 RWL_16 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x10T_1x8_magic
X10T_1x8_magic_97 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x62/WWL RWL_15 WBLb_24 WBL_24
+ WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29 WBLb_30
+ WBL_30 WBLb_31 WBL_31 x62/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_100 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x118/WWL RWL_13 WBLb_16
+ WBL_16 WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21
+ WBLb_22 WBL_22 WBLb_23 WBL_23 x118/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_53 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x73/WWL RWL_10 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x73/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_111 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x1/WWL RWL_8 WBLb_24 WBL_24
+ WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29 WBLb_30
+ WBL_30 WBLb_31 WBL_31 x1/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_123 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x31/WWL RWL_2 WBLb_24 WBL_24
+ WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29 WBLb_30
+ WBL_30 WBLb_31 WBL_31 x31/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_112 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x17/WWL RWL_7 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x17/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_32 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x54/WWL RWL_30 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x54/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_65 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x87/WWL RWL_30 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x87/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_21 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_25 RWL_25 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x10T_1x8_magic
X10T_1x8_magic_76 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x16/WWL RWL_25 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x16/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_43 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x123/WWL RWL_20 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_87 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x124/WWL RWL_20 WBLb_24
+ WBL_24 WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29
+ WBLb_30 WBL_30 WBLb_31 WBL_31 VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_98 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x116/WWL RWL_14 WBLb_16
+ WBL_16 WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21
+ WBLb_22 WBL_22 WBLb_23 WBL_23 x116/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_10 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_13 RWL_13 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x10T_1x8_magic
X10T_1x8_magic_101 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x56/WWL RWL_13 WBLb_24 WBL_24
+ WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29 WBLb_30
+ WBL_30 WBLb_31 WBL_31 x56/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_54 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x37/WWL RWL_9 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x37/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_124 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x91/WWL RWL_1 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x91/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_113 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x82/WWL RWL_7 WBLb_24 WBL_24
+ WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29 WBLb_30
+ WBL_30 WBLb_31 WBL_31 x82/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_33 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x92/WWL RWL_31 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x92/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_66 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x9/WWL RWL_30 WBLb_24 WBL_24
+ WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29 WBLb_30
+ WBL_30 WBLb_31 WBL_31 x9/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_22 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_26 RWL_26 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x10T_1x8_magic
X10T_1x8_magic_77 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x59/WWL RWL_24 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x59/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_44 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x50/WWL RWL_19 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x50/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_88 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x64/WWL RWL_19 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x64/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_99 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x5/WWL RWL_14 WBLb_24 WBL_24
+ WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29 WBLb_30
+ WBL_30 WBLb_31 WBL_31 x5/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_11 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_12 RWL_12 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x10T_1x8_magic
X10T_1x8_magic_102 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x38/WWL RWL_12 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x38/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_55 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x13/WWL RWL_8 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x13/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_12 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_11 RWL_11 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x10T_1x8_magic
X10T_1x8_magic_125 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x43/WWL RWL_1 WBLb_24 WBL_24
+ WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29 WBLb_30
+ WBL_30 WBLb_31 WBL_31 x43/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_114 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x30/WWL RWL_6 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x30/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_56 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x42/WWL RWL_7 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x42/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_67 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x15/WWL RWL_31 WBLb_24 WBL_24
+ WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29 WBLb_30
+ WBL_30 WBLb_31 WBL_31 x15/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_34 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x70/WWL RWL_28 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x70/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_78 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x80/WWL RWL_24 WBLb_24 WBL_24
+ WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29 WBLb_30
+ WBL_30 WBLb_31 WBL_31 x80/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_23 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_23 RWL_23 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x10T_1x8_magic
X10T_1x8_magic_89 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x108/WWL RWL_19 WBLb_24
+ WBL_24 WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29
+ WBLb_30 WBL_30 WBLb_31 WBL_31 x108/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_45 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x49/WWL RWL_17 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x49/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_103 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x53/WWL RWL_12 WBLb_24 WBL_24
+ WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29 WBLb_30
+ WBL_30 WBLb_31 WBL_31 x53/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_126 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x7/WWL RWL_0 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x7/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_115 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x26/WWL RWL_6 WBLb_24 WBL_24
+ WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29 WBLb_30
+ WBL_30 WBLb_31 WBL_31 x26/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_57 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x109/WWL RWL_6 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x109/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_35 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x25/WWL RWL_29 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x25/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_68 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x12/WWL RWL_29 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x12/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_79 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x119/WWL RWL_25 WBLb_24
+ WBL_24 WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29
+ WBLb_30 WBL_30 WBLb_31 WBL_31 x119/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_24 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_24 RWL_24 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x10T_1x8_magic
X10T_1x8_magic_46 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x93/WWL RWL_18 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x93/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_104 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x35/WWL RWL_11 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x35/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_13 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_10 RWL_10 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x10T_1x8_magic
X10T_1x8_magic_127 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x55/WWL RWL_0 WBLb_24 WBL_24
+ WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29 WBLb_30
+ WBL_30 WBLb_31 WBL_31 x55/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_116 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x69/WWL RWL_4 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x69/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_58 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x40/WWL RWL_5 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x40/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_69 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x58/WWL RWL_29 WBLb_24 WBL_24
+ WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29 WBLb_30
+ WBL_30 WBLb_31 WBL_31 x58/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_36 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x6/WWL RWL_26 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x6/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_25 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_21 RWL_21 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x10T_1x8_magic
X10T_1x8_magic_47 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x8/WWL RWL_16 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x8/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_105 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x90/WWL RWL_10 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x90/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_14 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_8 RWL_8 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x10T_1x8_magic
X10T_1x8_magic_59 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x34/WWL RWL_4 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x34/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_117 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x83/WWL RWL_5 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x83/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_37 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x46/WWL RWL_27 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x46/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_26 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_22 RWL_22 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x10T_1x8_magic
X10T_1x8_magic_48 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x101/WWL RWL_15 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x101/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_106 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x0/WWL RWL_11 WBLb_24 WBL_24
+ WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29 WBLb_30
+ WBL_30 WBLb_31 WBL_31 x0/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_15 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_9 RWL_9 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x10T_1x8_magic
X10T_1x8_magic_118 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x79/WWL RWL_5 WBLb_24 WBL_24
+ WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29 WBLb_30
+ WBL_30 WBLb_31 WBL_31 x79/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_16 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_31 RWL_31 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x10T_1x8_magic
X10T_1x8_magic_38 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x44/WWL RWL_24 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x44/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_27 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_19 RWL_19 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x10T_1x8_magic
X10T_1x8_magic_49 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x95/WWL RWL_14 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x95/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_107 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x68/WWL RWL_10 WBLb_24 WBL_24
+ WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29 WBLb_30
+ WBL_30 WBLb_31 WBL_31 x68/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_119 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x75/WWL RWL_4 WBLb_24 WBL_24
+ WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29 WBLb_30
+ WBL_30 WBLb_31 WBL_31 x75/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_17 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_29 RWL_29 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x10T_1x8_magic
X10T_1x8_magic_39 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x125/WWL RWL_23 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_28 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_20 RWL_20 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x10T_1x8_magic
X10T_1x8_magic_108 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x45/WWL RWL_9 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x45/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_18 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_30 RWL_30 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x10T_1x8_magic
X10T_1x8_magic_29 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_17 RWL_17 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x10T_1x8_magic
X10T_1x8_magic_109 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x51/WWL RWL_9 WBLb_24 WBL_24
+ WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29 WBLb_30
+ WBL_30 WBLb_31 WBL_31 x51/VDD VSUBS x10T_1x8_magic
X10T_1x8_magic_19 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_27 RWL_27 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x10T_1x8_magic
C195 x61/VDD VSUBS 7.76fF
C196 x48/VDD VSUBS 7.76fF
C197 x89/VDD VSUBS 7.76fF
C198 x100/VDD VSUBS 7.76fF
C199 x112/VDD VSUBS 7.76fF
C200 x96/VDD VSUBS 7.76fF
C201 x18/VDD VSUBS 2.19fF
C202 x97/VDD VSUBS 7.76fF
C203 x107/VDD VSUBS 7.76fF
C204 x85/VDD VSUBS 7.76fF
C205 x67/VDD VSUBS 7.76fF
C206 x32/VDD VSUBS 7.76fF
C207 x23/VDD VSUBS 7.77fF
C208 x117/VDD VSUBS 7.26fF
C209 x60/VDD VSUBS 7.76fF
C210 x63/VDD VSUBS 7.94fF
C211 x11/VDD VSUBS 7.76fF
C212 x29/VDD VSUBS 7.76fF
C213 x66/VDD VSUBS 7.76fF
C214 x33/VDD VSUBS 7.76fF
C215 x52/VDD VSUBS 7.76fF
C216 x24/VDD VSUBS 7.76fF
C217 x65/VDD VSUBS 7.76fF
C218 x98/VDD VSUBS 7.76fF
C219 x74/VDD VSUBS 7.76fF
C220 x47/VDD VSUBS 7.76fF
C221 x71/VDD VSUBS 7.76fF
C222 x99/VDD VSUBS 7.76fF
C223 x77/VDD VSUBS 7.76fF
C224 x10/VDD VSUBS 7.76fF
.ends

** hspice subcircuit dictionary
* x0	10T_1x8_magic_106
* x1	10T_1x8_magic_111
* x2	10T_1x8_magic_51
* x3	10T_1x8_magic_84
* x4	10T_1x8_magic_41
* x5	10T_1x8_magic_99
* x6	10T_1x8_magic_36
* x7	10T_1x8_magic_126
* x8	10T_1x8_magic_47
* x9	10T_1x8_magic_66
* x10	10T_1x8_magic_92/10T_toy_magic_7
* x11	10T_1x8_magic_113/10T_toy_magic_7
* x12	10T_1x8_magic_68
* x13	10T_1x8_magic_55
* x14	10T_1x8_magic_74
* x15	10T_1x8_magic_67
* x16	10T_1x8_magic_76
* x17	10T_1x8_magic_112
* x18	10T_1x8_magic_127/10T_toy_magic_7
* x19	10T_1x8_magic_60
* x20	10T_1x8_magic_96
* x21	10T_1x8_magic_64
* x22	10T_1x8_magic_110
* x23	10T_1x8_magic_67/10T_toy_magic_7
* x24	10T_1x8_magic_75/10T_toy_magic_7
* x25	10T_1x8_magic_35
* x26	10T_1x8_magic_115
* x27	10T_1x8_magic_122
* x28	10T_1x8_magic_83
* x29	10T_1x8_magic_101/10T_toy_magic_7
* x30	10T_1x8_magic_114
* x31	10T_1x8_magic_123
* x32	10T_1x8_magic_78/10T_toy_magic_7
* x33	10T_1x8_magic_111/10T_toy_magic_7
* x34	10T_1x8_magic_59
* x35	10T_1x8_magic_104
* x36	10T_1x8_magic_75
* x37	10T_1x8_magic_54
* x38	10T_1x8_magic_102
* x39	10T_1x8_magic_72
* x40	10T_1x8_magic_58
* x41	10T_1x8_magic_52
* x42	10T_1x8_magic_56
* x43	10T_1x8_magic_125
* x44	10T_1x8_magic_38
* x45	10T_1x8_magic_108
* x46	10T_1x8_magic_37
* x47	10T_1x8_magic_73/10T_toy_magic_7
* x48	10T_1x8_magic_119/10T_toy_magic_7
* x49	10T_1x8_magic_45
* x50	10T_1x8_magic_44
* x51	10T_1x8_magic_109
* x52	10T_1x8_magic_97/10T_toy_magic_7
* x53	10T_1x8_magic_103
* x54	10T_1x8_magic_32
* x55	10T_1x8_magic_127
* x56	10T_1x8_magic_101
* x57	10T_1x8_magic_70
* x58	10T_1x8_magic_69
* x59	10T_1x8_magic_77
* x60	10T_1x8_magic_99/10T_toy_magic_7
* x61	10T_1x8_magic_109/10T_toy_magic_7
* x62	10T_1x8_magic_97
* x63	10T_1x8_magic_66/10T_toy_magic_7
* x64	10T_1x8_magic_88
* x65	10T_1x8_magic_85/10T_toy_magic_7
* x66	10T_1x8_magic_123/10T_toy_magic_7
* x67	10T_1x8_magic_89/10T_toy_magic_7
* x68	10T_1x8_magic_107
* x69	10T_1x8_magic_116
* x70	10T_1x8_magic_34
* x71	10T_1x8_magic_83/10T_toy_magic_7
* x72	10T_1x8_magic_90
* x73	10T_1x8_magic_53
* x74	10T_1x8_magic_95/10T_toy_magic_7
* x75	10T_1x8_magic_119
* x76	10T_1x8_magic_62
* x77	10T_1x8_magic_71/10T_toy_magic_7
* x78	10T_1x8_magic_94
* x79	10T_1x8_magic_118
* x80	10T_1x8_magic_78
* x81	10T_1x8_magic_40
* x82	10T_1x8_magic_113
* x83	10T_1x8_magic_117
* x84	10T_1x8_magic_82
* x85	10T_1x8_magic_103/10T_toy_magic_7
* x86	10T_1x8_magic_71
* x87	10T_1x8_magic_65
* x88	10T_1x8_magic_95
* x89	10T_1x8_magic_107/10T_toy_magic_7
* x90	10T_1x8_magic_105
* x91	10T_1x8_magic_124
* x92	10T_1x8_magic_33
* x93	10T_1x8_magic_46
* x94	10T_1x8_magic_121
* x95	10T_1x8_magic_49
* x96	10T_1x8_magic_69/10T_toy_magic_7
* x97	10T_1x8_magic_79/10T_toy_magic_7
* x98	10T_1x8_magic_121/10T_toy_magic_7
* x99	10T_1x8_magic_93/10T_toy_magic_7
* x100	10T_1x8_magic_118/10T_toy_magic_7
* x101	10T_1x8_magic_48
* x102	10T_1x8_magic_61
* x103	10T_1x8_magic_73
* x104	10T_1x8_magic_92
* x105	10T_1x8_magic_91
* x106	10T_1x8_magic_50
* x107	10T_1x8_magic_115/10T_toy_magic_7
* x108	10T_1x8_magic_89
* x109	10T_1x8_magic_57
* x110	10T_1x8_magic_93
* x111	10T_1x8_magic_120
* x112	10T_1x8_magic_106/10T_toy_magic_7
* x113	10T_1x8_magic_85
* x114	10T_1x8_magic_42
* x115	10T_1x8_magic_63
* x116	10T_1x8_magic_98
* x117	10T_1x8_magic_125/10T_toy_magic_7
* x118	10T_1x8_magic_100
* x119	10T_1x8_magic_79
* x120	10T_1x8_magic_80
* x121	10T_1x8_magic_81
* x122	10T_1x8_magic_86
* x123	10T_1x8_magic_43
* x124	10T_1x8_magic_87
* x125	10T_1x8_magic_39
