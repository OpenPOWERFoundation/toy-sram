magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< pwell >>
rect 15 163 2283 817
<< mvnmos >>
rect 241 189 341 791
rect 397 189 497 791
rect 553 189 653 791
rect 709 189 809 791
rect 865 189 965 791
rect 1021 189 1121 791
rect 1177 189 1277 791
rect 1333 189 1433 791
rect 1489 189 1589 791
rect 1645 189 1745 791
rect 1801 189 1901 791
rect 1957 189 2057 791
<< mvndiff >>
rect 181 779 241 791
rect 181 745 196 779
rect 230 745 241 779
rect 181 711 241 745
rect 181 677 196 711
rect 230 677 241 711
rect 181 643 241 677
rect 181 609 196 643
rect 230 609 241 643
rect 181 575 241 609
rect 181 541 196 575
rect 230 541 241 575
rect 181 507 241 541
rect 181 473 196 507
rect 230 473 241 507
rect 181 439 241 473
rect 181 405 196 439
rect 230 405 241 439
rect 181 371 241 405
rect 181 337 196 371
rect 230 337 241 371
rect 181 303 241 337
rect 181 269 196 303
rect 230 269 241 303
rect 181 235 241 269
rect 181 201 196 235
rect 230 201 241 235
rect 181 189 241 201
rect 341 779 397 791
rect 341 745 352 779
rect 386 745 397 779
rect 341 711 397 745
rect 341 677 352 711
rect 386 677 397 711
rect 341 643 397 677
rect 341 609 352 643
rect 386 609 397 643
rect 341 575 397 609
rect 341 541 352 575
rect 386 541 397 575
rect 341 507 397 541
rect 341 473 352 507
rect 386 473 397 507
rect 341 439 397 473
rect 341 405 352 439
rect 386 405 397 439
rect 341 371 397 405
rect 341 337 352 371
rect 386 337 397 371
rect 341 303 397 337
rect 341 269 352 303
rect 386 269 397 303
rect 341 235 397 269
rect 341 201 352 235
rect 386 201 397 235
rect 341 189 397 201
rect 497 779 553 791
rect 497 745 508 779
rect 542 745 553 779
rect 497 711 553 745
rect 497 677 508 711
rect 542 677 553 711
rect 497 643 553 677
rect 497 609 508 643
rect 542 609 553 643
rect 497 575 553 609
rect 497 541 508 575
rect 542 541 553 575
rect 497 507 553 541
rect 497 473 508 507
rect 542 473 553 507
rect 497 439 553 473
rect 497 405 508 439
rect 542 405 553 439
rect 497 371 553 405
rect 497 337 508 371
rect 542 337 553 371
rect 497 303 553 337
rect 497 269 508 303
rect 542 269 553 303
rect 497 235 553 269
rect 497 201 508 235
rect 542 201 553 235
rect 497 189 553 201
rect 653 779 709 791
rect 653 745 664 779
rect 698 745 709 779
rect 653 711 709 745
rect 653 677 664 711
rect 698 677 709 711
rect 653 643 709 677
rect 653 609 664 643
rect 698 609 709 643
rect 653 575 709 609
rect 653 541 664 575
rect 698 541 709 575
rect 653 507 709 541
rect 653 473 664 507
rect 698 473 709 507
rect 653 439 709 473
rect 653 405 664 439
rect 698 405 709 439
rect 653 371 709 405
rect 653 337 664 371
rect 698 337 709 371
rect 653 303 709 337
rect 653 269 664 303
rect 698 269 709 303
rect 653 235 709 269
rect 653 201 664 235
rect 698 201 709 235
rect 653 189 709 201
rect 809 779 865 791
rect 809 745 820 779
rect 854 745 865 779
rect 809 711 865 745
rect 809 677 820 711
rect 854 677 865 711
rect 809 643 865 677
rect 809 609 820 643
rect 854 609 865 643
rect 809 575 865 609
rect 809 541 820 575
rect 854 541 865 575
rect 809 507 865 541
rect 809 473 820 507
rect 854 473 865 507
rect 809 439 865 473
rect 809 405 820 439
rect 854 405 865 439
rect 809 371 865 405
rect 809 337 820 371
rect 854 337 865 371
rect 809 303 865 337
rect 809 269 820 303
rect 854 269 865 303
rect 809 235 865 269
rect 809 201 820 235
rect 854 201 865 235
rect 809 189 865 201
rect 965 779 1021 791
rect 965 745 976 779
rect 1010 745 1021 779
rect 965 711 1021 745
rect 965 677 976 711
rect 1010 677 1021 711
rect 965 643 1021 677
rect 965 609 976 643
rect 1010 609 1021 643
rect 965 575 1021 609
rect 965 541 976 575
rect 1010 541 1021 575
rect 965 507 1021 541
rect 965 473 976 507
rect 1010 473 1021 507
rect 965 439 1021 473
rect 965 405 976 439
rect 1010 405 1021 439
rect 965 371 1021 405
rect 965 337 976 371
rect 1010 337 1021 371
rect 965 303 1021 337
rect 965 269 976 303
rect 1010 269 1021 303
rect 965 235 1021 269
rect 965 201 976 235
rect 1010 201 1021 235
rect 965 189 1021 201
rect 1121 779 1177 791
rect 1121 745 1132 779
rect 1166 745 1177 779
rect 1121 711 1177 745
rect 1121 677 1132 711
rect 1166 677 1177 711
rect 1121 643 1177 677
rect 1121 609 1132 643
rect 1166 609 1177 643
rect 1121 575 1177 609
rect 1121 541 1132 575
rect 1166 541 1177 575
rect 1121 507 1177 541
rect 1121 473 1132 507
rect 1166 473 1177 507
rect 1121 439 1177 473
rect 1121 405 1132 439
rect 1166 405 1177 439
rect 1121 371 1177 405
rect 1121 337 1132 371
rect 1166 337 1177 371
rect 1121 303 1177 337
rect 1121 269 1132 303
rect 1166 269 1177 303
rect 1121 235 1177 269
rect 1121 201 1132 235
rect 1166 201 1177 235
rect 1121 189 1177 201
rect 1277 779 1333 791
rect 1277 745 1288 779
rect 1322 745 1333 779
rect 1277 711 1333 745
rect 1277 677 1288 711
rect 1322 677 1333 711
rect 1277 643 1333 677
rect 1277 609 1288 643
rect 1322 609 1333 643
rect 1277 575 1333 609
rect 1277 541 1288 575
rect 1322 541 1333 575
rect 1277 507 1333 541
rect 1277 473 1288 507
rect 1322 473 1333 507
rect 1277 439 1333 473
rect 1277 405 1288 439
rect 1322 405 1333 439
rect 1277 371 1333 405
rect 1277 337 1288 371
rect 1322 337 1333 371
rect 1277 303 1333 337
rect 1277 269 1288 303
rect 1322 269 1333 303
rect 1277 235 1333 269
rect 1277 201 1288 235
rect 1322 201 1333 235
rect 1277 189 1333 201
rect 1433 779 1489 791
rect 1433 745 1444 779
rect 1478 745 1489 779
rect 1433 711 1489 745
rect 1433 677 1444 711
rect 1478 677 1489 711
rect 1433 643 1489 677
rect 1433 609 1444 643
rect 1478 609 1489 643
rect 1433 575 1489 609
rect 1433 541 1444 575
rect 1478 541 1489 575
rect 1433 507 1489 541
rect 1433 473 1444 507
rect 1478 473 1489 507
rect 1433 439 1489 473
rect 1433 405 1444 439
rect 1478 405 1489 439
rect 1433 371 1489 405
rect 1433 337 1444 371
rect 1478 337 1489 371
rect 1433 303 1489 337
rect 1433 269 1444 303
rect 1478 269 1489 303
rect 1433 235 1489 269
rect 1433 201 1444 235
rect 1478 201 1489 235
rect 1433 189 1489 201
rect 1589 779 1645 791
rect 1589 745 1600 779
rect 1634 745 1645 779
rect 1589 711 1645 745
rect 1589 677 1600 711
rect 1634 677 1645 711
rect 1589 643 1645 677
rect 1589 609 1600 643
rect 1634 609 1645 643
rect 1589 575 1645 609
rect 1589 541 1600 575
rect 1634 541 1645 575
rect 1589 507 1645 541
rect 1589 473 1600 507
rect 1634 473 1645 507
rect 1589 439 1645 473
rect 1589 405 1600 439
rect 1634 405 1645 439
rect 1589 371 1645 405
rect 1589 337 1600 371
rect 1634 337 1645 371
rect 1589 303 1645 337
rect 1589 269 1600 303
rect 1634 269 1645 303
rect 1589 235 1645 269
rect 1589 201 1600 235
rect 1634 201 1645 235
rect 1589 189 1645 201
rect 1745 779 1801 791
rect 1745 745 1756 779
rect 1790 745 1801 779
rect 1745 711 1801 745
rect 1745 677 1756 711
rect 1790 677 1801 711
rect 1745 643 1801 677
rect 1745 609 1756 643
rect 1790 609 1801 643
rect 1745 575 1801 609
rect 1745 541 1756 575
rect 1790 541 1801 575
rect 1745 507 1801 541
rect 1745 473 1756 507
rect 1790 473 1801 507
rect 1745 439 1801 473
rect 1745 405 1756 439
rect 1790 405 1801 439
rect 1745 371 1801 405
rect 1745 337 1756 371
rect 1790 337 1801 371
rect 1745 303 1801 337
rect 1745 269 1756 303
rect 1790 269 1801 303
rect 1745 235 1801 269
rect 1745 201 1756 235
rect 1790 201 1801 235
rect 1745 189 1801 201
rect 1901 779 1957 791
rect 1901 745 1912 779
rect 1946 745 1957 779
rect 1901 711 1957 745
rect 1901 677 1912 711
rect 1946 677 1957 711
rect 1901 643 1957 677
rect 1901 609 1912 643
rect 1946 609 1957 643
rect 1901 575 1957 609
rect 1901 541 1912 575
rect 1946 541 1957 575
rect 1901 507 1957 541
rect 1901 473 1912 507
rect 1946 473 1957 507
rect 1901 439 1957 473
rect 1901 405 1912 439
rect 1946 405 1957 439
rect 1901 371 1957 405
rect 1901 337 1912 371
rect 1946 337 1957 371
rect 1901 303 1957 337
rect 1901 269 1912 303
rect 1946 269 1957 303
rect 1901 235 1957 269
rect 1901 201 1912 235
rect 1946 201 1957 235
rect 1901 189 1957 201
rect 2057 779 2117 791
rect 2057 745 2068 779
rect 2102 745 2117 779
rect 2057 711 2117 745
rect 2057 677 2068 711
rect 2102 677 2117 711
rect 2057 643 2117 677
rect 2057 609 2068 643
rect 2102 609 2117 643
rect 2057 575 2117 609
rect 2057 541 2068 575
rect 2102 541 2117 575
rect 2057 507 2117 541
rect 2057 473 2068 507
rect 2102 473 2117 507
rect 2057 439 2117 473
rect 2057 405 2068 439
rect 2102 405 2117 439
rect 2057 371 2117 405
rect 2057 337 2068 371
rect 2102 337 2117 371
rect 2057 303 2117 337
rect 2057 269 2068 303
rect 2102 269 2117 303
rect 2057 235 2117 269
rect 2057 201 2068 235
rect 2102 201 2117 235
rect 2057 189 2117 201
<< mvndiffc >>
rect 196 745 230 779
rect 196 677 230 711
rect 196 609 230 643
rect 196 541 230 575
rect 196 473 230 507
rect 196 405 230 439
rect 196 337 230 371
rect 196 269 230 303
rect 196 201 230 235
rect 352 745 386 779
rect 352 677 386 711
rect 352 609 386 643
rect 352 541 386 575
rect 352 473 386 507
rect 352 405 386 439
rect 352 337 386 371
rect 352 269 386 303
rect 352 201 386 235
rect 508 745 542 779
rect 508 677 542 711
rect 508 609 542 643
rect 508 541 542 575
rect 508 473 542 507
rect 508 405 542 439
rect 508 337 542 371
rect 508 269 542 303
rect 508 201 542 235
rect 664 745 698 779
rect 664 677 698 711
rect 664 609 698 643
rect 664 541 698 575
rect 664 473 698 507
rect 664 405 698 439
rect 664 337 698 371
rect 664 269 698 303
rect 664 201 698 235
rect 820 745 854 779
rect 820 677 854 711
rect 820 609 854 643
rect 820 541 854 575
rect 820 473 854 507
rect 820 405 854 439
rect 820 337 854 371
rect 820 269 854 303
rect 820 201 854 235
rect 976 745 1010 779
rect 976 677 1010 711
rect 976 609 1010 643
rect 976 541 1010 575
rect 976 473 1010 507
rect 976 405 1010 439
rect 976 337 1010 371
rect 976 269 1010 303
rect 976 201 1010 235
rect 1132 745 1166 779
rect 1132 677 1166 711
rect 1132 609 1166 643
rect 1132 541 1166 575
rect 1132 473 1166 507
rect 1132 405 1166 439
rect 1132 337 1166 371
rect 1132 269 1166 303
rect 1132 201 1166 235
rect 1288 745 1322 779
rect 1288 677 1322 711
rect 1288 609 1322 643
rect 1288 541 1322 575
rect 1288 473 1322 507
rect 1288 405 1322 439
rect 1288 337 1322 371
rect 1288 269 1322 303
rect 1288 201 1322 235
rect 1444 745 1478 779
rect 1444 677 1478 711
rect 1444 609 1478 643
rect 1444 541 1478 575
rect 1444 473 1478 507
rect 1444 405 1478 439
rect 1444 337 1478 371
rect 1444 269 1478 303
rect 1444 201 1478 235
rect 1600 745 1634 779
rect 1600 677 1634 711
rect 1600 609 1634 643
rect 1600 541 1634 575
rect 1600 473 1634 507
rect 1600 405 1634 439
rect 1600 337 1634 371
rect 1600 269 1634 303
rect 1600 201 1634 235
rect 1756 745 1790 779
rect 1756 677 1790 711
rect 1756 609 1790 643
rect 1756 541 1790 575
rect 1756 473 1790 507
rect 1756 405 1790 439
rect 1756 337 1790 371
rect 1756 269 1790 303
rect 1756 201 1790 235
rect 1912 745 1946 779
rect 1912 677 1946 711
rect 1912 609 1946 643
rect 1912 541 1946 575
rect 1912 473 1946 507
rect 1912 405 1946 439
rect 1912 337 1946 371
rect 1912 269 1946 303
rect 1912 201 1946 235
rect 2068 745 2102 779
rect 2068 677 2102 711
rect 2068 609 2102 643
rect 2068 541 2102 575
rect 2068 473 2102 507
rect 2068 405 2102 439
rect 2068 337 2102 371
rect 2068 269 2102 303
rect 2068 201 2102 235
<< mvpsubdiff >>
rect 41 779 181 791
rect 41 201 60 779
rect 162 201 181 779
rect 41 189 181 201
rect 2117 779 2257 791
rect 2117 201 2136 779
rect 2238 201 2257 779
rect 2117 189 2257 201
<< mvpsubdiffcont >>
rect 60 201 162 779
rect 2136 201 2238 779
<< poly >>
rect 383 959 1915 980
rect 190 867 341 883
rect 190 833 206 867
rect 240 833 341 867
rect 383 857 418 959
rect 1880 857 1915 959
rect 383 841 1915 857
rect 1957 867 2108 883
rect 190 817 341 833
rect 241 791 341 817
rect 397 791 497 841
rect 553 791 653 841
rect 709 791 809 841
rect 865 791 965 841
rect 1021 791 1121 841
rect 1177 791 1277 841
rect 1333 791 1433 841
rect 1489 791 1589 841
rect 1645 791 1745 841
rect 1801 791 1901 841
rect 1957 833 2058 867
rect 2092 833 2108 867
rect 1957 817 2108 833
rect 1957 791 2057 817
rect 241 163 341 189
rect 190 147 341 163
rect 190 113 206 147
rect 240 113 341 147
rect 397 139 497 189
rect 553 139 653 189
rect 709 139 809 189
rect 865 139 965 189
rect 1021 139 1121 189
rect 1177 139 1277 189
rect 1333 139 1433 189
rect 1489 139 1589 189
rect 1645 139 1745 189
rect 1801 139 1901 189
rect 1957 163 2057 189
rect 1957 147 2108 163
rect 190 97 341 113
rect 383 123 1915 139
rect 383 21 418 123
rect 1880 21 1915 123
rect 1957 113 2058 147
rect 2092 113 2108 147
rect 1957 97 2108 113
rect 383 0 1915 21
<< polycont >>
rect 206 833 240 867
rect 418 857 1880 959
rect 2058 833 2092 867
rect 206 113 240 147
rect 418 21 1880 123
rect 2058 113 2092 147
<< locali >>
rect 385 961 1913 980
rect 190 867 256 883
rect 190 833 206 867
rect 240 833 256 867
rect 385 855 412 961
rect 1886 855 1913 961
rect 385 843 1913 855
rect 2042 867 2108 883
rect 190 817 256 833
rect 2042 833 2058 867
rect 2092 833 2108 867
rect 2042 817 2108 833
rect 190 795 230 817
rect 2068 795 2108 817
rect 41 779 230 795
rect 41 201 60 779
rect 162 745 196 779
rect 162 711 230 745
rect 162 677 196 711
rect 162 643 230 677
rect 162 609 196 643
rect 162 575 230 609
rect 162 541 196 575
rect 162 507 230 541
rect 162 473 196 507
rect 162 439 230 473
rect 162 405 196 439
rect 162 371 230 405
rect 162 337 196 371
rect 162 303 230 337
rect 162 269 196 303
rect 162 235 230 269
rect 162 201 196 235
rect 41 185 230 201
rect 352 779 386 795
rect 352 711 386 725
rect 352 643 386 653
rect 352 575 386 581
rect 352 507 386 509
rect 352 471 386 473
rect 352 399 386 405
rect 352 327 386 337
rect 352 255 386 269
rect 352 185 386 201
rect 508 779 542 795
rect 508 711 542 725
rect 508 643 542 653
rect 508 575 542 581
rect 508 507 542 509
rect 508 471 542 473
rect 508 399 542 405
rect 508 327 542 337
rect 508 255 542 269
rect 508 185 542 201
rect 664 779 698 795
rect 664 711 698 725
rect 664 643 698 653
rect 664 575 698 581
rect 664 507 698 509
rect 664 471 698 473
rect 664 399 698 405
rect 664 327 698 337
rect 664 255 698 269
rect 664 185 698 201
rect 820 779 854 795
rect 820 711 854 725
rect 820 643 854 653
rect 820 575 854 581
rect 820 507 854 509
rect 820 471 854 473
rect 820 399 854 405
rect 820 327 854 337
rect 820 255 854 269
rect 820 185 854 201
rect 976 779 1010 795
rect 976 711 1010 725
rect 976 643 1010 653
rect 976 575 1010 581
rect 976 507 1010 509
rect 976 471 1010 473
rect 976 399 1010 405
rect 976 327 1010 337
rect 976 255 1010 269
rect 976 185 1010 201
rect 1132 779 1166 795
rect 1132 711 1166 725
rect 1132 643 1166 653
rect 1132 575 1166 581
rect 1132 507 1166 509
rect 1132 471 1166 473
rect 1132 399 1166 405
rect 1132 327 1166 337
rect 1132 255 1166 269
rect 1132 185 1166 201
rect 1288 779 1322 795
rect 1288 711 1322 725
rect 1288 643 1322 653
rect 1288 575 1322 581
rect 1288 507 1322 509
rect 1288 471 1322 473
rect 1288 399 1322 405
rect 1288 327 1322 337
rect 1288 255 1322 269
rect 1288 185 1322 201
rect 1444 779 1478 795
rect 1444 711 1478 725
rect 1444 643 1478 653
rect 1444 575 1478 581
rect 1444 507 1478 509
rect 1444 471 1478 473
rect 1444 399 1478 405
rect 1444 327 1478 337
rect 1444 255 1478 269
rect 1444 185 1478 201
rect 1600 779 1634 795
rect 1600 711 1634 725
rect 1600 643 1634 653
rect 1600 575 1634 581
rect 1600 507 1634 509
rect 1600 471 1634 473
rect 1600 399 1634 405
rect 1600 327 1634 337
rect 1600 255 1634 269
rect 1600 185 1634 201
rect 1756 779 1790 795
rect 1756 711 1790 725
rect 1756 643 1790 653
rect 1756 575 1790 581
rect 1756 507 1790 509
rect 1756 471 1790 473
rect 1756 399 1790 405
rect 1756 327 1790 337
rect 1756 255 1790 269
rect 1756 185 1790 201
rect 1912 779 1946 795
rect 1912 711 1946 725
rect 1912 643 1946 653
rect 1912 575 1946 581
rect 1912 507 1946 509
rect 1912 471 1946 473
rect 1912 399 1946 405
rect 1912 327 1946 337
rect 1912 255 1946 269
rect 1912 185 1946 201
rect 2068 779 2257 795
rect 2102 745 2136 779
rect 2068 711 2136 745
rect 2102 677 2136 711
rect 2068 643 2136 677
rect 2102 609 2136 643
rect 2068 575 2136 609
rect 2102 541 2136 575
rect 2068 507 2136 541
rect 2102 473 2136 507
rect 2068 439 2136 473
rect 2102 405 2136 439
rect 2068 371 2136 405
rect 2102 337 2136 371
rect 2068 303 2136 337
rect 2102 269 2136 303
rect 2068 235 2136 269
rect 2102 201 2136 235
rect 2238 201 2257 779
rect 2068 185 2257 201
rect 190 163 230 185
rect 2068 163 2108 185
rect 190 147 256 163
rect 190 113 206 147
rect 240 113 256 147
rect 2042 147 2108 163
rect 190 97 256 113
rect 385 125 1913 137
rect 385 19 412 125
rect 1886 19 1913 125
rect 2042 113 2058 147
rect 2092 113 2108 147
rect 2042 97 2108 113
rect 385 0 1913 19
<< viali >>
rect 412 959 1886 961
rect 412 857 418 959
rect 418 857 1880 959
rect 1880 857 1886 959
rect 412 855 1886 857
rect 60 725 94 759
rect 60 653 94 687
rect 60 581 94 615
rect 60 509 94 543
rect 60 437 94 471
rect 60 365 94 399
rect 60 293 94 327
rect 60 221 94 255
rect 352 745 386 759
rect 352 725 386 745
rect 352 677 386 687
rect 352 653 386 677
rect 352 609 386 615
rect 352 581 386 609
rect 352 541 386 543
rect 352 509 386 541
rect 352 439 386 471
rect 352 437 386 439
rect 352 371 386 399
rect 352 365 386 371
rect 352 303 386 327
rect 352 293 386 303
rect 352 235 386 255
rect 352 221 386 235
rect 508 745 542 759
rect 508 725 542 745
rect 508 677 542 687
rect 508 653 542 677
rect 508 609 542 615
rect 508 581 542 609
rect 508 541 542 543
rect 508 509 542 541
rect 508 439 542 471
rect 508 437 542 439
rect 508 371 542 399
rect 508 365 542 371
rect 508 303 542 327
rect 508 293 542 303
rect 508 235 542 255
rect 508 221 542 235
rect 664 745 698 759
rect 664 725 698 745
rect 664 677 698 687
rect 664 653 698 677
rect 664 609 698 615
rect 664 581 698 609
rect 664 541 698 543
rect 664 509 698 541
rect 664 439 698 471
rect 664 437 698 439
rect 664 371 698 399
rect 664 365 698 371
rect 664 303 698 327
rect 664 293 698 303
rect 664 235 698 255
rect 664 221 698 235
rect 820 745 854 759
rect 820 725 854 745
rect 820 677 854 687
rect 820 653 854 677
rect 820 609 854 615
rect 820 581 854 609
rect 820 541 854 543
rect 820 509 854 541
rect 820 439 854 471
rect 820 437 854 439
rect 820 371 854 399
rect 820 365 854 371
rect 820 303 854 327
rect 820 293 854 303
rect 820 235 854 255
rect 820 221 854 235
rect 976 745 1010 759
rect 976 725 1010 745
rect 976 677 1010 687
rect 976 653 1010 677
rect 976 609 1010 615
rect 976 581 1010 609
rect 976 541 1010 543
rect 976 509 1010 541
rect 976 439 1010 471
rect 976 437 1010 439
rect 976 371 1010 399
rect 976 365 1010 371
rect 976 303 1010 327
rect 976 293 1010 303
rect 976 235 1010 255
rect 976 221 1010 235
rect 1132 745 1166 759
rect 1132 725 1166 745
rect 1132 677 1166 687
rect 1132 653 1166 677
rect 1132 609 1166 615
rect 1132 581 1166 609
rect 1132 541 1166 543
rect 1132 509 1166 541
rect 1132 439 1166 471
rect 1132 437 1166 439
rect 1132 371 1166 399
rect 1132 365 1166 371
rect 1132 303 1166 327
rect 1132 293 1166 303
rect 1132 235 1166 255
rect 1132 221 1166 235
rect 1288 745 1322 759
rect 1288 725 1322 745
rect 1288 677 1322 687
rect 1288 653 1322 677
rect 1288 609 1322 615
rect 1288 581 1322 609
rect 1288 541 1322 543
rect 1288 509 1322 541
rect 1288 439 1322 471
rect 1288 437 1322 439
rect 1288 371 1322 399
rect 1288 365 1322 371
rect 1288 303 1322 327
rect 1288 293 1322 303
rect 1288 235 1322 255
rect 1288 221 1322 235
rect 1444 745 1478 759
rect 1444 725 1478 745
rect 1444 677 1478 687
rect 1444 653 1478 677
rect 1444 609 1478 615
rect 1444 581 1478 609
rect 1444 541 1478 543
rect 1444 509 1478 541
rect 1444 439 1478 471
rect 1444 437 1478 439
rect 1444 371 1478 399
rect 1444 365 1478 371
rect 1444 303 1478 327
rect 1444 293 1478 303
rect 1444 235 1478 255
rect 1444 221 1478 235
rect 1600 745 1634 759
rect 1600 725 1634 745
rect 1600 677 1634 687
rect 1600 653 1634 677
rect 1600 609 1634 615
rect 1600 581 1634 609
rect 1600 541 1634 543
rect 1600 509 1634 541
rect 1600 439 1634 471
rect 1600 437 1634 439
rect 1600 371 1634 399
rect 1600 365 1634 371
rect 1600 303 1634 327
rect 1600 293 1634 303
rect 1600 235 1634 255
rect 1600 221 1634 235
rect 1756 745 1790 759
rect 1756 725 1790 745
rect 1756 677 1790 687
rect 1756 653 1790 677
rect 1756 609 1790 615
rect 1756 581 1790 609
rect 1756 541 1790 543
rect 1756 509 1790 541
rect 1756 439 1790 471
rect 1756 437 1790 439
rect 1756 371 1790 399
rect 1756 365 1790 371
rect 1756 303 1790 327
rect 1756 293 1790 303
rect 1756 235 1790 255
rect 1756 221 1790 235
rect 1912 745 1946 759
rect 1912 725 1946 745
rect 1912 677 1946 687
rect 1912 653 1946 677
rect 1912 609 1946 615
rect 1912 581 1946 609
rect 1912 541 1946 543
rect 1912 509 1946 541
rect 1912 439 1946 471
rect 1912 437 1946 439
rect 1912 371 1946 399
rect 1912 365 1946 371
rect 1912 303 1946 327
rect 1912 293 1946 303
rect 1912 235 1946 255
rect 1912 221 1946 235
rect 2204 725 2238 759
rect 2204 653 2238 687
rect 2204 581 2238 615
rect 2204 509 2238 543
rect 2204 437 2238 471
rect 2204 365 2238 399
rect 2204 293 2238 327
rect 2204 221 2238 255
rect 412 123 1886 125
rect 412 21 418 123
rect 418 21 1880 123
rect 1880 21 1886 123
rect 412 19 1886 21
<< metal1 >>
rect 381 961 1917 980
rect 381 855 412 961
rect 1886 855 1917 961
rect 381 843 1917 855
rect 41 759 100 771
rect 41 725 60 759
rect 94 725 100 759
rect 41 687 100 725
rect 41 653 60 687
rect 94 653 100 687
rect 41 615 100 653
rect 41 581 60 615
rect 94 581 100 615
rect 41 543 100 581
rect 41 509 60 543
rect 94 509 100 543
rect 41 471 100 509
rect 41 437 60 471
rect 94 437 100 471
rect 41 399 100 437
rect 41 365 60 399
rect 94 365 100 399
rect 41 327 100 365
rect 41 293 60 327
rect 94 293 100 327
rect 41 255 100 293
rect 41 221 60 255
rect 94 221 100 255
rect 41 209 100 221
rect 343 759 395 771
rect 343 725 352 759
rect 386 725 395 759
rect 343 687 395 725
rect 343 653 352 687
rect 386 653 395 687
rect 343 615 395 653
rect 343 581 352 615
rect 386 581 395 615
rect 343 543 395 581
rect 343 509 352 543
rect 386 509 395 543
rect 343 471 395 509
rect 343 459 352 471
rect 386 459 395 471
rect 343 399 395 407
rect 343 395 352 399
rect 386 395 395 399
rect 343 331 395 343
rect 343 267 395 279
rect 343 209 395 215
rect 499 765 551 771
rect 499 701 551 713
rect 499 637 551 649
rect 499 581 508 585
rect 542 581 551 585
rect 499 573 551 581
rect 499 509 508 521
rect 542 509 551 521
rect 499 471 551 509
rect 499 437 508 471
rect 542 437 551 471
rect 499 399 551 437
rect 499 365 508 399
rect 542 365 551 399
rect 499 327 551 365
rect 499 293 508 327
rect 542 293 551 327
rect 499 255 551 293
rect 499 221 508 255
rect 542 221 551 255
rect 499 209 551 221
rect 655 759 707 771
rect 655 725 664 759
rect 698 725 707 759
rect 655 687 707 725
rect 655 653 664 687
rect 698 653 707 687
rect 655 615 707 653
rect 655 581 664 615
rect 698 581 707 615
rect 655 543 707 581
rect 655 509 664 543
rect 698 509 707 543
rect 655 471 707 509
rect 655 459 664 471
rect 698 459 707 471
rect 655 399 707 407
rect 655 395 664 399
rect 698 395 707 399
rect 655 331 707 343
rect 655 267 707 279
rect 655 209 707 215
rect 811 765 863 771
rect 811 701 863 713
rect 811 637 863 649
rect 811 581 820 585
rect 854 581 863 585
rect 811 573 863 581
rect 811 509 820 521
rect 854 509 863 521
rect 811 471 863 509
rect 811 437 820 471
rect 854 437 863 471
rect 811 399 863 437
rect 811 365 820 399
rect 854 365 863 399
rect 811 327 863 365
rect 811 293 820 327
rect 854 293 863 327
rect 811 255 863 293
rect 811 221 820 255
rect 854 221 863 255
rect 811 209 863 221
rect 967 759 1019 771
rect 967 725 976 759
rect 1010 725 1019 759
rect 967 687 1019 725
rect 967 653 976 687
rect 1010 653 1019 687
rect 967 615 1019 653
rect 967 581 976 615
rect 1010 581 1019 615
rect 967 543 1019 581
rect 967 509 976 543
rect 1010 509 1019 543
rect 967 471 1019 509
rect 967 459 976 471
rect 1010 459 1019 471
rect 967 399 1019 407
rect 967 395 976 399
rect 1010 395 1019 399
rect 967 331 1019 343
rect 967 267 1019 279
rect 967 209 1019 215
rect 1123 765 1175 771
rect 1123 701 1175 713
rect 1123 637 1175 649
rect 1123 581 1132 585
rect 1166 581 1175 585
rect 1123 573 1175 581
rect 1123 509 1132 521
rect 1166 509 1175 521
rect 1123 471 1175 509
rect 1123 437 1132 471
rect 1166 437 1175 471
rect 1123 399 1175 437
rect 1123 365 1132 399
rect 1166 365 1175 399
rect 1123 327 1175 365
rect 1123 293 1132 327
rect 1166 293 1175 327
rect 1123 255 1175 293
rect 1123 221 1132 255
rect 1166 221 1175 255
rect 1123 209 1175 221
rect 1279 759 1331 771
rect 1279 725 1288 759
rect 1322 725 1331 759
rect 1279 687 1331 725
rect 1279 653 1288 687
rect 1322 653 1331 687
rect 1279 615 1331 653
rect 1279 581 1288 615
rect 1322 581 1331 615
rect 1279 543 1331 581
rect 1279 509 1288 543
rect 1322 509 1331 543
rect 1279 471 1331 509
rect 1279 459 1288 471
rect 1322 459 1331 471
rect 1279 399 1331 407
rect 1279 395 1288 399
rect 1322 395 1331 399
rect 1279 331 1331 343
rect 1279 267 1331 279
rect 1279 209 1331 215
rect 1435 765 1487 771
rect 1435 701 1487 713
rect 1435 637 1487 649
rect 1435 581 1444 585
rect 1478 581 1487 585
rect 1435 573 1487 581
rect 1435 509 1444 521
rect 1478 509 1487 521
rect 1435 471 1487 509
rect 1435 437 1444 471
rect 1478 437 1487 471
rect 1435 399 1487 437
rect 1435 365 1444 399
rect 1478 365 1487 399
rect 1435 327 1487 365
rect 1435 293 1444 327
rect 1478 293 1487 327
rect 1435 255 1487 293
rect 1435 221 1444 255
rect 1478 221 1487 255
rect 1435 209 1487 221
rect 1591 759 1643 771
rect 1591 725 1600 759
rect 1634 725 1643 759
rect 1591 687 1643 725
rect 1591 653 1600 687
rect 1634 653 1643 687
rect 1591 615 1643 653
rect 1591 581 1600 615
rect 1634 581 1643 615
rect 1591 543 1643 581
rect 1591 509 1600 543
rect 1634 509 1643 543
rect 1591 471 1643 509
rect 1591 459 1600 471
rect 1634 459 1643 471
rect 1591 399 1643 407
rect 1591 395 1600 399
rect 1634 395 1643 399
rect 1591 331 1643 343
rect 1591 267 1643 279
rect 1591 209 1643 215
rect 1747 765 1799 771
rect 1747 701 1799 713
rect 1747 637 1799 649
rect 1747 581 1756 585
rect 1790 581 1799 585
rect 1747 573 1799 581
rect 1747 509 1756 521
rect 1790 509 1799 521
rect 1747 471 1799 509
rect 1747 437 1756 471
rect 1790 437 1799 471
rect 1747 399 1799 437
rect 1747 365 1756 399
rect 1790 365 1799 399
rect 1747 327 1799 365
rect 1747 293 1756 327
rect 1790 293 1799 327
rect 1747 255 1799 293
rect 1747 221 1756 255
rect 1790 221 1799 255
rect 1747 209 1799 221
rect 1903 759 1955 771
rect 1903 725 1912 759
rect 1946 725 1955 759
rect 1903 687 1955 725
rect 1903 653 1912 687
rect 1946 653 1955 687
rect 1903 615 1955 653
rect 1903 581 1912 615
rect 1946 581 1955 615
rect 1903 543 1955 581
rect 1903 509 1912 543
rect 1946 509 1955 543
rect 1903 471 1955 509
rect 1903 459 1912 471
rect 1946 459 1955 471
rect 1903 399 1955 407
rect 1903 395 1912 399
rect 1946 395 1955 399
rect 1903 331 1955 343
rect 1903 267 1955 279
rect 1903 209 1955 215
rect 2198 759 2257 771
rect 2198 725 2204 759
rect 2238 725 2257 759
rect 2198 687 2257 725
rect 2198 653 2204 687
rect 2238 653 2257 687
rect 2198 615 2257 653
rect 2198 581 2204 615
rect 2238 581 2257 615
rect 2198 543 2257 581
rect 2198 509 2204 543
rect 2238 509 2257 543
rect 2198 471 2257 509
rect 2198 437 2204 471
rect 2238 437 2257 471
rect 2198 399 2257 437
rect 2198 365 2204 399
rect 2238 365 2257 399
rect 2198 327 2257 365
rect 2198 293 2204 327
rect 2238 293 2257 327
rect 2198 255 2257 293
rect 2198 221 2204 255
rect 2238 221 2257 255
rect 2198 209 2257 221
rect 381 125 1917 137
rect 381 19 412 125
rect 1886 19 1917 125
rect 381 0 1917 19
<< via1 >>
rect 343 437 352 459
rect 352 437 386 459
rect 386 437 395 459
rect 343 407 395 437
rect 343 365 352 395
rect 352 365 386 395
rect 386 365 395 395
rect 343 343 395 365
rect 343 327 395 331
rect 343 293 352 327
rect 352 293 386 327
rect 386 293 395 327
rect 343 279 395 293
rect 343 255 395 267
rect 343 221 352 255
rect 352 221 386 255
rect 386 221 395 255
rect 343 215 395 221
rect 499 759 551 765
rect 499 725 508 759
rect 508 725 542 759
rect 542 725 551 759
rect 499 713 551 725
rect 499 687 551 701
rect 499 653 508 687
rect 508 653 542 687
rect 542 653 551 687
rect 499 649 551 653
rect 499 615 551 637
rect 499 585 508 615
rect 508 585 542 615
rect 542 585 551 615
rect 499 543 551 573
rect 499 521 508 543
rect 508 521 542 543
rect 542 521 551 543
rect 655 437 664 459
rect 664 437 698 459
rect 698 437 707 459
rect 655 407 707 437
rect 655 365 664 395
rect 664 365 698 395
rect 698 365 707 395
rect 655 343 707 365
rect 655 327 707 331
rect 655 293 664 327
rect 664 293 698 327
rect 698 293 707 327
rect 655 279 707 293
rect 655 255 707 267
rect 655 221 664 255
rect 664 221 698 255
rect 698 221 707 255
rect 655 215 707 221
rect 811 759 863 765
rect 811 725 820 759
rect 820 725 854 759
rect 854 725 863 759
rect 811 713 863 725
rect 811 687 863 701
rect 811 653 820 687
rect 820 653 854 687
rect 854 653 863 687
rect 811 649 863 653
rect 811 615 863 637
rect 811 585 820 615
rect 820 585 854 615
rect 854 585 863 615
rect 811 543 863 573
rect 811 521 820 543
rect 820 521 854 543
rect 854 521 863 543
rect 967 437 976 459
rect 976 437 1010 459
rect 1010 437 1019 459
rect 967 407 1019 437
rect 967 365 976 395
rect 976 365 1010 395
rect 1010 365 1019 395
rect 967 343 1019 365
rect 967 327 1019 331
rect 967 293 976 327
rect 976 293 1010 327
rect 1010 293 1019 327
rect 967 279 1019 293
rect 967 255 1019 267
rect 967 221 976 255
rect 976 221 1010 255
rect 1010 221 1019 255
rect 967 215 1019 221
rect 1123 759 1175 765
rect 1123 725 1132 759
rect 1132 725 1166 759
rect 1166 725 1175 759
rect 1123 713 1175 725
rect 1123 687 1175 701
rect 1123 653 1132 687
rect 1132 653 1166 687
rect 1166 653 1175 687
rect 1123 649 1175 653
rect 1123 615 1175 637
rect 1123 585 1132 615
rect 1132 585 1166 615
rect 1166 585 1175 615
rect 1123 543 1175 573
rect 1123 521 1132 543
rect 1132 521 1166 543
rect 1166 521 1175 543
rect 1279 437 1288 459
rect 1288 437 1322 459
rect 1322 437 1331 459
rect 1279 407 1331 437
rect 1279 365 1288 395
rect 1288 365 1322 395
rect 1322 365 1331 395
rect 1279 343 1331 365
rect 1279 327 1331 331
rect 1279 293 1288 327
rect 1288 293 1322 327
rect 1322 293 1331 327
rect 1279 279 1331 293
rect 1279 255 1331 267
rect 1279 221 1288 255
rect 1288 221 1322 255
rect 1322 221 1331 255
rect 1279 215 1331 221
rect 1435 759 1487 765
rect 1435 725 1444 759
rect 1444 725 1478 759
rect 1478 725 1487 759
rect 1435 713 1487 725
rect 1435 687 1487 701
rect 1435 653 1444 687
rect 1444 653 1478 687
rect 1478 653 1487 687
rect 1435 649 1487 653
rect 1435 615 1487 637
rect 1435 585 1444 615
rect 1444 585 1478 615
rect 1478 585 1487 615
rect 1435 543 1487 573
rect 1435 521 1444 543
rect 1444 521 1478 543
rect 1478 521 1487 543
rect 1591 437 1600 459
rect 1600 437 1634 459
rect 1634 437 1643 459
rect 1591 407 1643 437
rect 1591 365 1600 395
rect 1600 365 1634 395
rect 1634 365 1643 395
rect 1591 343 1643 365
rect 1591 327 1643 331
rect 1591 293 1600 327
rect 1600 293 1634 327
rect 1634 293 1643 327
rect 1591 279 1643 293
rect 1591 255 1643 267
rect 1591 221 1600 255
rect 1600 221 1634 255
rect 1634 221 1643 255
rect 1591 215 1643 221
rect 1747 759 1799 765
rect 1747 725 1756 759
rect 1756 725 1790 759
rect 1790 725 1799 759
rect 1747 713 1799 725
rect 1747 687 1799 701
rect 1747 653 1756 687
rect 1756 653 1790 687
rect 1790 653 1799 687
rect 1747 649 1799 653
rect 1747 615 1799 637
rect 1747 585 1756 615
rect 1756 585 1790 615
rect 1790 585 1799 615
rect 1747 543 1799 573
rect 1747 521 1756 543
rect 1756 521 1790 543
rect 1790 521 1799 543
rect 1903 437 1912 459
rect 1912 437 1946 459
rect 1946 437 1955 459
rect 1903 407 1955 437
rect 1903 365 1912 395
rect 1912 365 1946 395
rect 1946 365 1955 395
rect 1903 343 1955 365
rect 1903 327 1955 331
rect 1903 293 1912 327
rect 1912 293 1946 327
rect 1946 293 1955 327
rect 1903 279 1955 293
rect 1903 255 1955 267
rect 1903 221 1912 255
rect 1912 221 1946 255
rect 1946 221 1955 255
rect 1903 215 1955 221
<< metal2 >>
rect 14 765 2284 771
rect 14 713 499 765
rect 551 713 811 765
rect 863 713 1123 765
rect 1175 713 1435 765
rect 1487 713 1747 765
rect 1799 713 2284 765
rect 14 701 2284 713
rect 14 649 499 701
rect 551 649 811 701
rect 863 649 1123 701
rect 1175 649 1435 701
rect 1487 649 1747 701
rect 1799 649 2284 701
rect 14 637 2284 649
rect 14 585 499 637
rect 551 585 811 637
rect 863 585 1123 637
rect 1175 585 1435 637
rect 1487 585 1747 637
rect 1799 585 2284 637
rect 14 573 2284 585
rect 14 521 499 573
rect 551 521 811 573
rect 863 521 1123 573
rect 1175 521 1435 573
rect 1487 521 1747 573
rect 1799 521 2284 573
rect 14 515 2284 521
rect 14 459 2284 465
rect 14 407 343 459
rect 395 407 655 459
rect 707 407 967 459
rect 1019 407 1279 459
rect 1331 407 1591 459
rect 1643 407 1903 459
rect 1955 407 2284 459
rect 14 395 2284 407
rect 14 343 343 395
rect 395 343 655 395
rect 707 343 967 395
rect 1019 343 1279 395
rect 1331 343 1591 395
rect 1643 343 1903 395
rect 1955 343 2284 395
rect 14 331 2284 343
rect 14 279 343 331
rect 395 279 655 331
rect 707 279 967 331
rect 1019 279 1279 331
rect 1331 279 1591 331
rect 1643 279 1903 331
rect 1955 279 2284 331
rect 14 267 2284 279
rect 14 215 343 267
rect 395 215 655 267
rect 707 215 967 267
rect 1019 215 1279 267
rect 1331 215 1591 267
rect 1643 215 1903 267
rect 1955 215 2284 267
rect 14 209 2284 215
<< labels >>
flabel metal1 s 1098 85 1195 120 0 FreeSans 200 0 0 0 GATE
port 2 nsew
flabel metal2 s 36 313 66 417 0 FreeSans 400 90 0 0 SOURCE
port 3 nsew
flabel metal2 s 35 602 70 699 0 FreeSans 400 270 0 0 DRAIN
port 1 nsew
flabel comment s 1617 490 1617 490 0 FreeSans 300 0 0 0 S
flabel comment s 1929 490 1929 490 0 FreeSans 300 0 0 0 S
flabel comment s 1773 490 1773 490 0 FreeSans 300 0 0 0 D
flabel comment s 1617 490 1617 490 0 FreeSans 300 0 0 0 S
flabel comment s 1461 490 1461 490 0 FreeSans 300 0 0 0 D
flabel comment s 1773 490 1773 490 0 FreeSans 300 0 0 0 S
flabel comment s 1461 490 1461 490 0 FreeSans 300 0 0 0 S
flabel comment s 993 490 993 490 0 FreeSans 300 0 0 0 S
flabel comment s 1149 490 1149 490 0 FreeSans 300 0 0 0 S
flabel comment s 1305 490 1305 490 0 FreeSans 300 0 0 0 S
flabel comment s 993 490 993 490 0 FreeSans 300 0 0 0 D
flabel comment s 1149 490 1149 490 0 FreeSans 300 0 0 0 S
flabel comment s 1305 490 1305 490 0 FreeSans 300 0 0 0 D
flabel comment s 681 490 681 490 0 FreeSans 300 0 0 0 S
flabel comment s 837 490 837 490 0 FreeSans 300 0 0 0 S
flabel comment s 681 490 681 490 0 FreeSans 300 0 0 0 S
flabel comment s 837 490 837 490 0 FreeSans 300 0 0 0 D
flabel comment s 369 490 369 490 0 FreeSans 300 0 0 0 S
flabel comment s 369 490 369 490 0 FreeSans 300 0 0 0 S
flabel comment s 525 490 525 490 0 FreeSans 300 0 0 0 S
flabel comment s 525 490 525 490 0 FreeSans 300 0 0 0 D
flabel comment s 2002 480 2002 480 0 FreeSans 400 90 0 0 dummy_poly
flabel comment s 286 493 286 493 0 FreeSans 400 90 0 0 dummy_poly
flabel metal1 s 2198 469 2257 499 0 FreeSans 200 90 0 0 SUBSTRATE
port 4 nsew
flabel metal1 s 41 466 100 496 0 FreeSans 200 90 0 0 SUBSTRATE
port 4 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 8765500
string GDS_START 8724470
<< end >>
