magic
tech sky130A
magscale 1 2
timestamp 1658880696
<< nwell >>
rect 98 125 251 221
<< pwell >>
rect -100 79 70 251
rect 282 79 452 251
rect -100 -19 452 79
<< nmos >>
rect 7 165 37 193
rect 315 165 345 193
rect -57 19 -27 61
rect 379 19 409 61
<< npd >>
rect 122 19 152 61
rect 200 19 230 61
<< npass >>
rect 29 19 59 47
rect 293 19 323 47
<< ppu >>
rect 122 155 152 183
rect 200 155 230 183
<< ndiff >>
rect -11 165 7 193
rect 37 165 55 193
rect 297 165 315 193
rect 345 165 364 193
rect -85 19 -57 61
rect -27 47 -2 61
rect 97 51 122 61
rect -27 19 29 47
rect 59 19 93 47
tri 107 44 114 51 ne
rect 114 19 122 51
rect 152 19 200 61
rect 230 51 255 61
rect 230 19 238 51
rect 354 47 379 61
rect 259 19 293 47
rect 323 19 379 47
rect 409 19 437 61
rect 66 -5 93 19
rect 160 -3 192 19
rect 160 -5 162 -3
rect 190 -5 192 -3
rect 259 -5 286 19
rect 66 -19 160 -5
rect 192 -19 286 -5
<< pdiff >>
rect 160 205 162 207
rect 190 205 192 207
rect 160 183 192 205
rect 113 155 122 183
rect 152 155 200 183
rect 230 155 239 183
tri 239 155 251 167 sw
<< ndiffc >>
rect -26 165 -11 193
rect 55 165 70 193
rect 282 165 297 193
rect 364 165 379 194
rect -100 19 -85 61
rect 97 44 107 51
tri 107 44 114 51 sw
rect 97 19 114 44
rect 238 19 255 51
rect 437 19 452 61
rect 160 -19 192 -5
<< pdiffc >>
rect 160 207 192 221
rect 98 155 113 183
rect 239 167 251 183
tri 239 155 251 167 ne
<< psubdiffcont >>
rect 162 -5 190 -3
<< nsubdiffcont >>
rect 162 205 190 207
<< poly >>
rect -100 221 452 251
rect 7 193 37 221
rect 122 183 152 205
rect 200 183 230 205
rect 315 193 345 221
rect 7 143 37 165
rect 122 122 152 155
rect -57 61 -27 83
rect 29 61 44 95
rect 122 61 152 88
rect 200 122 230 155
rect 315 143 345 165
rect 200 61 230 88
rect 308 61 323 95
rect 379 61 409 83
rect 29 47 59 61
rect 293 47 323 61
rect -57 -3 -27 19
rect 29 -3 59 19
rect 122 -3 152 19
rect 200 -3 230 19
rect 293 -3 323 19
rect 379 -3 409 19
<< polycont >>
rect -57 83 -27 117
rect 44 61 74 95
rect 122 88 152 122
rect 200 88 230 122
rect 278 61 308 95
rect 379 83 409 117
<< corelocali >>
rect -100 61 -85 251
tri -20 215 2 237 se
rect 2 230 17 251
tri 2 215 17 230 nw
rect 336 230 351 251
tri -26 209 -20 215 se
rect -20 209 -11 215
rect -26 193 -11 209
tri -11 202 2 215 nw
rect 143 207 160 221
rect 192 207 209 221
tri 336 215 351 230 ne
tri 351 215 373 237 sw
rect -26 157 -11 165
rect 55 193 115 207
rect 70 183 115 193
rect 70 165 98 183
tri -26 142 -11 157 ne
tri -11 142 11 164 sw
rect 55 155 98 165
rect 113 179 115 183
rect 237 193 297 207
tri 351 202 364 215 ne
rect 364 209 373 215
tri 373 209 379 215 sw
rect 237 183 282 193
rect 113 155 187 179
rect 55 151 187 155
tri 187 151 215 179 sw
rect 237 169 239 183
tri 237 167 239 169 ne
rect 251 165 282 183
rect 251 155 297 165
rect 364 194 379 209
tri -11 130 1 142 ne
rect 1 137 11 142
tri 11 137 16 142 sw
rect -100 -19 -85 19
rect 1 -19 16 137
rect 55 95 83 151
tri 175 133 193 151 ne
rect 193 131 215 151
tri 215 131 235 151 sw
tri 251 137 269 155 ne
rect 74 61 83 95
rect 117 122 159 123
rect 117 88 122 122
rect 152 88 159 122
rect 117 79 159 88
rect 193 122 235 131
rect 193 88 200 122
rect 230 88 235 122
rect 193 83 235 88
rect 269 95 297 155
tri 342 142 364 164 se
rect 364 157 379 165
tri 364 142 379 157 nw
tri 336 136 342 142 se
rect 342 136 351 142
rect 55 51 83 61
tri 83 51 107 75 sw
rect 55 19 97 51
tri 114 43 115 44 sw
rect 114 19 115 43
tri 117 42 154 79 ne
rect 154 51 159 79
tri 159 51 185 77 sw
rect 269 61 278 95
rect 269 51 297 61
rect 154 42 238 51
tri 154 23 173 42 ne
rect 173 23 238 42
rect 55 -3 115 19
rect 237 19 238 23
rect 255 19 297 51
rect 237 -3 297 19
rect 143 -19 160 -5
rect 192 -19 209 -5
rect 336 -19 351 136
tri 351 129 364 142 nw
rect 437 61 452 251
rect 437 -19 452 19
<< viali >>
rect 160 207 192 221
rect 160 -19 192 -5
<< metal1 >>
rect -100 207 160 221
rect 192 207 452 221
rect -100 -19 160 -5
rect 192 -19 452 -5
<< labels >>
rlabel poly -100 221 452 251 1 WWL
port 1 ew signal input
rlabel locali 379 83 409 117 1 RWL
port 2 ew signal input
rlabel locali -57 83 -27 117 1 RWL
port 3 ew signal input
rlabel locali 364 165 379 194 1 WBL
port 4 ns signal input
rlabel locali -26 165 -11 193 1 WBLb
port 5 ns signal input
rlabel locali 437 19 452 61 1 RBL0
port 6 ns signal output
rlabel locali -100 19 -85 61 1 RBL1
port 7 ns signal output
rlabel metal1 160 207 192 221 1 VDD
port 8 ew power bidirectional abutment
rlabel metal1 160 -19 192 -5 7 GND
port 9 ew ground bidirectional abutment
rlabel polycont 122 88 152 122 1 junc0
rlabel polycont 200 88 230 122 1 junc1
rlabel ndiff -27 19 29 47 1 RWL1_junc
rlabel ndiff 323 19 379 47 1 RWL0_junc
<< end >>
