VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO toysram_bit
  CLASS BLOCK ;
  FOREIGN toysram_bit ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.750 BY 2.500 ;
  PIN WWL
    ANTENNAGATEAREA 0.147000 ;
    PORT
      LAYER li1 ;
        RECT 0.110 1.940 0.450 2.280 ;
        RECT 0.110 0.400 0.450 0.740 ;
      LAYER mcon ;
        RECT 0.195 2.025 0.365 2.195 ;
        RECT 0.195 0.485 0.365 0.655 ;
      LAYER met1 ;
        RECT 0.110 1.940 0.450 2.280 ;
        RECT 0.110 0.400 0.450 0.740 ;
      LAYER via ;
        RECT 0.140 1.970 0.420 2.250 ;
        RECT 0.140 0.430 0.420 0.710 ;
      LAYER met2 ;
        RECT 0.000 1.940 0.560 2.280 ;
        RECT 0.110 0.400 0.450 1.940 ;
    END
  END WWL
  PIN WBL
    ANTENNADIFFAREA 0.181300 ;
    PORT
      LAYER li1 ;
        RECT 2.315 2.160 2.655 2.500 ;
      LAYER mcon ;
        RECT 2.400 2.245 2.570 2.415 ;
      LAYER met1 ;
        RECT 1.960 2.160 2.800 2.500 ;
    END
  END WBL
  PIN GND
    ANTENNADIFFAREA 0.380800 ;
    PORT
      LAYER li1 ;
        RECT 2.315 1.120 2.655 1.460 ;
        RECT 3.505 1.120 3.845 1.460 ;
      LAYER mcon ;
        RECT 2.400 1.205 2.570 1.375 ;
        RECT 3.590 1.205 3.760 1.375 ;
      LAYER met1 ;
        RECT 2.100 1.120 4.750 1.460 ;
    END
  END GND
  PIN VDD
    ANTENNADIFFAREA 0.142800 ;
    PORT
      LAYER li1 ;
        RECT 1.300 1.120 1.640 1.460 ;
      LAYER mcon ;
        RECT 1.385 1.205 1.555 1.375 ;
      LAYER met1 ;
        RECT 1.050 1.120 1.890 1.460 ;
    END
  END VDD
  PIN WBLb
    ANTENNADIFFAREA 0.196000 ;
    PORT
      LAYER li1 ;
        RECT 2.315 0.060 2.655 0.400 ;
      LAYER mcon ;
        RECT 2.400 0.145 2.570 0.315 ;
      LAYER met1 ;
        RECT 1.820 0.060 2.800 0.400 ;
    END
  END WBLb
  PIN RBL0
    ANTENNADIFFAREA 0.245700 ;
    PORT
      LAYER li1 ;
        RECT 3.505 2.160 3.845 2.500 ;
      LAYER mcon ;
        RECT 3.590 2.245 3.760 2.415 ;
      LAYER met1 ;
        RECT 3.220 2.160 4.130 2.500 ;
    END
  END RBL0
  PIN RBL1
    ANTENNADIFFAREA 0.239400 ;
    PORT
      LAYER li1 ;
        RECT 3.505 0.060 3.845 0.400 ;
      LAYER mcon ;
        RECT 3.590 0.145 3.760 0.315 ;
      LAYER met1 ;
        RECT 3.220 0.060 4.130 0.400 ;
    END
  END RBL1
  PIN RWL0
    ANTENNAGATEAREA 0.094500 ;
    PORT
      LAYER li1 ;
        RECT 4.410 1.895 4.750 2.235 ;
      LAYER mcon ;
        RECT 4.495 1.980 4.665 2.150 ;
      LAYER met1 ;
        RECT 4.410 1.895 4.750 2.235 ;
      LAYER via ;
        RECT 4.440 1.925 4.720 2.205 ;
      LAYER met2 ;
        RECT 4.410 1.895 4.750 2.235 ;
    END
  END RWL0
  PIN RWL1
    ANTENNAGATEAREA 0.094500 ;
    PORT
      LAYER li1 ;
        RECT 4.410 0.315 4.750 0.655 ;
      LAYER mcon ;
        RECT 4.495 0.400 4.665 0.570 ;
      LAYER met1 ;
        RECT 4.410 0.315 4.750 0.655 ;
      LAYER via ;
        RECT 4.440 0.345 4.720 0.625 ;
      LAYER met2 ;
        RECT 4.410 0.315 4.750 0.655 ;
    END
  END RWL1
  OBS
      LAYER pwell ;
        RECT 3.230 2.630 4.120 2.650 ;
      LAYER nwell ;
        RECT 1.050 0.445 1.890 2.105 ;
      LAYER pwell ;
        RECT 2.110 -0.110 4.120 2.630 ;
        RECT 2.110 -0.130 2.860 -0.110 ;
      LAYER li1 ;
        RECT 0.460 1.375 0.800 1.715 ;
        RECT 0.980 1.680 3.080 1.850 ;
        RECT 0.630 0.890 0.800 1.375 ;
        RECT 2.910 1.225 3.080 1.680 ;
        RECT 0.630 0.720 2.730 0.890 ;
        RECT 2.910 0.885 3.250 1.225 ;
  END
END toysram_bit
END LIBRARY

