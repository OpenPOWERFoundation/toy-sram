VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS

MACRO sky130_fd_sc_hdll__nand2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nand2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.990 1.075 1.375 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.277500 ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.055 0.430 1.325 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.085 0.395 0.885 ;
        RECT 0.000 -0.085 1.840 0.085 ;
      LAYER mcon ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.025 0.105 1.475 1.015 ;
        RECT 0.140 -0.085 0.310 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.635 1.840 2.805 ;
        RECT 0.085 1.495 0.365 2.635 ;
        RECT 1.135 1.495 1.395 2.635 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.491500 ;
    PORT
      LAYER li1 ;
        RECT 0.535 1.485 0.915 2.465 ;
        RECT 0.650 0.885 0.820 1.485 ;
        RECT 0.650 0.255 1.395 0.885 ;
    END
  END Y
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand2_1
MACRO local_eval
  CLASS BLOCK ;
  FOREIGN local_eval ;
  ORIGIN 0.270 0.150 ;
  SIZE 2.220 BY 3.200 ;
  OBS
      LAYER nwell ;
        RECT -0.270 1.395 1.950 3.000 ;
      LAYER pwell ;
        RECT -0.055 0.195 1.395 1.105 ;
        RECT 0.060 0.005 0.230 0.195 ;
      LAYER li1 ;
        RECT -0.080 2.725 1.760 2.895 ;
        RECT 0.005 1.585 0.285 2.725 ;
        RECT 0.455 1.575 0.835 2.555 ;
        RECT 1.055 1.585 1.315 2.725 ;
        RECT 0.015 1.145 0.350 1.415 ;
        RECT 0.570 0.975 0.740 1.575 ;
        RECT 0.910 1.165 1.295 1.415 ;
        RECT 0.005 0.175 0.315 0.975 ;
        RECT 0.570 0.345 1.315 0.975 ;
        RECT -0.080 0.005 1.760 0.175 ;
      LAYER mcon ;
        RECT 0.065 2.725 0.235 2.895 ;
        RECT 0.525 2.725 0.695 2.895 ;
        RECT 0.985 2.725 1.155 2.895 ;
        RECT 1.445 2.725 1.615 2.895 ;
        RECT 0.065 0.005 0.235 0.175 ;
        RECT 0.525 0.005 0.695 0.175 ;
        RECT 0.985 0.005 1.155 0.175 ;
        RECT 1.445 0.005 1.615 0.175 ;
      LAYER met1 ;
        RECT -0.080 2.570 1.760 3.050 ;
        RECT -0.080 -0.150 1.760 0.330 ;
  END
END local_eval
END LIBRARY

