magic
tech sky130A
magscale 1 2
timestamp 1656020757
<< error_s >>
rect 15 524 28 540
rect 117 538 130 540
rect 83 524 98 538
rect 107 524 137 538
rect 198 536 351 582
rect 180 524 372 536
rect 415 524 445 538
rect 451 524 464 540
rect 552 524 565 540
rect 595 524 608 540
rect 697 538 710 540
rect 663 524 678 538
rect 687 524 717 538
rect 778 536 931 582
rect 760 524 952 536
rect 995 524 1025 538
rect 1031 524 1044 540
rect 1132 524 1145 540
rect 1175 524 1188 540
rect 1277 538 1290 540
rect 1243 524 1258 538
rect 1267 524 1297 538
rect 1358 536 1511 582
rect 1340 524 1532 536
rect 1575 524 1605 538
rect 1611 524 1624 540
rect 1712 524 1725 540
rect 1755 524 1768 540
rect 1857 538 1870 540
rect 1823 524 1838 538
rect 1847 524 1877 538
rect 1938 536 2091 582
rect 1920 524 2112 536
rect 2155 524 2185 538
rect 2191 524 2204 540
rect 2292 524 2305 540
rect 2335 524 2348 540
rect 2437 538 2450 540
rect 2403 524 2418 538
rect 2427 524 2457 538
rect 2518 536 2671 582
rect 2500 524 2692 536
rect 2735 524 2765 538
rect 2771 524 2784 540
rect 2872 524 2885 540
rect 2915 524 2928 540
rect 3017 538 3030 540
rect 2983 524 2998 538
rect 3007 524 3037 538
rect 3098 536 3251 582
rect 3080 524 3272 536
rect 3315 524 3345 538
rect 3351 524 3364 540
rect 3452 524 3465 540
rect 3495 524 3508 540
rect 3597 538 3610 540
rect 3563 524 3578 538
rect 3587 524 3617 538
rect 3678 536 3831 582
rect 3660 524 3852 536
rect 3895 524 3925 538
rect 3931 524 3944 540
rect 4032 524 4045 540
rect 4075 524 4088 540
rect 4177 538 4190 540
rect 4143 524 4158 538
rect 4167 524 4197 538
rect 4258 536 4411 582
rect 4240 524 4432 536
rect 4475 524 4505 538
rect 4511 524 4524 540
rect 4612 524 4625 540
rect 0 510 4625 524
rect 15 406 28 510
rect 73 488 74 498
rect 89 488 102 498
rect 73 484 102 488
rect 107 484 137 510
rect 155 496 171 498
rect 243 496 296 510
rect 244 494 308 496
rect 351 494 366 510
rect 415 507 445 510
rect 415 504 451 507
rect 381 496 397 498
rect 155 484 170 488
rect 73 482 170 484
rect 198 482 366 494
rect 382 484 397 488
rect 415 485 454 504
rect 473 498 480 499
rect 479 491 480 498
rect 463 488 464 491
rect 479 488 492 491
rect 415 484 445 485
rect 454 484 460 485
rect 463 484 492 488
rect 382 483 492 484
rect 382 482 498 483
rect 57 474 108 482
rect 57 462 82 474
rect 89 462 108 474
rect 139 474 189 482
rect 139 466 155 474
rect 162 472 189 474
rect 198 472 419 482
rect 162 462 419 472
rect 448 474 498 482
rect 448 465 464 474
rect 57 454 108 462
rect 155 454 419 462
rect 445 462 464 465
rect 471 462 498 474
rect 445 454 498 462
rect 73 446 74 454
rect 89 446 102 454
rect 73 438 89 446
rect 70 431 89 434
rect 70 422 92 431
rect 43 412 92 422
rect 43 406 73 412
rect 92 407 97 412
rect 15 390 89 406
rect 107 398 137 454
rect 172 444 380 454
rect 415 450 460 454
rect 463 453 464 454
rect 479 453 492 454
rect 198 414 387 444
rect 213 411 387 414
rect 206 408 387 411
rect 15 388 28 390
rect 43 388 77 390
rect 15 372 89 388
rect 116 384 129 398
rect 144 384 160 400
rect 206 395 217 408
rect -1 350 0 366
rect 15 350 28 372
rect 43 350 73 372
rect 116 368 178 384
rect 206 377 217 393
rect 222 388 232 408
rect 242 388 256 408
rect 259 395 268 408
rect 284 395 293 408
rect 222 377 256 388
rect 259 377 268 393
rect 284 377 293 393
rect 300 388 310 408
rect 320 388 334 408
rect 335 395 346 408
rect 300 377 334 388
rect 335 377 346 393
rect 392 384 408 400
rect 415 398 445 450
rect 479 446 480 453
rect 464 438 480 446
rect 451 406 464 425
rect 479 406 509 422
rect 451 390 525 406
rect 451 388 464 390
rect 479 388 513 390
rect 116 366 129 368
rect 144 366 178 368
rect 116 350 178 366
rect 222 361 238 364
rect 300 361 330 372
rect 378 368 424 384
rect 451 372 525 388
rect 378 366 412 368
rect 377 350 424 366
rect 451 350 464 372
rect 479 350 509 372
rect 536 350 537 366
rect 552 350 565 510
rect 595 406 608 510
rect 653 488 654 498
rect 669 488 682 498
rect 653 484 682 488
rect 687 484 717 510
rect 735 496 751 498
rect 823 496 876 510
rect 824 494 888 496
rect 931 494 946 510
rect 995 507 1025 510
rect 995 504 1031 507
rect 961 496 977 498
rect 735 484 750 488
rect 653 482 750 484
rect 778 482 946 494
rect 962 484 977 488
rect 995 485 1034 504
rect 1053 498 1060 499
rect 1059 491 1060 498
rect 1043 488 1044 491
rect 1059 488 1072 491
rect 995 484 1025 485
rect 1034 484 1040 485
rect 1043 484 1072 488
rect 962 483 1072 484
rect 962 482 1078 483
rect 637 474 688 482
rect 637 462 662 474
rect 669 462 688 474
rect 719 474 769 482
rect 719 466 735 474
rect 742 472 769 474
rect 778 472 999 482
rect 742 462 999 472
rect 1028 474 1078 482
rect 1028 465 1044 474
rect 637 454 688 462
rect 735 454 999 462
rect 1025 462 1044 465
rect 1051 462 1078 474
rect 1025 454 1078 462
rect 653 446 654 454
rect 669 446 682 454
rect 653 438 669 446
rect 650 431 669 434
rect 650 422 672 431
rect 623 412 672 422
rect 623 406 653 412
rect 672 407 677 412
rect 595 390 669 406
rect 687 398 717 454
rect 752 444 960 454
rect 995 450 1040 454
rect 1043 453 1044 454
rect 1059 453 1072 454
rect 778 414 967 444
rect 793 411 967 414
rect 786 408 967 411
rect 595 388 608 390
rect 623 388 657 390
rect 595 372 669 388
rect 696 384 709 398
rect 724 384 740 400
rect 786 395 797 408
rect 579 350 580 366
rect 595 350 608 372
rect 623 350 653 372
rect 696 368 758 384
rect 786 377 797 393
rect 802 388 812 408
rect 822 388 836 408
rect 839 395 848 408
rect 864 395 873 408
rect 802 377 836 388
rect 839 377 848 393
rect 864 377 873 393
rect 880 388 890 408
rect 900 388 914 408
rect 915 395 926 408
rect 880 377 914 388
rect 915 377 926 393
rect 972 384 988 400
rect 995 398 1025 450
rect 1059 446 1060 453
rect 1044 438 1060 446
rect 1031 406 1044 425
rect 1059 406 1089 422
rect 1031 390 1105 406
rect 1031 388 1044 390
rect 1059 388 1093 390
rect 696 366 709 368
rect 724 366 758 368
rect 696 350 758 366
rect 802 361 818 364
rect 880 361 910 372
rect 958 368 1004 384
rect 1031 372 1105 388
rect 958 366 992 368
rect 957 350 1004 366
rect 1031 350 1044 372
rect 1059 350 1089 372
rect 1116 350 1117 366
rect 1132 350 1145 510
rect 1175 406 1188 510
rect 1233 488 1234 498
rect 1249 488 1262 498
rect 1233 484 1262 488
rect 1267 484 1297 510
rect 1315 496 1331 498
rect 1403 496 1456 510
rect 1404 494 1468 496
rect 1511 494 1526 510
rect 1575 507 1605 510
rect 1575 504 1611 507
rect 1541 496 1557 498
rect 1315 484 1330 488
rect 1233 482 1330 484
rect 1358 482 1526 494
rect 1542 484 1557 488
rect 1575 485 1614 504
rect 1633 498 1640 499
rect 1639 491 1640 498
rect 1623 488 1624 491
rect 1639 488 1652 491
rect 1575 484 1605 485
rect 1614 484 1620 485
rect 1623 484 1652 488
rect 1542 483 1652 484
rect 1542 482 1658 483
rect 1217 474 1268 482
rect 1217 462 1242 474
rect 1249 462 1268 474
rect 1299 474 1349 482
rect 1299 466 1315 474
rect 1322 472 1349 474
rect 1358 472 1579 482
rect 1322 462 1579 472
rect 1608 474 1658 482
rect 1608 465 1624 474
rect 1217 454 1268 462
rect 1315 454 1579 462
rect 1605 462 1624 465
rect 1631 462 1658 474
rect 1605 454 1658 462
rect 1233 446 1234 454
rect 1249 446 1262 454
rect 1233 438 1249 446
rect 1230 431 1249 434
rect 1230 422 1252 431
rect 1203 412 1252 422
rect 1203 406 1233 412
rect 1252 407 1257 412
rect 1175 390 1249 406
rect 1267 398 1297 454
rect 1332 444 1540 454
rect 1575 450 1620 454
rect 1623 453 1624 454
rect 1639 453 1652 454
rect 1358 414 1547 444
rect 1373 411 1547 414
rect 1366 408 1547 411
rect 1175 388 1188 390
rect 1203 388 1237 390
rect 1175 372 1249 388
rect 1276 384 1289 398
rect 1304 384 1320 400
rect 1366 395 1377 408
rect 1159 350 1160 366
rect 1175 350 1188 372
rect 1203 350 1233 372
rect 1276 368 1338 384
rect 1366 377 1377 393
rect 1382 388 1392 408
rect 1402 388 1416 408
rect 1419 395 1428 408
rect 1444 395 1453 408
rect 1382 377 1416 388
rect 1419 377 1428 393
rect 1444 377 1453 393
rect 1460 388 1470 408
rect 1480 388 1494 408
rect 1495 395 1506 408
rect 1460 377 1494 388
rect 1495 377 1506 393
rect 1552 384 1568 400
rect 1575 398 1605 450
rect 1639 446 1640 453
rect 1624 438 1640 446
rect 1611 406 1624 425
rect 1639 406 1669 422
rect 1611 390 1685 406
rect 1611 388 1624 390
rect 1639 388 1673 390
rect 1276 366 1289 368
rect 1304 366 1338 368
rect 1276 350 1338 366
rect 1382 361 1398 364
rect 1460 361 1490 372
rect 1538 368 1584 384
rect 1611 372 1685 388
rect 1538 366 1572 368
rect 1537 350 1584 366
rect 1611 350 1624 372
rect 1639 350 1669 372
rect 1696 350 1697 366
rect 1712 350 1725 510
rect 1755 406 1768 510
rect 1813 488 1814 498
rect 1829 488 1842 498
rect 1813 484 1842 488
rect 1847 484 1877 510
rect 1895 496 1911 498
rect 1983 496 2036 510
rect 1984 494 2048 496
rect 2091 494 2106 510
rect 2155 507 2185 510
rect 2155 504 2191 507
rect 2121 496 2137 498
rect 1895 484 1910 488
rect 1813 482 1910 484
rect 1938 482 2106 494
rect 2122 484 2137 488
rect 2155 485 2194 504
rect 2213 498 2220 499
rect 2219 491 2220 498
rect 2203 488 2204 491
rect 2219 488 2232 491
rect 2155 484 2185 485
rect 2194 484 2200 485
rect 2203 484 2232 488
rect 2122 483 2232 484
rect 2122 482 2238 483
rect 1797 474 1848 482
rect 1797 462 1822 474
rect 1829 462 1848 474
rect 1879 474 1929 482
rect 1879 466 1895 474
rect 1902 472 1929 474
rect 1938 472 2159 482
rect 1902 462 2159 472
rect 2188 474 2238 482
rect 2188 465 2204 474
rect 1797 454 1848 462
rect 1895 454 2159 462
rect 2185 462 2204 465
rect 2211 462 2238 474
rect 2185 454 2238 462
rect 1813 446 1814 454
rect 1829 446 1842 454
rect 1813 438 1829 446
rect 1810 431 1829 434
rect 1810 422 1832 431
rect 1783 412 1832 422
rect 1783 406 1813 412
rect 1832 407 1837 412
rect 1755 390 1829 406
rect 1847 398 1877 454
rect 1912 444 2120 454
rect 2155 450 2200 454
rect 2203 453 2204 454
rect 2219 453 2232 454
rect 1938 414 2127 444
rect 1953 411 2127 414
rect 1946 408 2127 411
rect 1755 388 1768 390
rect 1783 388 1817 390
rect 1755 372 1829 388
rect 1856 384 1869 398
rect 1884 384 1900 400
rect 1946 395 1957 408
rect 1739 350 1740 366
rect 1755 350 1768 372
rect 1783 350 1813 372
rect 1856 368 1918 384
rect 1946 377 1957 393
rect 1962 388 1972 408
rect 1982 388 1996 408
rect 1999 395 2008 408
rect 2024 395 2033 408
rect 1962 377 1996 388
rect 1999 377 2008 393
rect 2024 377 2033 393
rect 2040 388 2050 408
rect 2060 388 2074 408
rect 2075 395 2086 408
rect 2040 377 2074 388
rect 2075 377 2086 393
rect 2132 384 2148 400
rect 2155 398 2185 450
rect 2219 446 2220 453
rect 2204 438 2220 446
rect 2191 406 2204 425
rect 2219 406 2249 422
rect 2191 390 2265 406
rect 2191 388 2204 390
rect 2219 388 2253 390
rect 1856 366 1869 368
rect 1884 366 1918 368
rect 1856 350 1918 366
rect 1962 361 1978 364
rect 2040 361 2070 372
rect 2118 368 2164 384
rect 2191 372 2265 388
rect 2118 366 2152 368
rect 2117 350 2164 366
rect 2191 350 2204 372
rect 2219 350 2249 372
rect 2276 350 2277 366
rect 2292 350 2305 510
rect 2335 406 2348 510
rect 2393 488 2394 498
rect 2409 488 2422 498
rect 2393 484 2422 488
rect 2427 484 2457 510
rect 2475 496 2491 498
rect 2563 496 2616 510
rect 2564 494 2628 496
rect 2671 494 2686 510
rect 2735 507 2765 510
rect 2735 504 2771 507
rect 2701 496 2717 498
rect 2475 484 2490 488
rect 2393 482 2490 484
rect 2518 482 2686 494
rect 2702 484 2717 488
rect 2735 485 2774 504
rect 2793 498 2800 499
rect 2799 491 2800 498
rect 2783 488 2784 491
rect 2799 488 2812 491
rect 2735 484 2765 485
rect 2774 484 2780 485
rect 2783 484 2812 488
rect 2702 483 2812 484
rect 2702 482 2818 483
rect 2377 474 2428 482
rect 2377 462 2402 474
rect 2409 462 2428 474
rect 2459 474 2509 482
rect 2459 466 2475 474
rect 2482 472 2509 474
rect 2518 472 2739 482
rect 2482 462 2739 472
rect 2768 474 2818 482
rect 2768 465 2784 474
rect 2377 454 2428 462
rect 2475 454 2739 462
rect 2765 462 2784 465
rect 2791 462 2818 474
rect 2765 454 2818 462
rect 2393 446 2394 454
rect 2409 446 2422 454
rect 2393 438 2409 446
rect 2390 431 2409 434
rect 2390 422 2412 431
rect 2363 412 2412 422
rect 2363 406 2393 412
rect 2412 407 2417 412
rect 2335 390 2409 406
rect 2427 398 2457 454
rect 2492 444 2700 454
rect 2735 450 2780 454
rect 2783 453 2784 454
rect 2799 453 2812 454
rect 2518 414 2707 444
rect 2533 411 2707 414
rect 2526 408 2707 411
rect 2335 388 2348 390
rect 2363 388 2397 390
rect 2335 372 2409 388
rect 2436 384 2449 398
rect 2464 384 2480 400
rect 2526 395 2537 408
rect 2319 350 2320 366
rect 2335 350 2348 372
rect 2363 350 2393 372
rect 2436 368 2498 384
rect 2526 377 2537 393
rect 2542 388 2552 408
rect 2562 388 2576 408
rect 2579 395 2588 408
rect 2604 395 2613 408
rect 2542 377 2576 388
rect 2579 377 2588 393
rect 2604 377 2613 393
rect 2620 388 2630 408
rect 2640 388 2654 408
rect 2655 395 2666 408
rect 2620 377 2654 388
rect 2655 377 2666 393
rect 2712 384 2728 400
rect 2735 398 2765 450
rect 2799 446 2800 453
rect 2784 438 2800 446
rect 2771 406 2784 425
rect 2799 406 2829 422
rect 2771 390 2845 406
rect 2771 388 2784 390
rect 2799 388 2833 390
rect 2436 366 2449 368
rect 2464 366 2498 368
rect 2436 350 2498 366
rect 2542 361 2558 364
rect 2620 361 2650 372
rect 2698 368 2744 384
rect 2771 372 2845 388
rect 2698 366 2732 368
rect 2697 350 2744 366
rect 2771 350 2784 372
rect 2799 350 2829 372
rect 2856 350 2857 366
rect 2872 350 2885 510
rect 2915 406 2928 510
rect 2973 488 2974 498
rect 2989 488 3002 498
rect 2973 484 3002 488
rect 3007 484 3037 510
rect 3055 496 3071 498
rect 3143 496 3196 510
rect 3144 494 3208 496
rect 3251 494 3266 510
rect 3315 507 3345 510
rect 3315 504 3351 507
rect 3281 496 3297 498
rect 3055 484 3070 488
rect 2973 482 3070 484
rect 3098 482 3266 494
rect 3282 484 3297 488
rect 3315 485 3354 504
rect 3373 498 3380 499
rect 3379 491 3380 498
rect 3363 488 3364 491
rect 3379 488 3392 491
rect 3315 484 3345 485
rect 3354 484 3360 485
rect 3363 484 3392 488
rect 3282 483 3392 484
rect 3282 482 3398 483
rect 2957 474 3008 482
rect 2957 462 2982 474
rect 2989 462 3008 474
rect 3039 474 3089 482
rect 3039 466 3055 474
rect 3062 472 3089 474
rect 3098 472 3319 482
rect 3062 462 3319 472
rect 3348 474 3398 482
rect 3348 465 3364 474
rect 2957 454 3008 462
rect 3055 454 3319 462
rect 3345 462 3364 465
rect 3371 462 3398 474
rect 3345 454 3398 462
rect 2973 446 2974 454
rect 2989 446 3002 454
rect 2973 438 2989 446
rect 2970 431 2989 434
rect 2970 422 2992 431
rect 2943 412 2992 422
rect 2943 406 2973 412
rect 2992 407 2997 412
rect 2915 390 2989 406
rect 3007 398 3037 454
rect 3072 444 3280 454
rect 3315 450 3360 454
rect 3363 453 3364 454
rect 3379 453 3392 454
rect 3098 414 3287 444
rect 3113 411 3287 414
rect 3106 408 3287 411
rect 2915 388 2928 390
rect 2943 388 2977 390
rect 2915 372 2989 388
rect 3016 384 3029 398
rect 3044 384 3060 400
rect 3106 395 3117 408
rect 2899 350 2900 366
rect 2915 350 2928 372
rect 2943 350 2973 372
rect 3016 368 3078 384
rect 3106 377 3117 393
rect 3122 388 3132 408
rect 3142 388 3156 408
rect 3159 395 3168 408
rect 3184 395 3193 408
rect 3122 377 3156 388
rect 3159 377 3168 393
rect 3184 377 3193 393
rect 3200 388 3210 408
rect 3220 388 3234 408
rect 3235 395 3246 408
rect 3200 377 3234 388
rect 3235 377 3246 393
rect 3292 384 3308 400
rect 3315 398 3345 450
rect 3379 446 3380 453
rect 3364 438 3380 446
rect 3351 406 3364 425
rect 3379 406 3409 422
rect 3351 390 3425 406
rect 3351 388 3364 390
rect 3379 388 3413 390
rect 3016 366 3029 368
rect 3044 366 3078 368
rect 3016 350 3078 366
rect 3122 361 3138 364
rect 3200 361 3230 372
rect 3278 368 3324 384
rect 3351 372 3425 388
rect 3278 366 3312 368
rect 3277 350 3324 366
rect 3351 350 3364 372
rect 3379 350 3409 372
rect 3436 350 3437 366
rect 3452 350 3465 510
rect 3495 406 3508 510
rect 3553 488 3554 498
rect 3569 488 3582 498
rect 3553 484 3582 488
rect 3587 484 3617 510
rect 3635 496 3651 498
rect 3723 496 3776 510
rect 3724 494 3788 496
rect 3831 494 3846 510
rect 3895 507 3925 510
rect 3895 504 3931 507
rect 3861 496 3877 498
rect 3635 484 3650 488
rect 3553 482 3650 484
rect 3678 482 3846 494
rect 3862 484 3877 488
rect 3895 485 3934 504
rect 3953 498 3960 499
rect 3959 491 3960 498
rect 3943 488 3944 491
rect 3959 488 3972 491
rect 3895 484 3925 485
rect 3934 484 3940 485
rect 3943 484 3972 488
rect 3862 483 3972 484
rect 3862 482 3978 483
rect 3537 474 3588 482
rect 3537 462 3562 474
rect 3569 462 3588 474
rect 3619 474 3669 482
rect 3619 466 3635 474
rect 3642 472 3669 474
rect 3678 472 3899 482
rect 3642 462 3899 472
rect 3928 474 3978 482
rect 3928 465 3944 474
rect 3537 454 3588 462
rect 3635 454 3899 462
rect 3925 462 3944 465
rect 3951 462 3978 474
rect 3925 454 3978 462
rect 3553 446 3554 454
rect 3569 446 3582 454
rect 3553 438 3569 446
rect 3550 431 3569 434
rect 3550 422 3572 431
rect 3523 412 3572 422
rect 3523 406 3553 412
rect 3572 407 3577 412
rect 3495 390 3569 406
rect 3587 398 3617 454
rect 3652 444 3860 454
rect 3895 450 3940 454
rect 3943 453 3944 454
rect 3959 453 3972 454
rect 3678 414 3867 444
rect 3693 411 3867 414
rect 3686 408 3867 411
rect 3495 388 3508 390
rect 3523 388 3557 390
rect 3495 372 3569 388
rect 3596 384 3609 398
rect 3624 384 3640 400
rect 3686 395 3697 408
rect 3479 350 3480 366
rect 3495 350 3508 372
rect 3523 350 3553 372
rect 3596 368 3658 384
rect 3686 377 3697 393
rect 3702 388 3712 408
rect 3722 388 3736 408
rect 3739 395 3748 408
rect 3764 395 3773 408
rect 3702 377 3736 388
rect 3739 377 3748 393
rect 3764 377 3773 393
rect 3780 388 3790 408
rect 3800 388 3814 408
rect 3815 395 3826 408
rect 3780 377 3814 388
rect 3815 377 3826 393
rect 3872 384 3888 400
rect 3895 398 3925 450
rect 3959 446 3960 453
rect 3944 438 3960 446
rect 3931 406 3944 425
rect 3959 406 3989 422
rect 3931 390 4005 406
rect 3931 388 3944 390
rect 3959 388 3993 390
rect 3596 366 3609 368
rect 3624 366 3658 368
rect 3596 350 3658 366
rect 3702 361 3718 364
rect 3780 361 3810 372
rect 3858 368 3904 384
rect 3931 372 4005 388
rect 3858 366 3892 368
rect 3857 350 3904 366
rect 3931 350 3944 372
rect 3959 350 3989 372
rect 4016 350 4017 366
rect 4032 350 4045 510
rect 4075 406 4088 510
rect 4133 488 4134 498
rect 4149 488 4162 498
rect 4133 484 4162 488
rect 4167 484 4197 510
rect 4215 496 4231 498
rect 4303 496 4356 510
rect 4304 494 4368 496
rect 4411 494 4426 510
rect 4475 507 4505 510
rect 4475 504 4511 507
rect 4441 496 4457 498
rect 4215 484 4230 488
rect 4133 482 4230 484
rect 4258 482 4426 494
rect 4442 484 4457 488
rect 4475 485 4514 504
rect 4533 498 4540 499
rect 4539 491 4540 498
rect 4523 488 4524 491
rect 4539 488 4552 491
rect 4475 484 4505 485
rect 4514 484 4520 485
rect 4523 484 4552 488
rect 4442 483 4552 484
rect 4442 482 4558 483
rect 4117 474 4168 482
rect 4117 462 4142 474
rect 4149 462 4168 474
rect 4199 474 4249 482
rect 4199 466 4215 474
rect 4222 472 4249 474
rect 4258 472 4479 482
rect 4222 462 4479 472
rect 4508 474 4558 482
rect 4508 465 4524 474
rect 4117 454 4168 462
rect 4215 454 4479 462
rect 4505 462 4524 465
rect 4531 462 4558 474
rect 4505 454 4558 462
rect 4133 446 4134 454
rect 4149 446 4162 454
rect 4133 438 4149 446
rect 4130 431 4149 434
rect 4130 422 4152 431
rect 4103 412 4152 422
rect 4103 406 4133 412
rect 4152 407 4157 412
rect 4075 390 4149 406
rect 4167 398 4197 454
rect 4232 444 4440 454
rect 4475 450 4520 454
rect 4523 453 4524 454
rect 4539 453 4552 454
rect 4258 414 4447 444
rect 4273 411 4447 414
rect 4266 408 4447 411
rect 4075 388 4088 390
rect 4103 388 4137 390
rect 4075 372 4149 388
rect 4176 384 4189 398
rect 4204 384 4220 400
rect 4266 395 4277 408
rect 4059 350 4060 366
rect 4075 350 4088 372
rect 4103 350 4133 372
rect 4176 368 4238 384
rect 4266 377 4277 393
rect 4282 388 4292 408
rect 4302 388 4316 408
rect 4319 395 4328 408
rect 4344 395 4353 408
rect 4282 377 4316 388
rect 4319 377 4328 393
rect 4344 377 4353 393
rect 4360 388 4370 408
rect 4380 388 4394 408
rect 4395 395 4406 408
rect 4360 377 4394 388
rect 4395 377 4406 393
rect 4452 384 4468 400
rect 4475 398 4505 450
rect 4539 446 4540 453
rect 4524 438 4540 446
rect 4511 406 4524 425
rect 4539 406 4569 422
rect 4511 390 4585 406
rect 4511 388 4524 390
rect 4539 388 4573 390
rect 4176 366 4189 368
rect 4204 366 4238 368
rect 4176 350 4238 366
rect 4282 361 4298 364
rect 4360 361 4390 372
rect 4438 368 4484 384
rect 4511 372 4585 388
rect 4438 366 4472 368
rect 4437 350 4484 366
rect 4511 350 4524 372
rect 4539 350 4569 372
rect 4596 350 4597 366
rect 4612 350 4625 510
rect -7 342 34 350
rect -7 316 8 342
rect 15 316 34 342
rect 98 338 160 350
rect 172 338 247 350
rect 305 338 380 350
rect 392 338 423 350
rect 429 338 464 350
rect 98 336 260 338
rect -7 308 34 316
rect 116 312 129 336
rect 144 334 159 336
rect -1 298 0 308
rect 15 298 28 308
rect 43 298 73 312
rect 116 298 159 312
rect 183 309 190 316
rect 193 312 260 336
rect 292 336 464 338
rect 262 314 290 318
rect 292 314 372 336
rect 393 334 408 336
rect 262 312 372 314
rect 193 308 372 312
rect 166 298 196 308
rect 198 298 351 308
rect 359 298 389 308
rect 393 298 423 312
rect 451 298 464 336
rect 536 342 571 350
rect 536 316 537 342
rect 544 316 571 342
rect 479 298 509 312
rect 536 308 571 316
rect 573 342 614 350
rect 573 316 588 342
rect 595 316 614 342
rect 678 338 740 350
rect 752 338 827 350
rect 885 338 960 350
rect 972 338 1003 350
rect 1009 338 1044 350
rect 678 336 840 338
rect 573 308 614 316
rect 696 312 709 336
rect 724 334 739 336
rect 536 298 537 308
rect 552 298 565 308
rect 579 298 580 308
rect 595 298 608 308
rect 623 298 653 312
rect 696 298 739 312
rect 763 309 770 316
rect 773 312 840 336
rect 872 336 1044 338
rect 842 314 870 318
rect 872 314 952 336
rect 973 334 988 336
rect 842 312 952 314
rect 773 308 952 312
rect 746 298 776 308
rect 778 298 931 308
rect 939 298 969 308
rect 973 298 1003 312
rect 1031 298 1044 336
rect 1116 342 1151 350
rect 1116 316 1117 342
rect 1124 316 1151 342
rect 1059 298 1089 312
rect 1116 308 1151 316
rect 1153 342 1194 350
rect 1153 316 1168 342
rect 1175 316 1194 342
rect 1258 338 1320 350
rect 1332 338 1407 350
rect 1465 338 1540 350
rect 1552 338 1583 350
rect 1589 338 1624 350
rect 1258 336 1420 338
rect 1153 308 1194 316
rect 1276 312 1289 336
rect 1304 334 1319 336
rect 1116 298 1117 308
rect 1132 298 1145 308
rect 1159 298 1160 308
rect 1175 298 1188 308
rect 1203 298 1233 312
rect 1276 298 1319 312
rect 1343 309 1350 316
rect 1353 312 1420 336
rect 1452 336 1624 338
rect 1422 314 1450 318
rect 1452 314 1532 336
rect 1553 334 1568 336
rect 1422 312 1532 314
rect 1353 308 1532 312
rect 1326 298 1356 308
rect 1358 298 1511 308
rect 1519 298 1549 308
rect 1553 298 1583 312
rect 1611 298 1624 336
rect 1696 342 1731 350
rect 1696 316 1697 342
rect 1704 316 1731 342
rect 1639 298 1669 312
rect 1696 308 1731 316
rect 1733 342 1774 350
rect 1733 316 1748 342
rect 1755 316 1774 342
rect 1838 338 1900 350
rect 1912 338 1987 350
rect 2045 338 2120 350
rect 2132 338 2163 350
rect 2169 338 2204 350
rect 1838 336 2000 338
rect 1733 308 1774 316
rect 1856 312 1869 336
rect 1884 334 1899 336
rect 1696 298 1697 308
rect 1712 298 1725 308
rect 1739 298 1740 308
rect 1755 298 1768 308
rect 1783 298 1813 312
rect 1856 298 1899 312
rect 1923 309 1930 316
rect 1933 312 2000 336
rect 2032 336 2204 338
rect 2002 314 2030 318
rect 2032 314 2112 336
rect 2133 334 2148 336
rect 2002 312 2112 314
rect 1933 308 2112 312
rect 1906 298 1936 308
rect 1938 298 2091 308
rect 2099 298 2129 308
rect 2133 298 2163 312
rect 2191 298 2204 336
rect 2276 342 2311 350
rect 2276 316 2277 342
rect 2284 316 2311 342
rect 2219 298 2249 312
rect 2276 308 2311 316
rect 2313 342 2354 350
rect 2313 316 2328 342
rect 2335 316 2354 342
rect 2418 338 2480 350
rect 2492 338 2567 350
rect 2625 338 2700 350
rect 2712 338 2743 350
rect 2749 338 2784 350
rect 2418 336 2580 338
rect 2313 308 2354 316
rect 2436 312 2449 336
rect 2464 334 2479 336
rect 2276 298 2277 308
rect 2292 298 2305 308
rect 2319 298 2320 308
rect 2335 298 2348 308
rect 2363 298 2393 312
rect 2436 298 2479 312
rect 2503 309 2510 316
rect 2513 312 2580 336
rect 2612 336 2784 338
rect 2582 314 2610 318
rect 2612 314 2692 336
rect 2713 334 2728 336
rect 2582 312 2692 314
rect 2513 308 2692 312
rect 2486 298 2516 308
rect 2518 298 2671 308
rect 2679 298 2709 308
rect 2713 298 2743 312
rect 2771 298 2784 336
rect 2856 342 2891 350
rect 2856 316 2857 342
rect 2864 316 2891 342
rect 2799 298 2829 312
rect 2856 308 2891 316
rect 2893 342 2934 350
rect 2893 316 2908 342
rect 2915 316 2934 342
rect 2998 338 3060 350
rect 3072 338 3147 350
rect 3205 338 3280 350
rect 3292 338 3323 350
rect 3329 338 3364 350
rect 2998 336 3160 338
rect 2893 308 2934 316
rect 3016 312 3029 336
rect 3044 334 3059 336
rect 2856 298 2857 308
rect 2872 298 2885 308
rect 2899 298 2900 308
rect 2915 298 2928 308
rect 2943 298 2973 312
rect 3016 298 3059 312
rect 3083 309 3090 316
rect 3093 312 3160 336
rect 3192 336 3364 338
rect 3162 314 3190 318
rect 3192 314 3272 336
rect 3293 334 3308 336
rect 3162 312 3272 314
rect 3093 308 3272 312
rect 3066 298 3096 308
rect 3098 298 3251 308
rect 3259 298 3289 308
rect 3293 298 3323 312
rect 3351 298 3364 336
rect 3436 342 3471 350
rect 3436 316 3437 342
rect 3444 316 3471 342
rect 3379 298 3409 312
rect 3436 308 3471 316
rect 3473 342 3514 350
rect 3473 316 3488 342
rect 3495 316 3514 342
rect 3578 338 3640 350
rect 3652 338 3727 350
rect 3785 338 3860 350
rect 3872 338 3903 350
rect 3909 338 3944 350
rect 3578 336 3740 338
rect 3473 308 3514 316
rect 3596 312 3609 336
rect 3624 334 3639 336
rect 3436 298 3437 308
rect 3452 298 3465 308
rect 3479 298 3480 308
rect 3495 298 3508 308
rect 3523 298 3553 312
rect 3596 298 3639 312
rect 3663 309 3670 316
rect 3673 312 3740 336
rect 3772 336 3944 338
rect 3742 314 3770 318
rect 3772 314 3852 336
rect 3873 334 3888 336
rect 3742 312 3852 314
rect 3673 308 3852 312
rect 3646 298 3676 308
rect 3678 298 3831 308
rect 3839 298 3869 308
rect 3873 298 3903 312
rect 3931 298 3944 336
rect 4016 342 4051 350
rect 4016 316 4017 342
rect 4024 316 4051 342
rect 3959 298 3989 312
rect 4016 308 4051 316
rect 4053 342 4094 350
rect 4053 316 4068 342
rect 4075 316 4094 342
rect 4158 338 4220 350
rect 4232 338 4307 350
rect 4365 338 4440 350
rect 4452 338 4483 350
rect 4489 338 4524 350
rect 4158 336 4320 338
rect 4053 308 4094 316
rect 4176 312 4189 336
rect 4204 334 4219 336
rect 4016 298 4017 308
rect 4032 298 4045 308
rect 4059 298 4060 308
rect 4075 298 4088 308
rect 4103 298 4133 312
rect 4176 298 4219 312
rect 4243 309 4250 316
rect 4253 312 4320 336
rect 4352 336 4524 338
rect 4322 314 4350 318
rect 4352 314 4432 336
rect 4453 334 4468 336
rect 4322 312 4432 314
rect 4253 308 4432 312
rect 4226 298 4256 308
rect 4258 298 4411 308
rect 4419 298 4449 308
rect 4453 298 4483 312
rect 4511 298 4524 336
rect 4596 342 4631 350
rect 4596 316 4597 342
rect 4604 316 4631 342
rect 4539 298 4569 312
rect 4596 308 4631 316
rect 4596 298 4597 308
rect 4612 298 4625 308
rect -1 292 4625 298
rect 0 284 4625 292
rect 15 254 28 284
rect 43 266 73 284
rect 116 270 130 284
rect 166 270 386 284
rect 117 268 130 270
rect 83 256 98 268
rect 80 254 102 256
rect 107 254 137 268
rect 198 266 351 270
rect 180 254 372 266
rect 415 254 445 268
rect 451 254 464 284
rect 479 266 509 284
rect 552 254 565 284
rect 595 254 608 284
rect 623 266 653 284
rect 696 270 710 284
rect 746 270 966 284
rect 697 268 710 270
rect 663 256 678 268
rect 660 254 682 256
rect 687 254 717 268
rect 778 266 931 270
rect 760 254 952 266
rect 995 254 1025 268
rect 1031 254 1044 284
rect 1059 266 1089 284
rect 1132 254 1145 284
rect 1175 254 1188 284
rect 1203 266 1233 284
rect 1276 270 1290 284
rect 1326 270 1546 284
rect 1277 268 1290 270
rect 1243 256 1258 268
rect 1240 254 1262 256
rect 1267 254 1297 268
rect 1358 266 1511 270
rect 1340 254 1532 266
rect 1575 254 1605 268
rect 1611 254 1624 284
rect 1639 266 1669 284
rect 1712 254 1725 284
rect 1755 254 1768 284
rect 1783 266 1813 284
rect 1856 270 1870 284
rect 1906 270 2126 284
rect 1857 268 1870 270
rect 1823 256 1838 268
rect 1820 254 1842 256
rect 1847 254 1877 268
rect 1938 266 2091 270
rect 1920 254 2112 266
rect 2155 254 2185 268
rect 2191 254 2204 284
rect 2219 266 2249 284
rect 2292 254 2305 284
rect 2335 254 2348 284
rect 2363 266 2393 284
rect 2436 270 2450 284
rect 2486 270 2706 284
rect 2437 268 2450 270
rect 2403 256 2418 268
rect 2400 254 2422 256
rect 2427 254 2457 268
rect 2518 266 2671 270
rect 2500 254 2692 266
rect 2735 254 2765 268
rect 2771 254 2784 284
rect 2799 266 2829 284
rect 2872 254 2885 284
rect 2915 254 2928 284
rect 2943 266 2973 284
rect 3016 270 3030 284
rect 3066 270 3286 284
rect 3017 268 3030 270
rect 2983 256 2998 268
rect 2980 254 3002 256
rect 3007 254 3037 268
rect 3098 266 3251 270
rect 3080 254 3272 266
rect 3315 254 3345 268
rect 3351 254 3364 284
rect 3379 266 3409 284
rect 3452 254 3465 284
rect 3495 254 3508 284
rect 3523 266 3553 284
rect 3596 270 3610 284
rect 3646 270 3866 284
rect 3597 268 3610 270
rect 3563 256 3578 268
rect 3560 254 3582 256
rect 3587 254 3617 268
rect 3678 266 3831 270
rect 3660 254 3852 266
rect 3895 254 3925 268
rect 3931 254 3944 284
rect 3959 266 3989 284
rect 4032 254 4045 284
rect 4075 254 4088 284
rect 4103 266 4133 284
rect 4176 270 4190 284
rect 4226 270 4446 284
rect 4177 268 4190 270
rect 4143 256 4158 268
rect 4140 254 4162 256
rect 4167 254 4197 268
rect 4258 266 4411 270
rect 4240 254 4432 266
rect 4475 254 4505 268
rect 4511 254 4524 284
rect 4539 266 4569 284
rect 4612 254 4625 284
rect 0 240 4625 254
rect 15 136 28 240
rect 73 218 74 228
rect 89 218 102 228
rect 73 214 102 218
rect 107 214 137 240
rect 155 226 171 228
rect 243 226 296 240
rect 244 224 308 226
rect 155 214 170 218
rect 73 212 170 214
rect 57 204 108 212
rect 57 192 82 204
rect 89 192 108 204
rect 139 204 189 212
rect 139 196 155 204
rect 162 202 189 204
rect 198 204 213 208
rect 260 204 292 224
rect 351 212 366 240
rect 415 237 445 240
rect 415 234 451 237
rect 381 226 397 228
rect 382 214 397 218
rect 415 215 454 234
rect 473 228 480 229
rect 479 221 480 228
rect 463 218 464 221
rect 479 218 492 221
rect 415 214 445 215
rect 454 214 460 215
rect 463 214 492 218
rect 382 213 492 214
rect 382 212 498 213
rect 351 204 419 212
rect 198 202 267 204
rect 285 202 419 204
rect 162 198 234 202
rect 162 196 287 198
rect 162 192 234 196
rect 57 184 108 192
rect 155 188 234 192
rect 315 188 419 202
rect 448 204 498 212
rect 448 195 464 204
rect 155 184 419 188
rect 445 192 464 195
rect 471 192 498 204
rect 445 184 498 192
rect 73 176 74 184
rect 89 176 102 184
rect 73 168 89 176
rect 70 161 89 164
rect 70 152 92 161
rect 43 142 92 152
rect 43 136 73 142
rect 92 137 97 142
rect 15 120 89 136
rect 107 128 137 184
rect 172 174 380 184
rect 415 180 460 184
rect 463 183 464 184
rect 479 183 492 184
rect 339 170 387 174
rect 222 148 252 157
rect 315 150 330 157
rect 351 148 387 170
rect 198 144 387 148
rect 213 141 387 144
rect 206 138 387 141
rect 15 118 28 120
rect 43 118 77 120
rect 15 102 89 118
rect 116 114 129 128
rect 144 114 160 130
rect 206 125 217 138
rect -1 80 0 96
rect 15 80 28 102
rect 43 80 73 102
rect 116 98 178 114
rect 206 107 217 123
rect 222 118 232 138
rect 242 118 256 138
rect 259 125 268 138
rect 284 125 293 138
rect 222 107 256 118
rect 259 107 267 123
rect 284 107 293 123
rect 300 118 310 138
rect 320 118 334 138
rect 335 125 346 138
rect 300 107 334 118
rect 335 107 346 123
rect 392 114 408 130
rect 415 128 445 180
rect 479 176 480 183
rect 464 168 480 176
rect 451 136 464 155
rect 479 136 509 152
rect 451 120 525 136
rect 451 118 464 120
rect 479 118 513 120
rect 116 96 129 98
rect 144 96 178 98
rect 116 80 178 96
rect 222 91 235 94
rect 300 91 330 102
rect 378 98 424 114
rect 451 102 525 118
rect 378 96 412 98
rect 377 80 424 96
rect 451 80 464 102
rect 479 80 509 102
rect 536 80 537 96
rect 552 80 565 240
rect 595 136 608 240
rect 653 218 654 228
rect 669 218 682 228
rect 653 214 682 218
rect 687 214 717 240
rect 735 226 751 228
rect 823 226 876 240
rect 824 224 888 226
rect 735 214 750 218
rect 653 212 750 214
rect 637 204 688 212
rect 637 192 662 204
rect 669 192 688 204
rect 719 204 769 212
rect 719 196 735 204
rect 742 202 769 204
rect 778 204 793 208
rect 840 204 872 224
rect 931 212 946 240
rect 995 237 1025 240
rect 995 234 1031 237
rect 961 226 977 228
rect 962 214 977 218
rect 995 215 1034 234
rect 1053 228 1060 229
rect 1059 221 1060 228
rect 1043 218 1044 221
rect 1059 218 1072 221
rect 995 214 1025 215
rect 1034 214 1040 215
rect 1043 214 1072 218
rect 962 213 1072 214
rect 962 212 1078 213
rect 931 204 999 212
rect 778 202 847 204
rect 865 202 999 204
rect 742 198 814 202
rect 742 196 867 198
rect 742 192 814 196
rect 637 184 688 192
rect 735 188 814 192
rect 895 188 999 202
rect 1028 204 1078 212
rect 1028 195 1044 204
rect 735 184 999 188
rect 1025 192 1044 195
rect 1051 192 1078 204
rect 1025 184 1078 192
rect 653 176 654 184
rect 669 176 682 184
rect 653 168 669 176
rect 650 161 669 164
rect 650 152 672 161
rect 623 142 672 152
rect 623 136 653 142
rect 672 137 677 142
rect 595 120 669 136
rect 687 128 717 184
rect 752 174 960 184
rect 995 180 1040 184
rect 1043 183 1044 184
rect 1059 183 1072 184
rect 919 170 967 174
rect 802 148 832 157
rect 895 150 910 157
rect 931 148 967 170
rect 778 144 967 148
rect 793 141 967 144
rect 786 138 967 141
rect 595 118 608 120
rect 623 118 657 120
rect 595 102 669 118
rect 696 114 709 128
rect 724 114 740 130
rect 786 125 797 138
rect 579 80 580 96
rect 595 80 608 102
rect 623 80 653 102
rect 696 98 758 114
rect 786 107 797 123
rect 802 118 812 138
rect 822 118 836 138
rect 839 125 848 138
rect 864 125 873 138
rect 802 107 836 118
rect 839 107 847 123
rect 864 107 873 123
rect 880 118 890 138
rect 900 118 914 138
rect 915 125 926 138
rect 880 107 914 118
rect 915 107 926 123
rect 972 114 988 130
rect 995 128 1025 180
rect 1059 176 1060 183
rect 1044 168 1060 176
rect 1031 136 1044 155
rect 1059 136 1089 152
rect 1031 120 1105 136
rect 1031 118 1044 120
rect 1059 118 1093 120
rect 696 96 709 98
rect 724 96 758 98
rect 696 80 758 96
rect 802 91 815 94
rect 880 91 910 102
rect 958 98 1004 114
rect 1031 102 1105 118
rect 958 96 992 98
rect 957 80 1004 96
rect 1031 80 1044 102
rect 1059 80 1089 102
rect 1116 80 1117 96
rect 1132 80 1145 240
rect 1175 136 1188 240
rect 1233 218 1234 228
rect 1249 218 1262 228
rect 1233 214 1262 218
rect 1267 214 1297 240
rect 1315 226 1331 228
rect 1403 226 1456 240
rect 1404 224 1468 226
rect 1315 214 1330 218
rect 1233 212 1330 214
rect 1217 204 1268 212
rect 1217 192 1242 204
rect 1249 192 1268 204
rect 1299 204 1349 212
rect 1299 196 1315 204
rect 1322 202 1349 204
rect 1358 204 1373 208
rect 1420 204 1452 224
rect 1511 212 1526 240
rect 1575 237 1605 240
rect 1575 234 1611 237
rect 1541 226 1557 228
rect 1542 214 1557 218
rect 1575 215 1614 234
rect 1633 228 1640 229
rect 1639 221 1640 228
rect 1623 218 1624 221
rect 1639 218 1652 221
rect 1575 214 1605 215
rect 1614 214 1620 215
rect 1623 214 1652 218
rect 1542 213 1652 214
rect 1542 212 1658 213
rect 1511 204 1579 212
rect 1358 202 1427 204
rect 1445 202 1579 204
rect 1322 198 1394 202
rect 1322 196 1447 198
rect 1322 192 1394 196
rect 1217 184 1268 192
rect 1315 188 1394 192
rect 1475 188 1579 202
rect 1608 204 1658 212
rect 1608 195 1624 204
rect 1315 184 1579 188
rect 1605 192 1624 195
rect 1631 192 1658 204
rect 1605 184 1658 192
rect 1233 176 1234 184
rect 1249 176 1262 184
rect 1233 168 1249 176
rect 1230 161 1249 164
rect 1230 152 1252 161
rect 1203 142 1252 152
rect 1203 136 1233 142
rect 1252 137 1257 142
rect 1175 120 1249 136
rect 1267 128 1297 184
rect 1332 174 1540 184
rect 1575 180 1620 184
rect 1623 183 1624 184
rect 1639 183 1652 184
rect 1499 170 1547 174
rect 1382 148 1412 157
rect 1475 150 1490 157
rect 1511 148 1547 170
rect 1358 144 1547 148
rect 1373 141 1547 144
rect 1366 138 1547 141
rect 1175 118 1188 120
rect 1203 118 1237 120
rect 1175 102 1249 118
rect 1276 114 1289 128
rect 1304 114 1320 130
rect 1366 125 1377 138
rect 1159 80 1160 96
rect 1175 80 1188 102
rect 1203 80 1233 102
rect 1276 98 1338 114
rect 1366 107 1377 123
rect 1382 118 1392 138
rect 1402 118 1416 138
rect 1419 125 1428 138
rect 1444 125 1453 138
rect 1382 107 1416 118
rect 1419 107 1427 123
rect 1444 107 1453 123
rect 1460 118 1470 138
rect 1480 118 1494 138
rect 1495 125 1506 138
rect 1460 107 1494 118
rect 1495 107 1506 123
rect 1552 114 1568 130
rect 1575 128 1605 180
rect 1639 176 1640 183
rect 1624 168 1640 176
rect 1611 136 1624 155
rect 1639 136 1669 152
rect 1611 120 1685 136
rect 1611 118 1624 120
rect 1639 118 1673 120
rect 1276 96 1289 98
rect 1304 96 1338 98
rect 1276 80 1338 96
rect 1382 91 1395 94
rect 1460 91 1490 102
rect 1538 98 1584 114
rect 1611 102 1685 118
rect 1538 96 1572 98
rect 1537 80 1584 96
rect 1611 80 1624 102
rect 1639 80 1669 102
rect 1696 80 1697 96
rect 1712 80 1725 240
rect 1755 136 1768 240
rect 1813 218 1814 228
rect 1829 218 1842 228
rect 1813 214 1842 218
rect 1847 214 1877 240
rect 1895 226 1911 228
rect 1983 226 2036 240
rect 1984 224 2048 226
rect 1895 214 1910 218
rect 1813 212 1910 214
rect 1797 204 1848 212
rect 1797 192 1822 204
rect 1829 192 1848 204
rect 1879 204 1929 212
rect 1879 196 1895 204
rect 1902 202 1929 204
rect 1938 204 1953 208
rect 2000 204 2032 224
rect 2091 212 2106 240
rect 2155 237 2185 240
rect 2155 234 2191 237
rect 2121 226 2137 228
rect 2122 214 2137 218
rect 2155 215 2194 234
rect 2213 228 2220 229
rect 2219 221 2220 228
rect 2203 218 2204 221
rect 2219 218 2232 221
rect 2155 214 2185 215
rect 2194 214 2200 215
rect 2203 214 2232 218
rect 2122 213 2232 214
rect 2122 212 2238 213
rect 2091 204 2159 212
rect 1938 202 2007 204
rect 2025 202 2159 204
rect 1902 198 1974 202
rect 1902 196 2027 198
rect 1902 192 1974 196
rect 1797 184 1848 192
rect 1895 188 1974 192
rect 2055 188 2159 202
rect 2188 204 2238 212
rect 2188 195 2204 204
rect 1895 184 2159 188
rect 2185 192 2204 195
rect 2211 192 2238 204
rect 2185 184 2238 192
rect 1813 176 1814 184
rect 1829 176 1842 184
rect 1813 168 1829 176
rect 1810 161 1829 164
rect 1810 152 1832 161
rect 1783 142 1832 152
rect 1783 136 1813 142
rect 1832 137 1837 142
rect 1755 120 1829 136
rect 1847 128 1877 184
rect 1912 174 2120 184
rect 2155 180 2200 184
rect 2203 183 2204 184
rect 2219 183 2232 184
rect 2079 170 2127 174
rect 1962 148 1992 157
rect 2055 150 2070 157
rect 2091 148 2127 170
rect 1938 144 2127 148
rect 1953 141 2127 144
rect 1946 138 2127 141
rect 1755 118 1768 120
rect 1783 118 1817 120
rect 1755 102 1829 118
rect 1856 114 1869 128
rect 1884 114 1900 130
rect 1946 125 1957 138
rect 1739 80 1740 96
rect 1755 80 1768 102
rect 1783 80 1813 102
rect 1856 98 1918 114
rect 1946 107 1957 123
rect 1962 118 1972 138
rect 1982 118 1996 138
rect 1999 125 2008 138
rect 2024 125 2033 138
rect 1962 107 1996 118
rect 1999 107 2007 123
rect 2024 107 2033 123
rect 2040 118 2050 138
rect 2060 118 2074 138
rect 2075 125 2086 138
rect 2040 107 2074 118
rect 2075 107 2086 123
rect 2132 114 2148 130
rect 2155 128 2185 180
rect 2219 176 2220 183
rect 2204 168 2220 176
rect 2191 136 2204 155
rect 2219 136 2249 152
rect 2191 120 2265 136
rect 2191 118 2204 120
rect 2219 118 2253 120
rect 1856 96 1869 98
rect 1884 96 1918 98
rect 1856 80 1918 96
rect 1962 91 1975 94
rect 2040 91 2070 102
rect 2118 98 2164 114
rect 2191 102 2265 118
rect 2118 96 2152 98
rect 2117 80 2164 96
rect 2191 80 2204 102
rect 2219 80 2249 102
rect 2276 80 2277 96
rect 2292 80 2305 240
rect 2335 136 2348 240
rect 2393 218 2394 228
rect 2409 218 2422 228
rect 2393 214 2422 218
rect 2427 214 2457 240
rect 2475 226 2491 228
rect 2563 226 2616 240
rect 2564 224 2628 226
rect 2475 214 2490 218
rect 2393 212 2490 214
rect 2377 204 2428 212
rect 2377 192 2402 204
rect 2409 192 2428 204
rect 2459 204 2509 212
rect 2459 196 2475 204
rect 2482 202 2509 204
rect 2518 204 2533 208
rect 2580 204 2612 224
rect 2671 212 2686 240
rect 2735 237 2765 240
rect 2735 234 2771 237
rect 2701 226 2717 228
rect 2702 214 2717 218
rect 2735 215 2774 234
rect 2793 228 2800 229
rect 2799 221 2800 228
rect 2783 218 2784 221
rect 2799 218 2812 221
rect 2735 214 2765 215
rect 2774 214 2780 215
rect 2783 214 2812 218
rect 2702 213 2812 214
rect 2702 212 2818 213
rect 2671 204 2739 212
rect 2518 202 2587 204
rect 2605 202 2739 204
rect 2482 198 2554 202
rect 2482 196 2607 198
rect 2482 192 2554 196
rect 2377 184 2428 192
rect 2475 188 2554 192
rect 2635 188 2739 202
rect 2768 204 2818 212
rect 2768 195 2784 204
rect 2475 184 2739 188
rect 2765 192 2784 195
rect 2791 192 2818 204
rect 2765 184 2818 192
rect 2393 176 2394 184
rect 2409 176 2422 184
rect 2393 168 2409 176
rect 2390 161 2409 164
rect 2390 152 2412 161
rect 2363 142 2412 152
rect 2363 136 2393 142
rect 2412 137 2417 142
rect 2335 120 2409 136
rect 2427 128 2457 184
rect 2492 174 2700 184
rect 2735 180 2780 184
rect 2783 183 2784 184
rect 2799 183 2812 184
rect 2659 170 2707 174
rect 2542 148 2572 157
rect 2635 150 2650 157
rect 2671 148 2707 170
rect 2518 144 2707 148
rect 2533 141 2707 144
rect 2526 138 2707 141
rect 2335 118 2348 120
rect 2363 118 2397 120
rect 2335 102 2409 118
rect 2436 114 2449 128
rect 2464 114 2480 130
rect 2526 125 2537 138
rect 2319 80 2320 96
rect 2335 80 2348 102
rect 2363 80 2393 102
rect 2436 98 2498 114
rect 2526 107 2537 123
rect 2542 118 2552 138
rect 2562 118 2576 138
rect 2579 125 2588 138
rect 2604 125 2613 138
rect 2542 107 2576 118
rect 2579 107 2587 123
rect 2604 107 2613 123
rect 2620 118 2630 138
rect 2640 118 2654 138
rect 2655 125 2666 138
rect 2620 107 2654 118
rect 2655 107 2666 123
rect 2712 114 2728 130
rect 2735 128 2765 180
rect 2799 176 2800 183
rect 2784 168 2800 176
rect 2771 136 2784 155
rect 2799 136 2829 152
rect 2771 120 2845 136
rect 2771 118 2784 120
rect 2799 118 2833 120
rect 2436 96 2449 98
rect 2464 96 2498 98
rect 2436 80 2498 96
rect 2542 91 2555 94
rect 2620 91 2650 102
rect 2698 98 2744 114
rect 2771 102 2845 118
rect 2698 96 2732 98
rect 2697 80 2744 96
rect 2771 80 2784 102
rect 2799 80 2829 102
rect 2856 80 2857 96
rect 2872 80 2885 240
rect 2915 136 2928 240
rect 2973 218 2974 228
rect 2989 218 3002 228
rect 2973 214 3002 218
rect 3007 214 3037 240
rect 3055 226 3071 228
rect 3143 226 3196 240
rect 3144 224 3208 226
rect 3055 214 3070 218
rect 2973 212 3070 214
rect 2957 204 3008 212
rect 2957 192 2982 204
rect 2989 192 3008 204
rect 3039 204 3089 212
rect 3039 196 3055 204
rect 3062 202 3089 204
rect 3098 204 3113 208
rect 3160 204 3192 224
rect 3251 212 3266 240
rect 3315 237 3345 240
rect 3315 234 3351 237
rect 3281 226 3297 228
rect 3282 214 3297 218
rect 3315 215 3354 234
rect 3373 228 3380 229
rect 3379 221 3380 228
rect 3363 218 3364 221
rect 3379 218 3392 221
rect 3315 214 3345 215
rect 3354 214 3360 215
rect 3363 214 3392 218
rect 3282 213 3392 214
rect 3282 212 3398 213
rect 3251 204 3319 212
rect 3098 202 3167 204
rect 3185 202 3319 204
rect 3062 198 3134 202
rect 3062 196 3187 198
rect 3062 192 3134 196
rect 2957 184 3008 192
rect 3055 188 3134 192
rect 3215 188 3319 202
rect 3348 204 3398 212
rect 3348 195 3364 204
rect 3055 184 3319 188
rect 3345 192 3364 195
rect 3371 192 3398 204
rect 3345 184 3398 192
rect 2973 176 2974 184
rect 2989 176 3002 184
rect 2973 168 2989 176
rect 2970 161 2989 164
rect 2970 152 2992 161
rect 2943 142 2992 152
rect 2943 136 2973 142
rect 2992 137 2997 142
rect 2915 120 2989 136
rect 3007 128 3037 184
rect 3072 174 3280 184
rect 3315 180 3360 184
rect 3363 183 3364 184
rect 3379 183 3392 184
rect 3239 170 3287 174
rect 3122 148 3152 157
rect 3215 150 3230 157
rect 3251 148 3287 170
rect 3098 144 3287 148
rect 3113 141 3287 144
rect 3106 138 3287 141
rect 2915 118 2928 120
rect 2943 118 2977 120
rect 2915 102 2989 118
rect 3016 114 3029 128
rect 3044 114 3060 130
rect 3106 125 3117 138
rect 2899 80 2900 96
rect 2915 80 2928 102
rect 2943 80 2973 102
rect 3016 98 3078 114
rect 3106 107 3117 123
rect 3122 118 3132 138
rect 3142 118 3156 138
rect 3159 125 3168 138
rect 3184 125 3193 138
rect 3122 107 3156 118
rect 3159 107 3167 123
rect 3184 107 3193 123
rect 3200 118 3210 138
rect 3220 118 3234 138
rect 3235 125 3246 138
rect 3200 107 3234 118
rect 3235 107 3246 123
rect 3292 114 3308 130
rect 3315 128 3345 180
rect 3379 176 3380 183
rect 3364 168 3380 176
rect 3351 136 3364 155
rect 3379 136 3409 152
rect 3351 120 3425 136
rect 3351 118 3364 120
rect 3379 118 3413 120
rect 3016 96 3029 98
rect 3044 96 3078 98
rect 3016 80 3078 96
rect 3122 91 3135 94
rect 3200 91 3230 102
rect 3278 98 3324 114
rect 3351 102 3425 118
rect 3278 96 3312 98
rect 3277 80 3324 96
rect 3351 80 3364 102
rect 3379 80 3409 102
rect 3436 80 3437 96
rect 3452 80 3465 240
rect 3495 136 3508 240
rect 3553 218 3554 228
rect 3569 218 3582 228
rect 3553 214 3582 218
rect 3587 214 3617 240
rect 3635 226 3651 228
rect 3723 226 3776 240
rect 3724 224 3788 226
rect 3635 214 3650 218
rect 3553 212 3650 214
rect 3537 204 3588 212
rect 3537 192 3562 204
rect 3569 192 3588 204
rect 3619 204 3669 212
rect 3619 196 3635 204
rect 3642 202 3669 204
rect 3678 204 3693 208
rect 3740 204 3772 224
rect 3831 212 3846 240
rect 3895 237 3925 240
rect 3895 234 3931 237
rect 3861 226 3877 228
rect 3862 214 3877 218
rect 3895 215 3934 234
rect 3953 228 3960 229
rect 3959 221 3960 228
rect 3943 218 3944 221
rect 3959 218 3972 221
rect 3895 214 3925 215
rect 3934 214 3940 215
rect 3943 214 3972 218
rect 3862 213 3972 214
rect 3862 212 3978 213
rect 3831 204 3899 212
rect 3678 202 3747 204
rect 3765 202 3899 204
rect 3642 198 3714 202
rect 3642 196 3767 198
rect 3642 192 3714 196
rect 3537 184 3588 192
rect 3635 188 3714 192
rect 3795 188 3899 202
rect 3928 204 3978 212
rect 3928 195 3944 204
rect 3635 184 3899 188
rect 3925 192 3944 195
rect 3951 192 3978 204
rect 3925 184 3978 192
rect 3553 176 3554 184
rect 3569 176 3582 184
rect 3553 168 3569 176
rect 3550 161 3569 164
rect 3550 152 3572 161
rect 3523 142 3572 152
rect 3523 136 3553 142
rect 3572 137 3577 142
rect 3495 120 3569 136
rect 3587 128 3617 184
rect 3652 174 3860 184
rect 3895 180 3940 184
rect 3943 183 3944 184
rect 3959 183 3972 184
rect 3819 170 3867 174
rect 3702 148 3732 157
rect 3795 150 3810 157
rect 3831 148 3867 170
rect 3678 144 3867 148
rect 3693 141 3867 144
rect 3686 138 3867 141
rect 3495 118 3508 120
rect 3523 118 3557 120
rect 3495 102 3569 118
rect 3596 114 3609 128
rect 3624 114 3640 130
rect 3686 125 3697 138
rect 3479 80 3480 96
rect 3495 80 3508 102
rect 3523 80 3553 102
rect 3596 98 3658 114
rect 3686 107 3697 123
rect 3702 118 3712 138
rect 3722 118 3736 138
rect 3739 125 3748 138
rect 3764 125 3773 138
rect 3702 107 3736 118
rect 3739 107 3747 123
rect 3764 107 3773 123
rect 3780 118 3790 138
rect 3800 118 3814 138
rect 3815 125 3826 138
rect 3780 107 3814 118
rect 3815 107 3826 123
rect 3872 114 3888 130
rect 3895 128 3925 180
rect 3959 176 3960 183
rect 3944 168 3960 176
rect 3931 136 3944 155
rect 3959 136 3989 152
rect 3931 120 4005 136
rect 3931 118 3944 120
rect 3959 118 3993 120
rect 3596 96 3609 98
rect 3624 96 3658 98
rect 3596 80 3658 96
rect 3702 91 3715 94
rect 3780 91 3810 102
rect 3858 98 3904 114
rect 3931 102 4005 118
rect 3858 96 3892 98
rect 3857 80 3904 96
rect 3931 80 3944 102
rect 3959 80 3989 102
rect 4016 80 4017 96
rect 4032 80 4045 240
rect 4075 136 4088 240
rect 4133 218 4134 228
rect 4149 218 4162 228
rect 4133 214 4162 218
rect 4167 214 4197 240
rect 4215 226 4231 228
rect 4303 226 4356 240
rect 4304 224 4368 226
rect 4215 214 4230 218
rect 4133 212 4230 214
rect 4117 204 4168 212
rect 4117 192 4142 204
rect 4149 192 4168 204
rect 4199 204 4249 212
rect 4199 196 4215 204
rect 4222 202 4249 204
rect 4258 204 4273 208
rect 4320 204 4352 224
rect 4411 212 4426 240
rect 4475 237 4505 240
rect 4475 234 4511 237
rect 4441 226 4457 228
rect 4442 214 4457 218
rect 4475 215 4514 234
rect 4533 228 4540 229
rect 4539 221 4540 228
rect 4523 218 4524 221
rect 4539 218 4552 221
rect 4475 214 4505 215
rect 4514 214 4520 215
rect 4523 214 4552 218
rect 4442 213 4552 214
rect 4442 212 4558 213
rect 4411 204 4479 212
rect 4258 202 4327 204
rect 4345 202 4479 204
rect 4222 198 4294 202
rect 4222 196 4347 198
rect 4222 192 4294 196
rect 4117 184 4168 192
rect 4215 188 4294 192
rect 4375 188 4479 202
rect 4508 204 4558 212
rect 4508 195 4524 204
rect 4215 184 4479 188
rect 4505 192 4524 195
rect 4531 192 4558 204
rect 4505 184 4558 192
rect 4133 176 4134 184
rect 4149 176 4162 184
rect 4133 168 4149 176
rect 4130 161 4149 164
rect 4130 152 4152 161
rect 4103 142 4152 152
rect 4103 136 4133 142
rect 4152 137 4157 142
rect 4075 120 4149 136
rect 4167 128 4197 184
rect 4232 174 4440 184
rect 4475 180 4520 184
rect 4523 183 4524 184
rect 4539 183 4552 184
rect 4399 170 4447 174
rect 4282 148 4312 157
rect 4375 150 4390 157
rect 4411 148 4447 170
rect 4258 144 4447 148
rect 4273 141 4447 144
rect 4266 138 4447 141
rect 4075 118 4088 120
rect 4103 118 4137 120
rect 4075 102 4149 118
rect 4176 114 4189 128
rect 4204 114 4220 130
rect 4266 125 4277 138
rect 4059 80 4060 96
rect 4075 80 4088 102
rect 4103 80 4133 102
rect 4176 98 4238 114
rect 4266 107 4277 123
rect 4282 118 4292 138
rect 4302 118 4316 138
rect 4319 125 4328 138
rect 4344 125 4353 138
rect 4282 107 4316 118
rect 4319 107 4327 123
rect 4344 107 4353 123
rect 4360 118 4370 138
rect 4380 118 4394 138
rect 4395 125 4406 138
rect 4360 107 4394 118
rect 4395 107 4406 123
rect 4452 114 4468 130
rect 4475 128 4505 180
rect 4539 176 4540 183
rect 4524 168 4540 176
rect 4511 136 4524 155
rect 4539 136 4569 152
rect 4511 120 4585 136
rect 4511 118 4524 120
rect 4539 118 4573 120
rect 4176 96 4189 98
rect 4204 96 4238 98
rect 4176 80 4238 96
rect 4282 91 4295 94
rect 4360 91 4390 102
rect 4438 98 4484 114
rect 4511 102 4585 118
rect 4438 96 4472 98
rect 4437 80 4484 96
rect 4511 80 4524 102
rect 4539 80 4569 102
rect 4596 80 4597 96
rect 4612 80 4625 240
rect -7 72 34 80
rect -7 46 8 72
rect 15 46 34 72
rect 98 68 160 80
rect 172 68 247 80
rect 305 68 380 80
rect 392 68 423 80
rect 429 68 464 80
rect 98 66 260 68
rect -7 38 34 46
rect 116 38 129 66
rect 144 64 159 66
rect 183 39 190 46
rect 193 38 260 66
rect 292 66 464 68
rect 262 44 290 48
rect 292 44 372 66
rect 393 64 408 66
rect 262 42 372 44
rect 262 38 290 42
rect 292 38 372 42
rect -1 28 0 38
rect 15 28 28 38
rect 43 28 73 38
rect 116 28 159 38
rect 166 28 174 38
rect 193 30 196 38
rect 260 30 292 38
rect 193 28 359 30
rect 378 28 389 38
rect 393 28 423 38
rect 451 28 464 66
rect 536 72 571 80
rect 536 46 537 72
rect 544 46 571 72
rect 536 38 571 46
rect 573 72 614 80
rect 573 46 588 72
rect 595 46 614 72
rect 678 68 740 80
rect 752 68 827 80
rect 885 68 960 80
rect 972 68 1003 80
rect 1009 68 1044 80
rect 678 66 840 68
rect 573 38 614 46
rect 696 38 709 66
rect 724 64 739 66
rect 763 39 770 46
rect 773 38 840 66
rect 872 66 1044 68
rect 842 44 870 48
rect 872 44 952 66
rect 973 64 988 66
rect 842 42 952 44
rect 842 38 870 42
rect 872 38 952 42
rect 479 28 509 38
rect 536 28 537 38
rect 552 28 565 38
rect 579 28 580 38
rect 595 28 608 38
rect 623 28 653 38
rect 696 28 739 38
rect 746 28 754 38
rect 773 30 776 38
rect 840 30 872 38
rect 773 28 939 30
rect 958 28 969 38
rect 973 28 1003 38
rect 1031 28 1044 66
rect 1116 72 1151 80
rect 1116 46 1117 72
rect 1124 46 1151 72
rect 1116 38 1151 46
rect 1153 72 1194 80
rect 1153 46 1168 72
rect 1175 46 1194 72
rect 1258 68 1320 80
rect 1332 68 1407 80
rect 1465 68 1540 80
rect 1552 68 1583 80
rect 1589 68 1624 80
rect 1258 66 1420 68
rect 1153 38 1194 46
rect 1276 38 1289 66
rect 1304 64 1319 66
rect 1343 39 1350 46
rect 1353 38 1420 66
rect 1452 66 1624 68
rect 1422 44 1450 48
rect 1452 44 1532 66
rect 1553 64 1568 66
rect 1422 42 1532 44
rect 1422 38 1450 42
rect 1452 38 1532 42
rect 1059 28 1089 38
rect 1116 28 1117 38
rect 1132 28 1145 38
rect 1159 28 1160 38
rect 1175 28 1188 38
rect 1203 28 1233 38
rect 1276 28 1319 38
rect 1326 28 1334 38
rect 1353 30 1356 38
rect 1420 30 1452 38
rect 1353 28 1519 30
rect 1538 28 1549 38
rect 1553 28 1583 38
rect 1611 28 1624 66
rect 1696 72 1731 80
rect 1696 46 1697 72
rect 1704 46 1731 72
rect 1696 38 1731 46
rect 1733 72 1774 80
rect 1733 46 1748 72
rect 1755 46 1774 72
rect 1838 68 1900 80
rect 1912 68 1987 80
rect 2045 68 2120 80
rect 2132 68 2163 80
rect 2169 68 2204 80
rect 1838 66 2000 68
rect 1733 38 1774 46
rect 1856 38 1869 66
rect 1884 64 1899 66
rect 1923 39 1930 46
rect 1933 38 2000 66
rect 2032 66 2204 68
rect 2002 44 2030 48
rect 2032 44 2112 66
rect 2133 64 2148 66
rect 2002 42 2112 44
rect 2002 38 2030 42
rect 2032 38 2112 42
rect 1639 28 1669 38
rect 1696 28 1697 38
rect 1712 28 1725 38
rect 1739 28 1740 38
rect 1755 28 1768 38
rect 1783 28 1813 38
rect 1856 28 1899 38
rect 1906 28 1914 38
rect 1933 30 1936 38
rect 2000 30 2032 38
rect 1933 28 2099 30
rect 2118 28 2129 38
rect 2133 28 2163 38
rect 2191 28 2204 66
rect 2276 72 2311 80
rect 2276 46 2277 72
rect 2284 46 2311 72
rect 2276 38 2311 46
rect 2313 72 2354 80
rect 2313 46 2328 72
rect 2335 46 2354 72
rect 2418 68 2480 80
rect 2492 68 2567 80
rect 2625 68 2700 80
rect 2712 68 2743 80
rect 2749 68 2784 80
rect 2418 66 2580 68
rect 2313 38 2354 46
rect 2436 38 2449 66
rect 2464 64 2479 66
rect 2503 39 2510 46
rect 2513 38 2580 66
rect 2612 66 2784 68
rect 2582 44 2610 48
rect 2612 44 2692 66
rect 2713 64 2728 66
rect 2582 42 2692 44
rect 2582 38 2610 42
rect 2612 38 2692 42
rect 2219 28 2249 38
rect 2276 28 2277 38
rect 2292 28 2305 38
rect 2319 28 2320 38
rect 2335 28 2348 38
rect 2363 28 2393 38
rect 2436 28 2479 38
rect 2486 28 2494 38
rect 2513 30 2516 38
rect 2580 30 2612 38
rect 2513 28 2679 30
rect 2698 28 2709 38
rect 2713 28 2743 38
rect 2771 28 2784 66
rect 2856 72 2891 80
rect 2856 46 2857 72
rect 2864 46 2891 72
rect 2856 38 2891 46
rect 2893 72 2934 80
rect 2893 46 2908 72
rect 2915 46 2934 72
rect 2998 68 3060 80
rect 3072 68 3147 80
rect 3205 68 3280 80
rect 3292 68 3323 80
rect 3329 68 3364 80
rect 2998 66 3160 68
rect 2893 38 2934 46
rect 3016 38 3029 66
rect 3044 64 3059 66
rect 3083 39 3090 46
rect 3093 38 3160 66
rect 3192 66 3364 68
rect 3162 44 3190 48
rect 3192 44 3272 66
rect 3293 64 3308 66
rect 3162 42 3272 44
rect 3162 38 3190 42
rect 3192 38 3272 42
rect 2799 28 2829 38
rect 2856 28 2857 38
rect 2872 28 2885 38
rect 2899 28 2900 38
rect 2915 28 2928 38
rect 2943 28 2973 38
rect 3016 28 3059 38
rect 3066 28 3074 38
rect 3093 30 3096 38
rect 3160 30 3192 38
rect 3093 28 3259 30
rect 3278 28 3289 38
rect 3293 28 3323 38
rect 3351 28 3364 66
rect 3436 72 3471 80
rect 3436 46 3437 72
rect 3444 46 3471 72
rect 3436 38 3471 46
rect 3473 72 3514 80
rect 3473 46 3488 72
rect 3495 46 3514 72
rect 3578 68 3640 80
rect 3652 68 3727 80
rect 3785 68 3860 80
rect 3872 68 3903 80
rect 3909 68 3944 80
rect 3578 66 3740 68
rect 3473 38 3514 46
rect 3596 38 3609 66
rect 3624 64 3639 66
rect 3663 39 3670 46
rect 3673 38 3740 66
rect 3772 66 3944 68
rect 3742 44 3770 48
rect 3772 44 3852 66
rect 3873 64 3888 66
rect 3742 42 3852 44
rect 3742 38 3770 42
rect 3772 38 3852 42
rect 3379 28 3409 38
rect 3436 28 3437 38
rect 3452 28 3465 38
rect 3479 28 3480 38
rect 3495 28 3508 38
rect 3523 28 3553 38
rect 3596 28 3639 38
rect 3646 28 3654 38
rect 3673 30 3676 38
rect 3740 30 3772 38
rect 3673 28 3839 30
rect 3858 28 3869 38
rect 3873 28 3903 38
rect 3931 28 3944 66
rect 4016 72 4051 80
rect 4016 46 4017 72
rect 4024 46 4051 72
rect 4016 38 4051 46
rect 4053 72 4094 80
rect 4053 46 4068 72
rect 4075 46 4094 72
rect 4158 68 4220 80
rect 4232 68 4307 80
rect 4365 68 4440 80
rect 4452 68 4483 80
rect 4489 68 4524 80
rect 4158 66 4320 68
rect 4053 38 4094 46
rect 4176 38 4189 66
rect 4204 64 4219 66
rect 4243 39 4250 46
rect 4253 38 4320 66
rect 4352 66 4524 68
rect 4322 44 4350 48
rect 4352 44 4432 66
rect 4453 64 4468 66
rect 4322 42 4432 44
rect 4322 38 4350 42
rect 4352 38 4432 42
rect 3959 28 3989 38
rect 4016 28 4017 38
rect 4032 28 4045 38
rect 4059 28 4060 38
rect 4075 28 4088 38
rect 4103 28 4133 38
rect 4176 28 4219 38
rect 4226 28 4234 38
rect 4253 30 4256 38
rect 4320 30 4352 38
rect 4253 28 4419 30
rect 4438 28 4449 38
rect 4453 28 4483 38
rect 4511 28 4524 66
rect 4596 72 4631 80
rect 4596 46 4597 72
rect 4604 46 4631 72
rect 4596 38 4631 46
rect 4539 28 4569 38
rect 4596 28 4597 38
rect 4612 28 4625 38
rect -1 22 4625 28
rect 0 14 4625 22
rect 15 0 28 14
rect 43 -4 73 14
rect 116 0 129 14
rect 166 1 174 14
rect 207 1 345 14
rect 378 1 386 14
rect 243 0 294 1
rect 451 0 464 14
rect 244 -2 308 0
rect 479 -4 509 14
rect 552 0 565 14
rect 595 0 608 14
rect 623 -4 653 14
rect 696 0 709 14
rect 746 1 754 14
rect 787 1 925 14
rect 958 1 966 14
rect 823 0 874 1
rect 1031 0 1044 14
rect 824 -2 888 0
rect 1059 -4 1089 14
rect 1132 0 1145 14
rect 1175 0 1188 14
rect 1203 -4 1233 14
rect 1276 0 1289 14
rect 1326 1 1334 14
rect 1367 1 1505 14
rect 1538 1 1546 14
rect 1403 0 1454 1
rect 1611 0 1624 14
rect 1404 -2 1468 0
rect 1639 -4 1669 14
rect 1712 0 1725 14
rect 1755 0 1768 14
rect 1783 -4 1813 14
rect 1856 0 1869 14
rect 1906 1 1914 14
rect 1947 1 2085 14
rect 2118 1 2126 14
rect 1983 0 2034 1
rect 2191 0 2204 14
rect 1984 -2 2048 0
rect 2219 -4 2249 14
rect 2292 0 2305 14
rect 2335 0 2348 14
rect 2363 -4 2393 14
rect 2436 0 2449 14
rect 2486 1 2494 14
rect 2527 1 2665 14
rect 2698 1 2706 14
rect 2563 0 2614 1
rect 2771 0 2784 14
rect 2564 -2 2628 0
rect 2799 -4 2829 14
rect 2872 0 2885 14
rect 2915 0 2928 14
rect 2943 -4 2973 14
rect 3016 0 3029 14
rect 3066 1 3074 14
rect 3107 1 3245 14
rect 3278 1 3286 14
rect 3143 0 3194 1
rect 3351 0 3364 14
rect 3144 -2 3208 0
rect 3379 -4 3409 14
rect 3452 0 3465 14
rect 3495 0 3508 14
rect 3523 -4 3553 14
rect 3596 0 3609 14
rect 3646 1 3654 14
rect 3687 1 3825 14
rect 3858 1 3866 14
rect 3723 0 3774 1
rect 3931 0 3944 14
rect 3724 -2 3788 0
rect 3959 -4 3989 14
rect 4032 0 4045 14
rect 4075 0 4088 14
rect 4103 -4 4133 14
rect 4176 0 4189 14
rect 4226 1 4234 14
rect 4267 1 4405 14
rect 4438 1 4446 14
rect 4303 0 4354 1
rect 4511 0 4524 14
rect 4304 -2 4368 0
rect 4539 -4 4569 14
rect 4612 0 4625 14
<< pwell >>
rect 74 184 89 212
rect 464 184 479 213
rect 0 38 15 80
rect 537 38 552 80
rect 580 38 595 80
<< ndiffc >>
rect 74 184 89 212
rect 464 184 479 213
rect 654 184 669 212
rect 1044 184 1059 213
rect 1234 184 1249 212
rect 1624 184 1639 213
rect 1814 184 1829 212
rect 2204 184 2219 213
rect 2394 184 2409 212
rect 2784 184 2799 213
rect 2974 184 2989 212
rect 3364 184 3379 213
rect 3554 184 3569 212
rect 3944 184 3959 213
rect 4134 184 4149 212
rect 4524 184 4539 213
rect 0 38 15 80
rect 537 38 552 80
rect 580 38 595 80
rect 1117 38 1132 80
rect 1160 38 1175 80
rect 1697 38 1712 80
rect 1740 38 1755 80
rect 2277 38 2292 80
rect 2320 38 2335 80
rect 2857 38 2872 80
rect 2900 38 2915 80
rect 3437 38 3452 80
rect 3480 38 3495 80
rect 4017 38 4032 80
rect 4060 38 4075 80
rect 4597 38 4612 80
<< poly >>
rect 0 510 30 540
rect 0 240 30 270
<< metal1 >>
rect 0 496 15 510
rect 0 372 15 406
rect 0 270 15 284
rect 0 226 15 240
rect 0 102 15 136
rect 0 0 15 14
use 10T_1x8_magic  10T_1x8_magic_1
timestamp 1656019537
transform 1 0 0 0 1 0
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_0
timestamp 1656019537
transform 1 0 0 0 1 270
box -7 -4 4631 312
<< labels >>
rlabel locali 74 184 89 212 1 WBLb_0
port 21 ns signal input
rlabel locali 464 184 479 213 1 WBL_0
port 22 ns signal input
rlabel locali 0 38 15 80 1 RBL1_0
port 1 ns signal output
rlabel locali 537 38 552 80 1 RBL0_0
port 2 ns signal output
rlabel locali 654 184 669 212 1 WBLb_1
port 23 ns signal input
rlabel locali 1044 184 1059 213 1 WBL_1
port 24 ns signal input
rlabel locali 580 38 595 80 1 RBL1_1
port 3 ns signal output
rlabel locali 1117 38 1132 80 1 RBL0_1
port 4 ns signal output
rlabel locali 1234 184 1249 212 1 WBLb_2
port 25 ns signal input
rlabel locali 1624 184 1639 213 1 WBL_2
port 26 ns signal input
rlabel locali 1160 38 1175 80 1 RBL1_2
port 5 ns signal output
rlabel locali 1697 38 1712 80 1 RBL0_2
port 6 ns signal output
rlabel locali 1814 184 1829 212 1 WBLb_3
port 27 ns signal input
rlabel locali 2204 184 2219 213 1 WBL_3
port 28 ns signal input
rlabel locali 1740 38 1755 80 1 RBL1_3
port 7 ns signal output
rlabel locali 2277 38 2292 80 1 RBL0_3
port 8 ns signal output
rlabel locali 2394 184 2409 212 1 WBLb_4
port 29 ns signal input
rlabel locali 2784 184 2799 213 1 WBL_4
port 30 ns signal input
rlabel locali 2320 38 2335 80 1 RBL1_4
port 8 ns signal output
rlabel locali 2857 38 2872 80 1 RBL0_4
port 10 ns signal output
rlabel locali 2974 184 2989 212 1 WBLb_5
port 31 ns signal input
rlabel locali 3364 184 3379 213 1 WBL_5
port 32 ns signal input
rlabel locali 2900 38 2915 80 1 RBL1_5
port 11 ns signal output
rlabel locali 3437 38 3452 80 1 RBL0_5
port 12 ns signal output
rlabel locali 3554 184 3569 212 1 WBLb_6
port 33 ns signal input
rlabel locali 3944 184 3959 213 1 WBL_6
port 32 ns signal input
rlabel locali 3480 38 3495 80 1 RBL1_6
port 13 ns signal output
rlabel locali 4017 38 4032 80 1 RBL0_6
port 14 ns signal output
rlabel locali 4134 184 4149 212 1 WBLb_7
port 33 ns signal input
rlabel locali 4524 184 4539 213 1 WBL_7
port 34 ns signal input
rlabel locali 4060 38 4075 80 1 RBL1_7
port 15 ns signal output
rlabel locali 4597 38 4612 80 1 RBL0_7
port 16 ns signal output
rlabel poly 0 510 30 540 1 WWL_0
port 17 ew signal input
rlabel poly 0 240 30 270 1 WWL_1
port 18 ew signal input
rlabel metal1 0 372 15 406 1 RWL_0
port 19 ew signal input
rlabel metal1 0 102 15 136 1 RWL_1
port 20 ew signal input
rlabel metal1 0 496 15 510 1 VDD
port 35 ew power bidirectional abutment
rlabel metal1 0 226 15 240 1 VDD
rlabel metal1 0 270 15 284 1 GND
port 36 ew ground bidirectional abutment
rlabel metal1 0 0 15 14 1 GND
<< end >>
