magic
tech sky130A
magscale 1 2
timestamp 1656018194
<< error_s >>
rect 9 258 22 274
rect 111 272 124 322
rect 77 258 92 272
rect 101 258 131 272
rect 192 270 345 316
rect 174 258 366 270
rect 409 258 439 272
rect 445 258 458 322
rect 546 258 559 274
rect 589 258 602 274
rect 691 272 704 322
rect 657 258 672 272
rect 681 258 711 272
rect 772 270 925 316
rect 754 258 946 270
rect 989 258 1019 272
rect 1025 258 1038 322
rect 1126 258 1139 274
rect -54 244 1139 258
rect 9 140 22 244
rect 67 222 68 232
rect 88 230 96 232
rect 86 228 96 230
rect 83 222 96 228
rect 67 218 96 222
rect 101 218 131 244
rect 149 230 165 232
rect 237 230 288 244
rect 238 228 302 230
rect 345 228 360 244
rect 409 241 439 244
rect 409 238 445 241
rect 375 230 391 232
rect 149 218 164 222
rect 67 216 164 218
rect 192 216 360 228
rect 376 218 391 222
rect 409 219 448 238
rect 467 232 474 233
rect 473 225 474 232
rect 457 222 458 225
rect 473 222 486 225
rect 409 218 439 219
rect 448 218 454 219
rect 457 218 486 222
rect 376 217 486 218
rect 376 216 492 217
rect 51 208 102 216
rect 51 196 76 208
rect 83 196 102 208
rect 133 208 183 216
rect 133 200 149 208
rect 156 206 183 208
rect 192 206 413 216
rect 156 196 413 206
rect 442 208 492 216
rect 442 199 458 208
rect 51 188 102 196
rect 149 188 413 196
rect 439 196 458 199
rect 465 196 492 208
rect 439 188 492 196
rect 67 180 68 188
rect 83 180 96 188
rect 67 172 83 180
rect 64 165 83 168
rect 64 156 86 165
rect 37 146 86 156
rect 37 140 67 146
rect 86 141 91 146
rect 9 124 83 140
rect 101 132 131 188
rect 166 178 374 188
rect 409 184 454 188
rect 457 187 458 188
rect 473 187 486 188
rect 192 148 381 178
rect 207 145 381 148
rect 200 142 381 145
rect 9 122 22 124
rect 37 122 71 124
rect 9 106 83 122
rect 110 118 123 132
rect 138 118 154 134
rect 200 129 211 142
rect -7 84 -6 100
rect 9 84 22 106
rect 37 84 67 106
rect 110 102 172 118
rect 200 111 211 127
rect 216 122 226 142
rect 236 122 250 142
rect 253 129 262 142
rect 278 129 287 142
rect 216 111 250 122
rect 253 111 262 127
rect 278 111 287 127
rect 294 122 304 142
rect 314 122 328 142
rect 329 129 340 142
rect 294 111 328 122
rect 329 111 340 127
rect 386 118 402 134
rect 409 132 439 184
rect 473 180 474 187
rect 458 172 474 180
rect 445 140 458 159
rect 473 140 503 156
rect 445 124 519 140
rect 445 122 458 124
rect 473 122 507 124
rect 110 100 123 102
rect 138 100 172 102
rect 110 84 172 100
rect 216 95 232 98
rect 294 95 324 106
rect 372 102 418 118
rect 445 106 519 122
rect 372 100 406 102
rect 371 84 418 100
rect 445 84 458 106
rect 473 84 503 106
rect 530 84 531 100
rect 546 84 559 244
rect 589 140 602 244
rect 647 222 648 232
rect 668 230 676 232
rect 666 228 676 230
rect 663 222 676 228
rect 647 218 676 222
rect 681 218 711 244
rect 729 230 745 232
rect 817 230 868 244
rect 818 228 882 230
rect 925 228 940 244
rect 989 241 1019 244
rect 989 238 1025 241
rect 955 230 971 232
rect 729 218 744 222
rect 647 216 744 218
rect 772 216 940 228
rect 956 218 971 222
rect 989 219 1028 238
rect 1047 232 1054 233
rect 1053 225 1054 232
rect 1037 222 1038 225
rect 1053 222 1066 225
rect 989 218 1019 219
rect 1028 218 1034 219
rect 1037 218 1066 222
rect 956 217 1066 218
rect 956 216 1072 217
rect 631 208 682 216
rect 631 196 656 208
rect 663 196 682 208
rect 713 208 763 216
rect 713 200 729 208
rect 736 206 763 208
rect 772 206 993 216
rect 736 196 993 206
rect 1022 208 1072 216
rect 1022 199 1038 208
rect 631 188 682 196
rect 729 188 993 196
rect 1019 196 1038 199
rect 1045 196 1072 208
rect 1019 188 1072 196
rect 647 180 648 188
rect 663 180 676 188
rect 647 172 663 180
rect 644 165 663 168
rect 644 156 666 165
rect 617 146 666 156
rect 617 140 647 146
rect 666 141 671 146
rect 589 124 663 140
rect 681 132 711 188
rect 746 178 954 188
rect 989 184 1034 188
rect 1037 187 1038 188
rect 1053 187 1066 188
rect 772 148 961 178
rect 787 145 961 148
rect 780 142 961 145
rect 589 122 602 124
rect 617 122 651 124
rect 589 106 663 122
rect 690 118 703 132
rect 718 118 734 134
rect 780 129 791 142
rect 573 84 574 100
rect 589 84 602 106
rect 617 84 647 106
rect 690 102 752 118
rect 780 111 791 127
rect 796 122 806 142
rect 816 122 830 142
rect 833 129 842 142
rect 858 129 867 142
rect 796 111 830 122
rect 833 111 842 127
rect 858 111 867 127
rect 874 122 884 142
rect 894 122 908 142
rect 909 129 920 142
rect 874 111 908 122
rect 909 111 920 127
rect 966 118 982 134
rect 989 132 1019 184
rect 1053 180 1054 187
rect 1038 172 1054 180
rect 1025 140 1038 159
rect 1053 140 1083 156
rect 1025 124 1099 140
rect 1025 122 1038 124
rect 1053 122 1087 124
rect 690 100 703 102
rect 718 100 752 102
rect 690 84 752 100
rect 796 95 812 98
rect 874 95 904 106
rect 952 102 998 118
rect 1025 106 1099 122
rect 952 100 986 102
rect 951 84 998 100
rect 1025 84 1038 106
rect 1053 84 1083 106
rect 1110 84 1111 100
rect 1126 84 1139 244
rect -13 76 28 84
rect -13 50 2 76
rect 9 50 28 76
rect 92 72 154 84
rect 166 72 241 84
rect 299 72 374 84
rect 386 72 417 84
rect 423 72 458 84
rect 92 70 254 72
rect -13 42 28 50
rect 110 46 123 70
rect 138 68 153 70
rect 187 52 254 70
rect 286 70 458 72
rect 286 52 366 70
rect 387 68 402 70
rect -7 32 -6 42
rect 9 32 22 42
rect 37 32 67 46
rect 110 32 153 46
rect 177 43 184 50
rect 187 42 366 52
rect 160 32 190 42
rect 192 32 345 42
rect 353 32 383 42
rect 387 32 417 46
rect 445 32 458 70
rect 530 76 565 84
rect 530 50 531 76
rect 538 50 565 76
rect 473 32 503 46
rect 530 42 565 50
rect 567 76 608 84
rect 567 50 582 76
rect 589 50 608 76
rect 672 72 734 84
rect 746 72 821 84
rect 879 72 954 84
rect 966 72 997 84
rect 1003 72 1038 84
rect 672 70 834 72
rect 567 42 608 50
rect 690 46 703 70
rect 718 68 733 70
rect 767 52 834 70
rect 866 70 1038 72
rect 866 52 946 70
rect 967 68 982 70
rect 530 32 531 42
rect 546 32 559 42
rect 573 32 574 42
rect 589 32 602 42
rect 617 32 647 46
rect 690 32 733 46
rect 757 43 764 50
rect 767 42 946 52
rect 740 32 770 42
rect 772 32 925 42
rect 933 32 963 42
rect 967 32 997 46
rect 1025 32 1038 70
rect 1110 76 1145 84
rect 1110 50 1111 76
rect 1118 50 1145 76
rect 1053 32 1083 46
rect 1110 42 1145 50
rect 1110 32 1111 42
rect 1126 32 1139 42
rect -54 18 1139 32
rect 9 -12 22 18
rect 37 0 67 18
rect 110 4 124 18
rect 160 4 380 18
rect 111 2 124 4
rect 77 -10 92 2
rect 74 -12 96 -10
rect 101 -12 131 2
rect 192 0 345 4
rect 174 -12 366 0
rect 409 -12 439 2
rect 445 -12 458 18
rect 473 0 503 18
rect 546 -12 559 18
rect 589 -12 602 18
rect 617 0 647 18
rect 690 4 704 18
rect 740 4 960 18
rect 691 2 704 4
rect 657 -10 672 2
rect 654 -12 676 -10
rect 681 -12 711 2
rect 772 0 925 4
rect 754 -12 946 0
rect 989 -12 1019 2
rect 1025 -12 1038 18
rect 1053 0 1083 18
rect 1126 -12 1139 18
rect -54 -26 1139 -12
rect 9 -130 22 -26
rect 67 -48 68 -38
rect 88 -40 96 -38
rect 86 -42 96 -40
rect 83 -48 96 -42
rect 67 -52 96 -48
rect 101 -52 131 -26
rect 149 -40 165 -38
rect 237 -40 288 -26
rect 238 -42 302 -40
rect 149 -52 164 -48
rect 67 -54 164 -52
rect 51 -62 102 -54
rect 51 -74 76 -62
rect 83 -74 102 -62
rect 133 -62 183 -54
rect 133 -70 149 -62
rect 156 -64 183 -62
rect 192 -62 207 -58
rect 254 -62 286 -42
rect 345 -54 360 -26
rect 409 -29 439 -26
rect 409 -32 445 -29
rect 375 -40 391 -38
rect 376 -52 391 -48
rect 409 -51 448 -32
rect 467 -38 474 -37
rect 473 -45 474 -38
rect 457 -48 458 -45
rect 473 -48 486 -45
rect 409 -52 439 -51
rect 448 -52 454 -51
rect 457 -52 486 -48
rect 376 -53 486 -52
rect 376 -54 492 -53
rect 345 -62 413 -54
rect 192 -64 261 -62
rect 279 -64 413 -62
rect 156 -68 228 -64
rect 156 -70 281 -68
rect 156 -74 228 -70
rect 51 -82 102 -74
rect 149 -78 228 -74
rect 309 -78 413 -64
rect 442 -62 492 -54
rect 442 -71 458 -62
rect 149 -82 413 -78
rect 439 -74 458 -71
rect 465 -74 492 -62
rect 439 -82 492 -74
rect 67 -90 68 -82
rect 83 -90 96 -82
rect 67 -98 83 -90
rect 64 -105 83 -102
rect 64 -114 86 -105
rect 37 -124 86 -114
rect 37 -130 67 -124
rect 86 -129 91 -124
rect 9 -146 83 -130
rect 101 -138 131 -82
rect 166 -92 374 -82
rect 409 -86 454 -82
rect 457 -83 458 -82
rect 473 -83 486 -82
rect 333 -96 381 -92
rect 216 -118 246 -109
rect 309 -116 324 -109
rect 345 -118 381 -96
rect 192 -122 381 -118
rect 207 -125 381 -122
rect 200 -128 381 -125
rect 9 -148 22 -146
rect 37 -148 71 -146
rect 9 -164 83 -148
rect 110 -152 123 -138
rect 138 -152 154 -136
rect 200 -141 211 -128
rect -7 -186 -6 -170
rect 9 -186 22 -164
rect 37 -186 67 -164
rect 110 -168 172 -152
rect 200 -159 211 -143
rect 216 -148 226 -128
rect 236 -148 250 -128
rect 253 -141 262 -128
rect 278 -141 287 -128
rect 216 -159 250 -148
rect 253 -159 262 -143
rect 278 -159 287 -143
rect 294 -148 304 -128
rect 314 -148 328 -128
rect 329 -141 340 -128
rect 294 -159 328 -148
rect 329 -159 340 -143
rect 386 -152 402 -136
rect 409 -138 439 -86
rect 473 -90 474 -83
rect 458 -98 474 -90
rect 445 -130 458 -111
rect 473 -130 503 -114
rect 445 -146 519 -130
rect 445 -148 458 -146
rect 473 -148 507 -146
rect 110 -170 123 -168
rect 138 -170 172 -168
rect 110 -186 172 -170
rect 216 -175 232 -172
rect 294 -175 324 -164
rect 372 -168 418 -152
rect 445 -164 519 -148
rect 372 -170 406 -168
rect 371 -186 418 -170
rect 445 -186 458 -164
rect 473 -186 503 -164
rect 530 -186 531 -170
rect 546 -186 559 -26
rect 589 -130 602 -26
rect 647 -48 648 -38
rect 668 -40 676 -38
rect 666 -42 676 -40
rect 663 -48 676 -42
rect 647 -52 676 -48
rect 681 -52 711 -26
rect 729 -40 745 -38
rect 817 -40 868 -26
rect 818 -42 882 -40
rect 729 -52 744 -48
rect 647 -54 744 -52
rect 631 -62 682 -54
rect 631 -74 656 -62
rect 663 -74 682 -62
rect 713 -62 763 -54
rect 713 -70 729 -62
rect 736 -64 763 -62
rect 772 -62 787 -58
rect 834 -62 866 -42
rect 925 -54 940 -26
rect 989 -29 1019 -26
rect 989 -32 1025 -29
rect 955 -40 971 -38
rect 956 -52 971 -48
rect 989 -51 1028 -32
rect 1047 -38 1054 -37
rect 1053 -45 1054 -38
rect 1037 -48 1038 -45
rect 1053 -48 1066 -45
rect 989 -52 1019 -51
rect 1028 -52 1034 -51
rect 1037 -52 1066 -48
rect 956 -53 1066 -52
rect 956 -54 1072 -53
rect 925 -62 993 -54
rect 772 -64 841 -62
rect 859 -64 993 -62
rect 736 -68 808 -64
rect 736 -70 861 -68
rect 736 -74 808 -70
rect 631 -82 682 -74
rect 729 -78 808 -74
rect 889 -78 993 -64
rect 1022 -62 1072 -54
rect 1022 -71 1038 -62
rect 729 -82 993 -78
rect 1019 -74 1038 -71
rect 1045 -74 1072 -62
rect 1019 -82 1072 -74
rect 647 -90 648 -82
rect 663 -90 676 -82
rect 647 -98 663 -90
rect 644 -105 663 -102
rect 644 -114 666 -105
rect 617 -124 666 -114
rect 617 -130 647 -124
rect 666 -129 671 -124
rect 589 -146 663 -130
rect 681 -138 711 -82
rect 746 -92 954 -82
rect 989 -86 1034 -82
rect 1037 -83 1038 -82
rect 1053 -83 1066 -82
rect 913 -96 961 -92
rect 796 -118 826 -109
rect 889 -116 904 -109
rect 925 -118 961 -96
rect 772 -122 961 -118
rect 787 -125 961 -122
rect 780 -128 961 -125
rect 589 -148 602 -146
rect 617 -148 651 -146
rect 589 -164 663 -148
rect 690 -152 703 -138
rect 718 -152 734 -136
rect 780 -141 791 -128
rect 573 -186 574 -170
rect 589 -186 602 -164
rect 617 -186 647 -164
rect 690 -168 752 -152
rect 780 -159 791 -143
rect 796 -148 806 -128
rect 816 -148 830 -128
rect 833 -141 842 -128
rect 858 -141 867 -128
rect 796 -159 830 -148
rect 833 -159 842 -143
rect 858 -159 867 -143
rect 874 -148 884 -128
rect 894 -148 908 -128
rect 909 -141 920 -128
rect 874 -159 908 -148
rect 909 -159 920 -143
rect 966 -152 982 -136
rect 989 -138 1019 -86
rect 1053 -90 1054 -83
rect 1038 -98 1054 -90
rect 1025 -130 1038 -111
rect 1053 -130 1083 -114
rect 1025 -146 1099 -130
rect 1025 -148 1038 -146
rect 1053 -148 1087 -146
rect 690 -170 703 -168
rect 718 -170 752 -168
rect 690 -186 752 -170
rect 796 -175 812 -172
rect 874 -175 904 -164
rect 952 -168 998 -152
rect 1025 -164 1099 -148
rect 952 -170 986 -168
rect 951 -186 998 -170
rect 1025 -186 1038 -164
rect 1053 -186 1083 -164
rect 1110 -186 1111 -170
rect 1126 -186 1139 -26
rect -13 -194 28 -186
rect -13 -220 2 -194
rect 9 -220 28 -194
rect 92 -198 154 -186
rect 166 -198 241 -186
rect 299 -198 374 -186
rect 386 -198 417 -186
rect 423 -198 458 -186
rect 92 -200 254 -198
rect -13 -228 28 -220
rect 110 -228 123 -200
rect 138 -202 153 -200
rect 187 -218 254 -200
rect 286 -200 458 -198
rect 286 -218 366 -200
rect 387 -202 402 -200
rect 177 -227 184 -220
rect 187 -228 366 -218
rect -7 -238 -6 -228
rect 9 -238 22 -228
rect 37 -238 67 -228
rect 110 -238 153 -228
rect 160 -238 168 -228
rect 187 -236 190 -228
rect 254 -236 286 -228
rect 187 -238 353 -236
rect 372 -238 383 -228
rect 387 -238 417 -228
rect 445 -238 458 -200
rect 530 -194 565 -186
rect 530 -220 531 -194
rect 538 -220 565 -194
rect 530 -228 565 -220
rect 567 -194 608 -186
rect 567 -220 582 -194
rect 589 -220 608 -194
rect 672 -198 734 -186
rect 746 -198 821 -186
rect 879 -198 954 -186
rect 966 -198 997 -186
rect 1003 -198 1038 -186
rect 672 -200 834 -198
rect 567 -228 608 -220
rect 690 -228 703 -200
rect 718 -202 733 -200
rect 767 -218 834 -200
rect 866 -200 1038 -198
rect 866 -218 946 -200
rect 967 -202 982 -200
rect 757 -227 764 -220
rect 767 -228 946 -218
rect 473 -238 503 -228
rect 530 -238 531 -228
rect 546 -238 559 -228
rect 573 -238 574 -228
rect 589 -238 602 -228
rect 617 -238 647 -228
rect 690 -238 733 -228
rect 740 -238 748 -228
rect 767 -236 770 -228
rect 834 -236 866 -228
rect 767 -238 933 -236
rect 952 -238 963 -228
rect 967 -238 997 -228
rect 1025 -238 1038 -200
rect 1110 -194 1145 -186
rect 1110 -220 1111 -194
rect 1118 -220 1145 -194
rect 1110 -228 1145 -220
rect 1053 -238 1083 -228
rect 1110 -238 1111 -228
rect 1126 -238 1139 -228
rect -54 -252 1139 -238
rect 9 -314 22 -252
rect 37 -270 67 -252
rect 110 -266 123 -252
rect 160 -265 168 -252
rect 201 -265 339 -252
rect 372 -265 380 -252
rect 237 -266 288 -265
rect 445 -266 458 -252
rect 254 -268 286 -266
rect 473 -270 503 -252
rect 546 -314 559 -252
rect 589 -314 602 -252
rect 617 -270 647 -252
rect 690 -266 703 -252
rect 740 -265 748 -252
rect 781 -265 919 -252
rect 952 -265 960 -252
rect 817 -266 868 -265
rect 1025 -266 1038 -252
rect 834 -268 866 -266
rect 1053 -270 1083 -252
rect 1126 -314 1139 -252
<< nwell >>
rect 834 228 866 230
rect 834 -42 866 -40
<< pwell >>
rect 254 18 286 20
rect -6 4 164 18
rect 237 -266 303 -252
rect 546 -266 574 274
rect 834 18 866 20
rect 834 -252 866 -250
<< psubdiffcont >>
rect 254 18 286 20
rect 834 18 866 20
rect 254 -252 286 -250
rect 834 -252 866 -250
<< nsubdiffcont >>
rect 254 228 286 230
rect 834 228 866 230
rect 254 -42 286 -40
rect 834 -42 866 -40
<< poly >>
rect -54 244 -6 274
rect 546 244 574 274
rect -54 -26 -6 4
rect 546 -26 574 4
<< corelocali >>
rect 96 274 111 322
rect 430 274 445 322
rect 676 274 691 322
rect 1010 274 1025 322
rect -6 -314 9 -266
rect 531 -314 546 -266
rect 574 -314 589 -266
rect 1111 -314 1126 -266
<< viali >>
rect 37 106 67 140
rect 473 106 503 140
rect 617 106 647 140
rect 1053 106 1083 140
rect 37 -164 67 -130
rect 473 -164 503 -130
rect 617 -164 647 -130
rect 1053 -164 1083 -130
<< metal1 >>
rect -54 230 -6 244
rect 546 230 574 244
rect -54 106 37 140
rect 67 106 473 140
rect 503 106 617 140
rect 647 106 1053 140
rect 1083 106 1126 140
rect -54 4 -6 18
rect 546 4 574 18
rect -54 -40 -6 -26
rect 546 -40 574 -26
rect -54 -164 37 -130
rect 67 -164 473 -130
rect 503 -164 617 -130
rect 647 -164 1053 -130
rect 1083 -164 1126 -130
rect -54 -266 -6 -252
rect 546 -266 574 -252
use 10T_toy_magic  10T_toy_magic_1
timestamp 1655238822
transform 1 0 674 0 1 23
box -107 -23 471 293
use 10T_toy_magic  10T_toy_magic_2
timestamp 1655238822
transform 1 0 94 0 1 -247
box -107 -23 471 293
use 10T_toy_magic  10T_toy_magic_0
timestamp 1655238822
transform 1 0 94 0 1 23
box -107 -23 471 293
use 10T_toy_magic  10T_toy_magic_3
timestamp 1655238822
transform 1 0 674 0 1 -247
box -107 -23 471 293
<< labels >>
rlabel poly -54 244 -24 274 1 WWL_0
rlabel poly -54 -26 -24 4 1 WWL_1
rlabel metal1 -54 230 -24 244 1 VDD
rlabel metal1 -54 -40 -24 -26 1 VDD
rlabel metal1 -54 4 -24 18 1 GND
rlabel metal1 -54 -266 -24 -252 1 GND
rlabel corelocali -6 -314 9 -284 1 RBL1_0
rlabel corelocali 531 -314 546 -284 1 RBL0_0
rlabel corelocali 574 -314 589 -284 1 RBL1_1
rlabel corelocali 1111 -314 1126 -284 1 RBL0_1
rlabel metal1 -54 -164 -24 -130 1 RWL_1
rlabel metal1 -54 106 -24 140 1 RWL_0
<< end >>
