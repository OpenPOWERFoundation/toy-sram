* HSPICE file created from 10T_32x32_magic_flattened.ext - technology: sky130A
.lib /import/angmar1/repos/openpdk/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.subckt x10T_32x32_magic_flattened RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3
+ RBL0_3 RBL1_4 RBL0_4 RBL1_5 RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 RBL1_8 RBL0_8 RBL1_9
+ RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL0_11 RBL1_12 RBL0_12 RBL1_13 RBL0_13 RBL1_14 RBL0_14
+ RBL1_15 RBL0_15 WWL_0 RWL_0 WWL_1 RWL_1 WWL_2 RWL_2 WWL_3 RWL_3 WWL_4 RWL_4 WWL_5
+ RWL_5 WWL_6 RWL_6 WWL_7 RWL_7 WWL_8 RWL_8 WWL_9 RWL_9 WWL_10 RWL_10 WWL_11 RWL_11
+ WWL_12 RWL_12 WWL_13 RWL_13 WWL_14 RWL_14 WWL_15 RWL_15 WWL_16 RWL_16 WWL_17 RWL_17
+ WWL_18 RWL_18 WWL_19 RWL_19 WWL_20 RWL_20 WWL_21 RWL_21 WWL_22 RWL_22 WWL_23 RWL_23
+ WWL_24 RWL_24 WWL_25 RWL_25 WWL_26 RWL_26 WWL_27 RWL_27 WWL_28 RWL_28 WWL_29 RWL_29
+ WWL_30 RWL_30 WWL_31 RWL_31 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19
+ RBL0_19 RBL1_20 RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 RBL1_24
+ RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL0_27 RBL1_28 RBL0_28 RBL1_29
+ RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 WBL_0 WBLb_0 WBL_1 WBLb_1 WBL_2 WBLb_2 WBL_3
+ WBLb_19 WBL_4 WBLb_4 WBL_5 WBLb_5 WBL_22 WBLb_6 WBL_7 WBLb_23 WBL_24 WBLb_8 WBL_25
+ WBLb_9 WBL_26 WBLb_10 WBL_11 WBLb_11 WBL_12 WBLb_12 WBL_13 WBLb_13 WBL_14 WBLb_30
+ WBL_15 WBLb_15 VDD GND
M1000 GND x0/junc1 x0/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1001 x1/RWL0_junc x1/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1002 x2/junc1 WWL_22 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1003 x3/junc0 x3/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1004 x4/RWL1_junc RWL_16 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1005 x5/RWL0_junc x5/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1006 x6/junc1 WWL_18 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1007 x7/RWL1_junc RWL_1 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1008 RBL0_13 RWL_2 x8/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1009 WBL_14 WWL_12 x9/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1010 x10/RWL0_junc x10/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1011 WBL_5 WWL_20 x11/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1012 x12/junc0 x12/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1013 x13/junc0 x13/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1014 x14/RWL0_junc x14/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1015 x15/junc0 x15/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1016 GND x16/junc0 x16/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1017 x17/junc0 x17/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1018 GND x18/junc1 x18/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1019 VDD x19/junc0 x19/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1020 GND x20/junc1 x20/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1021 GND x21/junc1 x21/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1022 GND x22/junc0 x22/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1023 x23/RWL1_junc RWL_3 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1024 x24/RWL0_junc x24/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1025 x25/RWL0_junc x25/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1026 x26/RWL0_junc x26/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1027 x27/RWL0_junc x27/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1028 GND x28/junc0 x28/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1029 x29/junc0 x29/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1030 VDD x30/junc0 x30/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1031 VDD x31/junc0 x31/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1032 x32/junc1 WWL_19 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1033 RBL0_22 RWL_6 x33/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1034 GND x34/junc1 x34/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1035 WBL_23 WWL_16 x35/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1036 RBL0_7 RWL_20 x36/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1037 GND x37/junc1 x37/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1038 x38/junc0 x38/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1039 RBL0_11 RWL_16 x39/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1040 GND x40/junc0 x40/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1041 RBL0_15 RWL_24 x41/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1042 x42/junc0 x42/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1043 RBL0_0 RWL_17 x43/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1044 VDD x44/junc0 x44/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1045 x45/junc1 WWL_25 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1046 x46/junc0 x46/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1047 GND x47/junc1 x47/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1048 x48/RWL1_junc RWL_19 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1049 x49/RWL0_junc x49/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1050 GND WWL_30 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1051 x50/RWL1_junc RWL_24 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1052 x51/RWL0_junc x51/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1053 x52/junc1 WWL_15 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1054 VDD x53/junc0 x53/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1055 GND x54/junc1 x54/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1056 x55/junc1 WWL_23 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1057 VDD x56/junc0 x56/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1058 x57/RWL0_junc x57/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1059 x58/junc1 WWL_28 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1060 x59/RWL0_junc x59/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1061 x60/junc1 WWL_0 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1062 RBL0_13 x61/RWL1 x62/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1063 WBL_14 WWL_13 x63/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1064 x64/RWL0_junc x64/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1065 x65/RWL1_junc RWL_27 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1066 x66/junc0 x66/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1067 x67/junc0 x67/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1068 x68/junc0 x68/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1069 x69/junc0 x69/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1070 x70/junc0 x70/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1071 WBL_31 WWL_29 x71/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1072 RBL0_11 RWL_31 x72/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1073 x73/RWL1_junc RWL_0 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1074 GND x74/junc0 x74/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1075 x75/junc0 x75/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1076 RBL0_7 RWL_9 x76/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1077 GND x77/junc1 x77/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1078 GND x78/junc1 x78/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1079 GND x79/junc1 x79/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1080 x80/RWL0_junc x80/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1081 x81/RWL0_junc x81/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1082 GND x82/junc0 x82/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1083 GND x83/junc0 x83/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1084 x84/junc1 WWL_30 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1085 x85/junc0 x85/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1086 x86/junc0 x86/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1087 VDD x87/junc0 x87/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1088 VDD x88/junc0 x88/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1089 x89/junc1 WWL_20 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1090 GND x90/junc1 x90/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1091 WBL_27 WWL_25 x91/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1092 GND x92/junc1 x92/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1093 GND x93/junc0 x93/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1094 WBL_31 WWL_21 x94/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1095 x95/RWL1_junc RWL_20 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1096 RBL0_15 RWL_25 x96/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1097 x97/junc0 x97/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1098 x98/junc0 x98/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1099 x99/junc1 WWL_26 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1100 RBL0_0 RWL_18 x100/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1101 GND x101/junc1 x101/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1102 WBL_10 WWL_6 x102/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1103 x103/junc0 x103/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1104 GND x104/junc1 x104/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1105 x105/junc0 x105/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1106 x106/RWL0_junc x106/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1107 x107/RWL1_junc RWL_25 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1108 x108/junc1 WWL_16 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1109 x109/junc1 WWL_24 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1110 x110/RWL0_junc x110/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1111 VDD x111/junc0 x111/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1112 x112/junc0 x112/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1113 x113/junc0 x113/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1114 GND x114/junc0 x114/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1115 x115/RWL0_junc x115/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1116 x116/junc1 WWL_1 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1117 VDD x117/junc0 x117/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1118 GND x118/junc1 x118/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1119 x119/junc0 x119/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1120 x120/RWL0_junc x120/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1121 GND x121/junc0 x121/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1122 x122/junc0 x122/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1123 x123/junc0 x123/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1124 x124/junc0 x124/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1125 WBL_19 WWL_10 x15/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1126 GND x125/junc1 x125/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1127 RBL0_3 RWL_14 x126/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1128 x127/RWL1_junc RWL_1 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1129 RBL0_16 RWL_2 x128/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1130 x129/junc0 x129/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1131 x130/RWL0_junc x130/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1132 x131/RWL0_junc x131/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1133 RBL0_27 RWL_4 x132/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1134 GND x133/junc0 x133/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1135 x134/RWL1_junc RWL_9 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1136 GND x135/junc0 x135/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1137 x136/junc1 WWL_31 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1138 GND x137/junc0 x137/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1139 x138/RWL1_junc RWL_13 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1140 VDD x139/junc0 x139/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1141 WBL_1 WWL_17 x29/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1142 GND x140/junc1 x140/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1143 GND x141/junc0 x141/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1144 WBL_27 WWL_26 x142/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1145 RBL0_21 RWL_10 x143/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1146 GND x144/junc1 x144/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1147 x145/junc0 x145/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1148 RBL0_15 RWL_26 x146/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1149 x147/junc0 x147/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1150 RBL0_25 RWL_6 x148/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1151 GND x149/junc1 x149/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1152 x150/junc1 WWL_27 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1153 x151/junc0 x151/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1154 RBL0_0 RWL_19 x152/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1155 WBL_10 WWL_7 x46/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1156 GND x153/junc1 x153/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1157 x154/RWL1_junc RWL_17 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1158 VDD x155/junc0 x155/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1159 RBL0_14 RWL_28 x156/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1160 VDD x157/junc0 x157/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1161 x158/RWL1_junc RWL_26 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1162 x159/RWL0_junc x159/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1163 x160/junc0 x160/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1164 x161/junc0 x161/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1165 x162/junc0 x162/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1166 RBL0_7 RWL_31 x149/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1167 x163/junc1 WWL_25 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1168 VDD x164/junc0 x164/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1169 x165/junc0 x165/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1170 x166/junc0 x166/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1171 x167/RWL0_junc x167/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1172 GND x168/junc0 x168/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1173 x169/junc0 x169/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1174 x170/junc1 WWL_6 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1175 WBL_28 WWL_3 x69/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1176 RBL0_12 RWL_7 x87/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1177 x171/junc1 WWL_14 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1178 GND x172/junc1 x172/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1179 WBL_19 WWL_11 x70/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1180 RBL0_3 RWL_15 x173/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1181 RBL0_16 x61/RWL1 x61/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1182 x174/junc0 x174/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1183 x95/RWL0_junc x95/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1184 x175/RWL0_junc x175/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1185 GND x176/junc0 x176/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1186 x177/RWL0_junc x177/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1187 GND x178/junc0 x178/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1188 x179/RWL1_junc RWL_10 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1189 VDD x180/junc0 x180/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1190 RBL0_27 RWL_5 x181/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1191 VDD x182/junc0 x182/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1192 GND x183/junc1 x183/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1193 GND x184/junc1 x184/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1194 GND x185/junc0 x185/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1195 GND x186/junc0 x186/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1196 x187/junc0 x187/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1197 WBL_1 WWL_18 x86/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1198 x188/RWL1_junc RWL_30 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1199 x189/junc1 WWL_10 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1200 x190/junc0 x190/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1201 VDD x191/junc0 x191/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1202 x192/junc0 x192/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1203 x193/junc0 x193/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1204 WBL_27 WWL_27 x194/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1205 VDD x195/junc0 x195/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1206 RBL0_21 RWL_11 x196/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1207 WBL_10 WWL_8 x103/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1208 GND x197/junc0 x197/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1209 x198/RWL1_junc RWL_14 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1210 RBL0_10 RWL_30 x199/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1211 x6/RWL1_junc RWL_18 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1212 RBL0_14 RWL_29 x200/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1213 VDD x201/junc0 x201/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1214 x202/junc0 x202/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1215 x203/junc0 x203/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1216 x204/junc0 x204/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1217 GND x205/junc0 x205/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1218 WBL_13 WWL_6 x112/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1219 x206/junc0 x206/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1220 x0/junc0 x0/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1221 WBL_4 WWL_14 x113/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1222 GND x207/junc1 x207/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1223 x208/junc1 WWL_26 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1224 x134/RWL0_junc x134/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1225 VDD x209/junc0 x209/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1226 RBL0_29 RWL_27 x210/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1227 VDD x211/junc0 x211/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1228 x212/junc1 WWL_28 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1229 x213/RWL0_junc x213/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1230 GND x214/junc0 x214/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1231 x215/junc1 WWL_7 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1232 WBL_28 WWL_4 x124/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1233 RBL0_12 RWL_8 x139/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1234 RBL0_3 RWL_16 x216/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1235 x217/junc0 x217/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1236 GND x218/junc0 x218/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1237 GND x219/junc1 x219/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1238 x220/RWL1_junc RWL_11 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1239 x221/junc0 x221/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1240 GND x222/junc0 x222/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1241 x223/junc0 x223/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1242 x224/junc0 x224/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1243 RBL0_6 RWL_14 x225/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1244 x226/junc0 x226/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1245 RBL0_20 RWL_28 x227/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1246 VDD x228/junc0 x228/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1247 x229/junc1 WWL_15 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1248 VDD x230/junc0 x230/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1249 GND x231/junc1 x231/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1250 x232/RWL1_junc RWL_17 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1251 x233/RWL0_junc x233/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1252 x234/junc1 WWL_29 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1253 x235/junc0 x235/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1254 RBL0_30 RWL_4 x236/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1255 x237/junc1 WWL_11 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1256 VDD x238/junc0 x238/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1257 x239/junc0 x239/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1258 RBL0_21 RWL_12 x240/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1259 VDD x241/junc0 x241/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1260 WBL_15 WWL_5 x242/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1261 GND x243/junc0 x243/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1262 RBL0_3 RWL_31 x244/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1263 x245/RWL1_junc RWL_15 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1264 x246/junc1 WWL_22 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1265 x247/RWL1_junc RWL_19 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1266 x248/junc0 x248/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1267 x249/junc0 x249/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1268 x60/RWL1_junc RWL_0 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1269 x138/junc0 x138/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1270 x250/junc0 x250/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1271 x251/RWL1_junc RWL_31 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1272 x252/junc0 x252/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1273 GND x253/junc0 x253/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1274 x231/junc0 x231/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1275 VDD x254/junc0 x254/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1276 x54/junc0 x54/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1277 WBL_13 WWL_7 x161/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1278 x255/RWL0_junc x255/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1279 GND x256/junc1 x256/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1280 x257/junc1 WWL_27 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1281 GND x258/junc0 x258/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1282 WBL_24 WWL_9 x165/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1283 GND x259/junc1 x259/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1284 GND x260/junc0 x260/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1285 GND x261/junc0 x261/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1286 x262/junc1 WWL_8 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1287 GND x263/junc0 x263/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1288 GND x264/junc1 x264/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1289 GND x265/junc1 x265/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1290 x266/junc0 x266/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1291 GND x267/junc1 x267/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1292 WBL_18 WWL_15 x268/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1293 GND x269/junc0 x269/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1294 x270/junc1 WWL_6 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1295 x9/RWL1_junc RWL_12 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1296 x271/junc0 x271/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1297 x272/junc0 x272/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1298 x273/junc1 WWL_14 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1299 x274/junc0 x274/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1300 RBL0_6 RWL_15 x275/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1301 x276/RWL0_junc x276/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1302 GND x277/junc0 x277/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1303 RBL0_20 RWL_29 x278/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1304 x279/junc0 x279/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1305 x280/junc0 x280/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1306 VDD x281/junc0 x281/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1307 x282/junc1 WWL_16 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1308 GND x283/junc1 x283/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1309 x284/junc0 x284/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1310 x285/RWL1_junc RWL_18 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1311 RBL0_30 RWL_5 x286/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1312 GND x287/junc0 x287/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1313 VDD x288/junc0 x288/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1314 x289/junc0 x289/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1315 x290/RWL1_junc RWL_20 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1316 x291/junc1 WWL_23 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1317 x35/RWL1_junc RWL_16 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1318 x292/RWL0_junc x292/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1319 x84/RWL1_junc RWL_30 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1320 x116/RWL1_junc RWL_1 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1321 RBL0_8 RWL_2 x293/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1322 WBL_9 WWL_12 x202/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1323 x294/RWL0_junc x294/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1324 VDD x295/junc0 x295/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1325 WBL_13 WWL_8 x206/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1326 x296/RWL0_junc x296/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1327 RBL0_23 RWL_30 x297/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1328 GND x298/junc1 x298/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1329 GND x299/junc1 x299/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1330 GND x300/junc0 x300/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1331 x301/RWL0_junc x301/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1332 GND x297/junc1 x297/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1333 VDD x91/junc0 x91/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1334 GND x302/junc1 x302/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1335 GND x303/junc0 x303/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1336 VDD x304/junc0 x304/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1337 VDD x305/junc0 x305/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1338 x306/junc1 WWL_19 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1339 RBL0_17 RWL_6 x270/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1340 GND x307/junc1 x307/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1341 WBL_18 WWL_16 x217/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1342 x308/junc1 WWL_7 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1343 x210/RWL0_junc x210/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1344 RBL0_2 RWL_20 x241/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1345 x309/junc0 x309/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1346 x310/junc0 x310/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1347 x311/junc0 x311/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1348 RBL0_6 RWL_16 x312/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1349 GND x313/junc0 x313/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1350 GND x314/junc0 x314/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1351 x315/RWL1_junc RWL_9 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1352 VDD x316/junc0 x316/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1353 x317/junc1 WWL_9 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1354 RBL0_10 RWL_24 x34/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1355 x318/junc0 x318/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1356 GND x319/junc1 x319/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1357 VDD x320/junc0 x320/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1358 x321/junc0 x321/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1359 GND x322/junc1 x322/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1360 x323/RWL1_junc RWL_19 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1361 x324/RWL1_junc RWL_31 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1362 x325/RWL0_junc x325/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1363 x326/junc0 x326/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1364 VDD x327/junc0 x327/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1365 x328/junc1 WWL_15 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1366 x329/RWL0_junc x329/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1367 WBL_20 WWL_3 x147/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1368 x50/junc1 WWL_24 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1369 WBL_30 WWL_28 x117/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1370 x330/RWL0_junc x330/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1371 RBL0_8 x61/RWL1 x331/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1372 WBL_9 WWL_13 x138/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1373 x332/RWL0_junc x332/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1374 x333/junc0 x333/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1375 VDD x334/junc0 x334/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1376 x335/junc0 x335/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1377 x336/junc0 x336/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1378 x337/RWL1_junc RWL_0 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1379 RBL0_2 RWL_9 x338/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1380 GND x339/junc1 x339/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1381 GND x340/junc1 x340/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1382 GND x341/junc0 x341/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1383 GND x342/junc0 x342/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1384 GND x343/junc0 x343/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1385 VDD x344/junc0 x344/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1386 x345/junc1 WWL_12 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1387 x346/junc1 WWL_30 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1388 x82/junc0 x82/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1389 VDD x347/junc0 x347/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1390 VDD x348/junc0 x348/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1391 x349/junc1 WWL_20 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1392 x350/junc1 WWL_8 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1393 x351/junc0 x351/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1394 x352/junc0 x352/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1395 x353/junc0 x353/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1396 WBL_22 WWL_25 x354/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1397 x355/RWL1_junc RWL_2 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1398 x356/RWL1_junc RWL_6 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1399 GND x357/junc0 x357/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1400 GND x358/junc0 x358/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1401 WBL_26 WWL_21 x280/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1402 x359/junc0 x359/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1403 VDD x360/junc0 x360/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1404 RBL0_10 RWL_25 x90/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1405 x361/junc0 x361/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1406 x362/junc0 x362/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1407 GND x363/junc1 x363/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1408 GND x364/junc1 x364/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1409 WBL_5 WWL_6 x284/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1410 x365/junc0 x365/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1411 x366/RWL0_junc x366/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1412 x367/junc0 x367/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1413 VDD x368/junc0 x368/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1414 x369/junc1 WWL_16 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1415 x233/junc0 x233/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1416 RBL0_13 RWL_0 x370/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1417 WBL_20 WWL_4 x371/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1418 VDD x372/junc0 x372/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1419 x373/RWL0_junc x373/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1420 x374/junc0 x374/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1421 GND x375/junc0 x375/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1422 x376/junc0 x376/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1423 GND x377/junc1 x377/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1424 GND x378/junc1 x378/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1425 x379/RWL1_junc RWL_1 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1426 RBL0_11 RWL_2 x380/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1427 x381/RWL0_junc x381/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1428 x382/junc0 x382/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1429 GND x383/junc1 x383/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1430 x384/RWL0_junc x384/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1431 x385/junc0 x385/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1432 x386/RWL0_junc x386/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1433 x387/RWL0_junc x387/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1434 x388/junc0 x388/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1435 x389/junc1 WWL_3 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1436 RBL0_22 RWL_4 x390/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1437 GND x391/junc1 x391/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1438 GND x392/junc0 x392/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1439 GND x393/junc0 x393/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1440 x394/junc1 WWL_31 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1441 GND x395/junc0 x395/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1442 x396/RWL1_junc RWL_13 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1443 VDD x397/junc0 x397/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1444 VDD x398/junc0 x398/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1445 x399/junc1 WWL_13 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1446 GND x400/junc0 x400/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1447 x141/junc0 x141/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1448 WBL_22 WWL_26 x311/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1449 x401/junc0 x401/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1450 WBL_30 WWL_22 x310/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1451 x402/RWL0_junc x402/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1452 x69/RWL1_junc x389/RWL1 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1453 x212/RWL1_junc RWL_28 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1454 GND x403/junc1 x403/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1455 GND x404/junc0 x404/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1456 x405/junc0 x405/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1457 RBL0_10 RWL_26 x140/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1458 x406/junc0 x406/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1459 GND x407/junc1 x407/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1460 x408/junc0 x408/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1461 WBL_5 WWL_7 x321/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1462 VDD x409/junc0 x409/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1463 x410/RWL0_junc x410/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1464 x411/junc0 x411/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1465 x412/RWL0_junc x412/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1466 x413/junc0 x413/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1467 RBL0_13 RWL_1 x414/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1468 x257/RWL1_junc RWL_27 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1469 x415/junc1 WWL_25 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1470 VDD x416/junc0 x416/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1471 x417/RWL0_junc x417/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1472 x315/junc0 x315/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1473 x418/junc0 x418/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1474 GND x419/junc0 x419/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1475 WBL_23 WWL_3 x335/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1476 x420/junc0 x420/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1477 x421/junc1 WWL_6 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1478 x422/junc0 x422/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1479 GND x14/junc1 x14/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1480 RBL0_7 RWL_7 x347/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1481 GND x423/junc1 x423/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1482 RBL0_11 x61/RWL1 x424/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1483 x425/junc0 x425/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1484 x426/RWL0_junc x426/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1485 GND x427/junc0 x427/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1486 x428/junc0 x428/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1487 x429/RWL1_junc RWL_10 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1488 x430/junc0 x430/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1489 x431/junc0 x431/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1490 x432/junc1 WWL_4 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1491 RBL0_22 RWL_5 x433/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1492 VDD x434/junc0 x434/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1493 GND x26/junc1 x26/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1494 GND x27/junc1 x27/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1495 x112/RWL1_junc RWL_6 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1496 GND x435/junc1 x435/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1497 GND x436/junc0 x436/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1498 GND x437/junc0 x437/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1499 VDD x242/junc0 x242/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1500 WBL_23 WWL_29 x230/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1501 WBL_31 WWL_19 x352/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1502 x438/junc1 WWL_10 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1503 WBL_30 WWL_23 x351/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1504 VDD x42/junc0 x42/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1505 x439/junc0 x439/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1506 x440/junc0 x440/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1507 WBL_22 WWL_27 x353/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1508 x441/RWL1_junc RWL_29 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1509 x442/junc0 x442/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1510 WBL_14 WWL_0 x362/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1511 RBL0_29 RWL_31 x443/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1512 WBL_5 WWL_8 x365/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1513 GND x444/junc0 x444/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1514 x445/RWL1_junc RWL_14 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1515 x446/junc0 x446/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1516 VDD x447/junc0 x447/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1517 x448/RWL0_junc x448/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1518 x449/junc0 x449/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1519 x450/junc0 x450/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1520 GND x451/junc0 x451/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1521 x452/junc0 x452/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1522 GND x57/junc1 x57/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1523 GND x453/junc1 x453/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1524 x454/junc1 WWL_26 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1525 VDD x66/junc0 x66/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1526 RBL0_24 RWL_27 x455/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1527 VDD x456/junc0 x456/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1528 VDD x68/junc0 x68/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1529 x355/junc0 x355/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1530 RBL0_16 RWL_0 x457/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1531 x458/junc1 WWL_7 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1532 x459/junc0 x459/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1533 WBL_23 WWL_4 x376/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1534 RBL0_7 RWL_8 x398/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1535 GND x460/junc0 x460/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1536 x308/RWL1_junc RWL_7 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1537 GND x461/junc0 x461/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1538 GND x80/junc1 x80/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1539 x462/RWL1_junc RWL_11 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1540 x463/junc0 x463/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1541 WBL_16 WWL_22 x388/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1542 x464/junc0 x464/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1543 WBL_1 WWL_15 x465/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1544 GND x81/junc1 x81/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1545 x466/RWL0_junc x466/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1546 VDD x467/junc0 x467/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1547 x468/junc1 WWL_3 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1548 x1/RWL1_junc RWL_17 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1549 x118/RWL0_junc x118/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1550 x469/junc1 WWL_11 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1551 WBL_30 WWL_24 x401/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1552 WBL_31 WWL_20 x141/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1553 x470/junc0 x470/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1554 RBL0_25 RWL_4 x471/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1555 WBL_0 WWL_28 x288/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1556 WBL_10 WWL_5 x472/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1557 WBL_14 WWL_1 x408/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1558 x268/RWL1_junc RWL_15 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1559 x473/junc0 x473/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1560 x474/junc0 x474/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1561 x475/RWL1_junc RWL_28 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1562 x396/junc0 x396/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1563 x476/junc0 x476/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1564 GND x477/junc0 x477/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1565 VDD x478/junc0 x478/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1566 x479/RWL0_junc x479/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1567 GND x480/junc1 x480/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1568 x481/junc1 WWL_27 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1569 VDD x119/junc0 x119/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1570 x482/junc0 x482/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1571 x45/junc0 x45/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1572 GND x483/junc0 x483/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1573 x484/junc1 WWL_12 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1574 RBL0_6 RWL_28 x485/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1575 WBL_19 WWL_9 x315/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1576 GND x120/junc1 x120/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1577 GND x486/junc0 x486/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1578 GND x487/junc0 x487/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1579 RBL0_16 RWL_1 x38/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1580 x488/junc1 WWL_8 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1581 x489/RWL0_junc x489/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1582 GND x490/junc1 x490/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1583 x491/junc1 WWL_29 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1584 GND x492/junc0 x492/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1585 GND x130/junc1 x130/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1586 x350/RWL1_junc RWL_8 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1587 GND x131/junc1 x131/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1588 GND x493/junc0 x493/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1589 x202/RWL1_junc RWL_12 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1590 WBL_16 WWL_23 x430/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1591 RBL0_15 RWL_13 x264/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1592 x494/junc0 x494/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1593 RBL0_0 RWL_6 x495/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1594 WBL_1 WWL_16 x431/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1595 x126/junc1 WWL_14 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1596 x496/RWL0_junc x496/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1597 x497/RWL1_junc RWL_24 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1598 GND x498/junc0 x498/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1599 VDD x499/junc0 x499/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1600 x500/junc0 x500/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1601 x277/junc0 x277/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1602 VDD x501/junc0 x501/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1603 x502/RWL1_junc RWL_13 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1604 x132/junc1 WWL_4 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1605 x51/RWL1_junc RWL_18 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1606 RBL0_25 RWL_5 x503/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1607 VDD x504/junc0 x504/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1608 x505/junc0 x505/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1609 RBL0_28 RWL_17 x66/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1610 RBL0_20 RWL_21 x283/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1611 x506/RWL0_junc x506/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1612 x507/junc0 x507/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1613 VDD x160/junc0 x160/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1614 x346/RWL1_junc RWL_30 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1615 x508/junc0 x508/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1616 x217/RWL1_junc RWL_16 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1617 GND x509/junc0 x509/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1618 x491/RWL1_junc RWL_29 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1619 RBL0_3 RWL_2 x75/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1620 WBL_4 WWL_12 x449/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1621 x308/RWL0_junc x308/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1622 VDD x510/junc0 x510/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1623 x511/RWL0_junc x511/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1624 GND x512/junc0 x512/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1625 x513/junc0 x513/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1626 x514/junc1 WWL_5 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1627 x515/junc0 x515/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1628 RBL0_2 RWL_30 x516/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1629 WBL_28 WWL_2 x355/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1630 GND x517/junc1 x517/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1631 GND x518/junc1 x518/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1632 x519/junc1 WWL_13 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1633 RBL0_6 RWL_29 x145/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1634 GND x167/junc1 x167/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1635 GND x516/junc1 x516/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1636 x520/RWL0_junc x520/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1637 GND x521/junc0 x521/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1638 VDD x354/junc0 x354/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1639 x522/junc0 x522/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1640 x523/junc0 x523/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1641 WBL_27 WWL_14 x524/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1642 VDD x525/junc0 x525/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1643 GND x175/junc1 x175/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1644 GND x177/junc1 x177/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1645 x455/RWL0_junc x455/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1646 x526/junc0 x526/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1647 WBL_16 WWL_24 x463/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1648 x47/junc0 x47/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1649 x527/junc0 x527/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1650 x528/RWL0_junc x528/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1651 GND x529/junc0 x529/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1652 GND x530/junc0 x530/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1653 x531/RWL1_junc RWL_25 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1654 GND x532/junc0 x532/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1655 VDD x192/junc0 x192/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1656 x207/RWL0_junc x207/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1657 x533/junc1 WWL_9 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1658 VDD x193/junc0 x193/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1659 RBL0_5 RWL_24 x534/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1660 VDD x535/junc0 x535/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1661 x536/junc0 x536/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1662 x110/RWL1_junc RWL_19 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1663 x537/junc0 x537/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1664 x538/junc1 WWL_17 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1665 x539/RWL0_junc x539/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1666 x540/junc0 x540/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1667 VDD x541/junc0 x541/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1668 RBL0_28 RWL_18 x119/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1669 RBL0_29 RWL_14 x319/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1670 RBL0_20 RWL_22 x322/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1671 x542/junc0 x542/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1672 x543/RWL0_junc x543/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1673 WBL_9 WWL_28 x372/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1674 GND x544/junc0 x544/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1675 WBL_13 WWL_5 x545/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1676 x546/RWL1_junc RWL_21 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1677 x547/RWL0_junc x547/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1678 RBL0_3 RWL_3 x129/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1679 WBL_4 WWL_13 x396/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1680 x350/RWL0_junc x350/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1681 x548/junc0 x548/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1682 VDD x549/junc0 x549/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1683 x78/junc0 x78/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1684 GND x550/junc0 x550/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1685 GND x551/junc0 x551/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1686 WBL_12 WWL_17 x482/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1687 GND x552/junc1 x552/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1688 x553/RWL1_junc RWL_31 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1689 GND x213/junc1 x213/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1690 GND x554/junc1 x554/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1691 x555/RWL0_junc x555/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1692 VDD x556/junc0 x556/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1693 x557/RWL0_junc x557/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1694 GND x558/junc0 x558/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1695 x559/junc0 x559/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1696 x560/junc0 x560/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1697 x22/junc1 WWL_12 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1698 x342/junc0 x342/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1699 VDD x224/junc0 x224/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1700 x101/junc0 x101/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1701 x561/junc0 x561/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1702 GND x562/junc0 x562/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1703 x563/junc0 x563/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1704 WBL_17 WWL_25 x564/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1705 x565/junc1 WWL_28 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1706 GND x566/junc0 x566/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1707 x567/RWL1_junc RWL_2 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1708 x33/RWL1_junc RWL_6 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1709 x568/RWL1_junc RWL_26 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1710 GND x569/junc0 x569/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1711 x256/RWL0_junc x256/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1712 WBL_21 WWL_21 x277/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1713 RBL0_14 RWL_17 x570/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1714 x571/junc0 x571/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1715 VDD x235/junc0 x235/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1716 VDD x239/junc0 x239/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1717 RBL0_5 RWL_25 x572/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1718 x573/junc0 x573/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1719 x41/RWL1_junc RWL_24 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1720 x574/junc1 WWL_18 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1721 x575/junc1 WWL_14 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1722 x576/RWL0_junc x576/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1723 x577/junc0 x577/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1724 VDD x249/junc0 x249/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1725 RBL0_29 RWL_15 x363/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1726 RBL0_20 RWL_23 x364/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1727 RBL0_28 RWL_19 x166/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1728 RBL0_8 RWL_0 x578/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1729 WBL_5 WWL_30 x416/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1730 x310/RWL1_junc RWL_22 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1731 x579/RWL0_junc x579/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1732 x580/junc0 x580/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1733 x394/junc0 x394/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1734 x581/junc0 x581/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1735 GND x255/junc1 x255/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1736 x582/junc0 x582/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1737 WBL_8 WWL_22 x450/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1738 GND x583/junc0 x583/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1739 GND x584/junc0 x584/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1740 WBL_12 WWL_18 x513/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1741 RBL0_6 RWL_2 x187/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1742 GND x585/junc1 x585/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1743 x586/RWL0_junc x586/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1744 GND x587/junc1 x587/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1745 x588/RWL0_junc x588/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1746 VDD x589/junc0 x589/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1747 x590/junc0 x590/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1748 x591/junc0 x591/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1749 x43/RWL1_junc RWL_17 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1750 x74/junc1 WWL_3 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1751 RBL0_17 RWL_4 x193/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1752 x239/junc1 WWL_5 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1753 GND x592/junc0 x592/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1754 VDD x274/junc0 x274/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1755 x593/junc0 x593/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1756 x594/junc1 WWL_13 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1757 GND x595/junc0 x595/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1758 x596/RWL1_junc RWL_7 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1759 x24/junc1 WWL_30 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1760 x597/junc0 x597/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1761 x400/junc0 x400/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1762 WBL_17 WWL_26 x527/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1763 WBL_25 WWL_22 x47/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1764 x335/RWL1_junc x61/RWL1 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1765 x598/junc1 WWL_10 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1766 x599/junc1 WWL_21 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1767 GND x276/junc1 x276/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1768 x600/junc1 WWL_17 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1769 GND x601/junc0 x601/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1770 RBL0_14 RWL_18 x602/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1771 x603/junc0 x603/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1772 x604/junc0 x604/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1773 RBL0_5 RWL_26 x605/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1774 x606/junc0 x606/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1775 GND x334/junc0 x334/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1776 VDD x289/junc0 x289/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1777 x156/RWL0_junc x156/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1778 x607/junc0 x607/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1779 GND x608/junc1 x608/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1780 x227/RWL0_junc x227/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1781 x96/RWL1_junc RWL_25 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1782 x609/RWL0_junc x609/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1783 x610/RWL0_junc x610/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1784 RBL0_29 RWL_16 x407/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1785 WBL_5 WWL_31 x456/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1786 RBL0_8 RWL_1 x611/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1787 x481/RWL1_junc RWL_27 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1788 x612/junc1 WWL_25 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1789 x613/RWL1_junc RWL_31 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1790 x351/RWL1_junc RWL_23 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1791 x614/junc0 x614/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1792 x211/RWL0_junc x211/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1793 x615/junc0 x615/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1794 x114/junc1 WWL_6 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1795 WBL_18 WWL_3 x78/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1796 x616/junc0 x616/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1797 WBL_8 WWL_23 x476/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1798 GND x296/junc1 x296/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1799 RBL0_2 RWL_7 x224/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1800 x319/RWL0_junc x319/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1801 RBL0_6 RWL_3 x226/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1802 x617/RWL0_junc x617/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1803 VDD x618/junc0 x618/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1804 GND x619/junc0 x619/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1805 x620/RWL1_junc RWL_10 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1806 x621/junc0 x621/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1807 x100/RWL1_junc RWL_18 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1808 x622/junc1 WWL_4 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1809 VDD x623/junc0 x623/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1810 RBL0_17 RWL_5 x239/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1811 GND x301/junc1 x301/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1812 x233/RWL1_junc RWL_6 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1813 GND x624/junc0 x624/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1814 WBL_2 WWL_29 x467/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1815 x625/RWL1_junc RWL_0 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1816 x132/RWL1_junc RWL_4 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1817 x135/junc1 WWL_22 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1818 x626/RWL1_junc RWL_8 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1819 WBL_26 WWL_19 x561/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1820 x613/junc1 WWL_31 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1821 WBL_17 WWL_27 x563/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1822 WBL_25 WWL_23 x101/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1823 VDD x318/junc0 x318/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1824 x11/junc0 x11/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1825 x21/junc1 WWL_11 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1826 x18/junc1 WWL_18 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1827 RBL0_14 RWL_19 x627/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1828 x628/junc0 x628/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1829 WBL_9 WWL_0 x573/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1830 GND x629/junc0 x629/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1831 VDD x326/junc0 x326/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1832 x200/RWL0_junc x200/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1833 GND x630/junc1 x630/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1834 x278/RWL0_junc x278/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1835 x146/RWL1_junc RWL_26 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1836 x631/RWL0_junc x631/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1837 WBL_20 WWL_2 x98/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1838 x632/junc1 WWL_28 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1839 x633/junc0 x633/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1840 GND x634/junc1 x634/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1841 GND x329/junc1 x329/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1842 x254/junc1 WWL_22 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1843 x570/RWL0_junc x570/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1844 x635/junc1 WWL_26 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1845 VDD x333/junc0 x333/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1846 RBL0_19 RWL_27 x636/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1847 GND x330/junc1 x330/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1848 x567/junc0 x567/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1849 x637/junc0 x637/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1850 RBL0_11 RWL_0 x271/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1851 x638/junc1 WWL_7 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1852 WBL_8 WWL_24 x639/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1853 WBL_18 WWL_4 x582/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1854 RBL0_2 RWL_8 x274/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1855 x401/junc0 x401/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1856 x363/RWL0_junc x363/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1857 VDD x231/junc0 x231/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1858 x640/junc0 x640/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1859 x641/junc0 x641/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1860 GND x555/junc0 x555/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1861 x642/junc0 x642/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1862 GND x643/junc0 x643/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1863 GND x36/junc0 x36/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1864 x644/junc0 x644/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1865 x645/RWL1_junc RWL_11 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1866 x28/junc0 x28/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1867 WBL_11 WWL_22 x590/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1868 x152/RWL1_junc RWL_19 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1869 VDD x646/junc0 x646/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1870 GND x647/junc1 x647/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1871 x648/RWL0_junc x648/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1872 x649/junc0 x649/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1873 x650/RWL1_junc RWL_1 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1874 x186/junc1 WWL_3 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1875 x181/RWL1_junc RWL_5 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1876 x185/junc1 WWL_23 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1877 VDD x359/junc0 x359/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1878 WBL_25 WWL_24 x597/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1879 WBL_26 WWL_20 x400/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1880 WBL_29 WWL_29 x504/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1881 WBL_5 WWL_5 x153/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1882 WBL_9 WWL_1 x606/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1883 GND x651/junc0 x651/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1884 GND x652/junc1 x652/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1885 x653/junc1 WWL_30 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1886 x654/RWL0_junc x654/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1887 VDD x655/junc0 x655/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1888 GND x656/junc1 x656/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1889 x657/RWL0_junc x657/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1890 x658/RWL0_junc x658/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1891 x602/RWL0_junc x602/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1892 x92/junc1 WWL_27 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1893 x295/junc1 WWL_23 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1894 VDD x374/junc0 x374/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1895 x659/junc0 x659/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1896 GND x373/junc1 x373/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1897 GND x76/junc0 x76/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1898 GND x660/junc0 x660/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1899 x370/junc1 WWL_0 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1900 RBL0_11 RWL_1 x309/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1901 x661/junc1 WWL_8 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1902 x210/RWL1_junc RWL_27 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1903 x662/junc0 x662/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1904 x94/junc0 x94/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1905 x407/RWL0_junc x407/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1906 VDD x663/junc0 x663/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1907 x492/junc0 x492/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1908 GND x664/junc0 x664/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1909 x665/junc0 x665/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1910 x328/junc0 x328/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1911 x666/junc1 WWL_2 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1912 GND x667/junc0 x667/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1913 GND x384/junc1 x384/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1914 GND x386/junc1 x386/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1915 x668/RWL1_junc RWL_4 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1916 x669/junc0 x669/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1917 x449/RWL1_junc RWL_12 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1918 WBL_11 WWL_23 x621/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1919 RBL0_10 RWL_13 x490/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1920 GND x670/junc1 x670/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1921 GND x671/junc0 x671/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1922 x672/RWL0_junc x672/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1923 x673/RWL1_junc RWL_24 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1924 VDD x674/junc0 x674/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1925 x390/junc1 WWL_4 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1926 x497/junc1 WWL_24 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1927 VDD x405/junc0 x405/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1928 x575/RWL1_junc RWL_14 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1929 x13/junc0 x13/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1930 x15/junc0 x15/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1931 RBL0_23 RWL_17 x333/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1932 x675/junc0 x675/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1933 VDD x411/junc0 x411/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1934 x17/junc0 x17/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1935 x676/junc1 WWL_31 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1936 GND x410/junc1 x410/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1937 VDD x677/junc0 x677/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1938 x678/RWL0_junc x678/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1939 x565/RWL1_junc RWL_28 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1940 x463/junc0 x463/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1941 x679/junc0 x679/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1942 x627/RWL0_junc x627/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1943 x29/junc0 x29/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1944 x680/RWL0_junc x680/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1945 GND x211/junc0 x211/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1946 x334/junc1 WWL_24 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1947 x512/junc0 x512/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1948 GND x31/junc0 x31/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1949 x681/junc0 x681/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1950 x682/junc0 x682/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1951 x253/junc1 WWL_5 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1952 GND x417/junc1 x417/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1953 x683/junc0 x683/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1954 WBL_23 WWL_2 x567/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1955 GND x684/junc0 x684/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1956 GND x685/junc1 x685/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1957 GND x686/junc1 x686/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1958 x414/junc1 WWL_1 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1959 x687/junc0 x687/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1960 x688/junc0 x688/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1961 x521/junc0 x521/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1962 GND x44/junc0 x44/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1963 RBL0_12 RWL_28 x689/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1964 WBL_31 WWL_6 x640/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1965 WBL_30 WWL_10 x641/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1966 RBL0_15 RWL_10 x517/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1967 x46/junc0 x46/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1968 WBL_22 WWL_14 x642/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1969 GND x426/junc1 x426/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1970 VDD x250/junc0 x250/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1971 x545/RWL1_junc RWL_5 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1972 x690/junc0 x690/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1973 x636/RWL0_junc x636/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1974 GND x689/junc1 x689/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1975 x115/junc1 WWL_29 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1976 WBL_11 WWL_24 x28/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1977 x322/junc0 x322/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1978 x691/RWL0_junc x691/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1979 x600/RWL1_junc RWL_17 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1980 x598/RWL1_junc RWL_10 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1981 GND x53/junc0 x53/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1982 GND x56/junc0 x56/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1983 x692/RWL1_junc RWL_25 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1984 VDD x440/junc0 x440/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1985 x453/RWL0_junc x453/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1986 x693/junc1 WWL_9 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1987 VDD x439/junc0 x439/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1988 x694/junc0 x694/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1989 x67/junc0 x67/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1990 x695/RWL1_junc RWL_15 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1991 x696/junc1 WWL_17 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1992 x70/junc0 x70/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1993 x697/junc0 x697/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1994 VDD x698/junc0 x698/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M1995 RBL0_23 RWL_18 x374/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1996 RBL0_24 RWL_14 x699/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1997 GND x448/junc1 x448/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1998 x700/RWL1_junc RWL_21 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M1999 x701/RWL0_junc x701/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2000 VDD x4/junc0 x4/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2001 x24/RWL1_junc RWL_30 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2002 VDD x12/junc0 x12/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2003 x25/RWL1_junc RWL_29 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2004 x85/junc0 x85/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2005 x702/junc0 x702/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2006 x703/RWL0_junc x703/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2007 GND x87/junc0 x87/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2008 x704/RWL1_junc RWL_30 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2009 x86/junc0 x86/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2010 x551/junc0 x551/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2011 GND x88/junc0 x88/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2012 x550/junc0 x550/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2013 WBL_7 WWL_17 x659/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2014 GND x705/junc1 x705/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2015 GND x706/junc1 x706/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2016 VDD x707/junc0 x707/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2017 x708/junc0 x708/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2018 RBL0_8 RWL_30 x709/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2019 GND x387/junc0 x387/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2020 RBL0_12 RWL_29 x446/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2021 WBL_31 WWL_7 x492/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2022 WBL_30 WWL_11 x665/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2023 RBL0_15 RWL_11 x552/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2024 RBL0_0 RWL_4 x710/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2025 x103/junc0 x103/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2026 x300/junc1 WWL_12 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2027 WBL_11 WWL_30 x174/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2028 x711/RWL0_junc x711/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2029 x105/junc0 x105/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2030 GND x446/junc1 x446/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2031 x712/junc0 x712/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2032 x364/junc0 x364/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2033 x21/RWL1_junc RWL_11 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2034 GND x713/junc0 x713/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2035 x18/RWL1_junc RWL_18 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2036 GND x111/junc0 x111/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2037 x714/junc1 WWL_2 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2038 x20/RWL1_junc RWL_2 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2039 x715/RWL1_junc RWL_26 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2040 RBL0_9 RWL_17 x716/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2041 x480/RWL0_junc x480/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2042 x113/junc0 x113/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2043 VDD x470/junc0 x470/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2044 x717/junc0 x717/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2045 GND x117/junc0 x117/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2046 x34/RWL1_junc RWL_24 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2047 x37/RWL1_junc RWL_16 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2048 x124/junc0 x124/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2049 VDD x48/junc0 x48/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2050 x718/junc1 WWL_18 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2051 x219/junc1 WWL_14 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2052 x719/junc0 x719/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2053 VDD x474/junc0 x474/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2054 RBL0_23 RWL_19 x418/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2055 RBL0_24 RWL_15 x720/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2056 RBL0_3 RWL_0 x422/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2057 x47/RWL1_junc RWL_22 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2058 x721/RWL0_junc x721/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2059 WBL_15 WWL_28 x203/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2060 x383/junc0 x383/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2061 VDD x54/junc0 x54/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2062 GND x382/junc1 x382/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2063 x722/junc0 x722/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2064 x723/junc0 x723/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2065 GND x479/junc1 x479/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2066 GND x139/junc0 x139/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2067 WBL_21 WWL_28 x0/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2068 WBL_3 WWL_22 x679/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2069 x724/junc0 x724/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2070 GND x725/junc0 x725/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2071 WBL_1 WWL_3 x681/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2072 x584/junc0 x584/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2073 WBL_16 WWL_10 x512/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2074 WBL_7 WWL_18 x682/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2075 x317/RWL0_junc x317/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2076 GND x726/junc1 x726/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2077 x727/RWL0_junc x727/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2078 GND x728/junc1 x728/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2079 VDD x729/junc0 x729/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2080 x730/junc0 x730/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2081 WBL_27 WWL_12 x637/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2082 WBL_31 WWL_8 x521/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2083 RBL0_0 RWL_5 x731/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2084 RBL0_15 RWL_12 x585/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2085 x732/junc1 WWL_13 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2086 WBL_11 WWL_31 x72/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2087 x733/junc0 x733/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2088 x734/junc0 x734/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2089 x595/junc0 x595/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2090 VDD x735/junc0 x735/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2091 x79/RWL1_junc RWL_12 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2092 x77/RWL1_junc RWL_19 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2093 x259/junc1 WWL_17 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2094 x78/RWL1_junc x61/RWL1 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2095 x161/junc0 x161/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2096 x42/junc1 WWL_21 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2097 GND x736/junc0 x736/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2098 RBL0_9 RWL_18 x737/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2099 x162/junc0 x162/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2100 x738/junc0 x738/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2101 GND x549/junc0 x549/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2102 GND x164/junc0 x164/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2103 GND x739/junc0 x739/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2104 x357/junc1 WWL_15 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2105 VDD x505/junc0 x505/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2106 GND x740/junc1 x740/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2107 RBL0_20 RWL_20 x276/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2108 GND x741/junc1 x741/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2109 x90/RWL1_junc RWL_25 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2110 x742/RWL0_junc x742/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2111 x169/junc0 x169/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2112 VDD x508/junc0 x508/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2113 RBL0_24 RWL_16 x743/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2114 x337/junc1 WWL_0 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2115 RBL0_3 RWL_1 x459/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2116 x92/RWL1_junc RWL_27 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2117 x101/RWL1_junc RWL_23 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2118 WBL_17 WWL_30 x231/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2119 WBL_12 WWL_15 x340/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2120 WBL_3 WWL_23 x702/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2121 GND x511/junc1 x511/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2122 x699/RWL0_junc x699/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2123 WBL_1 WWL_4 x550/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2124 WBL_16 WWL_11 x551/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2125 x27/junc0 x27/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2126 x744/RWL0_junc x744/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2127 VDD x745/junc0 x745/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2128 GND x191/junc0 x191/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2129 VDD x522/junc0 x522/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2130 x746/junc0 x746/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2131 GND x747/junc1 x747/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2132 WBL_27 WWL_13 x336/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2133 x441/junc0 x441/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2134 x118/RWL1_junc RWL_6 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2135 x125/RWL1_junc RWL_0 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2136 x390/RWL1_junc RWL_4 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2137 x393/junc1 WWL_22 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2138 RBL0_20 RWL_9 x301/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2139 WBL_21 WWL_19 x712/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2140 x206/junc0 x206/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2141 x299/junc1 WWL_18 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2142 RBL0_9 RWL_19 x32/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2143 x748/junc0 x748/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2144 WBL_4 WWL_0 x717/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2145 GND x209/junc0 x209/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2146 x749/junc1 WWL_12 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2147 x404/junc1 WWL_16 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2148 VDD x540/junc0 x540/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2149 GND x385/junc1 x385/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2150 GND x750/junc1 x750/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2151 GND x515/junc1 x515/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2152 x140/RWL1_junc RWL_26 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2153 x751/RWL0_junc x751/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2154 x752/junc1 WWL_28 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2155 x379/junc1 WWL_1 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2156 GND x753/junc1 x753/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2157 GND x543/junc1 x543/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2158 x144/RWL1_junc RWL_20 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2159 x754/RWL0_junc x754/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2160 x716/RWL0_junc x716/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2161 VDD x158/junc0 x158/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2162 VDD x548/junc0 x548/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2163 x399/RWL0_junc x399/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2164 GND x547/junc1 x547/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2165 x20/junc0 x20/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2166 x755/junc0 x755/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2167 WBL_17 WWL_31 x663/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2168 WBL_12 WWL_16 x383/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2169 RBL0_6 RWL_0 x494/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2170 WBL_3 WWL_24 x723/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2171 x597/junc0 x597/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2172 x720/RWL0_junc x720/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2173 x756/junc0 x756/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2174 x757/junc0 x757/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2175 x81/junc0 x81/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2176 x758/junc0 x758/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2177 GND x759/junc0 x759/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2178 GND x270/junc0 x270/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2179 GND x238/junc0 x238/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2180 x760/RWL1_junc RWL_13 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2181 GND x241/junc0 x241/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2182 VDD x559/junc0 x559/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2183 x303/junc0 x303/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2184 GND x761/junc1 x761/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2185 WBL_6 WWL_22 x730/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2186 x762/RWL0_junc x762/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2187 x763/junc1 WWL_15 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2188 x172/RWL1_junc RWL_1 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2189 RBL0_29 RWL_2 x647/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2190 x433/RWL1_junc RWL_5 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2191 x437/junc1 WWL_19 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2192 RBL0_28 RWL_6 x507/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2193 x436/junc1 WWL_23 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2194 WBL_21 WWL_20 x595/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2195 VDD x571/junc0 x571/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2196 WBL_8 WWL_29 x764/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2197 x183/RWL1_junc RWL_9 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2198 WBL_4 WWL_1 x738/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2199 GND x765/junc0 x765/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2200 x766/junc0 x766/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2201 x767/junc1 WWL_13 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2202 VDD x768/junc0 x768/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2203 GND x769/junc1 x769/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2204 x402/junc1 WWL_30 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2205 x770/RWL0_junc x770/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2206 GND x618/junc0 x618/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2207 GND x771/junc1 x771/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2208 x772/RWL0_junc x772/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2209 VDD x580/junc0 x580/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2210 x773/RWL0_junc x773/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2211 x737/RWL0_junc x737/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2212 VDD x774/junc0 x774/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2213 VDD x581/junc0 x581/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2214 x775/junc0 x775/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2215 x776/junc0 x776/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2216 GND x579/junc1 x579/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2217 GND x338/junc0 x338/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2218 GND x555/junc1 x555/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2219 x578/junc1 WWL_0 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2220 RBL0_6 RWL_1 x526/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2221 x455/RWL1_junc RWL_27 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2222 x279/junc0 x279/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2223 x280/junc0 x280/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2224 x743/RWL0_junc x743/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2225 x664/junc0 x664/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2226 GND x281/junc0 x281/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2227 x777/junc0 x777/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2228 x778/junc0 x778/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2229 WBL_0 WWL_22 x27/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2230 x779/junc0 x779/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2231 x16/junc1 WWL_2 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2232 RBL0_1 RWL_17 x29/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2233 GND x780/junc0 x780/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2234 GND x588/junc1 x588/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2235 GND x781/junc0 x781/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2236 x782/junc0 x782/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2237 x207/RWL1_junc RWL_4 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2238 WBL_6 WWL_23 x746/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2239 RBL0_5 RWL_13 x519/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2240 GND x288/junc0 x288/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2241 GND x783/junc1 x783/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2242 x2/RWL0_junc x2/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2243 x784/RWL1_junc RWL_24 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2244 VDD x785/junc0 x785/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2245 RBL0_29 x389/RWL1 x670/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2246 x786/junc1 WWL_9 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2247 x190/junc1 WWL_20 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2248 x787/junc1 WWL_16 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2249 x673/junc1 WWL_24 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2250 GND x788/junc1 x788/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2251 VDD x603/junc0 x603/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2252 x219/RWL1_junc RWL_14 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2253 VDD x789/junc0 x789/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2254 x790/junc0 x790/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2255 RBL0_18 RWL_17 x548/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2256 x791/junc0 x791/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2257 VDD x792/junc0 x792/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2258 WBL_8 WWL_10 x793/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2259 VDD x244/junc0 x244/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2260 GND x794/junc1 x794/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2261 GND x609/junc1 x609/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2262 x387/junc1 WWL_31 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2263 GND x91/junc0 x91/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2264 VDD x614/junc0 x614/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2265 VDD x537/junc0 x537/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2266 x28/junc0 x28/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2267 x32/RWL0_junc x32/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2268 x795/RWL0_junc x795/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2269 GND x305/junc0 x305/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2270 x31/junc0 x31/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2271 x796/junc0 x796/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2272 WBL_18 WWL_2 x20/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2273 x477/junc1 WWL_5 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2274 x611/junc1 WWL_1 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2275 x797/junc0 x797/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2276 x40/junc0 x40/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2277 GND x316/junc0 x316/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2278 x798/junc0 x798/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2279 WBL_26 WWL_6 x756/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2280 x44/junc0 x44/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2281 GND x320/junc0 x320/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2282 x321/junc0 x321/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2283 WBL_25 WWL_10 x757/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2284 RBL0_10 RWL_10 x685/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2285 WBL_0 WWL_23 x81/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2286 GND x799/junc1 x799/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2287 RBL0_1 RWL_18 x86/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2288 WBL_17 WWL_14 x758/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2289 GND x617/junc1 x617/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2290 GND x671/junc1 x671/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2291 x256/RWL1_junc RWL_5 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2292 RBL0_14 RWL_6 x170/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2293 x800/junc0 x800/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2294 WBL_6 WWL_24 x303/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2295 GND x801/junc0 x801/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2296 x55/RWL0_junc x55/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2297 x259/RWL1_junc RWL_17 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2298 x802/RWL1_junc RWL_25 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2299 VDD x9/junc0 x9/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2300 VDD x11/junc0 x11/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2301 x264/RWL1_junc RWL_13 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2302 GND x803/junc1 x803/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2303 x267/RWL1_junc RWL_15 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2304 x804/junc1 WWL_17 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2305 RBL0_18 RWL_18 x581/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2306 RBL0_19 RWL_14 x805/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2307 RBL0_14 RWL_30 x188/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2308 x324/junc0 x324/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2309 WBL_8 WWL_11 x806/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2310 GND x807/junc1 x807/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2311 x647/RWL0_junc x647/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2312 GND x631/junc1 x631/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2313 GND x211/junc1 x211/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2314 x283/RWL1_junc RWL_21 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2315 VDD x35/junc0 x35/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2316 GND x142/junc0 x142/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2317 VDD x555/junc0 x555/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2318 x82/junc0 x82/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2319 x808/RWL0_junc x808/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2320 GND x347/junc0 x347/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2321 x88/junc0 x88/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2322 GND x348/junc0 x348/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2323 x495/RWL1_junc RWL_6 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2324 WBL_2 WWL_17 x775/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2325 x353/junc0 x353/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2326 x183/junc0 x183/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2327 x809/RWL1_junc RWL_28 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2328 x810/junc0 x810/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2329 x93/junc0 x93/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2330 GND x360/junc0 x360/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2331 x491/junc0 x491/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2332 x362/junc0 x362/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2333 x49/junc1 WWL_10 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2334 WBL_26 WWL_7 x664/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2335 WBL_25 WWL_11 x777/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2336 RBL0_10 RWL_11 x705/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2337 WBL_0 WWL_24 x778/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2338 GND x811/junc1 x811/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2339 x365/junc0 x365/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2340 RBL0_1 RWL_19 x724/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2341 x812/RWL0_junc x812/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2342 x813/junc0 x813/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2343 GND x814/junc1 x814/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2344 GND x815/junc0 x815/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2345 GND x368/junc0 x368/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2346 RBL0_24 RWL_28 x816/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2347 x299/RWL1_junc RWL_18 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2348 x133/junc1 WWL_2 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2349 x817/RWL1_junc RWL_26 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2350 RBL0_4 RWL_17 x818/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2351 GND x819/junc1 x819/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2352 VDD x63/junc0 x63/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2353 GND x820/junc1 x820/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2354 VDD x302/junc0 x302/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2355 x821/RWL0_junc x821/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2356 x822/junc1 WWL_29 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2357 GND x823/junc1 x823/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2358 GND x372/junc0 x372/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2359 x289/junc1 WWL_10 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2360 x534/RWL1_junc RWL_24 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2361 x307/RWL1_junc RWL_16 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2362 x80/junc1 WWL_14 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2363 x376/junc0 x376/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2364 VDD x323/junc0 x323/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2365 x824/junc1 WWL_18 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2366 RBL0_18 RWL_19 x615/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2367 RBL0_19 RWL_15 x229/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2368 x382/junc0 x382/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2369 x385/junc0 x385/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2370 x319/RWL1_junc RWL_14 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2371 x670/RWL0_junc x670/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2372 x322/RWL1_junc RWL_22 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2373 x587/junc0 x587/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2374 GND x658/junc1 x658/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2375 x137/junc0 x137/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2376 GND x397/junc0 x397/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2377 GND x398/junc0 x398/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2378 x506/junc1 WWL_30 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2379 GND x825/junc0 x825/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2380 WBL_11 WWL_10 x31/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2381 WBL_2 WWL_18 x796/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2382 x533/RWL0_junc x533/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2383 GND x387/junc1 x387/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2384 VDD x662/junc0 x662/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2385 x141/junc0 x141/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2386 VDD x102/junc0 x102/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2387 x822/RWL1_junc RWL_29 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2388 WBL_22 WWL_12 x797/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2389 x106/junc1 WWL_11 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2390 x408/junc0 x408/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2391 WBL_26 WWL_8 x44/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2392 RBL0_10 RWL_12 x726/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2393 RBL0_20 RWL_30 x562/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2394 RBL0_13 RWL_24 x489/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2395 GND x826/junc1 x826/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2396 RBL0_24 RWL_29 x234/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2397 x339/RWL1_junc RWL_19 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2398 x120/junc1 WWL_17 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2399 x413/junc0 x413/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2400 x604/RWL1_junc RWL_31 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2401 x163/RWL0_junc x163/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2402 RBL0_4 RWL_18 x827/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2403 GND x416/junc0 x416/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2404 GND x12/junc0 x12/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2405 VDD x15/junc0 x15/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2406 GND x828/junc0 x828/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2407 x566/junc1 WWL_15 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2408 GND x109/junc1 x109/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2409 x646/RWL0_junc x646/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2410 x170/RWL0_junc x170/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2411 x326/junc1 WWL_11 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2412 GND x58/junc1 x58/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2413 x572/RWL1_junc RWL_25 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2414 x420/junc0 x420/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2415 VDD x17/junc0 x17/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2416 RBL0_19 RWL_16 x282/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2417 x176/junc0 x176/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2418 x363/RWL1_junc RWL_15 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2419 x364/RWL1_junc RWL_23 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2420 x829/junc0 x829/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2421 x182/junc0 x182/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2422 x180/junc0 x180/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2423 GND x678/junc1 x678/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2424 WBL_7 WWL_15 x554/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2425 GND x242/junc0 x242/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2426 x607/junc1 WWL_31 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2427 x805/RWL0_junc x805/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2428 WBL_11 WWL_11 x88/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2429 GND x42/junc0 x42/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2430 WBL_27 WWL_28 x265/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2431 x830/junc0 x830/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2432 WBL_31 WWL_5 x831/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2433 VDD x46/junc0 x46/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2434 WBL_30 WWL_9 x183/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2435 GND x84/junc1 x84/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2436 GND x832/junc1 x832/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2437 WBL_22 WWL_13 x810/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2438 x833/RWL0_junc x833/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2439 x377/RWL1_junc RWL_2 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2440 x378/RWL1_junc RWL_0 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2441 x43/junc1 WWL_17 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2442 RBL0_13 RWL_25 x520/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2443 x592/junc1 WWL_22 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2444 WBL_29 WWL_21 x813/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2445 GND x834/junc1 x834/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2446 x452/junc0 x452/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2447 x167/junc1 WWL_18 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2448 x208/RWL0_junc x208/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2449 RBL0_4 RWL_19 x306/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2450 GND x66/junc0 x66/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2451 GND x68/junc0 x68/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2452 VDD x69/junc0 x69/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2453 x835/junc1 WWL_12 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2454 VDD x649/junc0 x649/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2455 x723/junc0 x723/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2456 GND x836/junc1 x836/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2457 x601/junc1 WWL_16 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2458 VDD x70/junc0 x70/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2459 x344/RWL0_junc x344/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2460 x214/junc0 x214/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2461 GND x837/junc1 x837/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2462 GND x683/junc1 x683/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2463 x605/RWL1_junc RWL_26 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2464 GND x838/junc1 x838/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2465 x243/RWL0_junc x243/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2466 RBL0_31 RWL_21 x94/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2467 x403/RWL1_junc RWL_20 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2468 GND x593/junc1 x593/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2469 x818/RWL0_junc x818/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2470 x407/RWL1_junc RWL_16 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2471 GND x701/junc1 x701/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2472 WBL_7 WWL_16 x587/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2473 x839/RWL0_junc x839/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2474 x734/junc0 x734/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2475 x229/RWL0_junc x229/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2476 x228/junc0 x228/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2477 x840/junc0 x840/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2478 GND x98/junc0 x98/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2479 GND x97/junc0 x97/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2480 x5/RWL1_junc RWL_13 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2481 VDD x103/junc0 x103/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2482 GND x841/junc1 x841/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2483 x842/RWL1_junc RWL_31 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2484 x246/RWL0_junc x246/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2485 x14/RWL1_junc x389/RWL1 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2486 VDD x112/junc0 x112/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2487 x843/junc1 WWL_15 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2488 x423/RWL1_junc RWL_1 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2489 RBL0_24 RWL_2 x666/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2490 RBL0_13 RWL_26 x557/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2491 x674/junc1 WWL_19 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2492 x100/junc1 WWL_18 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2493 VDD x113/junc0 x113/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2494 RBL0_23 RWL_6 x675/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2495 x624/junc1 WWL_23 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2496 x652/junc0 x652/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2497 GND x119/junc0 x119/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2498 x26/RWL1_junc RWL_9 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2499 x844/junc0 x844/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2500 GND x123/junc0 x123/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2501 RBL0_16 RWL_24 x463/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2502 x482/junc0 x482/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2503 VDD x124/junc0 x124/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2504 VDD x3/junc0 x3/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2505 x45/junc0 x45/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2506 x845/junc1 WWL_13 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2507 x656/junc0 x656/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2508 GND x846/junc1 x846/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2509 x261/junc0 x261/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2510 GND x847/junc1 x847/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2511 x260/junc0 x260/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2512 x258/junc0 x258/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2513 WBL_30 WWL_30 x537/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2514 GND x745/junc0 x745/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2515 GND x848/junc1 x848/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2516 x849/RWL0_junc x849/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2517 x287/RWL0_junc x287/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2518 x171/RWL0_junc x171/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2519 VDD x850/junc0 x850/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2520 VDD x13/junc0 x13/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2521 GND x71/junc1 x71/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2522 RBL0_31 RWL_22 x687/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2523 x827/RWL0_junc x827/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2524 x156/junc1 WWL_28 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2525 GND x721/junc1 x721/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2526 WBL_1 WWL_2 x180/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2527 WBL_16 WWL_9 x182/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2528 x422/junc1 WWL_0 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2529 x851/RWL0_junc x851/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2530 x500/junc0 x500/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2531 x277/junc0 x277/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2532 x282/RWL0_junc x282/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2533 x49/RWL1_junc RWL_10 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2534 x281/junc0 x281/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2535 x852/junc0 x852/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2536 x57/RWL1_junc RWL_6 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2537 GND x727/junc1 x727/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2538 GND x151/junc0 x151/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2539 GND x147/junc0 x147/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2540 x19/junc0 x19/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2541 x453/RWL1_junc RWL_4 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2542 GND x853/junc1 x853/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2543 RBL0_20 RWL_7 x588/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2544 x291/RWL0_junc x291/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2545 GND x160/junc0 x160/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2546 RBL0_24 x389/RWL1 x389/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2547 VDD x161/junc0 x161/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2548 x439/junc1 WWL_20 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2549 x39/junc1 WWL_16 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2550 x784/junc1 WWL_24 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2551 VDD x162/junc0 x162/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2552 x854/junc0 x854/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2553 x80/RWL1_junc RWL_14 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2554 WBL_28 WWL_25 x630/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2555 VDD x165/junc0 x165/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2556 GND x166/junc0 x166/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2557 RBL0_16 RWL_25 x85/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2558 x513/junc0 x513/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2559 VDD x169/junc0 x169/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2560 x99/junc0 x99/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2561 GND x855/junc1 x855/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2562 x856/junc0 x856/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2563 WBL_3 WWL_10 x214/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2564 GND x857/junc1 x857/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2565 GND x742/junc1 x742/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2566 VDD x858/junc0 x858/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2567 x632/junc0 x632/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2568 RBL0_27 RWL_27 x194/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2569 WBL_30 WWL_31 x555/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2570 GND x354/junc0 x354/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2571 x859/RWL0_junc x859/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2572 VDD x67/junc0 x67/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2573 x303/junc0 x303/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2574 x860/RWL0_junc x860/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2575 VDD x861/junc0 x861/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2576 RBL0_31 RWL_23 x708/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2577 x306/RWL0_junc x306/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2578 WBL_27 WWL_0 x218/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2579 x305/junc0 x305/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2580 x459/junc1 WWL_1 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2581 x862/junc0 x862/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2582 x863/junc0 x863/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2583 x314/junc0 x314/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2584 GND x192/junc0 x192/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2585 GND x193/junc0 x193/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2586 x106/RWL1_junc RWL_11 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2587 WBL_21 WWL_6 x228/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2588 x320/junc0 x320/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2589 x864/RWL0_junc x864/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2590 RBL0_5 RWL_10 x865/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2591 GND x866/junc1 x866/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2592 x480/RWL1_junc RWL_5 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2593 RBL0_9 RWL_6 x421/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2594 x867/junc0 x867/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2595 x667/junc1 WWL_3 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2596 x120/RWL1_junc RWL_17 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2597 RBL0_29 RWL_0 x799/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2598 RBL0_28 RWL_4 x124/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2599 RBL0_20 RWL_8 x617/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2600 VDD x202/junc0 x202/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2601 GND x204/junc0 x204/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2602 x490/RWL1_junc RWL_13 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2603 VDD x206/junc0 x206/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2604 x506/RWL1_junc RWL_30 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2605 x130/RWL1_junc RWL_7 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2606 VDD x105/junc0 x105/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2607 WBL_28 WWL_26 x652/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2608 x131/RWL1_junc RWL_15 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2609 x25/junc0 x25/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2610 RBL0_16 RWL_26 x722/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2611 x868/junc0 x868/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2612 WBL_12 WWL_3 x656/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2613 x869/junc0 x869/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2614 WBL_3 WWL_11 x261/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2615 GND x7/junc1 x7/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2616 x666/RWL0_junc x666/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2617 x778/junc0 x778/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2618 GND x751/junc1 x751/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2619 VDD x870/junc0 x870/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2620 x341/junc0 x341/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2621 VDD x217/junc0 x217/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2622 x871/junc0 x871/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2623 GND x311/junc0 x311/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2624 x345/RWL0_junc x345/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2625 VDD x122/junc0 x122/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2626 GND x221/junc0 x221/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2627 x342/junc0 x342/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2628 x872/RWL0_junc x872/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2629 GND x224/junc0 x224/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2630 WBL_27 WWL_1 x269/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2631 x348/junc0 x348/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2632 GND x873/junc1 x873/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2633 x563/junc0 x563/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2634 x26/junc0 x26/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2635 x874/junc0 x874/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2636 x358/junc0 x358/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2637 GND x235/junc0 x235/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2638 GND x239/junc0 x239/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2639 x684/junc1 WWL_6 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2640 x159/RWL1_junc RWL_12 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2641 x573/junc0 x573/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2642 x325/junc1 WWL_10 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2643 x875/RWL0_junc x875/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2644 WBL_21 WWL_7 x281/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2645 RBL0_5 RWL_11 x876/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2646 x877/RWL0_junc x877/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2647 RBL0_30 RWL_31 x555/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2648 x878/junc0 x878/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2649 x517/RWL1_junc RWL_10 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2650 GND x879/junc1 x879/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2651 GND x248/junc0 x248/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2652 x330/junc1 WWL_0 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2653 GND x249/junc0 x249/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2654 x167/RWL1_junc RWL_18 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2655 RBL0_29 RWL_1 x811/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2656 x236/junc1 WWL_4 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2657 RBL0_28 RWL_5 x169/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2658 x880/RWL0_junc x880/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2659 GND x881/junc1 x881/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2660 VDD x138/junc0 x138/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2661 GND x882/junc1 x882/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2662 x883/junc1 WWL_29 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2663 GND x252/junc0 x252/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2664 x175/RWL1_junc RWL_8 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2665 VDD x884/junc0 x884/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2666 WBL_28 WWL_27 x854/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2667 x177/RWL1_junc RWL_16 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2668 VDD x885/junc0 x885/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2669 x582/junc0 x582/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2670 VDD x110/junc0 x110/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2671 WBL_12 WWL_4 x856/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2672 x699/RWL1_junc RWL_14 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2673 x389/RWL0_junc x389/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2674 VDD x266/junc0 x266/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2675 x591/junc0 x591/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2676 x392/junc0 x392/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2677 x886/junc0 x886/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2678 x728/junc0 x728/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2679 GND x272/junc0 x272/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2680 x395/junc0 x395/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2681 GND x274/junc0 x274/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2682 WBL_6 WWL_10 x305/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2683 x593/junc0 x593/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2684 x693/RWL0_junc x693/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2685 RBL0_30 RWL_27 x887/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2686 VDD x279/junc0 x279/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2687 x400/junc0 x400/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2688 VDD x284/junc0 x284/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2689 WBL_17 WWL_12 x862/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2690 x61/junc1 WWL_3 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2691 x523/junc1 WWL_7 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2692 RBL0_14 RWL_4 x888/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2693 x366/junc1 WWL_11 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2694 x606/junc0 x606/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2695 WBL_21 WWL_8 x320/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2696 RBL0_5 RWL_12 x484/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2697 GND x289/junc0 x289/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2698 GND x889/junc1 x889/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2699 x115/junc0 x115/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2700 RBL0_8 RWL_24 x639/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2701 x552/RWL1_junc RWL_11 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2702 GND x890/junc1 x890/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2703 x373/junc1 WWL_1 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2704 x213/RWL1_junc RWL_19 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2705 GND x95/junc1 x95/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2706 x415/RWL0_junc x415/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2707 WBL_0 WWL_30 x649/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2708 x111/junc1 WWL_15 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2709 x891/RWL0_junc x891/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2710 x421/RWL0_junc x421/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2711 VDD x465/junc0 x465/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2712 x616/junc0 x616/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2713 VDD x892/junc0 x892/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2714 WBL_8 WWL_9 x694/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2715 x199/RWL1_junc RWL_30 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2716 x799/RWL0_junc x799/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2717 x427/junc0 x427/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2718 x720/RWL1_junc RWL_15 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2719 x893/junc0 x893/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2720 x201/junc0 x201/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2721 x434/junc0 x434/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2722 WBL_0 WWL_10 x871/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2723 WBL_15 WWL_17 x341/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2724 x710/RWL1_junc RWL_4 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2725 WBL_2 WWL_15 x706/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2726 RBL0_6 RWL_30 x346/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2727 x425/RWL0_junc x425/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2728 VDD x310/junc0 x310/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2729 x71/junc0 x71/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2730 WBL_6 WWL_11 x348/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2731 RBL0_26 RWL_31 x211/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2732 GND x318/junc0 x318/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2733 x894/junc0 x894/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2734 WBL_26 WWL_5 x895/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2735 VDD x321/junc0 x321/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2736 WBL_25 WWL_9 x26/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2737 GND x896/junc1 x896/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2738 WBL_17 WWL_13 x874/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2739 x410/junc1 WWL_4 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2740 RBL0_14 RWL_5 x514/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2741 x560/junc1 WWL_8 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2742 GND x134/junc1 x134/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2743 x897/junc0 x897/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2744 WBL_20 WWL_25 x500/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2745 GND x326/junc0 x326/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2746 x255/RWL1_junc RWL_2 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2747 WBL_24 WWL_21 x878/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2748 GND x898/junc1 x898/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2749 RBL0_8 RWL_25 x899/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2750 GND x900/junc1 x900/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2751 x585/RWL1_junc RWL_12 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2752 x227/RWL1_junc RWL_28 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2753 x454/RWL0_junc x454/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2754 WBL_0 WWL_31 x3/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2755 GND x333/junc0 x333/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2756 x901/junc0 x901/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2757 VDD x335/junc0 x335/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2758 x240/junc1 WWL_12 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2759 GND x154/junc1 x154/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2760 x736/junc1 WWL_16 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2761 GND x336/junc0 x336/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2762 x902/RWL0_junc x902/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2763 WBL_13 WWL_28 x13/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2764 GND x231/junc0 x231/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2765 x811/RWL0_junc x811/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2766 x641/junc0 x641/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2767 x278/junc1 WWL_29 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2768 RBL0_26 RWL_21 x280/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2769 x276/RWL1_junc RWL_20 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2770 x642/junc0 x642/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2771 x460/junc0 x460/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2772 x743/RWL1_junc RWL_16 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2773 WBL_15 WWL_18 x392/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2774 x731/RWL1_junc RWL_5 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2775 WBL_0 WWL_11 x886/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2776 x608/RWL1_junc RWL_24 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2777 RBL0_1 RWL_6 x258/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2778 WBL_2 WWL_16 x728/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2779 x903/RWL0_junc x903/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2780 VDD x351/junc0 x351/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2781 x761/junc0 x761/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2782 GND x359/junc0 x359/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2783 GND x361/junc0 x361/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2784 VDD x362/junc0 x362/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2785 x483/junc1 WWL_9 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2786 x292/RWL1_junc RWL_13 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2787 VDD x365/junc0 x365/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2788 GND x904/junc1 x904/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2789 GND x905/junc1 x905/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2790 x906/junc0 x906/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2791 WBL_20 WWL_26 x863/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2792 GND x367/junc0 x367/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2793 RBL0_4 RWL_31 x387/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2794 x296/RWL1_junc x389/RWL1 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2795 VDD x233/junc0 x233/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2796 x275/junc1 WWL_15 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2797 RBL0_19 RWL_2 x16/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2798 GND x907/junc1 x907/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2799 RBL0_8 RWL_26 x908/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2800 RBL0_18 RWL_6 x791/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2801 x278/RWL1_junc RWL_29 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2802 x769/junc0 x769/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2803 GND x821/junc1 x821/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2804 GND x374/junc0 x374/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2805 x909/RWL0_junc x909/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2806 x888/RWL0_junc x888/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2807 x301/RWL1_junc RWL_9 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2808 x789/junc1 WWL_9 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2809 RBL0_11 RWL_24 x28/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2810 x659/junc0 x659/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2811 VDD x376/junc0 x376/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2812 x910/junc1 WWL_13 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2813 x771/junc0 x771/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2814 GND x6/junc1 x6/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2815 x486/junc0 x486/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2816 x663/RWL1_junc RWL_31 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2817 x209/junc1 WWL_25 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2818 WBL_9 WWL_30 x67/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2819 x492/junc0 x492/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2820 x466/junc1 WWL_21 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2821 x665/junc0 x665/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2822 VDD x146/junc0 x146/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2823 x328/junc0 x328/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2824 RBL0_26 RWL_22 x40/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2825 x493/junc0 x493/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2826 RBL0_22 RWL_31 x654/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2827 WBL_11 WWL_9 x434/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2828 x630/RWL1_junc RWL_25 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2829 x911/RWL0_junc x911/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2830 VDD x401/junc0 x401/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2831 x325/RWL1_junc RWL_10 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2832 x783/junc0 x783/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2833 GND x405/junc0 x405/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2834 x329/RWL1_junc RWL_6 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2835 GND x406/junc0 x406/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2836 VDD x408/junc0 x408/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2837 GND x912/junc1 x912/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2838 GND x913/junc1 x913/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2839 x330/RWL1_junc RWL_0 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2840 WBL_29 WWL_19 x897/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2841 x238/junc1 WWL_15 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2842 WBL_20 WWL_27 x444/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2843 GND x411/junc0 x411/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2844 x744/junc1 WWL_30 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2845 VDD x413/junc0 x413/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2846 x312/junc1 WWL_16 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2847 RBL0_19 x61/RWL1 x74/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2848 WBL_19 WWL_28 x105/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2849 x914/junc0 x914/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2850 GND x163/junc1 x163/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2851 WBL_23 WWL_25 x750/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2852 x647/RWL1_junc RWL_2 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2853 VDD x315/junc0 x315/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2854 x915/RWL0_junc x915/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2855 x512/junc0 x512/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2856 GND x418/junc0 x418/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2857 x514/RWL0_junc x514/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2858 RBL0_11 RWL_25 x82/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2859 x682/junc0 x682/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2860 VDD x420/junc0 x420/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2861 x916/junc0 x916/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2862 GND x247/junc1 x247/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2863 GND x60/junc1 x60/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2864 x765/junc1 WWL_26 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2865 VDD x917/junc0 x917/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2866 WBL_9 WWL_31 x122/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2867 RBL0_22 RWL_27 x353/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2868 x521/junc0 x521/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2869 x918/junc0 x918/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2870 VDD x381/junc0 x381/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2871 RBL0_26 RWL_23 x93/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2872 x369/junc0 x369/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2873 WBL_22 WWL_0 x460/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2874 x652/RWL1_junc RWL_26 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2875 GND x440/junc0 x440/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2876 x754/junc1 WWL_28 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2877 GND x439/junc0 x439/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2878 x366/RWL1_junc RWL_11 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2879 x919/junc0 x919/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2880 WBL_14 WWL_22 x761/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2881 GND x920/junc1 x920/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2882 GND x89/junc1 x89/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2883 x836/RWL0_junc x836/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2884 GND x442/junc0 x442/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2885 x676/junc0 x676/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2886 RBL0_4 RWL_6 x114/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2887 GND x921/junc1 x921/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2888 x767/RWL0_junc x767/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2889 x922/RWL0_junc x922/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2890 x923/RWL0_junc x923/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2891 x924/junc0 x924/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2892 x373/RWL1_junc RWL_1 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2893 WBL_6 WWL_29 x145/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2894 x780/junc1 WWL_3 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2895 x781/junc1 WWL_16 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2896 RBL0_24 RWL_0 x121/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2897 VDD x449/junc0 x449/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2898 GND x833/junc1 x833/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2899 WBL_29 WWL_20 x906/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2900 RBL0_23 RWL_4 x376/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2901 GND x450/junc0 x450/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2902 x553/junc1 WWL_31 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2903 x519/RWL1_junc RWL_13 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2904 VDD x452/junc0 x452/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2905 x384/RWL1_junc RWL_7 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2906 VDD x355/junc0 x355/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2907 GND x208/junc1 x208/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2908 WBL_23 WWL_26 x769/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2909 x188/RWL0_junc x188/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2910 x670/RWL1_junc x389/RWL1 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2911 x925/junc0 x925/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2912 x551/junc0 x551/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2913 x562/RWL0_junc x562/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2914 x550/junc0 x550/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2915 x926/junc0 x926/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2916 RBL0_11 RWL_26 x137/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2917 WBL_7 WWL_3 x771/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2918 x927/junc0 x927/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2919 GND x116/junc1 x116/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2920 x16/RWL0_junc x16/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2921 x455/junc1 WWL_27 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2922 VDD x928/junc0 x928/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2923 RBL0_31 RWL_20 x141/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2924 x929/junc0 x929/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2925 GND x464/junc0 x464/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2926 WBL_22 WWL_1 x493/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2927 GND x930/junc1 x930/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2928 x91/junc1 WWL_25 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2929 x301/junc0 x301/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2930 x786/RWL0_junc x786/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2931 x410/RWL1_junc RWL_4 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2932 GND x470/junc0 x470/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2933 x102/junc1 WWL_6 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2934 x412/RWL1_junc RWL_12 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2935 RBL0_13 RWL_13 x399/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2936 x717/junc0 x717/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2937 x539/junc1 WWL_10 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2938 WBL_14 WWL_23 x783/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2939 x846/RWL0_junc x846/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2940 x931/junc0 x931/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2941 x816/RWL0_junc x816/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2942 x932/junc0 x932/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2943 x685/RWL1_junc RWL_10 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2944 GND x474/junc0 x474/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2945 GND x473/junc0 x473/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2946 x547/junc1 WWL_0 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2947 RBL0_24 RWL_1 x168/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2948 x471/junc1 WWL_4 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2949 RBL0_23 RWL_5 x420/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2950 x933/RWL0_junc x933/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2951 GND x246/junc1 x246/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2952 GND x934/junc1 x934/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2953 VDD x396/junc0 x396/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2954 GND x150/junc1 x150/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2955 GND x476/junc0 x476/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2956 x426/RWL1_junc RWL_8 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2957 RBL0_31 RWL_9 x176/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2958 VDD x935/junc0 x935/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2959 VDD x482/junc0 x482/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2960 WBL_23 WWL_27 x914/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2961 x634/junc0 x634/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2962 x583/junc0 x583/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2963 x584/junc0 x584/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2964 x936/junc1 WWL_30 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2965 WBL_7 WWL_4 x916/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2966 x74/RWL0_junc x74/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2967 VDD x937/junc0 x937/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2968 x938/junc0 x938/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2969 GND x171/junc1 x171/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2970 x83/RWL0_junc x83/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2971 x142/junc1 WWL_26 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2972 RBL0_25 RWL_27 x197/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2973 VDD x500/junc0 x500/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2974 x595/junc0 x595/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2975 x448/RWL1_junc RWL_5 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2976 x424/junc1 WWL_3 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2977 x46/junc1 WWL_7 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2978 x738/junc0 x738/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2979 RBL0_9 RWL_4 x205/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2980 x576/junc1 WWL_11 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2981 WBL_14 WWL_24 x919/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2982 x855/RWL0_junc x855/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2983 GND x505/junc0 x505/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2984 x939/junc0 x939/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M2985 GND x507/junc0 x507/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2986 GND x189/junc1 x189/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2987 x234/RWL0_junc x234/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2988 RBL0_3 RWL_24 x723/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2989 x705/RWL1_junc RWL_11 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2990 GND x508/junc0 x508/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2991 x579/junc1 WWL_1 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2992 GND x356/junc1 x356/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2993 x538/RWL0_junc x538/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2994 x732/junc0 x732/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2995 x251/RWL0_junc x251/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2996 GND x291/junc1 x291/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2997 x612/RWL0_junc x612/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2998 RBL0_27 RWL_14 x524/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M2999 VDD x446/junc0 x446/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3000 x940/RWL0_junc x940/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3001 x114/RWL0_junc x114/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3002 VDD x513/junc0 x513/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3003 WBL_3 WWL_9 x925/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3004 x121/RWL0_junc x121/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3005 x443/junc1 WWL_31 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3006 VDD x37/junc0 x37/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3007 x619/junc0 x619/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3008 GND x522/junc0 x522/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3009 x447/junc0 x447/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3010 GND x215/junc1 x215/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3011 x623/junc0 x623/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3012 WBL_10 WWL_17 x929/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3013 GND x860/junc1 x860/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3014 x764/junc0 x764/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3015 VDD x527/junc0 x527/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3016 VDD x47/junc0 x47/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3017 x135/RWL0_junc x135/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3018 x194/junc1 WWL_27 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3019 x941/junc0 x941/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3020 x942/junc0 x942/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3021 WBL_21 WWL_5 x943/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3022 GND x536/junc0 x536/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3023 RBL0_16 RWL_28 x565/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3024 x609/junc1 WWL_4 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3025 RBL0_9 RWL_5 x253/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3026 x103/junc1 WWL_8 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3027 x834/junc0 x834/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3028 GND x540/junc0 x540/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3029 x479/RWL1_junc RWL_2 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3030 x944/junc0 x944/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3031 x643/junc1 WWL_2 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3032 WBL_19 WWL_21 x931/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3033 RBL0_12 RWL_17 x482/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3034 GND x237/junc1 x237/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3035 RBL0_3 RWL_25 x45/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3036 x30/junc0 x30/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3037 x726/RWL1_junc RWL_12 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3038 RBL0_16 RWL_13 x260/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3039 x574/RWL0_junc x574/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3040 x635/RWL0_junc x635/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3041 GND x548/junc0 x548/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3042 VDD x77/junc0 x77/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3043 VDD x78/junc0 x78/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3044 VDD x79/junc0 x79/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3045 RBL0_27 RWL_15 x52/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3046 x755/junc0 x755/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3047 GND x810/junc0 x810/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3048 x23/RWL0_junc x23/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3049 WBL_12 WWL_2 x634/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3050 x168/RWL0_junc x168/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3051 x757/junc0 x757/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3052 RBL0_21 RWL_21 x277/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3053 x758/junc0 x758/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3054 x703/junc0 x703/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3055 x945/junc0 x945/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3056 x417/junc0 x417/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3057 GND x559/junc0 x559/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3058 x744/RWL1_junc RWL_30 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3059 WBL_10 WWL_18 x938/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3060 GND x262/junc1 x262/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3061 x740/RWL1_junc RWL_24 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3062 x882/RWL0_junc x882/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3063 GND x872/junc1 x872/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3064 x178/RWL0_junc x178/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3065 VDD x563/junc0 x563/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3066 VDD x101/junc0 x101/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3067 x841/junc0 x841/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3068 x185/RWL0_junc x185/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3069 GND x571/junc0 x571/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3070 x242/junc1 WWL_5 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3071 x946/junc0 x946/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3072 VDD x573/junc0 x573/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3073 x76/junc1 WWL_9 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3074 RBL0_12 RWL_30 x24/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3075 RBL0_16 RWL_29 x25/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3076 GND x273/junc1 x273/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3077 x324/RWL0_junc x324/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3078 x947/junc0 x947/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3079 x766/junc0 x766/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3080 GND x24/junc1 x24/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3081 GND x577/junc0 x577/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3082 x511/RWL1_junc x61/RWL1 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3083 x570/junc1 WWL_17 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3084 WBL_28 WWL_14 x939/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3085 VDD x118/junc0 x118/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3086 GND x768/junc0 x768/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3087 RBL0_12 RWL_18 x513/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3088 GND x948/junc1 x948/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3089 RBL0_3 RWL_26 x99/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3090 x847/junc0 x847/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3091 x949/RWL0_junc x949/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3092 GND x580/junc0 x580/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3093 GND x880/junc1 x880/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3094 GND x774/junc0 x774/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3095 x747/RWL1_junc RWL_21 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3096 GND x581/junc0 x581/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3097 x73/RWL0_junc x73/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3098 x205/RWL0_junc x205/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3099 x754/RWL1_junc RWL_28 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3100 RBL0_6 RWL_24 x303/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3101 VDD x950/junc0 x950/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3102 x775/junc0 x775/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3103 RBL0_27 RWL_16 x108/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3104 VDD x502/junc0 x502/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3105 VDD x582/junc0 x582/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3106 x848/junc0 x848/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3107 x660/junc0 x660/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3108 x68/junc1 WWL_25 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3109 x664/junc0 x664/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3110 VDD x591/junc0 x591/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3111 x648/junc1 WWL_21 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3112 RBL0_30 RWL_14 x313/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3113 x777/junc0 x777/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3114 RBL0_21 RWL_22 x314/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3115 x779/junc0 x779/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3116 RBL0_22 RWL_28 x59/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3117 WBL_15 WWL_15 x680/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3118 x951/junc0 x951/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3119 VDD x515/junc0 x515/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3120 WBL_6 WWL_9 x623/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3121 x750/RWL1_junc RWL_25 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3122 x222/RWL0_junc x222/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3123 VDD x597/junc0 x597/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3124 x539/RWL1_junc RWL_10 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3125 x853/junc0 x853/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3126 GND x603/junc0 x603/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3127 x128/junc1 WWL_2 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3128 x543/RWL1_junc RWL_6 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3129 WBL_13 WWL_17 x941/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3130 VDD x606/junc0 x606/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3131 GND x308/junc1 x308/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3132 GND x952/junc1 x952/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3133 x547/RWL1_junc RWL_0 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3134 x790/junc0 x790/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3135 WBL_24 WWL_19 x834/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3136 x230/junc0 x230/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3137 GND x792/junc0 x792/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3138 x602/junc1 WWL_18 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3139 VDD x953/junc0 x953/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3140 RBL0_12 RWL_19 x868/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3141 x855/junc0 x855/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3142 x65/junc0 x65/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3143 GND x614/junc0 x614/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3144 GND x537/junc0 x537/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3145 GND x415/junc1 x415/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3146 WBL_18 WWL_25 x837/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3147 x666/RWL1_junc RWL_2 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3148 x761/RWL1_junc RWL_22 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3149 x127/RWL0_junc x127/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3150 x31/junc0 x31/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3151 GND x615/junc0 x615/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3152 x535/junc0 x535/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3153 x253/RWL0_junc x253/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3154 x773/RWL1_junc RWL_29 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3155 RBL0_6 RWL_25 x342/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3156 x796/junc0 x796/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3157 VDD x616/junc0 x616/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3158 GND x632/junc1 x632/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3159 x954/junc0 x954/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3160 x123/junc1 WWL_26 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3161 VDD x955/junc0 x955/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3162 RBL0_17 RWL_27 x563/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3163 x44/junc0 x44/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3164 x155/junc0 x155/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3165 x157/junc0 x157/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3166 RBL0_30 RWL_15 x357/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3167 RBL0_21 RWL_23 x358/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3168 RBL0_22 RWL_29 x115/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3169 WBL_15 WWL_16 x703/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3170 WBL_17 WWL_0 x945/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3171 RBL0_1 RWL_4 x550/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3172 WBL_0 WWL_9 x417/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3173 WBL_15 WWL_30 x382/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3174 WBL_21 WWL_30 x385/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3175 x956/junc0 x956/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3176 x769/RWL1_junc RWL_26 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3177 GND x11/junc0 x11/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3178 x576/RWL1_junc RWL_11 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3179 x957/junc0 x957/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3180 WBL_9 WWL_22 x841/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3181 GND x958/junc1 x958/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3182 GND x349/junc1 x349/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3183 x154/RWL0_junc x154/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3184 GND x628/junc0 x628/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3185 WBL_13 WWL_18 x946/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3186 GND x350/junc1 x350/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3187 GND x959/junc1 x959/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3188 x845/RWL0_junc x845/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3189 x960/RWL0_junc x960/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3190 x579/RWL1_junc RWL_1 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3191 x147/junc1 WWL_3 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3192 GND x497/junc1 x497/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3193 RBL0_19 RWL_0 x375/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3194 RBL0_18 RWL_4 x582/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3195 WBL_24 WWL_20 x947/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3196 GND x679/junc0 x679/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3197 VDD x961/junc0 x961/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3198 x588/RWL1_junc RWL_7 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3199 x962/junc0 x962/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3200 VDD x567/junc0 x567/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3201 GND x454/junc1 x454/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3202 WBL_18 WWL_26 x847/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3203 x389/RWL1_junc x389/RWL1 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3204 GND x637/junc0 x637/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3205 x783/RWL1_junc RWL_23 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3206 x498/junc1 WWL_17 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3207 x88/junc0 x88/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3208 GND x653/junc1 x653/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3209 RBL0_6 RWL_26 x395/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3210 x195/junc0 x195/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3211 GND x504/junc1 x504/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3212 GND x401/junc0 x401/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3213 WBL_2 WWL_3 x848/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3214 x963/junc0 x963/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3215 VDD x641/junc0 x641/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3216 x166/junc1 WWL_19 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3217 x636/junc1 WWL_27 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3218 GND x334/junc1 x334/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3219 VDD x964/junc0 x964/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3220 x117/RWL0_junc x117/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3221 RBL0_26 RWL_20 x400/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3222 x965/junc0 x965/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3223 GND x644/junc0 x644/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3224 RBL0_30 RWL_16 x404/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3225 WBL_17 WWL_1 x951/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3226 GND x966/junc1 x966/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3227 WBL_15 WWL_31 x425/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3228 RBL0_1 RWL_5 x584/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3229 x194/RWL1_junc RWL_27 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3230 x354/junc1 WWL_25 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3231 x813/junc0 x813/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3232 WBL_21 WWL_31 x428/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3233 x967/junc0 x967/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3234 x609/RWL1_junc RWL_4 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3235 x610/RWL1_junc RWL_12 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3236 WBL_9 WWL_23 x853/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3237 RBL0_8 RWL_13 x594/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3238 x968/RWL0_junc x968/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3239 x6/RWL0_junc x6/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3240 x53/RWL0_junc x53/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3241 x865/RWL1_junc RWL_10 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3242 x701/junc1 WWL_0 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3243 x371/junc1 WWL_4 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3244 GND x531/junc1 x531/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3245 RBL0_19 RWL_1 x419/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3246 RBL0_18 RWL_5 x616/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3247 GND x702/junc0 x702/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3248 WBL_12 WWL_29 x446/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3249 x799/RWL1_junc RWL_0 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3250 x617/RWL1_junc RWL_8 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3251 x204/junc1 WWL_22 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3252 x133/junc0 x133/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3253 RBL0_26 RWL_9 x427/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3254 VDD x969/junc0 x969/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3255 VDD x659/junc0 x659/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3256 WBL_18 WWL_27 x65/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3257 x753/junc0 x753/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3258 x265/junc0 x265/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3259 x532/junc1 WWL_18 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3260 x725/junc0 x725/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3261 x709/junc1 WWL_30 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3262 GND x662/junc0 x662/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3263 WBL_2 WWL_4 x954/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3264 VDD x665/junc0 x665/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3265 x919/junc0 x919/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3266 x711/junc1 WWL_20 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3267 x164/RWL0_junc x164/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3268 GND x629/junc1 x629/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3269 x179/junc0 x179/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3270 x739/RWL0_junc x739/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3271 x970/junc0 x970/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3272 GND x669/junc0 x669/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3273 GND x8/junc1 x8/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3274 x254/junc0 x254/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3275 x343/RWL0_junc x343/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3276 x311/junc1 WWL_26 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3277 x971/junc0 x971/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3278 WBL_29 WWL_6 x956/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3279 RBL0_13 RWL_10 x849/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3280 WBL_20 WWL_14 x56/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3281 GND x432/junc1 x432/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3282 x631/RWL1_junc RWL_5 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3283 x226/junc1 WWL_3 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3284 RBL0_4 RWL_4 x451/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3285 x972/RWL0_junc x972/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3286 WBL_9 WWL_24 x957/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3287 x247/RWL0_junc x247/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3288 GND x15/junc0 x15/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3289 x198/junc0 x198/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3290 x713/RWL0_junc x713/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3291 GND x675/junc0 x675/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3292 GND x438/junc1 x438/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3293 VDD x973/junc0 x973/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3294 GND x17/junc0 x17/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3295 x876/RWL1_junc RWL_11 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3296 x721/junc1 WWL_1 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3297 GND x33/junc1 x33/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3298 GND x568/junc1 x568/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3299 x696/RWL0_junc x696/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3300 x864/junc1 WWL_28 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3301 x776/RWL1_junc RWL_31 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3302 RBL0_22 RWL_14 x642/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3303 x811/RWL1_junc RWL_1 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3304 x252/junc1 WWL_23 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3305 VDD x657/junc0 x657/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3306 x186/junc0 x186/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3307 x297/junc0 x297/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3308 VDD x682/junc0 x682/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3309 x375/RWL0_junc x375/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3310 VDD x307/junc0 x307/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3311 x671/junc1 WWL_31 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3312 GND x688/junc0 x688/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3313 x820/RWL1_junc RWL_27 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3314 x819/RWL1_junc RWL_13 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3315 x830/junc0 x830/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3316 GND x46/junc0 x46/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3317 x220/junc0 x220/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3318 GND x651/junc1 x651/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3319 GND x690/junc0 x690/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3320 GND x458/junc1 x458/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3321 WBL_5 WWL_17 x965/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3322 VDD x322/junc0 x322/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3323 GND x62/junc1 x62/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3324 x974/RWL0_junc x974/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3325 x975/RWL0_junc x975/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3326 x295/junc0 x295/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3327 x393/RWL0_junc x393/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3328 x353/junc1 WWL_27 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3329 x232/junc0 x232/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3330 x272/junc1 WWL_3 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3331 WBL_29 WWL_7 x967/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3332 RBL0_13 RWL_11 x859/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3333 x932/RWL1_junc RWL_31 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3334 GND x976/junc1 x976/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3335 GND x694/junc0 x694/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3336 x742/junc1 WWL_4 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3337 RBL0_4 RWL_5 x477/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3338 x749/RWL0_junc x749/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3339 x900/junc0 x900/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3340 GND x649/junc0 x649/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3341 GND x70/junc0 x70/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3342 x759/junc1 WWL_2 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3343 x214/junc0 x214/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3344 x245/junc0 x245/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3345 GND x767/junc1 x767/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3346 GND x922/junc1 x922/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3347 RBL0_7 RWL_17 x659/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3348 GND x469/junc1 x469/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3349 GND x923/junc1 x923/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3350 x484/RWL1_junc RWL_12 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3351 x304/junc0 x304/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3352 RBL0_11 RWL_13 x486/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3353 x718/RWL0_junc x718/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3354 x158/junc0 x158/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3355 RBL0_31 RWL_7 x492/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3356 VDD x339/junc0 x339/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3357 x699/junc1 WWL_14 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3358 RBL0_22 RWL_15 x328/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3359 x489/junc1 WWL_24 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3360 VDD x680/junc0 x680/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3361 x251/junc0 x251/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3362 WBL_7 WWL_2 x753/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3363 x419/RWL0_junc x419/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3364 x840/junc0 x840/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3365 x808/junc0 x808/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3366 WBL_25 WWL_29 x515/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3367 x327/junc0 x327/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3368 GND x103/junc0 x103/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3369 WBL_14 WWL_10 x179/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3370 WBL_5 WWL_18 x970/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3371 GND x488/junc1 x488/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3372 x109/RWL1_junc RWL_24 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3373 x150/RWL0_junc x150/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3374 x428/junc0 x428/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3375 VDD x364/junc0 x364/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3376 x905/junc0 x905/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3377 x763/RWL0_junc x763/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3378 x977/RWL0_junc x977/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3379 x436/RWL0_junc x436/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3380 GND x113/junc0 x113/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3381 x710/junc1 WWL_4 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3382 x472/junc1 WWL_5 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3383 WBL_29 WWL_8 x971/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3384 x200/junc0 x200/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3385 x285/junc0 x285/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3386 VDD x717/junc0 x717/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3387 x338/junc1 WWL_9 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3388 GND x786/junc1 x786/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3389 RBL0_13 RWL_12 x345/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3390 GND x126/junc1 x126/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3391 x907/junc0 x907/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3392 x844/junc0 x844/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3393 x290/junc0 x290/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3394 GND x124/junc0 x124/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3395 GND x719/junc0 x719/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3396 x716/junc1 WWL_17 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3397 RBL0_16 RWL_10 x512/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3398 x122/RWL1_junc RWL_31 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3399 WBL_23 WWL_14 x198/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3400 GND x132/junc1 x132/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3401 x261/junc0 x261/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3402 RBL0_7 RWL_18 x682/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3403 GND x978/junc1 x978/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3404 GND x933/junc1 x933/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3405 x979/RWL0_junc x979/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3406 GND x850/junc0 x850/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3407 x288/RWL0_junc x288/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3408 GND x13/junc0 x13/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3409 x832/RWL1_junc RWL_21 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3410 x498/RWL1_junc RWL_17 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3411 x774/junc0 x774/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3412 WBL_1 WWL_25 x107/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3413 x337/RWL0_junc x337/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3414 x451/RWL0_junc x451/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3415 RBL0_31 RWL_8 x521/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3416 VDD x980/junc0 x980/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3417 VDD x383/junc0 x383/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3418 RBL0_22 RWL_16 x369/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3419 x281/junc0 x281/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3420 RBL0_0 RWL_27 x529/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3421 x762/junc1 WWL_21 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3422 RBL0_25 RWL_14 x530/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3423 x852/junc0 x852/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3424 RBL0_1 RWL_28 x212/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3425 WBL_10 WWL_15 x795/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3426 VDD x683/junc0 x683/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3427 WBL_14 WWL_11 x220/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3428 x287/junc1 WWL_29 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3429 x356/RWL0_junc x356/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3430 x837/RWL1_junc RWL_25 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3431 x461/RWL0_junc x461/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3432 VDD x734/junc0 x734/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3433 x787/RWL0_junc x787/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3434 x263/RWL1_junc RWL_30 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3435 x913/junc0 x913/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3436 GND x161/junc0 x161/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3437 GND x162/junc0 x162/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3438 x380/junc1 WWL_2 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3439 VDD x738/junc0 x738/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3440 GND x173/junc1 x173/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3441 x854/junc0 x854/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3442 x701/RWL1_junc RWL_0 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3443 x361/junc1 WWL_22 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3444 x819/junc0 x819/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3445 WBL_19 WWL_19 x900/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3446 GND x169/junc0 x169/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3447 x467/junc0 x467/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3448 RBL0_24 RWL_30 x981/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3449 x856/junc0 x856/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3450 RBL0_16 RWL_11 x551/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3451 x737/junc1 WWL_18 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3452 GND x181/junc1 x181/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3453 x300/junc0 x300/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3454 RBL0_7 RWL_19 x926/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3455 GND x858/junc0 x858/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3456 x632/junc0 x632/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3457 VDD x14/junc0 x14/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3458 GND x67/junc0 x67/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3459 GND x538/junc1 x538/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3460 GND x861/junc0 x861/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3461 GND x612/junc1 x612/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3462 x532/RWL1_junc RWL_18 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3463 x801/RWL0_junc x801/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3464 GND x697/junc0 x697/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3465 GND x136/junc0 x136/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3466 x841/RWL1_junc RWL_22 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3467 x379/RWL0_junc x379/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3468 x477/RWL0_junc x477/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3469 x305/junc0 x305/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3470 WBL_1 WWL_26 x158/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3471 GND x752/junc1 x752/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3472 GND x940/junc1 x940/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3473 VDD x27/junc0 x27/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3474 x483/RWL0_junc x483/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3475 x524/junc1 WWL_14 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3476 x320/junc0 x320/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3477 RBL0_25 RWL_15 x566/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3478 x409/junc0 x409/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3479 x663/junc0 x663/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3480 RBL0_1 RWL_29 x441/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3481 WBL_10 WWL_16 x808/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3482 x920/junc0 x920/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3483 x847/RWL1_junc RWL_26 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3484 VDD x71/junc0 x71/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3485 x921/junc0 x921/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3486 x982/junc0 x982/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3487 WBL_4 WWL_22 x905/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3488 GND x206/junc0 x206/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3489 WBL_31 WWL_28 x593/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3490 x498/RWL0_junc x498/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3491 GND x748/junc0 x748/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3492 GND x105/junc0 x105/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3493 GND x216/junc1 x216/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3494 x910/RWL0_junc x910/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3495 x983/RWL0_junc x983/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3496 VDD x57/junc0 x57/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3497 x721/RWL1_junc RWL_1 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3498 RBL0_27 RWL_2 x714/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3499 WBL_28 WWL_12 x907/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3500 x405/junc1 WWL_15 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3501 GND x673/junc1 x673/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3502 x406/junc1 WWL_23 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3503 WBL_19 WWL_20 x290/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3504 x869/junc0 x869/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3505 RBL0_16 RWL_12 x583/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3506 GND x870/junc0 x870/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3507 x504/junc0 x504/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3508 x341/junc0 x341/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3509 VDD x984/junc0 x984/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3510 x871/junc0 x871/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3511 VDD x20/junc0 x20/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3512 x344/junc0 x344/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3513 GND x574/junc1 x574/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3514 GND x797/junc0 x797/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3515 GND x635/junc1 x635/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3516 x569/RWL1_junc RWL_19 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3517 x853/RWL1_junc RWL_23 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3518 x348/junc0 x348/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3519 GND x402/junc1 x402/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3520 WBL_1 WWL_27 x774/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3521 GND x764/junc1 x764/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3522 GND x597/junc0 x597/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3523 GND x23/junc1 x23/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3524 x273/RWL0_junc x273/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3525 VDD x757/junc0 x757/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3526 VDD x81/junc0 x81/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3527 x418/junc1 WWL_19 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3528 RBL0_21 RWL_20 x595/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3529 VDD x758/junc0 x758/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3530 RBL0_25 RWL_16 x601/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3531 RBL0_29 RWL_24 x334/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3532 x353/RWL1_junc RWL_27 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3533 x878/junc0 x878/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3534 x985/junc0 x985/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3535 x742/RWL1_junc RWL_4 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3536 WBL_27 WWL_30 x84/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3537 WBL_13 WWL_15 x912/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3538 WBL_4 WWL_23 x913/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3539 RBL0_3 RWL_13 x732/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3540 x986/RWL0_junc x986/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3541 x532/RWL0_junc x532/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3542 x987/RWL0_junc x987/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3543 GND x733/junc0 x733/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3544 GND x884/junc0 x884/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3545 GND x885/junc0 x885/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3546 VDD x988/junc0 x988/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3547 RBL0_27 x389/RWL1 x468/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3548 VDD x989/junc0 x989/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3549 x442/junc1 WWL_16 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3550 GND x692/junc1 x692/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3551 x534/junc1 WWL_24 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3552 GND x599/junc1 x599/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3553 WBL_28 WWL_13 x819/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3554 GND x251/junc0 x251/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3555 GND x352/junc0 x352/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3556 x121/RWL1_junc RWL_0 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3557 x866/RWL1_junc RWL_20 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3558 x392/junc0 x392/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3559 x735/junc0 x735/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3560 VDD x831/junc0 x831/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3561 x886/junc0 x886/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3562 x450/junc1 WWL_22 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3563 VDD x775/junc0 x775/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3564 RBL0_21 RWL_9 x619/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3565 GND x949/junc1 x949/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3566 x397/junc0 x397/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3567 x485/junc0 x485/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3568 x838/junc0 x838/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3569 x825/junc0 x825/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3570 GND x279/junc0 x279/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3571 VDD x777/junc0 x777/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3572 x957/junc0 x957/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3573 VDD x778/junc0 x778/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3574 x812/junc1 WWL_20 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3575 x952/RWL0_junc x952/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3576 x416/RWL0_junc x416/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3577 GND x924/junc1 x924/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3578 VDD x779/junc0 x779/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3579 x429/junc0 x429/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3580 GND x782/junc0 x782/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3581 GND x293/junc1 x293/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3582 RBL0_29 RWL_25 x629/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3583 x478/junc0 x478/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3584 x558/RWL0_junc x558/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3585 x990/junc0 x990/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3586 WBL_24 WWL_6 x920/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3587 RBL0_8 RWL_10 x793/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3588 GND x622/junc1 x622/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3589 x751/RWL1_junc RWL_5 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3590 RBL0_12 RWL_6 x30/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3591 WBL_27 WWL_31 x136/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3592 WBL_13 WWL_16 x921/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3593 x991/RWL0_junc x991/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3594 WBL_4 WWL_24 x982/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3595 x569/RWL0_junc x569/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3596 x356/junc0 x356/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3597 x445/junc0 x445/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3598 x873/RWL1_junc RWL_9 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3599 GND x388/junc0 x388/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3600 GND x465/junc0 x465/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3601 GND x791/junc0 x791/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3602 GND x892/junc0 x892/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3603 VDD x992/junc0 x992/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3604 VDD x993/junc0 x993/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3605 GND x715/junc1 x715/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3606 GND x994/junc1 x994/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3607 x804/RWL0_junc x804/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3608 RBL0_17 RWL_14 x758/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3609 x168/RWL1_junc RWL_1 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3610 x779/junc1 WWL_15 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3611 RBL0_30 RWL_2 x643/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3612 x499/junc0 x499/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3613 x476/junc1 WWL_23 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3614 x437/junc0 x437/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3615 x501/junc0 x501/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3616 x516/junc0 x516/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3617 VDD x796/junc0 x796/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3618 WBL_15 WWL_3 x344/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3619 x242/junc0 x242/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3620 x879/RWL1_junc RWL_17 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3621 VDD x177/junc0 x177/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3622 GND x798/junc0 x798/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3623 x881/RWL1_junc RWL_13 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3624 x882/RWL1_junc RWL_27 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3625 x894/junc0 x894/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3626 x959/RWL0_junc x959/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3627 GND x321/junc0 x321/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3628 x462/junc0 x462/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3629 VDD x755/junc0 x755/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3630 x188/junc1 WWL_30 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3631 GND x800/junc0 x800/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3632 GND x638/junc1 x638/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3633 GND x331/junc1 x331/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3634 x995/RWL0_junc x995/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3635 RBL0_29 RWL_26 x651/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3636 x510/junc0 x510/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3637 x592/RWL0_junc x592/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3638 WBL_24 WWL_7 x985/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3639 RBL0_8 RWL_11 x806/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3640 GND x925/junc0 x925/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3641 GND x996/junc1 x996/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3642 RBL0_15 RWL_31 x425/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3643 x835/RWL0_junc x835/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3644 x901/junc0 x901/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3645 GND x324/junc0 x324/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3646 x10/junc0 x10/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3647 x98/junc1 WWL_2 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3648 RBL0_2 RWL_17 x775/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3649 x268/junc0 x268/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3650 GND x845/junc1 x845/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3651 GND x960/junc1 x960/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3652 x334/RWL0_junc x334/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3653 GND x430/junc0 x430/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3654 GND x431/junc0 x431/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3655 x525/junc0 x525/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3656 GND x997/junc1 x997/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3657 RBL0_6 RWL_13 x660/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3658 x824/RWL0_junc x824/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3659 x507/junc1 WWL_6 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3660 x460/junc0 x460/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3661 RBL0_26 RWL_7 x664/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3662 VDD x213/junc0 x213/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3663 x805/junc1 WWL_14 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3664 VDD x766/junc0 x766/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3665 RBL0_17 RWL_15 x779/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3666 x816/junc1 WWL_28 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3667 x157/junc1 WWL_16 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3668 RBL0_30 x389/RWL1 x667/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3669 x639/junc1 WWL_24 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3670 x633/junc0 x633/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3671 WBL_15 WWL_4 x397/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3672 x889/RWL1_junc RWL_10 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3673 WBL_2 WWL_2 x838/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3674 x890/RWL1_junc RWL_18 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3675 x524/RWL1_junc RWL_14 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3676 VDD x183/junc0 x183/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3677 x936/junc0 x936/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3678 WBL_4 WWL_29 x683/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3679 x833/junc1 WWL_21 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3680 x872/junc0 x872/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3681 GND x362/junc0 x362/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3682 x541/junc0 x541/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3683 GND x365/junc0 x365/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3684 VDD x776/junc0 x776/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3685 GND x370/junc1 x370/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3686 WBL_9 WWL_10 x429/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3687 x998/junc1 WWL_31 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3688 GND x661/junc1 x661/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3689 VDD x813/junc0 x813/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3690 x906/junc0 x906/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3691 x843/RWL0_junc x843/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3692 WBL_20 WWL_12 x409/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3693 x624/RWL0_junc x624/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3694 WBL_24 WWL_8 x990/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3695 RBL0_8 RWL_12 x22/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3696 x704/RWL0_junc x704/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3697 GND x968/junc1 x968/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3698 x948/junc0 x948/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3699 x556/junc0 x556/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3700 GND x376/junc0 x376/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3701 x64/junc0 x64/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3702 RBL0_11 RWL_10 x31/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3703 x818/junc1 WWL_17 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3704 WBL_18 WWL_14 x445/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3705 GND x390/junc1 x390/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3706 x629/RWL0_junc x629/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3707 RBL0_2 RWL_18 x796/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3708 x999/junc1 WWL_29 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3709 x1000/RWL0_junc x1000/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3710 x896/RWL1_junc RWL_21 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3711 x839/junc1 WWL_7 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3712 VDD x585/junc0 x585/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3713 x493/junc0 x493/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3714 RBL0_26 RWL_8 x44/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3715 VDD x790/junc0 x790/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3716 VDD x1001/junc0 x1001/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3717 VDD x587/junc0 x587/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3718 RBL0_17 RWL_16 x157/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3719 x789/junc0 x789/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3720 x898/RWL1_junc RWL_11 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3721 x52/RWL1_junc RWL_15 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3722 x900/RWL1_junc RWL_19 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3723 x873/junc0 x873/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3724 x443/junc0 x443/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3725 GND x408/junc0 x408/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3726 WBL_5 WWL_15 x860/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3727 WBL_9 WWL_11 x462/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3728 GND x414/junc1 x414/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3729 x33/RWL0_junc x33/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3730 x36/RWL0_junc x36/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3731 WBL_29 WWL_5 x1002/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3732 x39/RWL0_junc x39/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3733 WBL_20 WWL_13 x447/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3734 GND x413/junc0 x413/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3735 x187/junc1 WWL_2 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3736 x41/RWL0_junc x41/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3737 GND x760/junc1 x760/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3738 x43/RWL0_junc x43/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3739 x914/junc0 x914/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3740 GND x972/junc1 x972/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3741 x881/junc0 x881/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3742 x589/junc0 x589/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3743 GND x420/junc0 x420/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3744 x849/junc1 WWL_10 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3745 x773/junc0 x773/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3746 x916/junc0 x916/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3747 RBL0_11 RWL_11 x88/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3748 x827/junc1 WWL_18 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3749 GND x433/junc1 x433/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3750 x651/RWL0_junc x651/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3751 RBL0_2 RWL_19 x195/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3752 GND x917/junc0 x917/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3753 x546/junc0 x546/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3754 x858/junc0 x858/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3755 x354/junc0 x354/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3756 VDD x296/junc0 x296/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3757 x577/junc1 WWL_12 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3758 GND x696/junc1 x696/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3759 GND x381/junc0 x381/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3760 x904/RWL1_junc RWL_14 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3761 GND x829/junc0 x829/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3762 x851/junc1 WWL_8 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3763 x905/RWL1_junc RWL_22 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3764 VDD x264/junc0 x264/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3765 VDD x324/junc0 x324/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3766 GND x815/junc1 x815/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3767 x76/RWL0_junc x76/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3768 x907/RWL1_junc RWL_12 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3769 x108/RWL1_junc RWL_16 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3770 VDD x830/junc0 x830/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3771 x642/junc1 WWL_14 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3772 x821/RWL1_junc RWL_24 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3773 WBL_5 WWL_16 x872/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3774 x924/junc0 x924/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3775 x958/junc0 x958/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3776 x221/junc1 WWL_2 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3777 VDD x491/junc0 x491/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3778 x959/junc0 x959/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3779 GND x974/junc1 x974/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3780 GND x975/junc1 x975/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3781 GND x452/junc0 x452/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3782 x96/RWL0_junc x96/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3783 x100/RWL0_junc x100/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3784 x998/junc0 x998/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3785 VDD x329/junc0 x329/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3786 x603/junc1 WWL_15 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3787 RBL0_22 RWL_2 x133/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3788 WBL_23 WWL_12 x948/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3789 GND x749/junc1 x749/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3790 GND x784/junc1 x784/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3791 x859/junc1 WWL_11 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3792 x927/junc0 x927/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3793 RBL0_11 RWL_12 x725/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3794 x816/RWL1_junc RWL_28 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3795 GND x928/junc0 x928/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3796 x870/junc0 x870/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3797 GND x136/junc1 x136/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3798 x929/junc0 x929/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3799 VDD x1003/junc0 x1003/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3800 x248/junc1 WWL_13 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3801 x902/junc0 x902/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3802 GND x718/junc1 x718/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3803 x912/RWL1_junc RWL_15 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3804 x63/junc0 x63/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3805 x913/RWL1_junc RWL_23 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3806 x553/RWL0_junc x553/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3807 GND x734/junc0 x734/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3808 x126/RWL0_junc x126/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3809 VDD x840/junc0 x840/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3810 x615/junc1 WWL_19 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3811 x128/RWL0_junc x128/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3812 GND x156/junc1 x156/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3813 WBL_14 WWL_9 x873/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3814 x163/RWL1_junc RWL_25 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3815 x132/RWL0_junc x132/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3816 RBL0_24 RWL_24 x549/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3817 x931/junc0 x931/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3818 x596/junc0 x596/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3819 WBL_1 WWL_29 x441/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3820 GND x763/junc1 x763/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3821 GND x977/junc1 x977/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3822 x143/RWL0_junc x143/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3823 VDD x652/junc0 x652/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3824 x148/RWL0_junc x148/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3825 x146/RWL0_junc x146/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3826 x152/RWL0_junc x152/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3827 GND x935/junc0 x935/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3828 GND x482/junc0 x482/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3829 x884/junc0 x884/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3830 x885/junc0 x885/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3831 VDD x656/junc0 x656/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3832 RBL0_22 x61/RWL1 x186/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3833 VDD x1004/junc0 x1004/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3834 x628/junc1 WWL_16 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3835 WBL_23 WWL_13 x881/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3836 GND x802/junc1 x802/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3837 GND x42/junc1 x42/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3838 x562/RWL1_junc RWL_30 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3839 x234/RWL1_junc RWL_29 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3840 GND x561/junc0 x561/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3841 WBL_31 WWL_17 x858/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3842 RBL0_15 RWL_21 x599/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3843 WBL_30 WWL_21 x546/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3844 x89/RWL1_junc RWL_20 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3845 x938/junc0 x938/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3846 VDD x895/junc0 x895/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3847 x679/junc1 WWL_22 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3848 RBL0_0 RWL_14 x191/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3849 GND x979/junc1 x979/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3850 x1005/junc0 x1005/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3851 x921/RWL1_junc RWL_16 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3852 GND x337/junc1 x337/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3853 x87/RWL0_junc x87/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3854 GND x500/junc0 x500/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3855 x833/RWL1_junc RWL_21 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3856 x637/junc1 WWL_12 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3857 WBL_13 WWL_30 x755/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3858 VDD x852/junc0 x852/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3859 x982/junc0 x982/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3860 x877/junc1 WWL_20 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3861 x173/RWL0_junc x173/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3862 x61/RWL0_junc x61/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3863 x620/junc0 x620/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3864 GND x200/junc1 x200/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3865 GND x19/junc0 x19/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3866 GND x75/junc1 x75/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3867 x208/RWL1_junc RWL_26 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3868 x181/RWL0_junc x181/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3869 x203/RWL0_junc x203/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3870 x939/junc0 x939/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3871 RBL0_24 RWL_25 x209/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3872 x655/junc0 x655/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3873 x625/junc0 x625/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3874 WBL_19 WWL_6 x958/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3875 x626/junc0 x626/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3876 RBL0_3 RWL_10 x214/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3877 x1006/junc0 x1006/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3878 RBL0_7 RWL_6 x304/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3879 GND x787/junc1 x787/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3880 x196/RWL0_junc x196/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3881 VDD x854/junc0 x854/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3882 x568/junc0 x568/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3883 RBL0_27 RWL_0 x218/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3884 GND x513/junc0 x513/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3885 x930/RWL1_junc RWL_9 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3886 GND x251/junc1 x251/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3887 GND x590/junc0 x590/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3888 VDD x856/junc0 x856/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3889 x465/junc0 x465/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3890 VDD x1007/junc0 x1007/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3891 GND x817/junc1 x817/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3892 GND x97/junc1 x97/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3893 WBL_23 WWL_28 x766/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3894 WBL_27 WWL_22 x556/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3895 VDD x377/junc0 x377/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3896 x613/RWL0_junc x613/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3897 RBL0_15 RWL_22 x994/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3898 WBL_31 WWL_18 x870/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3899 RBL0_25 RWL_2 x759/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3900 x702/junc1 WWL_23 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3901 x674/junc0 x674/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3902 RBL0_0 RWL_15 x238/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3903 RBL0_23 RWL_31 x251/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3904 WBL_10 WWL_3 x902/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3905 x472/junc0 x472/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3906 GND x379/junc1 x379/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3907 VDD x862/junc0 x862/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3908 GND x863/junc0 x863/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3909 x246/RWL1_junc RWL_22 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3910 x934/RWL1_junc RWL_13 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3911 x139/RWL0_junc x139/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3912 x150/RWL1_junc RWL_27 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3913 x689/junc0 x689/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3914 WBL_13 WWL_31 x776/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3915 x941/junc0 x941/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3916 x336/junc1 WWL_13 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3917 x942/junc0 x942/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3918 x216/RWL0_junc x216/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3919 x62/junc0 x62/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3920 x645/junc0 x645/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3921 GND x867/junc0 x867/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3922 x662/junc1 WWL_25 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3923 GND x129/junc1 x129/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3924 x250/RWL0_junc x250/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3925 x944/junc0 x944/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3926 x225/RWL0_junc x225/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3927 RBL0_24 RWL_26 x765/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3928 x677/junc0 x677/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3929 x650/junc0 x650/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3930 x865/junc1 WWL_10 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3931 WBL_19 WWL_7 x596/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3932 RBL0_3 RWL_11 x261/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3933 x236/RWL0_junc x236/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3934 x240/RWL0_junc x240/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3935 x1008/junc0 x1008/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3936 WBL_12 WWL_25 x531/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3937 RBL0_27 RWL_1 x269/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3938 x270/RWL1_junc RWL_6 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3939 GND x868/junc0 x868/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3940 GND x910/junc1 x910/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3941 GND x983/junc1 x983/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3942 x549/RWL0_junc x549/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3943 GND x621/junc0 x621/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3944 WBL_16 WWL_21 x884/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3945 VDD x869/junc0 x869/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3946 WBL_1 WWL_14 x885/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3947 GND x151/junc1 x151/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3948 GND x778/junc0 x778/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3949 WBL_19 WWL_30 x790/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3950 x675/junc1 WWL_6 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3951 VDD x871/junc0 x871/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3952 x945/junc0 x945/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3953 WBL_27 WWL_23 x589/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3954 RBL0_21 RWL_7 x281/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3955 VDD x844/junc0 x844/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3956 x646/junc0 x646/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3957 RBL0_15 RWL_23 x997/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3958 RBL0_25 x389/RWL1 x780/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3959 x723/junc1 WWL_24 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3960 RBL0_0 RWL_16 x781/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3961 WBL_10 WWL_4 x1005/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3962 GND x553/junc0 x553/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3963 x189/RWL1_junc RWL_10 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3964 GND x563/junc0 x563/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3965 x642/RWL1_junc RWL_14 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3966 VDD x26/junc0 x26/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3967 VDD x874/junc0 x874/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3968 x291/RWL1_junc RWL_23 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3969 x946/junc0 x946/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3970 GND x573/junc0 x573/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3971 x698/junc0 x698/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3972 x668/junc0 x668/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3973 WBL_4 WWL_10 x620/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3974 GND x578/junc1 x578/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3975 x687/junc1 WWL_22 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3976 x688/junc1 WWL_26 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3977 VDD x878/junc0 x878/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3978 RBL0_28 RWL_27 x854/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3979 x947/junc0 x947/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3980 x4/junc0 x4/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3981 x275/RWL0_junc x275/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3982 x690/junc1 WWL_3 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3983 WBL_28 WWL_0 x625/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3984 RBL0_12 RWL_4 x856/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3985 x876/junc1 WWL_11 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3986 x164/junc1 WWL_30 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3987 WBL_19 WWL_8 x626/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3988 RBL0_3 RWL_12 x300/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3989 GND x324/junc1 x324/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3990 x286/RWL0_junc x286/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3991 x978/junc0 x978/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M3992 x475/junc1 WWL_28 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3993 GND x640/junc0 x640/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3994 GND x986/junc1 x986/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3995 x215/RWL1_junc RWL_7 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3996 GND x950/junc0 x950/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3997 GND x582/junc0 x582/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3998 WBL_12 WWL_26 x568/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M3999 GND x987/junc1 x987/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4000 RBL0_6 RWL_10 x305/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4001 x809/RWL0_junc x809/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4002 x671/RWL0_junc x671/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4003 GND x190/junc1 x190/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4004 x209/RWL0_junc x209/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4005 GND x591/junc0 x591/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4006 WBL_19 WWL_31 x324/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4007 x293/RWL0_junc x293/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4008 x903/junc1 WWL_7 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4009 RBL0_30 RWL_0 x316/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4010 VDD x886/junc0 x886/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4011 WBL_27 WWL_24 x618/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4012 x951/junc0 x951/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4013 RBL0_21 RWL_8 x320/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4014 VDD x728/junc0 x728/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4015 x237/RWL1_junc RWL_11 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4016 x85/junc1 WWL_25 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4017 x165/junc0 x165/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4018 VDD x632/junc0 x632/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4019 x328/RWL1_junc RWL_15 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4020 x930/junc0 x930/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4021 x48/junc0 x48/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4022 GND x606/junc0 x606/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4023 x545/junc0 x545/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4024 WBL_13 WWL_3 x62/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4025 GND x611/junc1 x611/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4026 WBL_4 WWL_11 x645/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4027 x708/junc1 WWL_23 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4028 x270/RWL0_junc x270/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4029 x887/junc1 WWL_27 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4030 WBL_10 WWL_29 x491/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4031 x241/RWL0_junc x241/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4032 GND x180/junc0 x180/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4033 WBL_24 WWL_5 x976/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4034 GND x182/junc0 x182/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4035 x312/RWL0_junc x312/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4036 GND x953/junc0 x953/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4037 x888/junc1 WWL_4 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4038 WBL_28 WWL_1 x650/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4039 RBL0_12 RWL_5 x869/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4040 GND x223/junc1 x223/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4041 x741/junc0 x741/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4042 x211/junc1 WWL_31 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4043 x34/RWL0_junc x34/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4044 GND x5/junc1 x5/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4045 x65/junc0 x65/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4046 GND x991/junc1 x991/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4047 x934/junc0 x934/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4048 x262/RWL1_junc RWL_8 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4049 x981/RWL0_junc x981/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4050 GND x616/junc0 x616/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4051 x684/junc0 x684/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4052 x793/junc1 WWL_10 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4053 x954/junc0 x954/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4054 x822/RWL0_junc x822/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4055 WBL_12 WWL_27 x1008/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4056 RBL0_6 RWL_11 x348/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4057 x765/RWL0_junc x765/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4058 GND x955/junc0 x955/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4059 x700/junc0 x700/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4060 x917/junc0 x917/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4061 VDD x511/junc0 x511/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4062 x719/junc1 WWL_12 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4063 x564/junc0 x564/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4064 GND x804/junc1 x804/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4065 GND x201/junc0 x201/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4066 GND x893/junc0 x893/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4067 x273/RWL1_junc RWL_14 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4068 x331/RWL0_junc x331/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4069 RBL0_30 RWL_1 x360/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4070 x911/junc1 WWL_8 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4071 WBL_15 WWL_2 x646/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4072 x722/junc1 WWL_26 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4073 x338/RWL0_junc x338/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4074 x948/RWL1_junc RWL_12 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4075 VDD x894/junc0 x894/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4076 x724/junc1 WWL_19 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4077 x369/RWL1_junc RWL_16 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4078 RBL0_29 RWL_13 x815/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4079 RBL0_14 RWL_27 x368/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4080 x880/RWL1_junc RWL_24 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4081 VDD x897/junc0 x897/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4082 WBL_13 WWL_4 x668/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4083 x821/junc1 WWL_24 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4084 GND x49/junc1 x49/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4085 GND x995/junc1 x995/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4086 GND x681/junc0 x681/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4087 GND x961/junc0 x961/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4088 x90/RWL0_junc x90/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4089 VDD x901/junc0 x901/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4090 x962/junc0 x962/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4091 VDD x543/junc0 x543/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4092 x162/junc1 WWL_15 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4093 RBL0_17 RWL_2 x735/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4094 WBL_18 WWL_12 x978/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4095 GND x835/junc1 x835/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4096 x501/junc1 WWL_3 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4097 x806/junc1 WWL_11 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4098 x963/junc0 x963/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4099 RBL0_6 RWL_12 x825/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4100 x53/RWL1_junc RWL_28 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4101 x707/junc0 x707/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4102 GND x641/junc0 x641/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4103 GND x964/junc0 x964/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4104 x928/junc0 x928/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4105 x169/junc1 WWL_5 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4106 GND x289/junc1 x289/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4107 x529/RWL1_junc RWL_27 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4108 x965/junc0 x965/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4109 VDD x1009/junc0 x1009/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4110 x473/junc1 WWL_13 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4111 x23/junc0 x23/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4112 GND x824/junc1 x824/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4113 x952/RWL1_junc RWL_15 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4114 x138/junc0 x138/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4115 x967/junc0 x967/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4116 VDD x761/junc0 x761/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4117 x380/RWL0_junc x380/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4118 x713/junc1 WWL_29 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4119 x922/junc1 WWL_27 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4120 x923/junc1 WWL_20 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4121 WBL_9 WWL_9 x930/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4122 x415/RWL1_junc RWL_25 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4123 x390/RWL0_junc x390/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4124 RBL0_19 RWL_24 x12/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4125 VDD x906/junc0 x906/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4126 x266/junc0 x266/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4127 WBL_8 WWL_21 x411/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4128 GND x106/junc1 x106/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4129 GND x843/junc1 x843/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4130 RBL0_16 RWL_30 x744/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4131 VDD x769/junc0 x769/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4132 x140/RWL0_junc x140/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4133 x1010/RWL0_junc x1010/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4134 GND x969/junc0 x969/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4135 GND x659/junc0 x659/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4136 x935/junc0 x935/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4137 VDD x771/junc0 x771/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4138 x265/junc0 x265/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4139 RBL0_17 x61/RWL1 x501/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4140 VDD x1011/junc0 x1011/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4141 x748/junc1 WWL_16 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4142 WBL_18 WWL_13 x934/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4143 x193/junc1 WWL_4 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4144 x949/junc0 x949/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4145 x729/junc0 x729/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4146 x713/RWL1_junc RWL_29 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4147 x714/RWL1_junc RWL_2 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4148 GND x665/junc0 x665/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4149 x958/RWL1_junc RWL_6 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4150 x179/junc0 x179/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4151 GND x712/junc0 x712/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4152 WBL_26 WWL_17 x917/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4153 RBL0_10 RWL_21 x42/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4154 WBL_25 WWL_21 x700/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4155 x349/RWL1_junc RWL_20 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4156 x970/junc0 x970/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4157 VDD x943/junc0 x943/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4158 GND x326/junc1 x326/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4159 x104/junc0 x104/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4160 GND x1000/junc1 x1000/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4161 x117/RWL1_junc RWL_28 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4162 x959/RWL1_junc RWL_16 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4163 x875/junc0 x875/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4164 x347/RWL0_junc x347/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4165 x971/junc0 x971/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4166 x797/junc1 WWL_12 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4167 VDD x783/junc0 x783/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4168 x424/RWL0_junc x424/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4169 WBL_20 WWL_0 x440/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4170 RBL0_26 RWL_28 x754/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4171 x454/RWL1_junc RWL_26 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4172 x433/RWL0_junc x433/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4173 x739/junc1 WWL_29 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4174 RBL0_19 RWL_25 x68/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4175 x198/junc0 x198/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4176 x125/junc0 x125/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4177 GND x973/junc0 x973/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4178 x334/RWL1_junc RWL_24 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4179 RBL0_2 RWL_6 x525/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4180 GND x159/junc1 x159/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4181 GND x39/junc1 x39/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4182 x815/RWL0_junc x815/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4183 x368/RWL0_junc x368/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4184 VDD x914/junc0 x914/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4185 x715/junc0 x715/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4186 RBL0_22 RWL_0 x460/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4187 GND x43/junc1 x43/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4188 GND x657/junc0 x657/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4189 x297/junc0 x297/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4190 GND x730/junc0 x730/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4191 GND x682/junc0 x682/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4192 x966/RWL1_junc RWL_9 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4193 VDD x909/junc0 x909/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4194 VDD x916/junc0 x916/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4195 x536/junc1 WWL_9 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4196 x302/junc0 x302/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4197 VDD x1012/junc0 x1012/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4198 WBL_2 WWL_28 x844/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4199 x37/junc0 x37/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4200 x745/junc0 x745/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4201 WBL_22 WWL_22 x707/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4202 x144/junc0 x144/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4203 VDD x255/junc0 x255/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4204 GND x918/junc0 x918/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4205 x468/RWL1_junc x389/RWL1 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4206 x220/junc0 x220/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4207 x83/junc1 WWL_21 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4208 RBL0_10 RWL_22 x97/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4209 x785/junc0 x785/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4210 WBL_26 WWL_18 x928/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4211 GND x367/junc1 x367/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4212 x164/RWL1_junc RWL_30 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4213 WBL_5 WWL_3 x23/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4214 x153/junc0 x153/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4215 x739/RWL1_junc RWL_29 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4216 x457/RWL0_junc x457/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4217 x398/RWL0_junc x398/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4218 x232/junc0 x232/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4219 VDD x919/junc0 x919/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4220 x810/junc1 WWL_13 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4221 x331/junc0 x331/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4222 WBL_20 WWL_1 x470/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4223 RBL0_22 RWL_30 x770/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4224 RBL0_26 RWL_29 x773/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4225 x279/junc1 WWL_25 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4226 x813/junc1 WWL_21 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4227 x245/junc0 x245/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4228 RBL0_19 RWL_26 x123/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4229 x172/junc0 x172/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4230 GND x999/junc0 x999/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4231 GND x485/junc1 x485/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4232 x629/RWL1_junc RWL_25 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4233 x471/RWL0_junc x471/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4234 x79/junc0 x79/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4235 x77/junc0 x77/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4236 x121/junc1 WWL_0 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4237 x184/junc0 x184/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4238 WBL_7 WWL_25 x692/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4239 RBL0_22 RWL_1 x493/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4240 GND x100/junc1 x100/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4241 x8/RWL1_junc RWL_2 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4242 x12/RWL0_junc x12/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4243 GND x926/junc0 x926/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4244 GND x680/junc0 x680/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4245 GND x746/junc0 x746/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4246 WBL_11 WWL_21 x935/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4247 VDD x915/junc0 x915/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4248 VDD x927/junc0 x927/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4249 WBL_31 WWL_15 x695/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4250 x791/junc1 WWL_6 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4251 WBL_30 WWL_19 x949/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4252 VDD x929/junc0 x929/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4253 WBL_22 WWL_23 x729/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4254 x891/junc0 x891/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4255 x9/junc0 x9/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4256 RBL0_10 RWL_23 x151/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4257 WBL_29 WWL_28 x632/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4258 WBL_5 WWL_4 x104/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4259 GND x936/junc1 x936/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4260 x438/RWL1_junc RWL_10 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4261 VDD x301/junc0 x301/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4262 x38/RWL0_junc x38/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4263 x285/junc0 x285/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4264 GND x717/junc0 x717/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4265 x207/junc0 x207/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4266 GND x128/junc1 x128/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4267 GND x422/junc1 x422/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4268 x40/junc1 WWL_22 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4269 x798/junc1 WWL_26 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4270 VDD x931/junc0 x931/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4271 RBL0_23 RWL_27 x914/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4272 x290/junc0 x290/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4273 x495/RWL0_junc x495/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4274 x264/RWL0_junc x264/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4275 x35/junc0 x35/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4276 x800/junc1 WWL_3 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4277 WBL_23 WWL_0 x125/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4278 RBL0_7 RWL_4 x916/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4279 GND x145/junc1 x145/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4280 x651/RWL1_junc RWL_26 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4281 x503/RWL0_junc x503/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4282 x774/junc0 x774/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4283 GND x756/junc0 x756/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4284 GND x143/junc1 x143/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4285 x458/RWL1_junc RWL_7 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4286 GND x980/junc0 x980/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4287 x950/junc0 x950/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4288 x168/junc1 WWL_1 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4289 VDD x634/junc0 x634/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4290 x1013/RWL0_junc x1013/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4291 WBL_7 WWL_26 x715/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4292 x502/junc0 x502/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4293 GND x148/junc1 x148/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4294 GND x152/junc1 x152/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4295 x66/RWL0_junc x66/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4296 x62/RWL1_junc x61/RWL1 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4297 GND x439/junc1 x439/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4298 GND x703/junc0 x703/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4299 x68/RWL0_junc x68/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4300 WBL_16 WWL_29 x25/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4301 x75/RWL0_junc x75/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4302 x178/junc1 WWL_7 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4303 RBL0_15 RWL_20 x190/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4304 WBL_30 WWL_20 x144/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4305 VDD x938/junc0 x938/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4306 WBL_31 WWL_16 x37/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4307 RBL0_25 RWL_0 x192/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4308 WBL_22 WWL_24 x745/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4309 GND x553/junc1 x553/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4310 x922/RWL1_junc RWL_27 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4311 x767/RWL1_junc RWL_13 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4312 x469/RWL1_junc RWL_11 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4313 x82/junc1 WWL_25 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4314 x923/RWL1_junc RWL_20 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4315 x315/junc0 x315/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4316 x966/junc0 x966/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4317 x537/RWL0_junc x537/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4318 x323/junc0 x323/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4319 GND x738/junc0 x738/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4320 x256/junc0 x256/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4321 GND x61/junc1 x61/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4322 GND x459/junc1 x459/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4323 x93/junc1 WWL_23 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4324 VDD x939/junc0 x939/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4325 x197/junc1 WWL_27 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4326 x792/junc0 x792/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4327 WBL_19 WWL_5 x996/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4328 GND x434/junc0 x434/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4329 x205/junc1 WWL_4 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4330 x58/junc0 x58/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4331 WBL_23 WWL_1 x172/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4332 RBL0_7 RWL_5 x927/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4333 GND x464/junc1 x464/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4334 GND x292/junc1 x292/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4335 x534/RWL0_junc x534/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4336 x193/RWL1_junc RWL_4 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4337 GND x196/junc1 x196/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4338 x488/RWL1_junc RWL_8 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4339 RBL0_15 RWL_9 x223/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4340 x768/RWL0_junc x768/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4341 WBL_16 WWL_19 x77/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4342 RBL0_0 RWL_2 x221/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4343 x102/junc0 x102/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4344 x214/junc1 WWL_10 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4345 WBL_1 WWL_12 x79/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4346 x883/RWL0_junc x883/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4347 VDD x203/junc0 x203/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4348 WBL_7 WWL_27 x184/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4349 x119/RWL0_junc x119/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4350 x123/RWL0_junc x123/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4351 x59/junc1 WWL_28 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4352 x283/junc0 x283/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4353 x955/junc0 x955/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4354 x786/RWL1_junc RWL_9 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4355 GND x447/junc0 x447/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4356 x218/junc1 WWL_0 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4357 x126/RWL1_junc RWL_14 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4358 x129/RWL0_junc x129/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4359 RBL0_25 RWL_1 x235/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4360 x222/junc1 WWL_8 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4361 WBL_10 WWL_2 x891/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4362 x84/junc0 x84/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4363 x801/junc1 WWL_29 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4364 RBL0_20 RWL_17 x804/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4365 x355/junc0 x355/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4366 x137/junc1 WWL_26 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4367 VDD x941/junc0 x941/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4368 x978/RWL1_junc RWL_12 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4369 VDD x942/junc0 x942/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4370 RBL0_24 RWL_13 x248/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4371 RBL0_9 RWL_27 x249/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4372 x8/junc0 x8/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4373 x933/RWL1_junc RWL_24 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4374 VDD x834/junc0 x834/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4375 x880/junc1 WWL_24 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4376 VDD x944/junc0 x944/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4377 x298/junc0 x298/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4378 GND x30/junc0 x30/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4379 x644/junc1 WWL_9 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4380 GND x325/junc1 x325/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4381 GND x225/junc1 x225/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4382 WBL_22 WWL_29 x115/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4383 x572/RWL0_junc x572/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4384 x160/RWL0_junc x160/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4385 GND x984/junc0 x984/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4386 VDD x1014/junc0 x1014/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4387 WBL_27 WWL_10 x580/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4388 GND x236/junc1 x236/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4389 GND x240/junc1 x240/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4390 x239/RWL1_junc RWL_5 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4391 RBL0_0 RWL_3 x272/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4392 x261/junc1 WWL_11 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4393 VDD x174/junc0 x174/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4394 WBL_16 WWL_20 x950/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4395 WBL_1 WWL_13 x502/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4396 x803/junc0 x803/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4397 x166/RWL0_junc x166/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4398 GND x757/junc0 x757/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4399 x704/junc1 WWL_30 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4400 RBL0_19 RWL_31 x324/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4401 x83/RWL1_junc RWL_21 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4402 GND x758/junc0 x758/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4403 x578/RWL0_junc x578/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4404 x420/junc1 WWL_5 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4405 x964/junc0 x964/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4406 VDD x945/junc0 x945/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4407 VDD x417/junc0 x417/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4408 x173/RWL1_junc RWL_15 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4409 x269/junc1 WWL_1 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4410 x396/junc0 x396/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4411 x136/junc0 x136/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4412 x985/junc0 x985/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4413 RBL0_29 RWL_10 x289/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4414 VDD x841/junc0 x841/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4415 RBL0_28 RWL_14 x939/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4416 RBL0_20 RWL_18 x824/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4417 x187/RWL0_junc x187/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4418 x69/junc0 x69/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4419 x960/junc1 WWL_27 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4420 VDD x946/junc0 x946/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4421 x538/RWL1_junc RWL_17 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4422 WBL_4 WWL_9 x966/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4423 x612/RWL1_junc RWL_25 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4424 x193/RWL0_junc x193/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4425 VDD x947/junc0 x947/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4426 GND x988/junc0 x988/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4427 GND x989/junc0 x989/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4428 x340/junc0 x340/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4429 x669/junc1 WWL_2 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4430 VDD x0/junc0 x0/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4431 GND x523/junc1 x523/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4432 WBL_3 WWL_21 x792/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4433 GND x366/junc1 x366/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4434 GND x275/junc1 x275/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4435 VDD x847/junc0 x847/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4436 x605/RWL0_junc x605/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4437 x204/RWL0_junc x204/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4438 GND x831/junc0 x831/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4439 GND x775/junc0 x775/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4440 x397/junc0 x397/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4441 WBL_27 WWL_11 x614/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4442 x485/junc0 x485/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4443 x969/junc0 x969/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4444 VDD x848/junc0 x848/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4445 GND x286/junc1 x286/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4446 VDD x72/junc0 x72/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4447 x979/junc0 x979/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4448 x823/junc0 x823/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4449 GND x777/junc0 x777/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4450 x1015/junc1 WWL_31 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4451 x133/RWL1_junc RWL_2 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4452 GND x613/junc0 x613/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4453 x135/RWL1_junc RWL_22 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4454 GND x779/junc0 x779/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4455 x611/RWL0_junc x611/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4456 x429/junc0 x429/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4457 WBL_21 WWL_17 x955/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4458 VDD x951/junc0 x951/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4459 RBL0_5 RWL_21 x318/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4460 x112/junc0 x112/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4461 x372/RWL1_junc RWL_28 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4462 x216/RWL1_junc RWL_16 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4463 x968/junc1 WWL_10 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4464 x313/junc1 WWL_14 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4465 x224/RWL0_junc x224/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4466 x990/junc0 x990/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4467 RBL0_29 RWL_11 x326/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4468 VDD x853/junc0 x853/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4469 RBL0_20 RWL_19 x1000/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4470 RBL0_28 RWL_15 x944/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4471 x226/RWL0_junc x226/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4472 RBL0_5 RWL_28 x243/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4473 WBL_13 WWL_2 x8/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4474 x574/RWL1_junc RWL_18 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4475 VDD x764/junc0 x764/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4476 x635/RWL1_junc RWL_26 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4477 x828/junc1 WWL_29 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4478 x239/RWL0_junc x239/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4479 x445/junc0 x445/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4480 x378/junc0 x378/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4481 GND x992/junc0 x992/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4482 x1006/RWL1_junc RWL_31 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4483 GND x993/junc0 x993/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4484 WBL_12 WWL_14 x298/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4485 GND x560/junc1 x560/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4486 x549/RWL1_junc RWL_24 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4487 GND x412/junc1 x412/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4488 GND x312/junc1 x312/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4489 x248/RWL0_junc x248/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4490 x249/RWL0_junc x249/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4491 VDD x855/junc0 x855/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4492 VDD x65/junc0 x65/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4493 x391/junc0 x391/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4494 x817/junc0 x817/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4495 x252/RWL0_junc x252/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4496 RBL0_17 RWL_0 x945/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4497 GND x535/junc0 x535/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4498 x516/junc0 x516/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4499 GND x796/junc0 x796/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4500 x242/junc0 x242/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4501 x694/junc1 WWL_9 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4502 x145/junc0 x145/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4503 VDD x954/junc0 x954/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4504 x212/junc0 x212/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4505 x403/junc0 x403/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4506 x307/junc0 x307/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4507 x1016/junc0 x1016/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4508 WBL_17 WWL_22 x803/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4509 VDD x479/junc0 x479/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4510 x186/RWL1_junc x61/RWL1 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4511 x258/junc1 WWL_6 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4512 GND x155/junc0 x155/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4513 x185/RWL1_junc RWL_23 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4514 x341/junc1 WWL_17 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4515 GND x157/junc0 x157/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4516 x462/junc0 x462/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4517 x649/RWL0_junc x649/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4518 GND x755/junc0 x755/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4519 x343/junc1 WWL_21 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4520 WBL_21 WWL_18 x964/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4521 RBL0_14 RWL_14 x359/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4522 RBL0_5 RWL_22 x361/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4523 x828/RWL1_junc RWL_29 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4524 VDD x956/junc0 x956/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4525 x599/RWL1_junc RWL_21 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4526 x271/RWL0_junc x271/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4527 x972/junc1 WWL_11 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4528 x274/RWL0_junc x274/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4529 RBL0_29 RWL_12 x367/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4530 VDD x957/junc0 x957/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4531 RBL0_28 RWL_16 x4/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4532 x234/junc0 x234/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4533 RBL0_1 RWL_30 x506/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4534 RBL0_5 RWL_29 x287/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4535 x500/junc1 WWL_25 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4536 x949/RWL1_junc RWL_19 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4537 x10/junc0 x10/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4538 VDD x107/junc0 x107/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4539 x268/junc0 x268/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4540 x423/junc0 x423/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4541 WBL_8 WWL_19 x323/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4542 x289/RWL0_junc x289/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4543 x209/RWL1_junc RWL_25 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4544 x371/RWL0_junc x371/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4545 VDD x962/junc0 x962/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4546 GND x766/junc0 x766/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4547 x339/junc0 x339/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4548 x191/RWL1_junc RWL_14 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4549 x375/junc1 WWL_0 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4550 x435/junc0 x435/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4551 WBL_2 WWL_25 x802/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4552 RBL0_17 RWL_1 x951/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4553 x293/RWL1_junc RWL_2 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4554 GND x195/junc0 x195/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4555 x735/junc1 WWL_2 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4556 WBL_6 WWL_21 x969/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4557 VDD x963/junc0 x963/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4558 x218/RWL1_junc RWL_0 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4559 x622/RWL1_junc RWL_4 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4560 x936/junc0 x936/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4561 WBL_26 WWL_15 x267/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4562 WBL_17 WWL_23 x823/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4563 WBL_25 WWL_19 x979/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4564 VDD x965/junc0 x965/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4565 RBL0_1 RWL_27 x774/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4566 x940/junc0 x940/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4567 x975/junc1 WWL_7 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4568 x1015/junc0 x1015/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4569 x392/junc1 WWL_18 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4570 x974/junc1 WWL_14 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4571 x202/junc0 x202/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4572 RBL0_14 RWL_15 x405/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4573 RBL0_5 RWL_23 x406/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4574 WBL_8 WWL_28 x752/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4575 GND x709/junc1 x709/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4576 GND x813/junc0 x813/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4577 VDD x967/junc0 x967/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4578 GND x466/junc1 x466/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4579 x994/RWL1_junc RWL_22 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4580 x309/RWL0_junc x309/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4581 GND x380/junc1 x380/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4582 x394/RWL1_junc RWL_31 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4583 x314/junc1 WWL_22 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4584 x59/RWL1_junc RWL_28 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4585 x863/junc1 WWL_26 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4586 RBL0_18 RWL_27 x65/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4587 x842/RWL0_junc x842/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4588 x490/RWL0_junc x490/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4589 x64/junc0 x64/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4590 x217/junc0 x217/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4591 WBL_18 WWL_0 x378/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4592 x867/junc1 WWL_3 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4593 WBL_8 WWL_20 x17/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4594 RBL0_2 RWL_4 x954/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4595 x326/RWL0_junc x326/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4596 WBL_31 WWL_30 x924/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4597 x745/junc0 x745/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4598 x987/junc0 x987/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4599 x850/junc0 x850/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4600 RBL0_18 RWL_28 x864/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4601 x765/RWL1_junc RWL_26 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4602 x1017/RWL0_junc x1017/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4603 GND x228/junc0 x228/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4604 GND x790/junc0 x790/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4605 GND x1001/junc0 x1001/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4606 x638/RWL1_junc RWL_7 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4607 GND x230/junc0 x230/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4608 WBL_0 WWL_21 x391/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4609 x980/junc0 x980/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4610 x238/RWL1_junc RWL_15 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4611 x419/junc1 WWL_1 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4612 VDD x753/junc0 x753/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4613 WBL_2 WWL_26 x817/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4614 GND x1010/junc1 x1010/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4615 x333/RWL0_junc x333/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4616 x331/RWL1_junc x61/RWL1 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4617 GND x864/junc1 x864/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4618 GND x919/junc0 x919/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4619 x269/RWL1_junc RWL_1 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4620 x996/RWL1_junc RWL_5 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4621 VDD x179/junc0 x179/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4622 x868/junc1 WWL_19 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4623 GND x489/junc1 x489/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4624 RBL0_10 RWL_20 x439/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4625 WBL_25 WWL_20 x403/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4626 VDD x970/junc0 x970/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4627 WBL_26 WWL_16 x307/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4628 WBL_17 WWL_24 x1016/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4629 x607/RWL1_junc RWL_31 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4630 x977/junc1 WWL_8 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4631 RBL0_14 RWL_16 x442/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4632 GND x254/junc0 x254/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4633 x960/RWL1_junc RWL_27 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4634 x845/RWL1_junc RWL_13 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4635 VDD x971/junc0 x971/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4636 x342/junc1 WWL_25 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4637 GND x496/junc1 x496/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4638 x997/RWL1_junc RWL_23 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4639 x517/RWL0_junc x517/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4640 GND x424/junc1 x424/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4641 x359/RWL0_junc x359/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4642 x358/junc1 WWL_23 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4643 x897/junc1 WWL_19 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4644 VDD x198/junc0 x198/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4645 x115/RWL1_junc RWL_29 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4646 x444/junc1 WWL_27 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4647 GND x623/junc0 x623/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4648 x451/junc1 WWL_4 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4649 WBL_18 WWL_1 x423/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4650 RBL0_2 RWL_5 x963/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4651 x367/RWL0_junc x367/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4652 x546/junc0 x546/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4653 x858/junc0 x858/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4654 WBL_31 WWL_31 x932/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4655 x354/junc0 x354/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4656 x14/junc0 x14/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4657 x130/junc0 x130/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4658 x861/junc0 x861/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4659 RBL0_18 RWL_29 x875/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4660 x370/RWL1_junc RWL_0 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4661 x661/RWL1_junc RWL_8 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4662 RBL0_10 RWL_9 x464/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4663 WBL_11 WWL_19 x339/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4664 x284/junc0 x284/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4665 WBL_2 WWL_27 x435/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4666 x781/RWL1_junc RWL_16 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4667 GND x875/junc1 x875/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4668 x374/RWL0_junc x374/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4669 GND x830/junc0 x830/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4670 x460/junc1 WWL_0 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4671 VDD x220/junc0 x220/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4672 x461/junc1 WWL_20 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4673 GND x520/junc1 x520/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4674 WBL_5 WWL_2 x940/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4675 x968/RWL1_junc RWL_10 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4676 x346/junc0 x346/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4677 x591/junc1 WWL_25 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4678 GND x455/junc1 x455/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4679 GND x295/junc0 x295/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4680 x633/RWL1_junc RWL_31 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4681 x567/junc0 x567/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4682 x395/junc1 WWL_26 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4683 VDD x232/junc0 x232/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4684 RBL0_4 RWL_27 x474/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4685 GND x528/junc1 x528/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4686 RBL0_19 RWL_13 x473/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4687 GND x457/junc1 x457/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4688 x293/junc0 x293/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4689 VDD x900/junc0 x900/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4690 x710/RWL0_junc x710/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4691 x552/RWL0_junc x552/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4692 x405/RWL0_junc x405/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4693 x933/junc1 WWL_24 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4694 x906/junc1 WWL_20 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4695 VDD x245/junc0 x245/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4696 x57/junc0 x57/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4697 x518/junc0 x518/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4698 GND x646/junc0 x646/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4699 GND x304/junc0 x304/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4700 GND x539/junc1 x539/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4701 x870/junc0 x870/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4702 x311/junc0 x311/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4703 x310/junc0 x310/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4704 x984/junc0 x984/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4705 GND x1003/junc0 x1003/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4706 WBL_30 WWL_6 x987/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4707 x175/junc0 x175/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4708 WBL_22 WWL_10 x850/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4709 GND x471/junc1 x471/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4710 x475/junc0 x475/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4711 x414/RWL1_junc RWL_1 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4712 WBL_11 WWL_20 x980/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4713 x418/RWL0_junc x418/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4714 GND x840/junc0 x840/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4715 x343/RWL1_junc RWL_21 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4716 x422/RWL0_junc x422/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4717 x616/junc1 WWL_5 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4718 VDD x808/junc0 x808/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4719 GND x327/junc0 x327/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4720 x493/junc1 WWL_1 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4721 VDD x265/junc0 x265/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4722 GND x557/junc1 x557/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4723 x809/junc1 WWL_28 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4724 x972/RWL1_junc RWL_11 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4725 x394/junc0 x394/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4726 x893/junc1 WWL_26 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4727 x596/junc0 x596/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4728 RBL0_24 RWL_10 x505/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4729 VDD x905/junc0 x905/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4730 RBL0_23 RWL_14 x198/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4731 x335/junc0 x335/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4732 x983/junc1 WWL_27 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4733 VDD x285/junc0 x285/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4734 RBL0_16 RWL_31 x553/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4735 GND x38/junc1 x38/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4736 x696/RWL1_junc RWL_17 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4737 VDD x907/junc0 x907/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4738 VDD x290/junc0 x290/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4739 GND x842/junc0 x842/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4740 x815/RWL1_junc RWL_13 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4741 x731/RWL0_junc x731/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4742 x585/RWL0_junc x585/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4743 x884/junc0 x884/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4744 x110/junc0 x110/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4745 x442/RWL0_junc x442/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4746 x885/junc0 x885/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4747 x989/junc0 x989/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4748 GND x1004/junc0 x1004/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4749 x988/junc0 x988/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4750 x554/junc0 x554/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4751 x782/junc1 WWL_2 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4752 GND x495/junc1 x495/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4753 GND x344/junc0 x344/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4754 GND x46/junc1 x46/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4755 GND x576/junc1 x576/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4756 x352/junc0 x352/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4757 x351/junc0 x351/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4758 GND x895/junc0 x895/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4759 WBL_31 WWL_3 x14/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4760 x831/junc0 x831/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4761 WBL_30 WWL_7 x130/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4762 RBL0_15 RWL_7 x523/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4763 RBL0_0 RWL_0 x522/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4764 x1005/junc0 x1005/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4765 WBL_22 WWL_11 x861/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4766 GND x503/junc1 x503/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4767 x1000/junc0 x1000/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4768 x975/RWL1_junc RWL_7 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4769 GND x852/junc0 x852/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4770 x974/RWL1_junc RWL_14 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4771 x393/RWL1_junc RWL_22 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4772 x459/RWL0_junc x459/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4773 x620/junc0 x620/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4774 VDD x297/junc0 x297/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4775 x233/junc0 x233/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4776 x981/junc1 WWL_30 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4777 x749/RWL1_junc RWL_12 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4778 x625/junc0 x625/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4779 x986/junc1 WWL_10 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4780 x529/junc1 WWL_27 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4781 x530/junc1 WWL_14 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4782 x626/junc0 x626/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4783 RBL0_24 RWL_11 x540/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4784 VDD x913/junc0 x913/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4785 RBL0_23 RWL_15 x245/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4786 GND x854/junc0 x854/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4787 x718/RWL1_junc RWL_18 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4788 GND x194/junc1 x194/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4789 VDD x819/junc0 x819/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4790 x159/junc0 x159/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4791 x388/junc0 x388/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4792 x892/junc0 x892/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4793 GND x856/junc0 x856/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4794 x465/junc0 x465/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4795 x992/junc0 x992/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4796 GND x1007/junc0 x1007/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4797 x993/junc0 x993/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4798 WBL_16 WWL_6 x57/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4799 WBL_7 WWL_14 x518/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4800 GND x103/junc1 x103/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4801 GND x610/junc1 x610/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4802 x473/RWL0_junc x473/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4803 x474/RWL0_junc x474/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4804 VDD x247/junc0 x247/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4805 GND x534/junc1 x534/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4806 WBL_31 WWL_4 x984/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4807 RBL0_0 RWL_1 x559/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4808 x472/junc0 x472/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4809 WBL_30 WWL_8 x175/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4810 RBL0_15 RWL_8 x560/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4811 x925/junc1 WWL_9 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4812 GND x613/junc1 x613/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4813 x276/junc0 x276/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4814 x177/junc0 x177/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4815 x689/junc0 x689/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4816 x977/RWL1_junc RWL_8 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4817 x763/RWL1_junc RWL_15 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4818 GND x409/junc0 x409/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4819 x436/RWL1_junc RWL_23 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4820 x929/junc1 WWL_17 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4821 x645/junc0 x645/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4822 x558/junc1 WWL_21 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4823 RBL0_9 RWL_14 x571/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4824 VDD x251/junc0 x251/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4825 x604/junc1 WWL_31 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4826 VDD x920/junc0 x920/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4827 RBL0_12 RWL_31 x613/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4828 x42/RWL1_junc RWL_21 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4829 x494/RWL0_junc x494/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4830 x650/junc0 x650/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4831 x991/junc1 WWL_11 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4832 VDD x921/junc0 x921/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4833 RBL0_24 RWL_12 x577/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4834 VDD x982/junc0 x982/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4835 RBL0_23 RWL_16 x35/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4836 x713/junc0 x713/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4837 RBL0_27 RWL_24 x618/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4838 x979/RWL1_junc RWL_19 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4839 x1008/junc0 x1008/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4840 x760/junc0 x760/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4841 x430/junc0 x430/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4842 WBL_3 WWL_19 x110/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4843 x431/junc0 x431/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4844 GND x869/junc0 x869/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4845 x505/RWL0_junc x505/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4846 VDD x208/junc0 x208/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4847 WBL_1 WWL_0 x988/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4848 WBL_16 WWL_7 x989/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4849 VDD x200/junc0 x200/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4850 x507/RWL0_junc x507/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4851 x54/junc1 WWL_29 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4852 x508/RWL0_junc x508/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4853 GND x871/junc0 x871/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4854 VDD x1018/junc0 x1018/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4855 GND x844/junc0 x844/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4856 WBL_27 WWL_9 x266/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4857 x213/junc0 x213/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4858 GND x570/junc1 x570/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4859 GND x572/junc1 x572/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4860 x75/RWL1_junc RWL_2 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4861 x460/RWL1_junc RWL_0 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4862 x461/RWL1_junc RWL_20 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4863 WBL_21 WWL_15 x131/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4864 x446/junc0 x446/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4865 x787/RWL1_junc RWL_16 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4866 x668/junc0 x668/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4867 x938/junc1 WWL_18 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4868 x995/junc1 WWL_14 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4869 x449/junc0 x449/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4870 RBL0_9 RWL_15 x603/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4871 GND x878/junc0 x878/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4872 x918/junc1 WWL_12 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4873 x630/junc0 x630/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4874 VDD x985/junc0 x985/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4875 GND x648/junc1 x648/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4876 x97/RWL1_junc RWL_22 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4877 x526/RWL0_junc x526/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4878 GND x187/junc1 x187/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4879 RBL0_27 RWL_25 x91/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4880 VDD x246/junc0 x246/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4881 x536/RWL0_junc x536/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4882 x519/RWL0_junc x519/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4883 WBL_12 WWL_12 x159/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4884 WBL_3 WWL_20 x892/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4885 x540/RWL0_junc x540/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4886 VDD x257/junc0 x257/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4887 WBL_16 WWL_8 x992/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4888 x1016/junc0 x1016/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4889 WBL_1 WWL_1 x993/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4890 x148/junc0 x148/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4891 x146/junc0 x146/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4892 x1019/junc0 x1019/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4893 x152/junc0 x152/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4894 GND x735/junc0 x735/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4895 x483/RWL1_junc RWL_9 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4896 GND x886/junc0 x886/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4897 GND x467/junc0 x467/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4898 x1001/junc0 x1001/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4899 GND x602/junc1 x602/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4900 VDD x838/junc0 x838/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4901 GND x605/junc1 x605/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4902 x548/RWL0_junc x548/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4903 x129/RWL1_junc RWL_3 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4904 GND x632/junc0 x632/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4905 GND x957/junc0 x957/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4906 x981/RWL1_junc RWL_30 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4907 x493/RWL1_junc RWL_1 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4908 x680/junc1 WWL_15 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4909 RBL0_28 RWL_2 x355/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4910 RBL0_20 RWL_6 x1010/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4911 VDD x429/junc0 x429/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4912 GND x639/junc1 x639/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4913 x926/junc1 WWL_19 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4914 WBL_21 WWL_16 x177/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4915 RBL0_8 RWL_31 x671/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4916 RBL0_5 RWL_20 x11/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4917 x545/junc0 x545/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4918 RBL0_9 RWL_16 x628/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4919 x542/RWL1_junc RWL_31 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4920 GND x478/junc0 x478/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4921 x176/junc1 WWL_9 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4922 x983/RWL1_junc RWL_27 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4923 x910/RWL1_junc RWL_13 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4924 x829/junc1 WWL_13 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4925 VDD x990/junc0 x990/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4926 GND x672/junc1 x672/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4927 x151/RWL1_junc RWL_23 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4928 x741/junc0 x741/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4929 GND x188/junc1 x188/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4930 x685/RWL0_junc x685/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4931 GND x226/junc1 x226/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4932 VDD x356/junc0 x356/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4933 x571/RWL0_junc x571/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4934 RBL0_27 RWL_26 x142/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4935 VDD x291/junc0 x291/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4936 VDD x445/junc0 x445/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4937 WBL_12 WWL_13 x760/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4938 x577/RWL0_junc x577/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4939 RBL0_30 RWL_24 x401/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4940 x700/junc0 x700/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4941 x917/junc0 x917/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4942 x564/junc0 x564/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4943 x296/junc0 x296/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4944 x381/junc0 x381/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4945 WBL_15 WWL_25 x96/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4946 x384/junc0 x384/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4947 x1020/junc0 x1020/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4948 x386/junc0 x386/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4949 GND x501/junc0 x501/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4950 GND x499/junc0 x499/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4951 x578/RWL1_junc RWL_0 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4952 RBL0_5 RWL_9 x644/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4953 WBL_6 WWL_19 x213/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4954 GND x627/junc1 x627/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4955 x581/RWL0_junc x581/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4956 GND x504/junc0 x504/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4957 GND x894/junc0 x894/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4958 x584/junc1 WWL_5 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4959 x583/junc1 WWL_12 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4960 x703/junc1 WWL_16 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4961 RBL0_28 x389/RWL1 x69/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4962 VDD x462/junc0 x462/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4963 GND x816/junc1 x816/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4964 x36/junc1 WWL_20 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4965 GND x498/junc1 x498/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4966 GND x899/junc1 x899/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4967 x986/RWL1_junc RWL_10 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4968 x987/RWL1_junc RWL_6 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4969 GND x636/junc1 x636/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4970 GND x510/junc0 x510/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4971 x190/RWL1_junc RWL_20 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4972 x20/junc0 x20/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4973 VDD x1/junc0 x1/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4974 GND x691/junc1 x691/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4975 WBL_8 WWL_6 x233/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4976 x565/junc0 x565/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4977 GND x271/junc1 x271/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4978 x515/junc0 x515/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4979 GND x901/junc0 x901/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4980 VDD x10/junc0 x10/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4981 x705/RWL0_junc x705/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4982 x603/RWL0_junc x603/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4983 x382/RWL0_junc x382/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4984 VDD x50/junc0 x50/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4985 VDD x268/junc0 x268/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4986 x329/junc0 x329/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4987 x686/junc0 x686/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4988 GND x525/junc0 x525/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4989 RBL0_30 RWL_25 x662/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4990 x928/junc0 x928/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4991 x776/RWL0_junc x776/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4992 x527/junc0 x527/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4993 x47/junc0 x47/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4994 x1003/junc0 x1003/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4995 GND x1009/junc0 x1009/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4996 WBL_25 WWL_6 x148/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4997 x426/junc0 x426/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M4998 WBL_15 WWL_26 x146/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M4999 WBL_0 WWL_19 x152/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5000 WBL_17 WWL_10 x1019/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5001 RBL0_1 RWL_14 x885/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5002 GND x371/junc1 x371/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5003 x611/RWL1_junc RWL_1 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5004 RBL0_14 RWL_2 x669/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5005 WBL_6 WWL_20 x1001/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5006 x615/RWL0_junc x615/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5007 x558/RWL1_junc RWL_21 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5008 WBL_23 WWL_30 x297/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5009 x223/RWL1_junc RWL_9 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5010 VDD x872/junc0 x872/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5011 GND x541/junc0 x541/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5012 x260/junc1 WWL_13 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5013 GND x234/junc1 x234/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5014 GND x532/junc1 x532/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5015 GND x908/junc1 x908/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5016 x1013/junc1 WWL_28 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5017 GND x906/junc0 x906/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5018 x991/RWL1_junc RWL_11 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5019 RBL0_19 RWL_10 x15/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5020 GND x711/junc1 x711/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5021 RBL0_18 RWL_14 x445/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5022 x78/junc0 x78/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5023 x24/junc0 x24/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5024 VDD x51/junc0 x51/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5025 WBL_8 WWL_7 x413/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5026 GND x309/junc1 x309/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5027 x804/RWL1_junc RWL_17 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5028 VDD x948/junc0 x948/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5029 GND x556/junc0 x556/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5030 x248/RWL1_junc RWL_13 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5031 VDD x64/junc0 x64/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5032 x726/RWL0_junc x726/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5033 x935/junc0 x935/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5034 x628/RWL0_junc x628/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5035 x1004/junc0 x1004/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5036 GND x1011/junc0 x1011/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5037 x221/RWL1_junc RWL_2 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5038 x706/junc0 x706/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5039 x19/junc1 WWL_2 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5040 x937/junc0 x937/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5041 RBL0_30 RWL_26 x688/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5042 x561/junc0 x561/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5043 x101/junc0 x101/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5044 x895/junc0 x895/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5045 GND x943/junc0 x943/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5046 x30/junc1 WWL_6 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5047 WBL_26 WWL_3 x296/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5048 WBL_25 WWL_7 x384/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5049 RBL0_10 RWL_7 x46/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5050 WBL_15 WWL_27 x381/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5051 WBL_0 WWL_20 x386/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5052 x104/junc0 x104/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5053 WBL_17 WWL_11 x1020/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5054 RBL0_1 RWL_15 x465/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5055 GND x1017/junc1 x1017/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5056 RBL0_14 x61/RWL1 x690/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5057 x1021/junc0 x1021/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5058 GND x789/junc0 x789/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5059 x995/RWL1_junc RWL_14 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5060 VDD x873/junc0 x873/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5061 GND x317/junc1 x317/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5062 x59/junc0 x59/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5063 x592/RWL1_junc RWL_22 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5064 WBL_23 WWL_31 x251/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5065 VDD x516/junc0 x516/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5066 GND x569/junc1 x569/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5067 x956/junc1 WWL_6 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5068 x143/junc1 WWL_10 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5069 x835/RWL1_junc RWL_12 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5070 x125/junc0 x125/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5071 x56/junc1 WWL_14 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5072 RBL0_19 RWL_11 x70/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5073 RBL0_18 RWL_15 x268/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5074 x613/junc0 x613/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5075 WBL_8 WWL_8 x452/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5076 GND x842/junc1 x842/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5077 x289/RWL1_junc RWL_10 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5078 GND x914/junc0 x914/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5079 x824/RWL1_junc RWL_18 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5080 VDD x881/junc0 x881/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5081 GND x353/junc1 x353/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5082 GND x589/junc0 x589/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5083 x412/junc0 x412/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5084 WBL_14 WWL_29 x200/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5085 x590/junc0 x590/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5086 GND x909/junc0 x909/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5087 GND x916/junc0 x916/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5088 x122/RWL0_junc x122/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5089 WBL_11 WWL_6 x329/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5090 x1007/junc0 x1007/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5091 GND x1012/junc0 x1012/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5092 x272/RWL1_junc RWL_3 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5093 WBL_2 WWL_14 x686/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5094 VDD x546/junc0 x546/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5095 x144/junc0 x144/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5096 x377/junc0 x377/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5097 x199/junc1 WWL_30 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5098 x87/junc1 WWL_7 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5099 WBL_26 WWL_4 x1003/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5100 WBL_25 WWL_8 x426/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5101 RBL0_10 RWL_8 x103/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5102 x153/junc0 x153/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5103 x263/RWL0_junc x263/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5104 RBL0_1 RWL_16 x431/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5105 x1022/junc0 x1022/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5106 GND x699/junc1 x699/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5107 x843/RWL1_junc RWL_15 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5108 x624/RWL1_junc RWL_23 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5109 x94/RWL0_junc x94/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5110 RBL0_4 RWL_14 x113/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5111 VDD x633/junc0 x633/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5112 VDD x958/junc0 x958/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5113 x669/RWL0_junc x669/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5114 x967/junc1 WWL_7 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5115 x318/RWL1_junc RWL_21 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5116 x172/junc0 x172/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5117 x196/junc1 WWL_11 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5118 VDD x936/junc0 x936/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5119 VDD x959/junc0 x959/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5120 RBL0_19 RWL_12 x719/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5121 RBL0_18 RWL_16 x217/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5122 RBL0_22 RWL_24 x745/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5123 x326/RWL1_junc RWL_11 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5124 x183/junc0 x183/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5125 x227/junc1 WWL_28 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5126 x1000/RWL1_junc RWL_19 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5127 x810/junc0 x810/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5128 x184/junc0 x184/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5129 x5/junc0 x5/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5130 GND x710/junc1 x710/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5131 x621/junc0 x621/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5132 GND x915/junc0 x915/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5133 GND x927/junc0 x927/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5134 x15/RWL0_junc x15/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5135 VDD x454/junc0 x454/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5136 WBL_11 WWL_7 x1004/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5137 x653/junc0 x653/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5138 x675/RWL0_junc x675/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5139 GND x929/junc0 x929/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5140 x747/junc0 x747/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5141 VDD x902/junc0 x902/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5142 WBL_30 WWL_5 x286/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5143 WBL_22 WWL_9 x937/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5144 GND x716/junc1 x716/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5145 GND x63/junc0 x63/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5146 x1006/junc1 WWL_31 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5147 x139/junc1 WWL_8 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5148 GND x399/junc1 x399/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5149 x463/RWL0_junc x463/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5150 x29/RWL0_junc x29/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5151 WBL_29 WWL_17 x1021/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5152 RBL0_13 RWL_21 x160/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5153 x36/RWL1_junc RWL_20 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5154 GND x720/junc1 x720/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5155 x39/RWL1_junc RWL_16 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5156 x225/junc1 WWL_14 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5157 x207/junc0 x207/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5158 x687/RWL0_junc x687/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5159 RBL0_4 RWL_15 x162/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5160 GND x931/junc0 x931/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5161 x750/junc0 x750/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5162 x155/junc1 WWL_12 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5163 VDD x596/junc0 x596/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5164 WBL_20 WWL_29 x278/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5165 x118/junc0 x118/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5166 GND x762/junc1 x762/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5167 x690/RWL0_junc x690/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5168 x971/junc1 WWL_8 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5169 x361/RWL1_junc RWL_22 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5170 VDD x443/junc0 x443/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5171 RBL0_31 RWL_17 x858/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5172 GND x212/junc1 x212/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5173 RBL0_22 RWL_25 x354/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5174 x640/junc0 x640/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5175 x367/RWL1_junc RWL_12 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5176 VDD x96/junc0 x96/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5177 x950/junc0 x950/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5178 WBL_7 WWL_12 x412/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5179 GND x731/junc1 x731/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5180 x70/RWL0_junc x70/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5181 VDD x481/junc0 x481/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5182 WBL_11 WWL_8 x1007/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5183 x1010/junc0 x1010/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5184 x676/junc0 x676/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5185 x140/junc0 x140/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5186 GND x938/junc0 x938/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5187 x76/RWL1_junc RWL_9 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5188 WBL_31 WWL_2 x377/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5189 VDD x1005/junc0 x1005/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5190 GND x737/junc1 x737/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5191 x85/RWL0_junc x85/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5192 x86/RWL0_junc x86/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5193 x768/RWL1_junc RWL_30 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5194 GND x982/junc0 x982/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5195 x191/junc1 WWL_14 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5196 VDD x620/junc0 x620/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5197 RBL0_13 RWL_22 x204/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5198 x195/junc1 WWL_19 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5199 WBL_29 WWL_18 x1022/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5200 x795/junc1 WWL_15 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5201 RBL0_23 RWL_2 x567/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5202 GND x723/junc1 x723/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5203 x194/RWL0_junc x194/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5204 GND x743/junc1 x743/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5205 x256/junc0 x256/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5206 x496/junc0 x496/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5207 x708/RWL0_junc x708/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5208 RBL0_4 RWL_16 x748/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5209 GND x939/junc0 x939/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5210 GND x655/junc0 x655/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5211 VDD x625/junc0 x625/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5212 x427/junc1 WWL_9 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5213 x792/junc0 x792/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5214 x201/junc1 WWL_13 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5215 VDD x626/junc0 x626/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5216 GND x524/junc1 x524/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5217 x953/junc0 x953/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5218 x182/junc0 x182/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5219 GND x2/junc1 x2/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5220 x180/junc0 x180/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5221 x406/RWL1_junc RWL_23 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5222 x58/junc0 x58/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5223 RBL0_30 RWL_28 x117/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5224 x865/RWL0_junc x865/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5225 VDD x568/junc0 x568/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5226 VDD x33/junc0 x33/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5227 GND x441/junc1 x441/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5228 RBL0_31 RWL_18 x870/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5229 x113/RWL0_junc x113/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5230 RBL0_22 RWL_26 x311/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5231 GND x203/junc0 x203/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5232 WBL_16 WWL_5 x448/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5233 x1013/RWL1_junc RWL_28 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5234 WBL_7 WWL_13 x5/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5235 x124/RWL0_junc x124/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5236 x719/RWL0_junc x719/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5237 RBL0_25 RWL_24 x597/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5238 x283/junc0 x283/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5239 x955/junc0 x955/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5240 x511/junc0 x511/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5241 x588/junc0 x588/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5242 x586/junc0 x586/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5243 WBL_10 WWL_25 x90/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5244 x128/RWL1_junc RWL_2 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5245 GND x674/junc0 x674/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5246 x422/RWL1_junc RWL_0 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5247 WBL_14 WWL_21 x747/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5248 VDD x472/junc0 x472/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5249 x84/junc0 x84/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5250 GND x32/junc1 x32/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5251 RBL0_3 RWL_28 x53/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5252 x722/RWL0_junc x722/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5253 VDD x145/junc0 x145/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5254 x724/RWL0_junc x724/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5255 GND x941/junc0 x941/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5256 WBL_6 WWL_28 x485/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5257 GND x942/junc0 x942/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5258 VDD x62/junc0 x62/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5259 x725/junc1 WWL_12 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5260 RBL0_13 RWL_23 x252/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5261 x808/junc1 WWL_16 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5262 RBL0_23 x61/RWL1 x335/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5263 VDD x645/junc0 x645/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5264 x241/junc1 WWL_20 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5265 GND x45/junc1 x45/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5266 x143/RWL1_junc RWL_10 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5267 x537/RWL1_junc RWL_30 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5268 x528/junc0 x528/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5269 GND x944/junc0 x944/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5270 x148/RWL1_junc RWL_6 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5271 GND x677/junc0 x677/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5272 RBL0_16 RWL_21 x884/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5273 x439/RWL1_junc RWL_20 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5274 x298/junc0 x298/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5275 VDD x650/junc0 x650/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5276 x679/junc0 x679/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5277 GND x52/junc1 x52/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5278 x794/junc0 x794/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5279 GND x55/junc1 x55/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5280 x681/junc0 x681/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5281 WBL_3 WWL_6 x118/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5282 x961/junc0 x961/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5283 GND x494/junc1 x494/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5284 x683/junc0 x683/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5285 RBL0_26 RWL_30 x164/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5286 GND x1014/junc0 x1014/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5287 x161/RWL0_junc x161/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5288 x876/RWL0_junc x876/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5289 RBL0_30 RWL_29 x739/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5290 VDD x294/junc0 x294/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5291 VDD x1008/junc0 x1008/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5292 RBL0_31 RWL_19 x352/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5293 x162/RWL0_junc x162/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5294 x543/junc0 x543/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5295 GND x174/junc0 x174/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5296 GND x250/junc0 x250/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5297 x883/RWL1_junc RWL_29 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5298 x169/RWL0_junc x169/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5299 GND x475/junc1 x475/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5300 RBL0_25 RWL_25 x279/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5301 x322/junc0 x322/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5302 x964/junc0 x964/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5303 GND x945/junc0 x945/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5304 x87/RWL1_junc RWL_7 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5305 x1009/junc0 x1009/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5306 x617/junc0 x617/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5307 WBL_10 WWL_26 x140/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5308 x61/RWL1_junc x61/RWL1 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5309 x459/RWL1_junc RWL_1 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5310 RBL0_9 RWL_2 x782/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5311 RBL0_3 RWL_29 x713/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5312 x557/junc0 x557/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5313 RBL0_28 RWL_0 x625/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5314 RBL0_20 RWL_4 x371/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5315 WBL_2 WWL_30 x516/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5316 x464/RWL1_junc RWL_9 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5317 GND x946/junc0 x946/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5318 GND x698/junc0 x698/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5319 VDD x668/junc0 x668/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5320 x486/junc1 WWL_13 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5321 GND x99/junc1 x99/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5322 x830/junc1 WWL_25 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5323 GND x947/junc0 x947/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5324 x196/RWL1_junc RWL_11 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5325 x608/junc0 x608/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5326 WBL_28 WWL_22 x496/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5327 GND x812/junc1 x812/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5328 GND x4/junc0 x4/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5329 GND x0/junc0 x0/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5330 RBL0_16 RWL_22 x388/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5331 x340/junc0 x340/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5332 x887/RWL0_junc x887/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5333 x702/junc0 x702/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5334 GND x108/junc1 x108/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5335 x807/junc0 x807/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5336 WBL_3 WWL_7 x953/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5337 GND x526/junc1 x526/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5338 VDD x575/junc0 x575/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5339 VDD x978/junc0 x978/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5340 x495/junc0 x495/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5341 GND x707/junc0 x707/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5342 x206/RWL0_junc x206/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5343 VDD x332/junc0 x332/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5344 x484/RWL0_junc x484/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5345 x969/junc0 x969/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5346 x748/RWL0_junc x748/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5347 x1011/junc0 x1011/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5348 x639/RWL0_junc x639/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5349 GND x519/junc1 x519/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5350 GND x346/junc1 x346/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5351 x134/junc0 x134/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5352 GND x491/junc1 x491/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5353 RBL0_25 RWL_26 x798/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5354 x712/junc0 x712/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5355 GND x951/junc0 x951/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5356 x139/RWL1_junc RWL_8 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5357 x364/junc0 x364/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5358 x943/junc0 x943/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5359 x304/junc1 WWL_6 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5360 WBL_21 WWL_3 x511/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5361 RBL0_5 RWL_7 x321/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5362 WBL_10 WWL_27 x586/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5363 x973/RWL0_junc x973/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5364 RBL0_9 x61/RWL1 x800/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5365 x814/junc0 x814/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5366 GND x165/junc0 x165/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5367 x225/RWL1_junc RWL_14 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5368 x316/junc1 WWL_0 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5369 x820/junc0 x820/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5370 WBL_13 WWL_25 x520/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5371 RBL0_28 RWL_1 x650/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5372 RBL0_20 RWL_5 x1017/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5373 VDD x930/junc0 x930/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5374 GND x533/junc1 x533/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5375 WBL_2 WWL_31 x633/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5376 GND x48/junc0 x48/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5377 VDD x545/junc0 x545/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5378 WBL_29 WWL_30 x936/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5379 GND x50/junc0 x50/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5380 x236/RWL1_junc RWL_4 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5381 x327/junc1 WWL_26 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5382 VDD x600/junc0 x600/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5383 VDD x598/junc0 x598/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5384 x240/RWL1_junc RWL_12 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5385 WBL_28 WWL_23 x528/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5386 RBL0_27 RWL_13 x336/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5387 x378/junc0 x378/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5388 RBL0_12 RWL_27 x1008/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5389 VDD x689/junc0 x689/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5390 GND x54/junc0 x54/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5391 x72/junc0 x72/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5392 RBL0_16 RWL_23 x430/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5393 x383/junc0 x383/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5394 WBL_12 WWL_0 x794/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5395 WBL_3 WWL_8 x961/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5396 x505/RWL1_junc RWL_10 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5397 GND x65/junc0 x65/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5398 x391/junc0 x391/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5399 VDD x695/junc0 x695/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5400 x657/junc0 x657/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5401 VDD x934/junc0 x934/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5402 x658/junc0 x658/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5403 GND x729/junc0 x729/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5404 x610/junc0 x610/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5405 x730/junc0 x730/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5406 GND x954/junc0 x954/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5407 WBL_6 WWL_6 x543/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5408 x1012/junc0 x1012/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5409 x212/junc0 x212/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5410 GND x170/junc1 x170/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5411 x899/RWL0_junc x899/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5412 x752/junc0 x752/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5413 VDD x564/junc0 x564/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5414 VDD x700/junc0 x700/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5415 x403/junc0 x403/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5416 x255/junc0 x255/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5417 x344/junc1 WWL_3 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5418 RBL0_14 RWL_0 x362/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5419 x347/junc1 WWL_7 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5420 WBL_21 WWL_4 x1009/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5421 RBL0_5 RWL_8 x365/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5422 x487/RWL0_junc x487/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5423 x999/RWL0_junc x999/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5424 x443/junc0 x443/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5425 x826/junc0 x826/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5426 x523/RWL1_junc RWL_7 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5427 GND x805/junc1 x805/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5428 x360/junc1 WWL_1 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5429 WBL_13 WWL_26 x557/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5430 x275/RWL1_junc RWL_15 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5431 x280/RWL0_junc x280/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5432 RBL0_0 RWL_28 x288/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5433 WBL_29 WWL_31 x443/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5434 GND x107/junc0 x107/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5435 x782/RWL0_junc x782/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5436 x286/RWL1_junc RWL_5 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5437 VDD x21/junc0 x21/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5438 x368/junc1 WWL_27 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5439 WBL_28 WWL_24 x608/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5440 VDD x18/junc0 x18/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5441 x423/junc0 x423/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5442 VDD x216/junc0 x216/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5443 WBL_8 WWL_5 x256/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5444 x932/RWL0_junc x932/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5445 WBL_12 WWL_1 x807/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5446 RBL0_17 RWL_24 x1016/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5447 GND x962/junc0 x962/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5448 x540/RWL1_junc RWL_11 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5449 x564/junc1 WWL_25 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5450 x26/junc0 x26/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5451 x27/junc0 x27/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5452 x874/junc0 x874/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5453 x435/junc0 x435/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5454 WBL_0 WWL_6 x495/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5455 x678/junc0 x678/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5456 x680/junc0 x680/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5457 x522/RWL1_junc RWL_0 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5458 x292/junc0 x292/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5459 x509/RWL0_junc x509/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5460 x746/junc0 x746/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5461 GND x963/junc0 x963/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5462 x441/junc0 x441/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5463 VDD x635/junc0 x635/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5464 WBL_6 WWL_7 x1011/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5465 x402/junc0 x402/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5466 x908/RWL0_junc x908/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5467 x791/RWL0_junc x791/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5468 GND x965/junc0 x965/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5469 WBL_26 WWL_29 x773/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5470 x832/junc0 x832/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5471 VDD x23/junc0 x23/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5472 WBL_25 WWL_5 x503/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5473 WBL_17 WWL_9 x134/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5474 GND x818/junc1 x818/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5475 GND x138/junc0 x138/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5476 x457/junc1 WWL_0 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5477 RBL0_14 RWL_1 x408/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5478 x397/junc1 WWL_4 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5479 x398/junc1 WWL_8 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5480 x28/RWL0_junc x28/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5481 GND x594/junc1 x594/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5482 GND x967/junc0 x967/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5483 VDD x382/junc0 x382/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5484 WBL_24 WWL_17 x814/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5485 GND x839/junc1 x839/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5486 x770/junc1 WWL_30 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5487 RBL0_8 RWL_21 x411/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5488 x241/RWL1_junc RWL_20 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5489 GND x229/junc1 x229/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5490 x560/RWL1_junc RWL_8 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5491 WBL_13 WWL_27 x820/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5492 x312/RWL1_junc RWL_16 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5493 x40/RWL0_junc x40/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5494 x149/junc0 x149/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5495 x836/junc0 x836/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5496 RBL0_0 RWL_29 x801/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5497 x837/junc0 x837/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5498 GND x266/junc0 x266/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5499 x409/junc1 WWL_12 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5500 GND x158/junc0 x158/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5501 x800/RWL0_junc x800/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5502 x850/junc0 x850/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5503 RBL0_26 RWL_17 x917/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5504 RBL0_17 RWL_25 x564/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5505 x756/junc0 x756/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5506 x577/RWL1_junc RWL_12 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5507 x527/junc1 WWL_26 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5508 x81/junc0 x81/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5509 x980/junc0 x980/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5510 RBL0_30 RWL_13 x829/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5511 WBL_15 WWL_14 x657/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5512 x559/RWL1_junc RWL_1 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5513 WBL_0 WWL_7 x658/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5514 RBL0_1 RWL_2 x180/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5515 WBL_2 WWL_12 x610/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5516 x544/RWL0_junc x544/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5517 x618/RWL1_junc RWL_24 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5518 VDD x741/junc0 x741/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5519 VDD x949/junc0 x949/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5520 VDD x92/junc0 x92/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5521 WBL_6 WWL_8 x1012/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5522 x387/junc0 x387/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5523 x605/junc0 x605/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5524 GND x179/junc0 x179/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5525 GND x970/junc0 x970/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5526 x869/junc1 WWL_5 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5527 x338/RWL1_junc RWL_9 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5528 WBL_26 WWL_2 x255/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5529 VDD x104/junc0 x104/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5530 GND x849/junc1 x849/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5531 GND x827/junc1 x827/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5532 x38/junc1 WWL_1 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5533 GND x270/junc1 x270/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5534 x407/junc0 x407/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5535 x82/RWL0_junc x82/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5536 WBL_20 WWL_22 x322/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5537 GND x971/junc0 x971/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5538 VDD x425/junc0 x425/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5539 GND x851/junc1 x851/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5540 x654/junc1 WWL_31 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5541 RBL0_8 RWL_22 x450/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5542 WBL_24 WWL_18 x826/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5543 RBL0_18 RWL_2 x20/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5544 x353/RWL0_junc x353/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5545 GND x282/junc1 x282/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5546 x672/junc0 x672/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5547 x13/RWL1_junc RWL_28 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5548 x93/RWL0_junc x93/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5549 x136/RWL0_junc x136/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5550 GND x198/junc0 x198/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5551 x362/RWL0_junc x362/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5552 x846/junc0 x846/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5553 x1002/junc1 WWL_5 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5554 VDD x125/junc0 x125/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5555 x619/junc1 WWL_9 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5556 GND x642/junc1 x642/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5557 x447/junc1 WWL_13 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5558 x434/junc0 x434/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5559 RBL0_9 RWL_28 x372/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5560 x66/junc1 WWL_17 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5561 x130/junc0 x130/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5562 x861/junc0 x861/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5563 VDD x715/junc0 x715/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5564 VDD x994/junc0 x994/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5565 RBL0_26 RWL_18 x928/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5566 RBL0_17 RWL_26 x527/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5567 x697/junc1 WWL_29 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5568 x563/junc1 WWL_27 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5569 WBL_11 WWL_5 x631/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5570 WBL_0 WWL_8 x678/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5571 x466/RWL1_junc RWL_21 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5572 RBL0_1 RWL_3 x681/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5573 VDD x385/junc0 x385/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5574 x91/RWL1_junc RWL_25 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5575 WBL_2 WWL_13 x292/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5576 x376/RWL0_junc x376/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5577 VDD x144/junc0 x144/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5578 x627/junc0 x627/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5579 GND x776/junc0 x776/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5580 x727/junc0 x727/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5581 WBL_5 WWL_25 x572/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5582 GND x220/junc0 x220/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5583 x380/RWL1_junc RWL_2 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5584 GND x785/junc0 x785/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5585 WBL_9 WWL_21 x832/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5586 VDD x153/junc0 x153/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5587 GND x859/junc1 x859/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5588 x346/junc0 x346/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5589 GND x306/junc1 x306/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5590 WBL_29 WWL_15 x363/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5591 x137/RWL0_junc x137/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5592 x244/junc0 x244/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5593 WBL_20 WWL_23 x364/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5594 GND x232/junc0 x232/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5595 VDD x331/junc0 x331/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5596 x825/junc1 WWL_12 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5597 RBL0_8 RWL_23 x476/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5598 RBL0_18 x61/RWL1 x78/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5599 x141/RWL0_junc x141/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5600 x67/RWL1_junc RWL_30 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5601 x691/junc0 x691/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5602 x697/RWL1_junc RWL_29 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5603 GND x94/junc1 x94/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5604 x1010/RWL1_junc RWL_6 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5605 GND x245/junc0 x245/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5606 x408/RWL0_junc x408/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5607 RBL0_11 RWL_21 x935/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5608 x11/RWL1_junc RWL_20 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5609 x518/junc0 x518/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5610 VDD x172/junc0 x172/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5611 x857/junc0 x857/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5612 GND x328/junc1 x328/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5613 GND x932/junc0 x932/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5614 x478/junc1 WWL_22 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5615 RBL0_5 RWL_30 x416/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5616 x456/RWL0_junc x456/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5617 x822/junc0 x822/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5618 x489/RWL1_junc RWL_24 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5619 x984/junc0 x984/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5620 RBL0_9 RWL_29 x828/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5621 x119/junc1 WWL_18 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5622 x175/junc0 x175/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5623 VDD x997/junc0 x997/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5624 x797/junc0 x797/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5625 VDD x184/junc0 x184/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5626 RBL0_26 RWL_19 x561/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5627 x475/junc0 x475/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5628 x496/RWL1_junc RWL_22 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5629 VDD x428/junc0 x428/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5630 x142/RWL1_junc RWL_26 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5631 x420/RWL0_junc x420/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5632 x347/RWL1_junc RWL_7 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5633 x866/junc0 x866/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5634 VDD x891/junc0 x891/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5635 WBL_5 WWL_26 x605/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5636 GND x666/junc1 x666/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5637 GND x9/junc0 x9/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5638 x424/RWL1_junc x61/RWL1 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5639 GND x265/junc0 x265/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5640 RBL0_4 RWL_2 x19/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5641 x176/RWL0_junc x176/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5642 GND x345/junc1 x345/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5643 x105/RWL1_junc RWL_28 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5644 x506/junc0 x506/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5645 x499/junc1 WWL_12 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5646 x908/junc0 x908/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5647 GND x463/junc1 x463/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5648 RBL0_13 RWL_20 x508/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5649 GND x29/junc1 x29/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5650 WBL_29 WWL_16 x407/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5651 RBL0_23 RWL_0 x125/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5652 WBL_20 WWL_24 x734/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5653 GND x285/junc0 x285/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5654 x644/RWL1_junc RWL_9 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5655 VDD x207/junc0 x207/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5656 x3/RWL0_junc x3/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5657 x660/junc1 WWL_13 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5658 WBL_12 WWL_28 x689/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5659 VDD x875/junc0 x875/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5660 x894/junc1 WWL_25 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5661 GND x290/junc0 x290/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5662 x740/junc0 x740/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5663 GND x687/junc1 x687/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5664 WBL_23 WWL_22 x672/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5665 x733/junc1 WWL_29 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5666 x989/junc0 x989/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5667 x160/junc1 WWL_21 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5668 GND x877/junc1 x877/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5669 GND x35/junc0 x35/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5670 x988/junc0 x988/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5671 x554/junc0 x554/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5672 RBL0_11 RWL_22 x590/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5673 x197/RWL0_junc x197/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5674 GND x369/junc1 x369/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5675 x7/junc0 x7/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5676 x510/junc1 WWL_23 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5677 VDD x219/junc0 x219/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5678 x520/RWL1_junc RWL_25 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5679 x831/junc0 x831/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5680 VDD x41/junc0 x41/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5681 x491/junc0 x491/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5682 GND x122/junc0 x122/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5683 x723/RWL0_junc x723/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5684 x528/RWL1_junc RWL_23 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5685 x457/RWL1_junc RWL_0 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5686 x398/RWL1_junc RWL_8 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5687 RBL0_13 RWL_9 x536/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5688 WBL_14 WWL_19 x627/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5689 x525/junc1 WWL_6 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5690 GND x389/junc1 x389/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5691 GND x297/junc0 x297/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5692 WBL_5 WWL_27 x727/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5693 x524/RWL0_junc x524/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5694 GND x302/junc0 x302/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5695 GND x565/junc1 x565/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5696 RBL0_4 RWL_3 x867/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5697 x733/RWL1_junc RWL_29 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5698 GND x59/junc1 x59/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5699 x879/junc0 x879/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5700 x607/junc0 x607/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5701 GND x315/junc0 x315/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5702 x192/junc1 WWL_0 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5703 x882/junc0 x882/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5704 GND x85/junc1 x85/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5705 x535/junc1 WWL_13 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5706 RBL0_23 RWL_1 x172/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5707 VDD x966/junc0 x966/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5708 GND x693/junc1 x693/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5709 GND x86/junc1 x86/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5710 GND x323/junc0 x323/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5711 VDD x256/junc0 x256/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5712 x471/RWL1_junc RWL_4 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5713 WBL_8 WWL_30 x709/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5714 x541/junc1 WWL_26 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5715 VDD x259/junc0 x259/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5716 GND x708/junc1 x708/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5717 WBL_23 WWL_23 x691/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5718 x892/junc0 x892/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5719 RBL0_22 RWL_13 x810/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5720 RBL0_7 RWL_27 x184/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5721 x992/junc0 x992/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5722 x993/junc0 x993/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5723 RBL0_11 RWL_23 x621/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5724 x587/junc0 x587/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5725 WBL_7 WWL_0 x857/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5726 RBL0_0 RWL_24 x778/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5727 x549/junc1 WWL_24 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5728 VDD x267/junc0 x267/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5729 x557/RWL1_junc RWL_26 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5730 x772/junc0 x772/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5731 x770/RWL1_junc RWL_30 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5732 GND x102/junc0 x102/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5733 GND x865/junc1 x865/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5734 GND x421/junc1 x421/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5735 x482/RWL0_junc x482/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5736 x45/RWL0_junc x45/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5737 x556/junc1 WWL_22 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5738 VDD x283/junc0 x283/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5739 x276/junc0 x276/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5740 x260/RWL0_junc x260/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5741 x479/junc0 x479/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5742 x258/RWL0_junc x258/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5743 RBL0_18 RWL_30 x704/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5744 x38/RWL1_junc RWL_1 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5745 x902/junc1 WWL_3 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5746 RBL0_9 RWL_0 x573/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5747 x224/junc1 WWL_7 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5748 WBL_14 WWL_20 x866/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5749 x608/junc0 x608/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5750 x52/RWL0_junc x52/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5751 GND x25/junc1 x25/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5752 x889/junc0 x889/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5753 GND x704/junc1 x704/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5754 GND x115/junc1 x115/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5755 x890/junc0 x890/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5756 GND x355/junc0 x355/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5757 x46/RWL1_junc RWL_7 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5758 x235/junc1 WWL_1 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5759 VDD x8/junc0 x8/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5760 GND x714/junc1 x714/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5761 x925/junc0 x925/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5762 GND x722/junc1 x722/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5763 GND x724/junc1 x724/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5764 x277/RWL0_junc x277/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5765 RBL0_27 RWL_10 x580/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5766 WBL_8 WWL_31 x671/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5767 x107/junc0 x107/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5768 x19/RWL0_junc x19/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5769 x503/RWL1_junc RWL_5 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5770 RBL0_31 RWL_6 x640/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5771 x249/junc1 WWL_27 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5772 VDD x299/junc0 x299/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5773 VDD x298/junc0 x298/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5774 WBL_23 WWL_24 x740/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5775 RBL0_16 RWL_20 x950/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5776 WBL_3 WWL_5 x480/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5777 VDD x749/junc0 x749/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5778 WBL_7 WWL_1 x7/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5779 GND x456/junc0 x456/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5780 x563/RWL1_junc RWL_27 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5781 GND x1018/junc0 x1018/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5782 RBL0_0 RWL_25 x591/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5783 x301/junc0 x301/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5784 x795/junc0 x795/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5785 WBL_25 WWL_28 x741/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5786 GND x876/junc1 x876/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5787 VDD x803/junc0 x803/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5788 x513/RWL0_junc x513/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5789 x99/RWL0_junc x99/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5790 x589/junc1 WWL_23 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5791 x896/junc0 x896/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5792 GND x396/junc0 x396/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5793 x271/junc1 WWL_0 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5794 RBL0_9 RWL_1 x606/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5795 x1005/junc1 WWL_4 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5796 x274/junc1 WWL_8 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5797 x156/junc0 x156/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5798 x303/RWL0_junc x303/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5799 GND x732/junc1 x732/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5800 x630/junc0 x630/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5801 x108/RWL0_junc x108/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5802 GND x985/junc0 x985/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5803 x898/junc0 x898/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5804 WBL_19 WWL_17 x879/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5805 GND x69/junc0 x69/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5806 GND x903/junc1 x903/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5807 RBL0_3 RWL_21 x792/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5808 x634/junc0 x634/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5809 x103/RWL1_junc RWL_8 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5810 RBL0_16 RWL_9 x182/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5811 GND x468/junc1 x468/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5812 GND x3/junc0 x3/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5813 x313/RWL0_junc x313/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5814 x314/RWL0_junc x314/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5815 RBL0_27 RWL_11 x614/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5816 GND x937/junc0 x937/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5817 x867/RWL0_junc x867/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5818 VDD x340/junc0 x340/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5819 GND x257/junc0 x257/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5820 x1019/junc0 x1019/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5821 RBL0_21 RWL_17 x955/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5822 VDD x767/junc0 x767/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5823 x585/junc0 x585/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5824 GND x887/junc1 x887/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5825 x228/junc0 x228/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5826 RBL0_25 RWL_13 x201/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5827 RBL0_0 RWL_26 x893/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5828 x1001/junc0 x1001/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5829 WBL_10 WWL_14 x772/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5830 GND x888/junc1 x888/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5831 x745/RWL1_junc RWL_24 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5832 GND x484/junc1 x484/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5833 VDD x58/junc0 x58/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5834 VDD x823/junc0 x823/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5835 VDD x979/junc0 x979/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5836 x243/junc1 WWL_28 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5837 x868/RWL0_junc x868/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5838 x618/junc1 WWL_24 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5839 GND x429/junc0 x429/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5840 x904/junc0 x904/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5841 x927/junc1 WWL_5 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5842 WBL_21 WWL_2 x479/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5843 GND x112/junc0 x112/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5844 GND x793/junc1 x793/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5845 GND x663/junc1 x663/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5846 x199/junc0 x199/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5847 x309/junc1 WWL_1 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5848 x743/junc0 x743/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5849 x652/junc0 x652/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5850 x342/RWL0_junc x342/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5851 GND x990/junc0 x990/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5852 WBL_28 WWL_10 x889/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5853 x318/junc1 WWL_21 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5854 WBL_19 WWL_18 x890/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5855 RBL0_12 RWL_14 x298/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5856 GND x911/junc1 x911/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5857 RBL0_3 RWL_22 x679/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5858 x656/junc0 x656/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5859 x563/RWL0_junc x563/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5860 VDD x84/junc0 x84/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5861 x2/junc0 x2/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5862 x357/RWL0_junc x357/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5863 x358/RWL0_junc x358/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5864 x263/junc1 WWL_30 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5865 x570/RWL1_junc RWL_17 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5866 GND x445/junc0 x445/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5867 x573/RWL0_junc x573/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5868 VDD x378/junc0 x378/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5869 VDD x786/junc0 x786/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5870 RBL0_27 RWL_12 x637/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5871 VDD x787/junc0 x787/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5872 x623/junc0 x623/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5873 RBL0_30 RWL_10 x641/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5874 x381/junc0 x381/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5875 VDD x391/junc0 x391/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5876 x333/junc1 WWL_17 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5877 x384/junc0 x384/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5878 x1020/junc0 x1020/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5879 VDD x817/junc0 x817/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5880 x386/junc0 x386/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5881 RBL0_21 RWL_18 x964/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5882 x264/junc0 x264/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5883 WBL_6 WWL_5 x751/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5884 GND x514/junc1 x514/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5885 x648/RWL1_junc RWL_21 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5886 x354/RWL1_junc RWL_25 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5887 x582/RWL0_junc x582/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5888 VDD x403/junc0 x403/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5889 VDD x1016/junc0 x1016/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5890 x32/junc0 x32/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5891 GND x462/junc0 x462/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5892 x187/RWL1_junc RWL_2 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5893 x912/junc0 x912/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5894 x646/junc1 WWL_2 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5895 VDD x593/junc0 x593/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5896 WBL_4 WWL_21 x896/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5897 GND x806/junc1 x806/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5898 x1006/junc0 x1006/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5899 WBL_24 WWL_15 x720/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5900 x395/RWL0_junc x395/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5901 GND x1/junc0 x1/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5902 x359/junc1 WWL_14 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5903 VDD x129/junc0 x129/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5904 WBL_28 WWL_11 x898/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5905 x565/junc0 x565/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5906 RBL0_12 RWL_15 x340/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5907 RBL0_3 RWL_23 x702/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5908 WBL_18 WWL_29 x875/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5909 x400/RWL0_junc x400/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5910 x55/junc0 x55/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5911 x404/RWL0_junc x404/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5912 GND x10/junc0 x10/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5913 VDD x136/junc0 x136/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5914 GND x280/junc1 x280/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5915 x542/junc1 WWL_31 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5916 x602/RWL1_junc RWL_18 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5917 GND x268/junc0 x268/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5918 x417/junc0 x417/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5919 x606/RWL0_junc x606/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5920 RBL0_6 RWL_21 x969/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5921 x686/junc0 x686/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5922 VDD x423/junc0 x423/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5923 x60/junc0 x60/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5924 x655/junc1 WWL_22 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5925 x883/junc0 x883/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5926 x639/RWL1_junc RWL_24 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5927 x1003/junc0 x1003/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5928 RBL0_30 RWL_11 x665/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5929 x374/junc1 WWL_18 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5930 x594/RWL0_junc x594/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5931 x426/junc0 x426/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5932 x862/junc0 x862/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5933 VDD x435/junc0 x435/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5934 RBL0_21 RWL_19 x712/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5935 WBL_15 WWL_12 x585/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5936 RBL0_1 RWL_0 x988/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5937 WBL_0 WWL_5 x731/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5938 RBL0_15 RWL_28 x203/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5939 GND x776/junc1 x776/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5940 x672/RWL1_junc RWL_22 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5941 x311/RWL1_junc RWL_26 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5942 x616/RWL0_junc x616/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5943 x224/RWL1_junc RWL_7 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5944 x89/junc0 x89/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5945 VDD x940/junc0 x940/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5946 GND x16/junc1 x16/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5947 GND x202/junc0 x202/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5948 x226/RWL1_junc RWL_3 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5949 WBL_13 WWL_14 x904/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5950 GND x193/junc1 x193/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5951 x427/RWL0_junc x427/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5952 GND x22/junc1 x22/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5953 RBL0_18 RWL_0 x378/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5954 GND x28/junc1 x28/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5955 RBL0_8 RWL_20 x17/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5956 WBL_24 WWL_16 x743/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5957 GND x502/junc0 x502/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5958 x24/junc0 x24/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5959 GND x51/junc0 x51/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5960 x25/junc0 x25/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5961 RBL0_12 RWL_16 x383/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5962 VDD x453/junc0 x453/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5963 x108/junc0 x108/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5964 x942/junc1 WWL_25 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5965 x109/junc0 x109/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5966 GND x40/junc1 x40/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5967 WBL_18 WWL_22 x2/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5968 GND x64/junc0 x64/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5969 GND x932/junc1 x932/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5970 x627/RWL1_junc RWL_19 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5971 x1004/junc0 x1004/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5972 x411/junc1 WWL_21 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5973 GND x217/junc0 x217/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5974 RBL0_6 RWL_22 x730/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5975 x706/junc0 x706/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5976 x444/RWL0_junc x444/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5977 x116/junc0 x116/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5978 VDD x987/junc0 x987/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5979 x944/junc1 WWL_15 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5980 x677/junc1 WWL_23 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5981 VDD x80/junc0 x80/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5982 x899/RWL1_junc RWL_25 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5983 x243/RWL1_junc RWL_28 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5984 x895/junc0 x895/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5985 RBL0_30 RWL_12 x918/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5986 WBL_15 WWL_13 x264/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5987 RBL0_1 RWL_1 x993/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5988 x636/RWL1_junc RWL_27 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5989 x1021/junc0 x1021/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5990 RBL0_15 RWL_29 x250/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5991 x670/junc0 x670/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M5992 x691/RWL1_junc RWL_23 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5993 x59/junc0 x59/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5994 x271/RWL1_junc RWL_0 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5995 x274/RWL1_junc RWL_8 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5996 RBL0_8 RWL_9 x694/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5997 WBL_9 WWL_19 x32/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5998 GND x516/junc0 x516/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M5999 GND x74/junc1 x74/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6000 x642/RWL0_junc x642/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6001 GND x239/junc1 x239/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6002 x440/junc1 WWL_0 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6003 GND x83/junc1 x83/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6004 GND x82/junc1 x82/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6005 RBL0_18 RWL_1 x423/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6006 GND x110/junc0 x110/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6007 VDD x480/junc0 x480/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6008 x371/RWL1_junc RWL_4 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6009 x698/junc1 WWL_26 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6010 VDD x120/junc0 x120/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6011 RBL0_2 RWL_27 x435/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6012 GND x93/junc1 x93/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6013 WBL_18 WWL_23 x55/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6014 RBL0_17 RWL_13 x874/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6015 x758/junc1 WWL_14 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6016 x1007/junc0 x1007/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6017 RBL0_6 RWL_23 x746/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6018 x728/junc0 x728/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6019 VDD x234/junc0 x234/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6020 GND x546/junc0 x546/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6021 WBL_2 WWL_0 x60/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6022 VDD x130/junc0 x130/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6023 x4/junc1 WWL_16 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6024 GND x813/junc1 x813/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6025 x170/junc0 x170/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6026 x12/junc1 WWL_24 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6027 VDD x131/junc0 x131/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6028 GND x122/junc1 x122/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6029 x908/RWL1_junc RWL_26 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6030 x171/junc0 x171/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6031 GND x284/junc0 x284/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6032 x287/RWL1_junc RWL_29 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6033 GND x114/junc1 x114/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6034 x711/RWL1_junc RWL_20 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6035 x1022/junc0 x1022/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6036 x659/RWL0_junc x659/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6037 x707/junc1 WWL_22 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6038 x1023/junc0 x1023/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6039 x486/RWL0_junc x486/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6040 WBL_20 WWL_10 x840/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6041 GND x121/junc1 x121/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6042 x278/junc0 x278/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6043 x309/RWL1_junc RWL_1 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6044 x115/junc0 x115/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6045 RBL0_4 RWL_0 x717/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6046 x492/RWL0_junc x492/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6047 WBL_9 WWL_20 x89/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6048 x740/junc0 x740/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6049 x328/RWL0_junc x328/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6050 x443/RWL1_junc RWL_31 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6051 x189/junc0 x189/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6052 RBL0_28 RWL_28 x809/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6053 GND x567/junc0 x567/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6054 GND x936/junc0 x936/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6055 x321/RWL1_junc RWL_7 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6056 x470/junc1 WWL_1 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6057 VDD x293/junc0 x293/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6058 GND x133/junc1 x133/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6059 GND x137/junc1 x137/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6060 GND x135/junc1 x135/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6061 GND x809/junc1 x809/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6062 RBL0_22 RWL_10 x850/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6063 GND x41/junc0 x41/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6064 GND x141/junc1 x141/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6065 VDD x517/junc0 x517/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6066 x48/junc1 WWL_19 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6067 x1017/RWL1_junc RWL_5 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6068 RBL0_26 RWL_6 x756/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6069 x474/junc1 WWL_27 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6070 VDD x167/junc0 x167/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6071 VDD x518/junc0 x518/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6072 WBL_18 WWL_24 x109/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6073 RBL0_11 RWL_20 x980/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6074 x208/junc0 x208/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6075 VDD x835/junc0 x835/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6076 x653/junc0 x653/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6077 GND x310/junc0 x310/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6078 WBL_2 WWL_1 x116/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6079 x317/RWL1_junc RWL_9 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6080 x336/RWL1_junc RWL_13 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6081 x747/junc0 x747/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6082 VDD x175/junc0 x175/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6083 x215/junc0 x215/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6084 GND x254/junc1 x254/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6085 WBL_4 WWL_28 x58/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6086 x860/junc0 x860/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6087 x512/RWL0_junc x512/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6088 x897/junc0 x897/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6089 x682/RWL0_junc x682/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6090 x729/junc1 WWL_23 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6091 WBL_29 WWL_3 x670/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6092 x1002/junc0 x1002/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6093 RBL0_13 RWL_7 x161/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6094 WBL_20 WWL_11 x852/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6095 GND x168/junc1 x168/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6096 x494/junc1 WWL_0 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6097 RBL0_4 RWL_1 x738/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6098 x521/RWL0_junc x521/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6099 x750/junc0 x750/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6100 x369/RWL0_junc x369/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6101 GND x596/junc0 x596/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6102 GND x176/junc1 x176/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6103 x237/junc0 x237/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6104 RBL0_28 RWL_29 x822/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6105 GND x335/junc0 x335/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6106 GND x178/junc1 x178/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6107 x365/RWL1_junc RWL_8 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6108 x753/junc0 x753/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6109 RBL0_11 RWL_9 x434/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6110 GND x186/junc1 x186/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6111 GND x981/junc1 x981/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6112 GND x185/junc1 x185/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6113 x529/RWL0_junc x529/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6114 x530/RWL0_junc x530/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6115 GND x822/junc1 x822/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6116 x973/junc1 WWL_28 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6117 x246/junc0 x246/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6118 x505/junc1 WWL_10 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6119 RBL0_22 RWL_11 x861/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6120 GND x96/junc0 x96/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6121 VDD x552/junc0 x552/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6122 x508/junc1 WWL_20 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6123 VDD x554/junc0 x554/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6124 GND x456/junc1 x456/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6125 GND x481/junc0 x481/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6126 x744/junc0 x744/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6127 x257/junc0 x257/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6128 WBL_31 WWL_25 x163/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6129 VDD x845/junc0 x845/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6130 x726/junc0 x726/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6131 GND x197/junc1 x197/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6132 GND x351/junc0 x351/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6133 x761/junc0 x761/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6134 GND x1005/junc0 x1005/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6135 x262/junc0 x262/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6136 GND x295/junc1 x295/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6137 WBL_14 WWL_6 x170/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6138 WBL_5 WWL_14 x171/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6139 GND x205/junc1 x205/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6140 VDD x1000/junc0 x1000/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6141 x551/RWL0_junc x551/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6142 x550/RWL0_junc x550/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6143 x926/RWL0_junc x926/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6144 x745/junc1 WWL_24 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6145 GND x620/junc0 x620/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6146 x676/RWL1_junc RWL_31 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6147 x522/junc1 WWL_0 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6148 WBL_29 WWL_4 x1023/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6149 x273/junc0 x273/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6150 x963/junc1 WWL_5 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6151 RBL0_13 RWL_8 x206/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6152 GND x233/junc0 x233/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6153 GND x214/junc1 x214/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6154 x526/junc1 WWL_1 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6155 x282/junc0 x282/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6156 GND x625/junc0 x625/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6157 x769/junc0 x769/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6158 GND x626/junc0 x626/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6159 WBL_23 WWL_10 x189/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6160 GND x3/junc1 x3/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6161 GND x218/junc1 x218/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6162 x953/junc0 x953/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6163 RBL0_7 RWL_14 x518/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6164 GND x222/junc1 x222/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6165 x754/junc0 x754/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6166 x771/junc0 x771/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6167 x566/RWL0_junc x566/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6168 x487/junc1 WWL_30 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6169 x716/RWL1_junc RWL_17 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6170 x291/junc0 x291/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6171 x717/RWL0_junc x717/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6172 RBL0_31 RWL_4 x984/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6173 x540/junc1 WWL_11 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6174 VDD x159/junc0 x159/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6175 VDD x39/junc0 x39/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6176 RBL0_22 RWL_12 x797/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6177 GND x146/junc0 x146/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6178 x399/RWL1_junc RWL_13 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6179 x372/RWL0_junc x372/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6180 x553/junc0 x553/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6181 WBL_31 WWL_26 x208/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6182 RBL0_25 RWL_10 x757/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6183 x586/junc0 x586/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6184 x548/junc1 WWL_17 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6185 x588/junc0 x588/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6186 x490/junc0 x490/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6187 x783/junc0 x783/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6188 GND x472/junc0 x472/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6189 WBL_14 WWL_7 x215/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6190 x714/RWL0_junc x714/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6191 GND x253/junc1 x253/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6192 x762/RWL1_junc RWL_21 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6193 VDD x276/junc0 x276/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6194 x583/RWL0_junc x583/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6195 x584/RWL0_junc x584/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6196 x306/junc0 x306/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6197 GND x645/junc0 x645/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6198 x559/junc1 WWL_1 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6199 x891/junc1 WWL_2 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6200 VDD x475/junc0 x475/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6201 x952/junc0 x952/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6202 GND x260/junc1 x260/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6203 GND x258/junc1 x258/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6204 GND x261/junc1 x261/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6205 x317/junc0 x317/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6206 WBL_19 WWL_15 x229/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6207 GND x650/junc0 x650/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6208 x244/RWL1_junc RWL_31 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6209 x794/junc0 x794/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6210 RBL0_16 RWL_7 x989/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6211 WBL_23 WWL_11 x237/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6212 x571/junc1 WWL_14 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6213 GND x269/junc1 x269/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6214 x961/junc0 x961/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6215 RBL0_7 RWL_15 x554/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6216 x770/junc0 x770/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6217 x595/RWL0_junc x595/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6218 x601/RWL0_junc x601/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6219 GND x294/junc0 x294/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6220 GND x1008/junc0 x1008/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6221 x149/junc1 WWL_31 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6222 GND x277/junc1 x277/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6223 x758/RWL1_junc RWL_14 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6224 x50/junc0 x50/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6225 x737/RWL1_junc RWL_18 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6226 x738/RWL0_junc x738/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6227 RBL0_31 RWL_5 x831/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6228 WBL_1 WWL_22 x246/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6229 VDD x760/junc0 x760/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6230 x828/RWL0_junc x828/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6231 x580/junc1 WWL_10 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6232 WBL_31 WWL_27 x257/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6233 x723/RWL1_junc RWL_24 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6234 x1009/junc0 x1009/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6235 RBL0_25 RWL_11 x777/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6236 x581/junc1 WWL_18 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6237 x732/RWL0_junc x732/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6238 x617/junc0 x617/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6239 WBL_10 WWL_12 x726/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6240 x428/RWL1_junc RWL_31 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6241 WBL_14 WWL_8 x262/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6242 x468/RWL0_junc x468/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6243 x2/RWL1_junc RWL_22 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6244 x345/junc0 x345/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6245 VDD x441/junc0 x441/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6246 x349/junc0 x349/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6247 GND x668/junc0 x668/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6248 WBL_1 WWL_28 x212/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6249 GND x449/junc0 x449/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6250 x619/RWL0_junc x619/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6251 GND x300/junc1 x300/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6252 VDD x630/junc0 x630/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6253 x785/junc1 WWL_19 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6254 WBL_19 WWL_16 x282/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6255 GND x303/junc1 x303/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6256 RBL0_3 RWL_20 x892/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6257 x807/junc0 x807/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6258 RBL0_16 RWL_8 x992/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6259 RBL0_7 RWL_16 x587/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6260 x654/junc0 x654/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6261 GND x575/junc0 x575/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6262 VDD x330/junc0 x330/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6263 GND x313/junc1 x313/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6264 GND x332/junc0 x332/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6265 GND x314/junc1 x314/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6266 x779/RWL1_junc RWL_15 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6267 x32/RWL1_junc RWL_19 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6268 x1011/junc0 x1011/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6269 WBL_24 WWL_29 x234/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6270 WBL_1 WWL_23 x291/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6271 x792/junc1 WWL_21 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6272 RBL0_0 RWL_13 x535/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6273 GND x1016/junc0 x1016/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6274 x793/RWL0_junc x793/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6275 VDD x148/junc0 x148/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6276 VDD x152/junc0 x152/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6277 x245/junc1 WWL_15 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6278 VDD x1019/junc0 x1019/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6279 x30/RWL0_junc x30/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6280 x614/junc1 WWL_11 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6281 x45/RWL1_junc RWL_25 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6282 x943/junc0 x943/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6283 RBL0_25 RWL_12 x155/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6284 x562/junc1 WWL_30 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6285 WBL_10 WWL_13 x490/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6286 RBL0_28 RWL_24 x608/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6287 x814/junc0 x814/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6288 x389/junc0 x389/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6289 x55/RWL1_junc RWL_23 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6290 x819/junc0 x819/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6291 x820/junc0 x820/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6292 x494/RWL1_junc RWL_0 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6293 x399/junc0 x399/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6294 RBL0_3 RWL_9 x925/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6295 WBL_4 WWL_19 x306/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6296 GND x545/junc0 x545/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6297 x758/RWL0_junc x758/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6298 x643/RWL0_junc x643/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6299 x71/junc1 WWL_29 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6300 GND x600/junc0 x600/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6301 GND x598/junc0 x598/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6302 x531/junc0 x531/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6303 VDD x61/junc0 x61/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6304 x9/junc1 WWL_12 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6305 GND x689/junc0 x689/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6306 WBL_28 WWL_9 x317/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6307 GND x343/junc1 x343/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6308 x11/junc1 WWL_20 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6309 GND x341/junc1 x341/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6310 GND x342/junc1 x342/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6311 GND x695/junc0 x695/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6312 x657/junc0 x657/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6313 VDD x373/junc0 x373/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6314 x658/junc0 x658/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6315 WBL_27 WWL_21 x901/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6316 GND x357/junc1 x357/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6317 x909/junc0 x909/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6318 GND x358/junc1 x358/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6319 x157/RWL1_junc RWL_16 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6320 x1012/junc0 x1012/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6321 WBL_1 WWL_24 x50/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6322 x752/junc0 x752/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6323 GND x700/junc0 x700/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6324 GND x564/junc0 x564/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6325 VDD x384/junc0 x384/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6326 x806/RWL0_junc x806/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6327 VDD x386/junc0 x386/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6328 x35/junc1 WWL_16 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6329 VDD x1020/junc0 x1020/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6330 x421/junc0 x421/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6331 GND x506/junc1 x506/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6332 x99/RWL1_junc RWL_26 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6333 x842/junc1 WWL_31 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6334 x812/RWL1_junc RWL_20 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6335 RBL0_28 RWL_25 x630/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6336 RBL0_29 RWL_21 x813/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6337 x826/junc0 x826/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6338 x775/RWL0_junc x775/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6339 x973/RWL1_junc RWL_28 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6340 x432/junc0 x432/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6341 x660/RWL0_junc x660/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6342 GND x375/junc1 x375/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6343 x526/RWL1_junc RWL_1 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6344 RBL0_12 RWL_2 x634/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6345 WBL_13 WWL_12 x345/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6346 x664/RWL0_junc x664/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6347 WBL_4 WWL_20 x349/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6348 x109/junc0 x109/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6349 x779/RWL0_junc x779/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6350 x667/RWL0_junc x667/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6351 x438/junc0 x438/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6352 RBL0_7 RWL_28 x1013/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6353 GND x21/junc0 x21/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6354 GND x18/junc0 x18/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6355 GND x20/junc0 x20/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6356 VDD x410/junc0 x410/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6357 GND x446/junc0 x446/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6358 x63/junc1 WWL_13 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6359 VDD x75/junc0 x75/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6360 GND x393/junc1 x393/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6361 GND x392/junc1 x392/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6362 GND x395/junc1 x395/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6363 GND x1013/junc1 x1013/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6364 RBL0_17 RWL_10 x1019/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6365 GND x400/junc1 x400/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6366 GND x37/junc0 x37/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6367 x678/junc0 x678/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6368 x323/junc1 WWL_19 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6369 x680/junc0 x680/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6370 RBL0_21 RWL_6 x228/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6371 RBL0_6 RWL_20 x1001/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6372 GND x404/junc1 x404/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6373 VDD x686/junc0 x686/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6374 x915/junc0 x915/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6375 x454/junc0 x454/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6376 VDD x240/junc0 x240/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6377 x402/junc0 x402/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6378 x533/RWL1_junc RWL_9 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6379 x764/junc0 x764/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6380 GND x47/junc0 x47/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6381 GND x527/junc0 x527/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6382 RBL0_14 RWL_24 x919/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6383 x810/RWL1_junc RWL_13 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6384 VDD x426/junc0 x426/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6385 x22/RWL0_junc x22/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6386 RBL0_30 RWL_30 x537/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6387 x832/junc0 x832/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6388 x458/junc0 x458/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6389 RBL0_31 RWL_31 x932/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6390 GND x382/junc0 x382/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6391 x31/RWL0_junc x31/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6392 x94/junc1 WWL_21 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6393 x487/RWL1_junc RWL_30 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6394 RBL0_28 RWL_26 x652/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6395 RBL0_29 RWL_22 x254/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6396 x834/junc0 x834/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6397 x796/RWL0_junc x796/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6398 x999/RWL1_junc RWL_29 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6399 x976/junc0 x976/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6400 WBL_24 WWL_3 x389/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6401 RBL0_8 RWL_7 x413/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6402 x3/RWL1_junc RWL_31 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6403 GND x419/junc1 x419/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6404 RBL0_12 x61/RWL1 x656/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6405 WBL_13 WWL_13 x399/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6406 x44/RWL0_junc x44/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6407 x836/junc0 x836/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6408 x837/junc0 x837/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6409 x157/RWL0_junc x157/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6410 x468/junc0 x468/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6411 RBL0_3 RWL_30 x768/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6412 GND x427/junc1 x427/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6413 x469/junc0 x469/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6414 RBL0_7 RWL_29 x883/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6415 x170/RWL1_junc RWL_6 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6416 GND x77/junc0 x77/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6417 GND x78/junc0 x78/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6418 GND x79/junc0 x79/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6419 x838/junc0 x838/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6420 VDD x448/junc0 x448/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6421 WBL_6 WWL_30 x346/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6422 RBL0_6 RWL_9 x623/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6423 GND x437/junc1 x437/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6424 GND x436/junc1 x436/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6425 x56/RWL0_junc x56/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6426 GND x883/junc1 x883/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6427 x15/junc1 WWL_10 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6428 x778/RWL1_junc RWL_24 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6429 RBL0_17 RWL_11 x1020/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6430 x862/junc1 WWL_12 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6431 x17/junc1 WWL_20 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6432 x703/junc0 x703/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6433 VDD x706/junc0 x706/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6434 WBL_15 WWL_0 x909/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6435 GND x741/junc0 x741/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6436 x580/RWL1_junc RWL_10 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6437 GND x92/junc0 x92/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6438 x805/RWL1_junc RWL_14 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6439 x481/junc0 x481/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6440 WBL_26 WWL_25 x415/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6441 VDD x910/junc0 x910/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6442 GND x444/junc1 x444/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6443 GND x101/junc0 x101/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6444 x484/junc0 x484/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6445 x29/junc1 WWL_17 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6446 RBL0_14 RWL_25 x830/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6447 x841/junc0 x841/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6448 GND x104/junc0 x104/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6449 x488/junc0 x488/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6450 WBL_9 WWL_6 x421/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6451 GND x451/junc1 x451/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6452 VDD x1021/junc0 x1021/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6453 x647/junc0 x647/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6454 x88/RWL0_junc x88/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6455 WBL_10 WWL_28 x475/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6456 RBL0_29 RWL_23 x295/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6457 x195/RWL0_junc x195/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6458 GND x199/junc1 x199/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6459 WBL_24 WWL_4 x432/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6460 RBL0_8 RWL_8 x452/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6461 RBL0_9 RWL_31 x122/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6462 GND x118/junc0 x118/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6463 x846/junc0 x846/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6464 GND x125/junc0 x125/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6465 x847/junc0 x847/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6466 x132/junc0 x132/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6467 WBL_18 WWL_10 x438/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6468 GND x461/junc1 x461/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6469 GND x460/junc1 x460/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6470 x813/RWL0_junc x813/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6471 RBL0_2 RWL_14 x686/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6472 WBL_6 WWL_31 x394/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6473 x848/junc0 x848/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6474 x111/RWL0_junc x111/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6475 x818/RWL1_junc RWL_17 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6476 x69/junc1 WWL_3 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6477 x591/RWL1_junc RWL_25 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6478 RBL0_26 RWL_4 x1003/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6479 x70/junc1 WWL_11 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6480 VDD x412/junc0 x412/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6481 VDD x312/junc0 x312/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6482 RBL0_17 RWL_12 x862/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6483 x594/RWL1_junc RWL_13 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6484 x874/junc1 WWL_13 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6485 GND x385/junc0 x385/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6486 WBL_15 WWL_1 x915/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6487 GND x515/junc0 x515/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6488 RBL0_27 RWL_31 x136/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6489 GND x144/junc0 x144/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6490 x839/RWL1_junc RWL_7 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6491 x614/RWL1_junc RWL_11 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6492 WBL_26 WWL_26 x454/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6493 x229/RWL1_junc RWL_15 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6494 x727/junc0 x727/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6495 GND x227/junc1 x227/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6496 GND x906/junc1 x906/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6497 x86/junc1 WWL_18 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6498 x519/junc0 x519/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6499 RBL0_14 RWL_26 x327/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6500 x853/junc0 x853/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6501 GND x153/junc0 x153/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6502 WBL_9 WWL_7 x458/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6503 x133/RWL0_junc x133/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6504 GND x477/junc1 x477/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6505 VDD x1022/junc0 x1022/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6506 x725/RWL0_junc x725/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6507 WBL_20 WWL_9 x301/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6508 GND x483/junc1 x483/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6509 GND x486/junc1 x486/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6510 x919/RWL0_junc x919/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6511 x174/RWL0_junc x174/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6512 GND x492/junc1 x492/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6513 x533/junc0 x533/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6514 x855/junc0 x855/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6515 GND x172/junc0 x172/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6516 x112/junc1 WWL_6 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6517 x181/junc0 x181/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6518 x857/junc0 x857/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6519 RBL0_11 RWL_7 x1004/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6520 WBL_18 WWL_11 x469/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6521 x113/junc1 WWL_14 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6522 GND x493/junc1 x493/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6523 x254/RWL0_junc x254/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6524 RBL0_2 RWL_15 x706/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6525 x538/junc0 x538/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6526 x1014/junc0 x1014/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6527 GND x183/junc0 x183/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6528 x849/RWL1_junc RWL_10 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6529 x736/RWL0_junc x736/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6530 GND x184/junc0 x184/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6531 x124/junc1 WWL_4 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6532 VDD x223/junc0 x223/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6533 x893/RWL1_junc RWL_26 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6534 x827/RWL1_junc RWL_18 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6535 RBL0_26 RWL_5 x895/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6536 GND x789/junc1 x789/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6537 VDD x5/junc0 x5/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6538 VDD x24/junc0 x24/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6539 x851/RWL1_junc RWL_8 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6540 x637/RWL1_junc RWL_12 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6541 x956/junc0 x956/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6542 x850/junc1 WWL_10 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6543 WBL_26 WWL_27 x481/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6544 VDD x747/junc0 x747/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6545 x866/junc0 x866/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6546 x282/RWL1_junc RWL_16 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6547 GND x278/junc1 x278/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6548 x53/junc1 WWL_28 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6549 WBL_5 WWL_12 x484/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6550 x0/RWL0_junc x0/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6551 WBL_9 WWL_8 x488/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6552 x506/junc0 x506/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6553 RBL0_5 RWL_31 x456/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6554 x555/junc0 x555/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6555 x186/RWL0_junc x186/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6556 x709/junc0 x709/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6557 WBL_29 WWL_2 x647/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6558 GND x512/junc1 x512/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6559 x22/junc0 x22/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6560 GND x207/junc0 x207/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6561 x599/RWL0_junc x599/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6562 x830/RWL0_junc x830/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6563 x191/RWL0_junc x191/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6564 VDD x750/junc0 x750/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6565 GND x521/junc1 x521/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6566 x161/junc1 WWL_7 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6567 x7/junc0 x7/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6568 RBL0_11 RWL_8 x1007/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6569 x295/RWL0_junc x295/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6570 RBL0_2 RWL_16 x728/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6571 GND x219/junc0 x219/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6572 x575/junc0 x575/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6573 x574/junc0 x574/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6574 VDD x547/junc0 x547/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6575 x165/junc1 WWL_9 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6576 RBL0_0 RWL_30 x649/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6577 GND x529/junc1 x529/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6578 GND x530/junc1 x530/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6579 x873/junc0 x873/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6580 x859/RWL1_junc RWL_11 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6581 WBL_3 WWL_29 x713/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6582 x306/RWL1_junc RWL_19 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6583 RBL0_0 RWL_31 x3/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6584 VDD x613/junc0 x613/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6585 x214/RWL0_junc x214/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6586 VDD x1010/junc0 x1010/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6587 VDD x140/junc0 x140/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6588 x268/junc1 WWL_15 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6589 x864/junc0 x864/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6590 x304/RWL0_junc x304/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6591 x861/junc1 WWL_11 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6592 WBL_14 WWL_5 x514/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6593 x94/RWL1_junc RWL_21 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6594 WBL_5 WWL_13 x519/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6595 x218/RWL0_junc x218/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6596 x231/RWL0_junc x231/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6597 RBL0_23 RWL_24 x740/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6598 x879/junc0 x879/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6599 x54/RWL0_junc x54/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6600 x74/junc0 x74/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6601 x117/junc1 WWL_28 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6602 x881/junc0 x881/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6603 x882/junc0 x882/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6604 x671/junc0 x671/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6605 GND x551/junc1 x551/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6606 x594/junc0 x594/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6607 GND x550/junc1 x550/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6608 GND x256/junc0 x256/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6609 VDD x496/junc0 x496/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6610 x671/junc0 x671/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6611 x759/RWL0_junc x759/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6612 x327/RWL0_junc x327/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6613 x50/junc0 x50/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6614 x994/RWL0_junc x994/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6615 x238/RWL0_junc x238/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6616 GND x259/junc0 x259/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6617 x598/junc0 x598/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6618 x600/junc0 x600/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6619 x692/junc0 x692/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6620 VDD x424/junc0 x424/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6621 WBL_23 WWL_9 x533/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6622 x202/junc1 WWL_12 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6623 GND x929/junc1 x929/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6624 GND x558/junc1 x558/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6625 GND x264/junc0 x264/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6626 x206/junc1 WWL_8 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6627 GND x267/junc0 x267/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6628 x695/junc0 x695/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6629 RBL0_15 RWL_17 x341/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6630 WBL_30 WWL_17 x538/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6631 x772/junc0 x772/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6632 VDD x579/junc0 x579/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6633 RBL0_0 RWL_10 x871/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6634 WBL_22 WWL_21 x1014/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6635 GND x566/junc1 x566/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6636 x73/junc0 x73/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6637 x345/RWL1_junc RWL_12 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6638 x463/RWL1_junc RWL_24 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6639 GND x283/junc0 x283/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6640 x29/RWL1_junc RWL_17 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6641 x261/RWL0_junc x261/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6642 VDD x588/junc0 x588/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6643 VDD x586/junc0 x586/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6644 x217/junc1 WWL_16 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6645 RBL0_1 RWL_31 x607/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6646 x114/junc0 x114/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6647 x544/junc1 WWL_29 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6648 x687/RWL1_junc RWL_22 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6649 x269/RWL0_junc x269/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6650 x889/junc0 x889/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6651 RBL0_24 RWL_21 x878/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6652 x877/RWL1_junc RWL_20 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6653 VDD x653/junc0 x653/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6654 RBL0_23 RWL_25 x750/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6655 x890/junc0 x890/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6656 x622/junc0 x622/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6657 RBL0_7 RWL_2 x753/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6658 GND x584/junc1 x584/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6659 GND x583/junc1 x583/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6660 x281/RWL0_junc x281/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6661 VDD x528/junc0 x528/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6662 x542/RWL0_junc x542/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6663 x135/junc0 x135/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6664 x780/RWL0_junc x780/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6665 x107/junc0 x107/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6666 x997/RWL0_junc x997/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6667 x781/RWL0_junc x781/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6668 GND x298/junc0 x298/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6669 GND x299/junc0 x299/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6670 x18/junc0 x18/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6671 VDD x794/junc0 x794/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6672 x21/junc0 x21/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6673 VDD x609/junc0 x609/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6674 x138/junc1 WWL_13 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6675 GND x592/junc1 x592/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6676 GND x938/junc1 x938/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6677 x755/RWL1_junc RWL_30 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6678 GND x595/junc1 x595/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6679 GND x307/junc0 x307/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6680 RBL0_15 RWL_18 x392/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6681 WBL_30 WWL_18 x574/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6682 WBL_31 WWL_14 x575/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6683 RBL0_0 RWL_11 x886/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6684 x110/junc1 WWL_19 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6685 x795/junc0 x795/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6686 GND x601/junc1 x601/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6687 x127/junc0 x127/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6688 x854/RWL0_junc x854/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6689 x635/junc0 x635/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6690 x85/RWL1_junc RWL_25 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6691 x693/RWL1_junc RWL_9 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6692 GND x322/junc0 x322/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6693 x86/RWL1_junc RWL_18 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6694 x856/RWL0_junc x856/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6695 x266/junc1 WWL_9 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6696 RBL0_9 RWL_30 x67/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6697 RBL0_9 RWL_24 x957/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6698 VDD x617/junc0 x617/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6699 x300/RWL0_junc x300/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6700 x896/junc0 x896/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6701 x638/junc0 x638/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6702 x156/junc0 x156/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6703 x708/RWL1_junc RWL_23 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6704 x280/junc1 WWL_21 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6705 x305/RWL0_junc x305/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6706 x898/junc0 x898/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6707 VDD x557/junc0 x557/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6708 RBL0_23 RWL_26 x769/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6709 RBL0_24 RWL_22 x478/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6710 x900/junc0 x900/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6711 x387/junc0 x387/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6712 VDD x676/junc0 x676/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6713 x996/junc0 x996/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6714 x284/junc1 WWL_6 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6715 WBL_19 WWL_3 x74/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6716 RBL0_3 RWL_7 x953/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6717 RBL0_7 RWL_3 x771/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6718 x316/RWL0_junc x316/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6719 x320/RWL0_junc x320/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6720 VDD x608/junc0 x608/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6721 x766/RWL1_junc RWL_28 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6722 x287/junc0 x287/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6723 x185/junc0 x185/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6724 x735/RWL1_junc RWL_2 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6725 GND x619/junc1 x619/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6726 x158/junc0 x158/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6727 GND x340/junc0 x340/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6728 x421/RWL1_junc RWL_6 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6729 GND x339/junc0 x339/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6730 WBL_16 WWL_17 x600/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6731 VDD x807/junc0 x807/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6732 WBL_1 WWL_10 x598/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6733 VDD x631/junc0 x631/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6734 GND x674/junc1 x674/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6735 RBL0_13 RWL_28 x13/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6736 GND x624/junc1 x624/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6737 x394/RWL0_junc x394/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6738 VDD x495/junc0 x495/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6739 RBL0_19 RWL_28 x105/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6740 VDD x25/junc0 x25/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6741 WBL_27 WWL_19 x855/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6742 WBL_16 WWL_28 x565/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6743 VDD x115/junc0 x115/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6744 RBL0_15 RWL_19 x437/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6745 RBL0_0 RWL_12 x499/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6746 x230/junc1 WWL_29 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6747 x892/junc1 WWL_20 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6748 x808/junc0 x808/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6749 WBL_10 WWL_0 x73/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6750 GND x58/junc0 x58/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6751 x850/RWL1_junc RWL_10 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6752 x92/junc0 x92/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6753 WBL_21 WWL_25 x612/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6754 VDD x134/junc0 x134/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6755 x722/RWL1_junc RWL_26 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6756 GND x364/junc0 x364/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6757 x724/RWL1_junc RWL_19 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6758 x869/RWL0_junc x869/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6759 x904/junc0 x904/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6760 RBL0_9 RWL_25 x894/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6761 x905/junc0 x905/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6762 x370/junc0 x370/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6763 WBL_4 WWL_6 x114/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6764 x661/junc0 x661/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6765 x199/junc0 x199/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6766 x200/junc0 x200/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6767 x310/junc1 WWL_22 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6768 VDD x814/junc0 x814/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6769 RBL0_20 RWL_27 x444/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6770 x666/junc0 x666/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6771 x348/RWL0_junc x348/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6772 x907/junc0 x907/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6773 VDD x820/junc0 x820/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6774 RBL0_24 RWL_23 x510/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6775 x604/RWL0_junc x604/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6776 RBL0_12 RWL_0 x794/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6777 x321/junc1 WWL_7 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6778 WBL_19 WWL_4 x622/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6779 RBL0_3 RWL_8 x961/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6780 x607/RWL0_junc x607/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6781 GND x84/junc0 x84/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6782 x360/RWL0_junc x360/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6783 x790/RWL1_junc RWL_30 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6784 GND x377/junc0 x377/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6785 x230/RWL1_junc RWL_29 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6786 GND x378/junc0 x378/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6787 x497/junc0 x497/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6788 WBL_12 WWL_22 x135/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6789 VDD x128/junc0 x128/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6790 GND x643/junc1 x643/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6791 GND x36/junc1 x36/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6792 GND x383/junc0 x383/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6793 x501/RWL1_junc x61/RWL1 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6794 x878/RWL0_junc x878/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6795 WBL_1 WWL_11 x21/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6796 WBL_16 WWL_18 x18/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6797 GND x391/junc0 x391/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6798 RBL0_13 RWL_29 x697/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6799 x335/junc1 WWL_3 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6800 VDD x658/junc0 x658/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6801 RBL0_19 RWL_29 x733/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6802 WBL_12 WWL_30 x24/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6803 WBL_27 WWL_20 x962/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6804 RBL0_21 RWL_4 x1009/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6805 VDD x610/junc0 x610/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6806 x732/RWL1_junc RWL_13 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6807 WBL_10 WWL_1 x127/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6808 x903/RWL1_junc RWL_7 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6809 GND x683/junc0 x683/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6810 GND x403/junc0 x403/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6811 x861/RWL1_junc RWL_11 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6812 x96/junc1 WWL_25 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6813 x288/junc1 WWL_28 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6814 WBL_21 WWL_26 x635/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6815 x912/junc0 x912/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6816 GND x593/junc0 x593/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6817 RBL0_9 RWL_26 x541/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6818 x913/junc0 x913/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6819 x414/junc0 x414/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6820 WBL_4 WWL_7 x638/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6821 x352/junc1 WWL_19 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6822 x735/RWL0_junc x735/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6823 x351/junc1 WWL_23 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6824 RBL0_29 RWL_20 x906/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6825 VDD x826/junc0 x826/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6826 x825/RWL0_junc x825/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6827 x362/junc1 WWL_0 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6828 RBL0_12 RWL_1 x807/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6829 x365/junc1 WWL_8 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6830 GND x76/junc1 x76/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6831 x887/RWL1_junc RWL_27 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6832 GND x660/junc1 x660/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6833 x957/RWL0_junc x957/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6834 WBL_22 WWL_28 x59/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6835 GND x744/junc1 x744/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6836 GND x14/junc0 x14/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6837 GND x664/junc1 x664/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6838 x693/junc0 x693/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6839 GND x770/junc1 x770/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6840 x888/RWL1_junc RWL_4 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6841 x633/RWL0_junc x633/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6842 GND x423/junc0 x423/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6843 x646/junc0 x646/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6844 x233/junc1 WWL_6 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6845 x60/junc0 x60/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6846 GND x667/junc1 x667/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6847 WBL_12 WWL_23 x185/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6848 RBL0_6 RWL_7 x1011/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6849 x478/RWL0_junc x478/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6850 x696/junc0 x696/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6851 x788/junc0 x788/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6852 GND x26/junc0 x26/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6853 x793/RWL1_junc RWL_10 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6854 GND x27/junc0 x27/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6855 GND x874/junc0 x874/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6856 GND x435/junc0 x435/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6857 x376/junc1 WWL_4 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6858 VDD x678/junc0 x678/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6859 RBL0_21 RWL_5 x943/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6860 WBL_12 WWL_31 x613/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6861 VDD x292/junc0 x292/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6862 x388/junc1 WWL_22 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6863 x920/junc0 x920/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6864 x911/RWL1_junc RWL_8 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6865 RBL0_29 RWL_9 x789/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6866 x797/RWL1_junc RWL_12 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6867 x146/junc1 WWL_26 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6868 VDD x832/junc0 x832/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6869 x465/junc1 WWL_15 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6870 WBL_21 WWL_27 x92/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6871 x89/junc0 x89/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6872 RBL0_28 RWL_13 x819/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6873 x921/junc0 x921/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6874 GND x71/junc0 x71/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6875 WBL_13 WWL_0 x370/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6876 WBL_4 WWL_8 x661/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6877 GND x754/junc1 x754/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6878 x401/junc1 WWL_24 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6879 x141/junc1 WWL_20 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6880 x501/RWL0_junc x501/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6881 WBL_24 WWL_2 x666/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6882 GND x57/junc0 x57/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6883 GND x31/junc1 x31/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6884 x408/junc1 WWL_1 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6885 GND x453/junc0 x453/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6886 GND x684/junc1 x684/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6887 x42/RWL0_junc x42/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6888 x894/RWL0_junc x894/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6889 VDD x836/junc0 x836/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6890 VDD x837/junc0 x837/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6891 x714/junc0 x714/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6892 GND x44/junc1 x44/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6893 x514/RWL1_junc RWL_5 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6894 x344/junc0 x344/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6895 x413/junc1 WWL_7 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6896 WBL_12 WWL_24 x497/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6897 x116/junc0 x116/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6898 RBL0_6 RWL_8 x1012/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6899 x510/RWL0_junc x510/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6900 GND x394/junc0 x394/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6901 GND x80/junc0 x80/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6902 x718/junc0 x718/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6903 x219/junc0 x219/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6904 VDD x701/junc0 x701/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6905 x315/junc1 WWL_9 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6906 RBL0_1 RWL_24 x50/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6907 x806/RWL1_junc RWL_11 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6908 GND x81/junc0 x81/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6909 GND x56/junc1 x56/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6910 x930/junc0 x930/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6911 VDD x605/junc0 x605/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6912 x525/RWL0_junc x525/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6913 x381/junc1 WWL_27 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6914 x430/junc1 WWL_23 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6915 x431/junc1 WWL_16 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6916 WBL_9 WWL_5 x253/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6917 WBL_25 WWL_30 x653/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6918 x280/RWL1_junc RWL_21 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6919 x460/RWL0_junc x460/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6920 VDD x407/junc0 x407/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6921 WBL_13 WWL_1 x414/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6922 RBL0_18 RWL_24 x109/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6923 VDD x752/junc0 x752/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6924 GND x773/junc1 x773/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6925 x372/junc1 WWL_28 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6926 x934/junc0 x934/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6927 WBL_8 WWL_17 x232/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6928 GND x87/junc1 x87/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6929 GND x88/junc1 x88/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6930 x265/RWL0_junc x265/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6931 GND x607/junc0 x607/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6932 GND x480/junc0 x480/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6933 VDD x672/junc0 x672/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6934 x188/junc0 x188/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6935 x97/RWL0_junc x97/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6936 x98/RWL0_junc x98/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6937 x541/RWL0_junc x541/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6938 VDD x846/junc0 x846/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6939 GND x120/junc0 x120/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6940 x259/junc0 x259/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6941 VDD x226/junc0 x226/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6942 x449/junc1 WWL_12 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6943 x802/junc0 x802/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6944 WBL_18 WWL_9 x693/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6945 x906/RWL0_junc x906/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6946 x945/junc1 WWL_0 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6947 x452/junc1 WWL_8 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6948 x247/junc0 x247/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6949 GND x130/junc0 x130/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6950 x16/RWL1_junc RWL_2 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6951 GND x131/junc0 x131/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6952 x267/junc0 x267/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6953 x355/junc1 WWL_2 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6954 WBL_17 WWL_21 x788/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6955 RBL0_10 RWL_17 x929/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6956 WBL_25 WWL_17 x696/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6957 x171/junc0 x171/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6958 VDD x721/junc0 x721/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6959 GND x967/junc1 x967/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6960 RBL0_1 RWL_25 x107/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6961 x337/junc0 x337/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6962 GND x111/junc1 x111/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6963 x22/RWL1_junc RWL_12 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6964 RBL0_14 RWL_13 x63/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6965 x28/RWL1_junc RWL_24 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6966 x1023/junc0 x1023/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6967 VDD x627/junc0 x627/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6968 VDD x727/junc0 x727/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6969 x463/junc1 WWL_24 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6970 x816/junc0 x816/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6971 x40/RWL1_junc RWL_22 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6972 WBL_25 WWL_31 x676/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6973 x493/RWL0_junc x493/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6974 x189/junc0 x189/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6975 RBL0_19 RWL_21 x931/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6976 VDD x402/junc0 x402/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6977 RBL0_18 RWL_25 x837/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6978 x416/junc1 WWL_30 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6979 x356/junc0 x356/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6980 WBL_8 WWL_18 x285/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6981 RBL0_2 RWL_2 x838/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6982 GND x139/junc1 x139/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6983 x789/RWL0_junc x789/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6984 GND x725/junc1 x725/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6985 x302/RWL0_junc x302/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6986 VDD x691/junc0 x691/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6987 x998/junc0 x998/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6988 x393/junc0 x393/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6989 x147/RWL0_junc x147/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6990 GND x517/junc0 x517/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6991 x151/RWL0_junc x151/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6992 GND x167/junc0 x167/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6993 GND x518/junc0 x518/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6994 x299/junc0 x299/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6995 x535/RWL1_junc RWL_13 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6996 VDD x857/junc0 x857/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6997 x545/junc1 WWL_5 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M6998 VDD x742/junc0 x742/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M6999 x396/junc1 WWL_13 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7000 x951/junc1 WWL_1 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7001 x749/junc0 x749/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7002 x404/junc0 x404/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7003 x1018/junc0 x1018/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7004 GND x175/junc0 x175/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7005 x74/RWL1_junc x61/RWL1 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7006 x215/junc0 x215/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7007 x482/junc1 WWL_17 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7008 GND x177/junc0 x177/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7009 RBL0_10 RWL_18 x938/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7010 WBL_25 WWL_18 x718/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7011 x860/junc0 x860/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7012 WBL_26 WWL_14 x219/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7013 GND x971/junc1 x971/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7014 RBL0_1 RWL_26 x158/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7015 x914/RWL0_junc x914/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7016 GND x736/junc1 x736/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7017 x379/junc0 x379/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7018 GND x549/junc1 x549/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7019 x82/RWL1_junc RWL_25 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7020 x916/RWL0_junc x916/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7021 x1002/junc0 x1002/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7022 x937/junc1 WWL_9 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7023 x999/junc0 x999/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7024 RBL0_4 RWL_24 x982/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7025 VDD x866/junc0 x866/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7026 x93/RWL1_junc RWL_23 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7027 x277/junc1 WWL_21 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7028 x1021/junc1 WWL_17 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7029 x237/junc0 x237/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7030 VDD x908/junc0 x908/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7031 VDD x387/junc0 x387/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7032 RBL0_18 RWL_26 x847/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7033 RBL0_19 RWL_22 x655/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7034 x456/junc1 WWL_31 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7035 RBL0_2 RWL_3 x848/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7036 VDD x924/junc0 x924/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7037 x813/RWL1_junc RWL_21 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7038 x190/RWL0_junc x190/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7039 x192/RWL0_junc x192/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7040 VDD x740/junc0 x740/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7041 x436/junc0 x436/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7042 GND x191/junc1 x191/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7043 GND x552/junc0 x552/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7044 GND x554/junc0 x554/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7045 x114/RWL1_junc RWL_6 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7046 GND x213/junc0 x213/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7047 WBL_11 WWL_17 x259/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7048 VDD x7/junc0 x7/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7049 VDD x751/junc0 x751/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7050 x744/junc0 x744/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7051 x257/junc0 x257/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7052 x767/junc0 x767/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7053 WBL_30 WWL_15 x357/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7054 WBL_22 WWL_19 x247/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7055 x513/junc1 WWL_18 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7056 x262/junc0 x262/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7057 x467/junc1 WWL_29 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7058 RBL0_10 RWL_19 x674/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7059 x872/junc0 x872/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7060 WBL_5 WWL_0 x337/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7061 GND x209/junc1 x209/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7062 x137/RWL1_junc RWL_26 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7063 x927/RWL0_junc x927/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7064 x211/junc0 x211/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7065 RBL0_4 RWL_25 x942/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7066 x273/junc0 x273/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7067 x578/junc0 x578/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7068 x141/RWL1_junc RWL_20 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7069 x47/junc1 WWL_22 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7070 VDD x879/junc0 x879/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7071 RBL0_15 RWL_30 x382/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7072 x221/RWL0_junc x221/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7073 x223/RWL0_junc x223/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7074 x63/RWL0_junc x63/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7075 x16/junc0 x16/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7076 x1022/junc1 WWL_18 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7077 x948/junc0 x948/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7078 VDD x882/junc0 x882/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7079 RBL0_19 RWL_23 x677/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7080 RBL0_7 RWL_0 x857/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7081 x754/junc0 x754/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7082 x998/RWL1_junc RWL_31 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7083 VDD x932/junc0 x932/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7084 x254/RWL1_junc RWL_22 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7085 x235/RWL0_junc x235/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7086 GND x255/junc0 x255/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7087 x787/junc0 x787/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7088 x786/junc0 x786/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7089 x673/junc0 x673/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7090 WBL_7 WWL_22 x393/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7091 VDD x380/junc0 x380/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7092 GND x759/junc1 x759/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7093 GND x238/junc1 x238/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7094 GND x585/junc0 x585/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7095 GND x241/junc1 x241/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7096 GND x587/junc0 x587/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7097 x931/RWL0_junc x931/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7098 WBL_11 WWL_18 x299/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7099 x544/junc0 x544/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7100 x78/junc1 WWL_3 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7101 WBL_31 WWL_12 x749/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7102 WBL_30 WWL_16 x404/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7103 VDD x772/junc0 x772/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7104 WBL_22 WWL_20 x1018/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7105 WBL_5 WWL_1 x379/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7106 x176/RWL1_junc RWL_9 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7107 x178/RWL1_junc RWL_7 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7108 GND x276/junc0 x276/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7109 VDD x822/junc0 x822/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7110 x90/junc1 WWL_25 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7111 GND x765/junc1 x765/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7112 GND x475/junc0 x475/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7113 x952/junc0 x952/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7114 x416/RWL1_junc RWL_30 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7115 RBL0_4 RWL_26 x698/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7116 x611/junc0 x611/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7117 GND x608/junc0 x608/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7118 VDD x889/junc0 x889/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7119 x561/junc1 WWL_19 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7120 GND x618/junc1 x618/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7121 x101/junc1 WWL_23 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7122 VDD x890/junc0 x890/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7123 RBL0_24 RWL_20 x947/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7124 x272/RWL0_junc x272/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7125 x1/junc0 x1/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7126 x573/junc1 WWL_0 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7127 x770/junc0 x770/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7128 RBL0_7 RWL_1 x7/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7129 GND x338/junc1 x338/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7130 x197/RWL1_junc RWL_27 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7131 x773/junc0 x773/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7132 x982/RWL0_junc x982/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7133 x295/RWL1_junc RWL_23 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7134 x945/RWL1_junc RWL_0 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7135 GND x296/junc0 x296/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7136 GND x281/junc1 x281/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7137 x205/RWL1_junc RWL_4 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7138 WBL_16 WWL_15 x763/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7139 x891/junc0 x891/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7140 x118/junc1 WWL_6 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7141 GND x780/junc1 x780/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7142 WBL_7 WWL_23 x436/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7143 GND x781/junc1 x781/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7144 x939/RWL0_junc x939/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7145 x655/RWL0_junc x655/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7146 x804/junc0 x804/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7147 GND x301/junc0 x301/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7148 x214/RWL1_junc RWL_10 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7149 GND x1006/junc1 x1006/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7150 VDD x795/junc0 x795/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7151 WBL_31 WWL_13 x767/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7152 x582/junc1 WWL_4 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7153 x654/junc0 x654/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7154 x590/junc1 WWL_22 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7155 x958/junc0 x958/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7156 x222/RWL1_junc RWL_8 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7157 RBL0_24 RWL_9 x165/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7158 x140/junc1 WWL_26 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7159 VDD x896/junc0 x896/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7160 RBL0_23 RWL_13 x881/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7161 x349/junc0 x349/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7162 GND x491/junc0 x491/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7163 x959/junc0 x959/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7164 GND x630/junc0 x630/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7165 GND x243/junc1 x243/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7166 x497/junc0 x497/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7167 VDD x898/junc0 x898/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7168 GND x91/junc1 x91/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7169 x597/junc1 WWL_24 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7170 x400/junc1 WWL_20 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7171 x49/junc0 x49/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7172 x51/junc0 x51/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7173 GND x634/junc0 x634/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7174 x153/junc1 WWL_5 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7175 x502/junc0 x502/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7176 WBL_19 WWL_2 x16/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7177 GND x329/junc0 x329/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7178 GND x305/junc1 x305/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7179 x606/junc1 WWL_1 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7180 GND x102/junc1 x102/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7181 x941/RWL0_junc x941/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7182 x318/RWL0_junc x318/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7183 GND x330/junc0 x330/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7184 x942/RWL0_junc x942/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7185 VDD x154/junc0 x154/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7186 WBL_27 WWL_6 x356/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7187 GND x316/junc1 x316/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7188 GND x320/junc1 x320/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7189 RBL0_28 RWL_30 x263/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7190 x951/RWL1_junc RWL_1 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7191 x253/RWL1_junc RWL_5 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7192 x902/junc0 x902/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7193 RBL0_15 RWL_6 x684/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7194 x953/junc1 WWL_7 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7195 WBL_1 WWL_9 x786/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7196 WBL_16 WWL_16 x787/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7197 WBL_7 WWL_24 x673/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7198 x944/RWL0_junc x944/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7199 x677/RWL0_junc x677/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7200 GND x1019/junc0 x1019/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7201 GND x263/junc1 x263/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7202 x482/RWL1_junc RWL_17 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7203 x824/junc0 x824/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7204 x80/junc0 x80/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7205 x258/RWL1_junc RWL_6 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7206 x260/RWL1_junc RWL_13 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7207 x261/RWL1_junc RWL_11 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7208 x966/junc0 x966/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7209 RBL0_28 RWL_10 x889/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7210 RBL0_20 RWL_14 x56/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7211 x621/junc1 WWL_23 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7212 VDD x904/junc0 x904/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7213 x586/junc1 WWL_27 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7214 WBL_4 WWL_5 x477/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7215 WBL_4 WWL_30 x402/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7216 x277/RWL1_junc RWL_21 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7217 x945/RWL0_junc x945/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7218 VDD x743/junc0 x743/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7219 GND x287/junc1 x287/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7220 GND x652/junc0 x652/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7221 x531/junc0 x531/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7222 x106/junc0 x106/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7223 GND x142/junc1 x142/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7224 WBL_3 WWL_17 x1/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7225 GND x656/junc0 x656/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7226 GND x347/junc1 x347/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7227 GND x348/junc1 x348/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7228 VDD x2/junc0 x2/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7229 GND x542/junc0 x542/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7230 x361/RWL0_junc x361/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7231 x946/RWL0_junc x946/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7232 GND x373/junc0 x373/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7233 x698/RWL0_junc x698/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7234 VDD x6/junc0 x6/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7235 x909/junc0 x909/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7236 WBL_27 WWL_7 x10/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7237 x120/junc0 x120/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7238 GND x360/junc1 x360/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7239 GND x394/junc1 x394/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7240 x947/RWL0_junc x947/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7241 x961/junc1 WWL_8 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7242 x569/junc0 x569/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7243 x4/RWL0_junc x4/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7244 GND x384/junc0 x384/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7245 GND x1020/junc0 x1020/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7246 GND x386/junc0 x386/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7247 x513/RWL1_junc RWL_18 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7248 x131/junc0 x131/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7249 x567/junc1 WWL_2 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7250 GND x368/junc1 x368/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7251 x174/junc1 WWL_30 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7252 RBL0_5 RWL_17 x965/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7253 x8/junc0 x8/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7254 x300/RWL1_junc RWL_12 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7255 RBL0_9 RWL_13 x138/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7256 x640/junc1 WWL_6 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7257 x641/junc1 WWL_10 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7258 x303/RWL1_junc RWL_24 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7259 x432/junc0 x432/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7260 RBL0_29 RWL_7 x967/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7261 VDD x32/junc0 x32/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7262 RBL0_28 RWL_11 x898/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7263 x13/RWL0_junc x13/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7264 RBL0_20 RWL_15 x111/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7265 x28/junc1 WWL_24 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7266 VDD x912/junc0 x912/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7267 x313/RWL1_junc RWL_14 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7268 x53/junc0 x53/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7269 WBL_4 WWL_31 x387/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7270 x314/RWL1_junc RWL_22 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7271 x951/RWL0_junc x951/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7272 x438/junc0 x438/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7273 x568/junc0 x568/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7274 GND x410/junc0 x410/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7275 GND x607/junc1 x607/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7276 WBL_12 WWL_10 x49/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7277 GND x397/junc1 x397/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7278 WBL_3 WWL_18 x51/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7279 GND x398/junc1 x398/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7280 x165/RWL0_junc x165/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7281 GND x825/junc1 x825/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7282 VDD x163/junc0 x163/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7283 VDD x156/junc0 x156/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7284 VDD x55/junc0 x55/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7285 x43/junc0 x43/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7286 x0/junc1 WWL_28 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7287 x592/junc0 x592/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7288 x48/RWL0_junc x48/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7289 GND x417/junc0 x417/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7290 x406/RWL0_junc x406/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7291 GND x686/junc0 x686/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7292 x915/junc0 x915/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7293 x256/junc1 WWL_5 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7294 WBL_27 WWL_8 x64/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7295 x167/junc0 x167/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7296 VDD x60/junc0 x60/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7297 x835/junc0 x835/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7298 x164/junc0 x164/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7299 x601/junc0 x601/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7300 x95/junc0 x95/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7301 GND x426/junc0 x426/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7302 GND x862/junc0 x862/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7303 x868/RWL1_junc RWL_19 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7304 x458/junc0 x458/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7305 RBL0_14 RWL_10 x179/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7306 x659/junc1 WWL_17 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7307 WBL_21 WWL_14 x80/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7308 x72/junc1 WWL_31 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7309 RBL0_5 RWL_18 x970/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7310 x62/junc0 x62/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7311 x65/RWL0_junc x65/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7312 GND x12/junc1 x12/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7313 x341/RWL1_junc RWL_17 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7314 x492/junc1 WWL_7 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7315 x665/junc1 WWL_11 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7316 x67/RWL0_junc x67/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7317 x342/RWL1_junc RWL_25 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7318 x954/RWL0_junc x954/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7319 RBL0_29 RWL_8 x971/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7320 x976/junc0 x976/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7321 RBL0_28 RWL_12 x907/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7322 x697/RWL0_junc x697/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7323 VDD x89/junc0 x89/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7324 RBL0_20 RWL_16 x736/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7325 x357/RWL1_junc RWL_15 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7326 x358/RWL1_junc RWL_23 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7327 VDD x833/junc0 x833/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7328 x469/junc0 x469/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7329 VDD x99/junc0 x99/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7330 GND x604/junc0 x604/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7331 WBL_8 WWL_15 x952/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7332 GND x448/junc0 x448/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7333 WBL_12 WWL_11 x106/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7334 GND x242/junc1 x242/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7335 VDD x199/junc0 x199/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7336 x878/RWL1_junc RWL_21 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7337 x439/RWL0_junc x439/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7338 x440/RWL0_junc x440/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7339 VDD x108/junc0 x108/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7340 x96/junc0 x96/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7341 VDD x109/junc0 x109/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7342 x871/RWL1_junc RWL_10 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7343 x100/junc0 x100/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7344 x624/junc0 x624/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7345 GND x706/junc0 x706/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7346 WBL_6 WWL_17 x120/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7347 VDD x116/junc0 x116/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7348 x481/junc0 x481/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7349 x105/RWL0_junc x105/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7350 x375/RWL1_junc RWL_0 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7351 x211/junc0 x211/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7352 x845/junc0 x845/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7353 WBL_17 WWL_19 x569/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7354 WBL_25 WWL_15 x566/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7355 x681/junc1 WWL_3 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7356 x512/junc1 WWL_10 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7357 x657/junc1 WWL_14 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7358 x488/junc0 x488/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7359 RBL0_14 RWL_11 x220/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7360 x682/junc1 WWL_18 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7361 RBL0_5 RWL_19 x785/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7362 x654/RWL1_junc RWL_31 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7363 WBL_28 WWL_29 x822/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7364 GND x1021/junc0 x1021/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7365 VDD x670/junc0 x670/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7366 GND x66/junc1 x66/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7367 GND x68/junc1 x68/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7368 x392/RWL1_junc RWL_18 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7369 x521/junc1 WWL_8 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7370 x395/RWL1_junc RWL_26 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7371 x963/RWL0_junc x963/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7372 GND x563/junc1 x563/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7373 x400/RWL1_junc RWL_20 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7374 x322/junc1 WWL_22 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7375 x464/RWL0_junc x464/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7376 x404/RWL1_junc RWL_16 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7377 x138/RWL0_junc x138/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7378 x132/junc0 x132/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7379 x978/junc0 x978/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7380 VDD x150/junc0 x150/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7381 WBL_8 WWL_16 x959/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7382 RBL0_2 RWL_0 x60/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7383 x967/RWL0_junc x967/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7384 WBL_1 WWL_30 x506/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7385 x33/junc0 x33/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7386 VDD x1006/junc0 x1006/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7387 x478/RWL1_junc RWL_22 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7388 x470/RWL0_junc x470/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7389 GND x479/junc0 x479/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7390 x886/RWL1_junc RWL_11 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7391 GND x633/junc0 x633/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7392 WBL_0 WWL_17 x43/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7393 x39/junc0 x39/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7394 x784/junc0 x784/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7395 WBL_2 WWL_22 x592/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7396 VDD x187/junc0 x187/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7397 GND x98/junc1 x98/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7398 GND x728/junc0 x728/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7399 WBL_6 WWL_18 x167/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7400 x419/RWL1_junc RWL_1 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7401 VDD x170/junc0 x170/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7402 WBL_26 WWL_12 x835/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7403 x733/RWL0_junc x733/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7404 x340/junc1 WWL_15 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7405 WBL_25 WWL_16 x601/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7406 VDD x171/junc0 x171/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7407 WBL_17 WWL_20 x95/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7408 x550/junc1 WWL_4 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7409 x551/junc1 WWL_11 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7410 RBL0_14 RWL_12 x9/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7411 x651/junc0 x651/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7412 GND x1022/junc0 x1022/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7413 x427/RWL1_junc RWL_9 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7414 VDD x1023/junc0 x1023/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7415 VDD x883/junc0 x883/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7416 GND x119/junc1 x119/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7417 GND x123/junc1 x123/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7418 x437/RWL1_junc RWL_19 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7419 GND x740/junc0 x740/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7420 x179/RWL0_junc x179/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7421 VDD x189/junc0 x189/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7422 x712/junc1 WWL_19 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7423 x363/junc1 WWL_15 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7424 GND x745/junc1 x745/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7425 x364/junc1 WWL_23 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7426 RBL0_19 RWL_20 x290/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7427 x181/junc0 x181/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7428 x203/RWL1_junc RWL_28 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7429 x717/junc1 WWL_0 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7430 RBL0_2 RWL_1 x116/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7431 x971/RWL0_junc x971/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7432 x538/junc0 x538/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7433 x444/RWL1_junc RWL_27 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7434 WBL_1 WWL_31 x607/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7435 x1014/junc0 x1014/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7436 x667/junc0 x667/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7437 x294/junc0 x294/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7438 x510/RWL1_junc RWL_23 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7439 GND x511/junc0 x511/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7440 x451/RWL1_junc RWL_4 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7441 RBL0_11 RWL_28 x973/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7442 WBL_0 WWL_18 x100/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7443 WBL_11 WWL_15 x843/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7444 x940/junc0 x940/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7445 x499/RWL1_junc RWL_12 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7446 WBL_2 WWL_23 x624/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7447 RBL0_1 RWL_13 x502/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7448 GND x147/junc1 x147/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7449 GND x24/junc0 x24/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7450 x198/RWL0_junc x198/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7451 x250/junc1 WWL_29 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7452 GND x747/junc0 x747/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7453 VDD x215/junc0 x215/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7454 x383/junc1 WWL_16 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7455 GND x160/junc1 x160/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7456 VDD x860/junc0 x860/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7457 WBL_26 WWL_13 x845/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7458 x210/junc0 x210/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7459 WBL_29 WWL_25 x629/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7460 GND x897/junc0 x897/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7461 VDD x1002/junc0 x1002/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7462 x709/junc0 x709/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7463 x730/junc1 WWL_22 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7464 RBL0_19 RWL_9 x315/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7465 GND x166/junc1 x166/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7466 RBL0_18 RWL_13 x934/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7467 GND x750/junc0 x750/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7468 x522/RWL0_junc x522/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7469 x523/RWL0_junc x523/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7470 x220/RWL0_junc x220/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7471 VDD x237/junc0 x237/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7472 x673/junc0 x673/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7473 x595/junc1 WWL_20 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7474 x407/junc1 WWL_16 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7475 GND x354/junc1 x354/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7476 x734/junc1 WWL_24 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7477 x325/junc0 x325/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7478 x174/RWL1_junc RWL_30 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7479 GND x753/junc0 x753/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7480 x250/RWL1_junc RWL_29 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7481 GND x543/junc0 x543/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7482 x738/junc1 WWL_1 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7483 x906/RWL1_junc RWL_20 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7484 x575/junc0 x575/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7485 x707/junc0 x707/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7486 x574/junc0 x574/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7487 x330/junc0 x330/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7488 GND x547/junc0 x547/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7489 x236/junc0 x236/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7490 x332/junc0 x332/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7491 WBL_22 WWL_6 x33/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7492 GND x192/junc1 x192/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7493 RBL0_7 RWL_30 x487/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7494 x739/junc0 x739/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7495 x477/RWL1_junc RWL_5 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7496 RBL0_10 RWL_6 x102/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7497 RBL0_11 RWL_29 x999/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7498 x23/junc0 x23/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7499 WBL_11 WWL_16 x39/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7500 WBL_2 WWL_24 x784/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7501 x245/RWL0_junc x245/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7502 x659/RWL1_junc RWL_17 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7503 x864/junc0 x864/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7504 GND x487/junc1 x487/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7505 VDD x726/junc0 x726/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7506 GND x761/junc0 x761/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7507 x486/RWL1_junc RWL_13 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7508 VDD x262/junc0 x262/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7509 GND x204/junc1 x204/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7510 x492/RWL1_junc RWL_7 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7511 WBL_29 WWL_26 x651/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7512 x27/junc1 WWL_22 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7513 RBL0_23 RWL_10 x189/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7514 x0/RWL1_junc RWL_28 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7515 x746/junc1 WWL_23 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7516 VDD x273/junc0 x273/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7517 VDD x282/junc0 x282/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7518 x789/RWL1_junc RWL_9 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7519 GND x769/junc0 x769/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7520 x559/RWL0_junc x559/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7521 x560/RWL0_junc x560/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7522 x598/junc0 x598/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7523 x9/RWL0_junc x9/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7524 x600/junc0 x600/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7525 RBL0_17 RWL_28 x509/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7526 x692/junc0 x692/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7527 x61/junc0 x61/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7528 x366/junc0 x366/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7529 GND x311/junc1 x311/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7530 GND x221/junc1 x221/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7531 WBL_14 WWL_28 x156/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7532 VDD x278/junc0 x278/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7533 GND x771/junc0 x771/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7534 GND x224/junc1 x224/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7535 x695/junc0 x695/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7536 x729/junc0 x729/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7537 x949/junc0 x949/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7538 GND x579/junc0 x579/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7539 x373/junc0 x373/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7540 WBL_30 WWL_3 x667/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7541 x286/junc0 x286/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7542 x73/junc0 x73/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7543 WBL_22 WWL_7 x294/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7544 GND x235/junc1 x235/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7545 x290/RWL0_junc x290/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7546 x35/RWL0_junc x35/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7547 GND x588/junc0 x588/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7548 x512/RWL1_junc RWL_10 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7549 GND x586/junc0 x586/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7550 x875/junc0 x875/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7551 x682/RWL1_junc RWL_18 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7552 GND x248/junc1 x248/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7553 VDD x490/junc0 x490/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7554 x20/junc1 WWL_2 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7555 GND x249/junc1 x249/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7556 x618/RWL0_junc x618/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7557 GND x783/junc0 x783/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7558 x293/junc0 x293/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7559 GND x252/junc1 x252/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7560 RBL0_4 RWL_13 x396/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7561 x774/RWL0_junc x774/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7562 x521/RWL1_junc RWL_8 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7563 GND x653/junc0 x653/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7564 x756/junc1 WWL_6 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7565 x757/junc1 WWL_10 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7566 x81/junc1 WWL_23 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7567 x622/junc0 x622/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7568 RBL0_24 RWL_7 x985/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7569 RBL0_23 RWL_11 x237/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7570 WBL_29 WWL_27 x210/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7571 VDD x306/junc0 x306/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7572 x54/RWL1_junc RWL_29 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7573 x303/junc1 WWL_24 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7574 VDD x952/junc0 x952/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7575 x425/junc0 x425/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7576 x530/RWL1_junc RWL_14 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7577 VDD x317/junc0 x317/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7578 x18/junc0 x18/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7579 x216/junc0 x216/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7580 GND x794/junc0 x794/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7581 x21/junc0 x21/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7582 x715/junc0 x715/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7583 x410/junc0 x410/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7584 GND x609/junc0 x609/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7585 RBL0_17 RWL_29 x544/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7586 WBL_10 WWL_30 x199/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7587 WBL_7 WWL_10 x325/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7588 GND x272/junc1 x272/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7589 GND x1005/junc1 x1005/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7590 GND x542/junc1 x542/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7591 GND x274/junc1 x274/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7592 x315/RWL0_junc x315/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7593 RBL0_31 RWL_27 x257/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7594 VDD x415/junc0 x415/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7595 x37/junc0 x37/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7596 WBL_31 WWL_0 x330/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7597 RBL0_15 RWL_4 x397/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7598 x127/junc0 x127/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7599 WBL_30 WWL_4 x236/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7600 x480/junc1 WWL_5 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7601 WBL_22 WWL_8 x332/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7602 RBL0_28 RWL_31 x542/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7603 x240/junc0 x240/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7604 x736/junc0 x736/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7605 x550/RWL1_junc RWL_4 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7606 GND x617/junc0 x617/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7607 x551/RWL1_junc RWL_11 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7608 x926/RWL1_junc RWL_19 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7609 x775/junc1 WWL_17 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7610 x638/junc0 x638/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7611 RBL0_9 RWL_10 x429/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7612 x91/RWL0_junc x91/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7613 x331/junc0 x331/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7614 x929/RWL1_junc RWL_17 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7615 x664/junc1 WWL_7 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7616 x777/junc1 WWL_11 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7617 VDD x345/junc0 x345/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7618 x996/junc0 x996/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7619 RBL0_24 RWL_8 x990/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7620 WBL_20 WWL_28 x227/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7621 x778/junc1 WWL_24 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7622 VDD x349/junc0 x349/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7623 RBL0_23 RWL_12 x948/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7624 GND x562/junc1 x562/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7625 x566/RWL1_junc RWL_15 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7626 x741/RWL0_junc x741/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7627 x483/junc0 x483/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7628 x77/junc0 x77/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7629 x79/junc0 x79/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7630 WBL_3 WWL_15 x173/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7631 GND x807/junc0 x807/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7632 GND x631/junc0 x631/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7633 VDD x687/junc0 x687/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7634 WBL_16 WWL_3 x61/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7635 x448/junc0 x448/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7636 WBL_10 WWL_31 x1006/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7637 WBL_7 WWL_11 x366/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7638 x355/RWL0_junc x355/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7639 GND x472/junc1 x472/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7640 x11/RWL0_junc x11/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7641 VDD x369/junc0 x369/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7642 x90/junc0 x90/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7643 WBL_27 WWL_5 x181/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7644 GND x318/junc1 x318/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7645 WBL_31 WWL_1 x373/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7646 RBL0_15 RWL_5 x242/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7647 x92/junc0 x92/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7648 x910/junc0 x910/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7649 x583/RWL1_junc RWL_12 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7650 x370/junc0 x370/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7651 x584/RWL1_junc RWL_5 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7652 x31/junc1 WWL_10 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7653 x772/junc1 WWL_14 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7654 x661/junc0 x661/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7655 RBL0_9 RWL_11 x462/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7656 x796/junc1 WWL_18 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7657 x142/RWL0_junc x142/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7658 WBL_7 WWL_29 x883/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7659 GND x814/junc0 x814/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7660 RBL0_6 RWL_31 x394/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7661 x466/junc0 x466/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7662 VDD x389/junc0 x389/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7663 GND x820/junc0 x820/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7664 GND x333/junc1 x333/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7665 GND x819/junc0 x819/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7666 x938/RWL1_junc RWL_18 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7667 x44/junc1 WWL_8 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7668 x401/RWL0_junc x401/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7669 GND x336/junc1 x336/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7670 VDD x399/junc0 x399/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7671 x768/junc1 WWL_30 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7672 x595/RWL1_junc RWL_20 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7673 RBL0_27 RWL_21 x901/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7674 x644/RWL0_junc x644/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7675 GND x604/junc1 x604/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7676 x385/RWL0_junc x385/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7677 x515/RWL0_junc x515/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7678 VDD x531/junc0 x531/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7679 x601/RWL1_junc RWL_16 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7680 x396/RWL0_junc x396/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7681 x801/junc0 x801/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7682 WBL_3 WWL_16 x216/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7683 x985/RWL0_junc x985/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7684 VDD x708/junc0 x708/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7685 WBL_16 WWL_4 x410/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7686 x994/junc0 x994/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7687 x69/RWL0_junc x69/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7688 x270/junc0 x270/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7689 GND x658/junc0 x658/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7690 x312/junc0 x312/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7691 GND x359/junc1 x359/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7692 GND x361/junc1 x361/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7693 RBL0_20 RWL_2 x98/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7694 VDD x421/junc0 x421/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7695 WBL_21 WWL_12 x240/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7696 VDD x485/junc0 x485/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7697 x554/junc1 WWL_15 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7698 x414/junc0 x414/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7699 x88/junc1 WWL_11 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7700 RBL0_9 RWL_12 x202/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7701 x765/junc0 x765/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7702 GND x826/junc0 x826/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7703 x831/junc1 WWL_5 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7704 x183/junc1 WWL_9 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7705 x619/RWL1_junc RWL_9 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7706 RBL0_12 RWL_24 x497/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7707 VDD x432/junc0 x432/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7708 GND x374/junc1 x374/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7709 x704/junc0 x704/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7710 x674/RWL1_junc RWL_19 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7711 x760/junc0 x760/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7712 x662/RWL0_junc x662/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7713 GND x109/junc0 x109/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7714 x429/RWL0_junc x429/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7715 x244/junc1 WWL_31 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7716 VDD x722/junc0 x722/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7717 VDD x438/junc0 x438/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7718 RBL0_27 RWL_22 x556/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7719 VDD x724/junc0 x724/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7720 x112/RWL0_junc x112/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7721 x537/junc1 WWL_30 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7722 WBL_12 WWL_9 x483/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7723 x990/RWL0_junc x990/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7724 x696/junc0 x696/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7725 VDD x821/junc0 x821/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7726 x788/junc0 x788/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7727 GND x633/junc1 x633/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7728 x997/junc0 x997/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7729 x780/junc0 x780/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7730 x308/junc0 x308/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7731 x781/junc0 x781/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7732 x30/RWL1_junc RWL_6 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7733 GND x678/junc0 x678/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7734 WBL_6 WWL_15 x275/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7735 GND x405/junc1 x405/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7736 GND x406/junc1 x406/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7737 x445/RWL0_junc x445/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7738 RBL0_2 RWL_31 x633/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7739 GND x832/junc0 x832/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7740 x585/junc1 WWL_12 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7741 x520/junc0 x520/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7742 RBL0_20 x61/RWL1 x147/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7743 VDD x458/junc0 x458/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7744 x587/junc1 WWL_16 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7745 GND x411/junc1 x411/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7746 WBL_21 WWL_13 x910/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7747 x455/junc0 x455/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7748 WBL_24 WWL_25 x209/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7749 x643/RWL1_junc RWL_2 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7750 GND x834/junc0 x834/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7751 WBL_28 WWL_21 x466/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7752 VDD x976/junc0 x976/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7753 RBL0_12 RWL_25 x531/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7754 GND x418/junc1 x418/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7755 x1015/junc0 x1015/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7756 x688/RWL0_junc x688/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7757 GND x836/junc0 x836/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7758 GND x837/junc0 x837/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7759 VDD x468/junc0 x468/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7760 x46/RWL0_junc x46/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7761 x462/RWL0_junc x462/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7762 VDD x922/junc0 x922/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7763 VDD x469/junc0 x469/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7764 x784/junc0 x784/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7765 RBL0_27 RWL_23 x589/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7766 VDD x923/junc0 x923/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7767 x539/junc0 x539/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7768 GND x838/junc0 x838/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7769 x555/junc1 WWL_31 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7770 RBL0_30 RWL_21 x546/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7771 x947/RWL1_junc RWL_20 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7772 x219/junc0 x219/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7773 x803/junc0 x803/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7774 x718/junc0 x718/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7775 x547/junc0 x547/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7776 GND x701/junc0 x701/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7777 x41/junc0 x41/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7778 x471/junc0 x471/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7779 x350/junc0 x350/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7780 WBL_15 WWL_22 x994/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7781 WBL_0 WWL_15 x238/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7782 WBL_17 WWL_6 x270/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7783 RBL0_1 RWL_10 x598/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7784 GND x440/junc1 x440/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7785 x828/junc0 x828/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7786 RBL0_5 RWL_6 x284/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7787 WBL_6 WWL_16 x312/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7788 GND x442/junc1 x442/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7789 x268/RWL0_junc x268/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7790 x775/RWL1_junc RWL_17 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7791 VDD x484/junc0 x484/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7792 GND x841/junc0 x841/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7793 x180/junc1 WWL_2 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7794 x182/junc1 WWL_9 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7795 x660/RWL1_junc RWL_13 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7796 x264/junc1 WWL_13 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7797 VDD x488/junc0 x488/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7798 GND x758/junc1 x758/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7799 GND x450/junc1 x450/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7800 x302/junc1 WWL_29 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7801 x664/RWL1_junc RWL_7 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7802 VDD x647/junc0 x647/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7803 GND x752/junc0 x752/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7804 WBL_24 WWL_26 x765/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7805 RBL0_18 RWL_10 x438/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7806 x667/RWL1_junc x389/RWL1 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7807 RBL0_12 RWL_26 x568/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7808 VDD x126/junc0 x126/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7809 WBL_8 WWL_3 x331/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7810 x142/junc0 x142/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7811 x188/junc0 x188/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7812 GND x846/junc0 x846/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7813 x165/RWL1_junc RWL_9 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7814 GND x847/junc0 x847/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7815 VDD x132/junc0 x132/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7816 x103/RWL0_junc x103/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7817 x202/RWL0_junc x202/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7818 x259/junc0 x259/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7819 x802/junc0 x802/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7820 x424/junc0 x424/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7821 x576/junc0 x576/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7822 GND x848/junc0 x848/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7823 x630/junc1 WWL_25 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7824 RBL0_30 RWL_22 x310/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7825 x267/junc0 x267/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7826 x823/junc0 x823/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7827 x979/junc0 x979/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7828 x579/junc0 x579/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7829 GND x721/junc0 x721/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7830 x297/RWL1_junc RWL_30 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7831 WBL_25 WWL_3 x780/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7832 x503/junc0 x503/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7833 WBL_15 WWL_23 x997/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7834 WBL_0 WWL_16 x781/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7835 x337/junc0 x337/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7836 WBL_17 WWL_7 x308/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7837 RBL0_1 RWL_11 x21/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7838 GND x470/junc1 x470/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7839 x31/RWL1_junc RWL_10 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7840 x1015/RWL1_junc RWL_31 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7841 x217/RWL0_junc x217/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7842 GND x727/junc0 x727/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7843 RBL0_13 RWL_30 x755/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7844 x796/RWL1_junc RWL_18 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7845 RBL0_19 RWL_30 x790/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7846 GND x473/junc1 x473/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7847 VDD x519/junc0 x519/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7848 x684/RWL1_junc RWL_6 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7849 GND x474/junc1 x474/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7850 x745/RWL0_junc x745/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7851 GND x853/junc0 x853/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7852 WBL_16 WWL_30 x744/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7853 GND x779/junc1 x779/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7854 x816/junc0 x816/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7855 GND x476/junc1 x476/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7856 x228/junc1 WWL_6 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7857 x44/RWL1_junc RWL_8 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7858 GND x402/junc0 x402/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7859 x840/junc1 WWL_10 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7860 GND x764/junc0 x764/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7861 WBL_24 WWL_27 x455/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7862 RBL0_19 RWL_7 x596/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7863 RBL0_18 RWL_11 x469/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7864 GND x53/junc1 x53/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7865 VDD x173/junc0 x173/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7866 WBL_8 WWL_4 x207/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7867 x194/junc0 x194/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7868 x56/RWL1_junc RWL_14 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7869 VDD x533/junc0 x533/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7870 GND x855/junc0 x855/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7871 x299/junc0 x299/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7872 GND x857/junc0 x857/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7873 VDD x181/junc0 x181/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7874 x817/junc0 x817/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7875 x609/junc0 x609/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7876 GND x742/junc0 x742/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7877 WBL_2 WWL_10 x539/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7878 x652/junc1 WWL_26 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7879 VDD x538/junc0 x538/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7880 RBL0_26 RWL_27 x481/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7881 VDD x612/junc0 x612/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7882 x1018/junc0 x1018/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7883 x643/junc0 x643/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7884 x307/junc0 x307/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7885 VDD x773/junc0 x773/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7886 RBL0_30 RWL_23 x351/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7887 x656/junc1 WWL_3 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7888 WBL_26 WWL_28 x754/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7889 WBL_26 WWL_0 x547/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7890 WBL_25 WWL_4 x471/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7891 RBL0_10 RWL_4 x1005/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7892 WBL_15 WWL_24 x41/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7893 x379/junc0 x379/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7894 WBL_17 WWL_8 x350/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7895 RBL0_1 RWL_12 x79/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7896 x319/junc0 x319/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7897 GND x956/junc0 x956/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7898 GND x505/junc1 x505/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7899 GND x866/junc0 x866/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7900 x88/RWL1_junc RWL_11 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7901 GND x507/junc1 x507/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7902 x195/RWL1_junc RWL_19 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7903 RBL0_4 RWL_10 x620/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7904 GND x508/junc1 x508/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7905 x858/RWL0_junc x858/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7906 x354/RWL0_junc x354/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7907 WBL_16 WWL_31 x553/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7908 GND x157/junc1 x157/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7909 x234/junc0 x234/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7910 x670/junc1 WWL_3 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7911 x965/RWL1_junc RWL_17 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7912 x281/junc1 WWL_7 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7913 x852/junc1 WWL_11 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7914 VDD x22/junc0 x22/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7915 RBL0_19 RWL_8 x626/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7916 RBL0_18 RWL_12 x978/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7917 x649/junc1 WWL_30 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7918 GND x713/junc1 x713/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7919 GND x924/junc0 x924/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7920 x967/RWL1_junc RWL_7 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7921 x937/junc0 x937/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7922 x111/RWL1_junc RWL_15 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7923 GND x117/junc1 x117/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7924 x76/junc0 x76/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7925 GND x522/junc1 x522/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7926 x339/junc0 x339/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7927 GND x7/junc0 x7/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7928 x631/junc0 x631/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7929 GND x751/junc0 x751/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7930 VDD x40/junc0 x40/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7931 WBL_11 WWL_3 x424/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7932 WBL_2 WWL_11 x576/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7933 x567/RWL0_junc x567/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7934 x854/junc1 WWL_27 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7935 VDD x574/junc0 x574/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7936 x570/junc0 x570/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7937 x572/junc0 x572/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7938 WBL_22 WWL_5 x433/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7939 GND x873/junc0 x873/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7940 WBL_22 WWL_30 x770/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7941 x856/junc1 WWL_4 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7942 WBL_26 WWL_1 x579/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7943 GND x536/junc1 x536/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7944 RBL0_10 RWL_5 x472/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7945 x363/junc0 x363/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7946 RBL0_13 RWL_17 x941/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7947 GND x540/junc1 x540/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7948 WBL_20 WWL_21 x283/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7949 x305/junc1 WWL_10 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7950 x725/RWL1_junc RWL_12 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7951 x578/junc0 x578/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7952 RBL0_4 RWL_11 x645/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7953 x870/RWL0_junc x870/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7954 x311/RWL0_junc x311/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7955 GND x879/junc0 x879/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7956 x648/junc0 x648/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7957 VDD x74/junc0 x74/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7958 GND x882/junc0 x882/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7959 GND x548/junc1 x548/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7960 GND x881/junc0 x881/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7961 x1023/junc1 WWL_4 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7962 x970/RWL1_junc RWL_18 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7963 x320/junc1 WWL_8 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7964 VDD x594/junc0 x594/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7965 x597/RWL0_junc x597/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7966 GND x810/junc1 x810/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7967 x3/junc1 WWL_31 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7968 RBL0_22 RWL_21 x1014/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7969 x377/junc0 x377/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7970 x971/RWL1_junc RWL_8 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7971 x987/junc0 x987/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7972 GND x164/junc1 x164/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7973 VDD x599/junc0 x599/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7974 x736/RWL1_junc RWL_16 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7975 VDD x692/junc0 x692/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7976 x128/junc0 x128/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7977 GND x739/junc1 x739/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7978 x13/junc1 WWL_28 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7979 GND x559/junc1 x559/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7980 x596/RWL0_junc x596/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7981 VDD x93/junc0 x93/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7982 WBL_11 WWL_4 x609/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7983 x593/RWL0_junc x593/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7984 x97/junc0 x97/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7985 x335/RWL0_junc x335/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7986 GND x772/junc0 x772/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7987 x602/junc0 x602/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7988 VDD x73/junc0 x73/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7989 WBL_30 WWL_2 x643/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7990 GND x571/junc1 x571/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7991 WBL_22 WWL_31 x654/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7992 x884/RWL0_junc x884/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7993 x885/RWL0_junc x885/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7994 x871/junc1 WWL_10 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7995 VDD x114/junc0 x114/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M7996 RBL0_13 RWL_18 x946/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7997 x706/junc1 WWL_15 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7998 WBL_29 WWL_14 x319/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M7999 GND x577/junc1 x577/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8000 x611/junc0 x611/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8001 x348/junc1 WWL_11 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8002 RBL0_4 RWL_12 x449/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8003 x123/junc0 x123/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8004 x352/RWL0_junc x352/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8005 GND x889/junc0 x889/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8006 GND x890/junc0 x890/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8007 x895/junc1 WWL_5 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8008 x26/junc1 WWL_9 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8009 RBL0_7 RWL_24 x673/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8010 x1/junc0 x1/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8011 VDD x622/junc0 x622/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8012 GND x580/junc1 x580/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8013 GND x774/junc1 x774/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8014 x129/junc0 x129/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8015 GND x581/junc1 x581/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8016 x785/RWL1_junc RWL_19 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8017 x5/junc0 x5/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8018 x279/RWL0_junc x279/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8019 VDD x135/junc0 x135/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8020 x878/junc1 WWL_21 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8021 x620/RWL0_junc x620/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8022 VDD x137/junc0 x137/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8023 RBL0_31 RWL_14 x575/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8024 x809/junc0 x809/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8025 RBL0_22 RWL_22 x707/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8026 x14/junc0 x14/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8027 VDD x709/junc0 x709/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8028 x67/junc1 WWL_30 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8029 WBL_7 WWL_9 x76/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8030 x625/RWL0_junc x625/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8031 x626/RWL0_junc x626/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8032 x84/RWL0_junc x84/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8033 VDD x880/junc0 x880/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8034 x804/junc0 x804/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8035 x71/RWL0_junc x71/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8036 x147/junc0 x147/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8037 x151/junc0 x151/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8038 GND x795/junc0 x795/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8039 x304/RWL1_junc RWL_6 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8040 WBL_14 WWL_17 x570/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8041 VDD x127/junc0 x127/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8042 GND x603/junc1 x603/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8043 x388/RWL0_junc x388/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8044 x465/RWL0_junc x465/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8045 GND x896/junc0 x896/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8046 x899/junc0 x899/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8047 x886/junc1 WWL_11 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8048 x726/junc1 WWL_12 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8049 RBL0_13 RWL_19 x48/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8050 VDD x638/junc0 x638/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8051 x728/junc1 WWL_16 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8052 GND x792/junc1 x792/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8053 x166/junc0 x166/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8054 x636/junc0 x636/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8055 WBL_19 WWL_25 x68/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8056 x759/RWL1_junc RWL_2 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8057 GND x898/junc0 x898/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8058 x49/junc0 x49/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8059 GND x900/junc0 x900/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8060 RBL0_16 RWL_17 x600/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8061 VDD x864/junc0 x864/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8062 WBL_23 WWL_21 x648/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8063 x51/junc0 x51/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8064 VDD x996/junc0 x996/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8065 GND x614/junc1 x614/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8066 x105/junc1 WWL_28 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8067 RBL0_7 RWL_25 x692/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8068 x57/junc0 x57/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8069 GND x615/junc1 x615/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8070 x453/junc0 x453/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8071 x288/RWL1_junc RWL_28 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8072 x798/RWL0_junc x798/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8073 x1016/RWL1_junc RWL_24 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8074 GND x154/junc0 x154/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8075 x321/RWL0_junc x321/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8076 VDD x186/junc0 x186/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8077 x645/RWL0_junc x645/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8078 x981/junc0 x981/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8079 VDD x960/junc0 x960/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8080 VDD x185/junc0 x185/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8081 RBL0_31 RWL_15 x695/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8082 RBL0_22 RWL_23 x729/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8083 VDD x671/junc0 x671/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8084 x122/junc1 WWL_31 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8085 WBL_16 WWL_2 x128/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8086 x650/RWL0_junc x650/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8087 RBL0_25 RWL_21 x700/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8088 x824/junc0 x824/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8089 x80/junc0 x80/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8090 x701/junc0 x701/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8091 x34/junc0 x34/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8092 x371/junc0 x371/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8093 RBL0_24 RWL_31 x604/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8094 WBL_10 WWL_22 x97/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8095 GND x11/junc1 x11/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8096 GND x808/junc0 x808/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8097 WBL_14 WWL_18 x602/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8098 x336/RWL0_junc x336/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8099 x1008/RWL0_junc x1008/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8100 GND x628/junc1 x628/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8101 x204/junc0 x204/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8102 x430/RWL0_junc x430/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8103 RBL0_20 RWL_0 x440/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8104 x431/RWL0_junc x431/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8105 GND x904/junc0 x904/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8106 GND x905/junc0 x905/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8107 VDD x370/junc0 x370/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8108 x434/junc1 WWL_9 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8109 x490/junc1 WWL_13 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8110 VDD x661/junc0 x661/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8111 GND x679/junc1 x679/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8112 x145/junc1 WWL_29 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8113 x281/RWL1_junc RWL_7 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8114 x711/junc0 x711/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8115 VDD x666/junc0 x666/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8116 GND x288/junc1 x288/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8117 WBL_19 WWL_26 x123/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8118 GND x907/junc0 x907/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8119 x780/RWL1_junc x389/RWL1 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8120 x106/junc0 x106/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8121 RBL0_16 RWL_18 x18/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8122 GND x637/junc1 x637/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8123 RBL0_7 RWL_26 x715/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8124 x110/junc0 x110/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8125 GND x821/junc0 x821/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8126 WBL_3 WWL_3 x129/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8127 x480/junc0 x480/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8128 x801/RWL1_junc RWL_29 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8129 VDD x968/junc0 x968/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8130 GND x401/junc1 x401/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8131 RBL0_27 RWL_20 x962/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8132 x564/RWL1_junc RWL_25 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8133 GND x6/junc0 x6/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8134 x668/RWL0_junc x668/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8135 VDD x390/junc0 x390/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8136 x365/RWL0_junc x365/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8137 x449/RWL0_junc x449/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8138 x604/junc0 x604/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8139 VDD x497/junc0 x497/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8140 x120/junc0 x120/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8141 RBL0_31 RWL_16 x37/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8142 x226/junc0 x226/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8143 GND x644/junc1 x644/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8144 x750/junc1 WWL_25 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8145 x901/junc1 WWL_21 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8146 RBL0_25 RWL_22 x47/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8147 x131/junc0 x131/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8148 x856/RWL1_junc RWL_4 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8149 x1000/junc0 x1000/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8150 x721/junc0 x721/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8151 x1017/junc0 x1017/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8152 WBL_10 WWL_23 x151/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8153 x305/RWL1_junc RWL_10 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8154 x252/junc0 x252/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8155 x250/junc0 x250/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8156 RBL0_20 RWL_1 x470/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8157 x54/junc0 x54/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8158 x136/junc0 x136/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8159 GND x912/junc0 x912/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8160 x102/RWL1_junc RWL_6 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8161 x1016/RWL0_junc x1016/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8162 GND x913/junc0 x913/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8163 VDD x414/junc0 x414/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8164 x53/junc0 x53/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8165 GND x702/junc1 x702/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8166 x316/RWL1_junc RWL_0 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8167 x761/junc1 WWL_22 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8168 VDD x258/junc0 x258/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8169 x320/RWL1_junc RWL_8 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8170 RBL0_27 RWL_9 x266/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8171 RBL0_29 RWL_28 x632/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8172 WBL_28 WWL_19 x166/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8173 WBL_19 WWL_27 x636/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8174 GND x801/junc1 x801/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8175 x159/junc0 x159/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8176 RBL0_16 RWL_19 x77/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8177 GND x163/junc0 x163/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8178 WBL_3 WWL_4 x453/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8179 GND x156/junc0 x156/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8180 x425/RWL1_junc RWL_31 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8181 x41/junc0 x41/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8182 VDD x972/junc0 x972/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8183 x43/junc0 x43/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8184 VDD x693/junc0 x693/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8185 x517/junc0 x517/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8186 GND x662/junc1 x662/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8187 x272/junc0 x272/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8188 x527/RWL1_junc RWL_26 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8189 GND x247/junc0 x247/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8190 x545/RWL0_junc x545/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8191 x167/junc0 x167/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8192 GND x60/junc0 x60/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8193 VDD x433/junc0 x433/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8194 x742/junc0 x742/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8195 GND x669/junc1 x669/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8196 RBL0_20 RWL_31 x842/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8197 x411/RWL0_junc x411/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8198 x164/junc0 x164/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8199 x769/junc1 WWL_26 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8200 VDD x788/junc0 x788/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8201 VDD x696/junc0 x696/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8202 RBL0_21 RWL_27 x92/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8203 x95/junc0 x95/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8204 x759/junc0 x759/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8205 VDD x287/junc0 x287/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8206 RBL0_25 RWL_23 x101/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8207 x177/junc0 x177/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8208 x869/RWL1_junc RWL_5 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8209 x771/junc1 WWL_3 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8210 WBL_21 WWL_0 x701/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8211 RBL0_5 RWL_4 x104/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8212 WBL_10 WWL_24 x34/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8213 x699/junc0 x699/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8214 GND x920/junc0 x920/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8215 GND x15/junc1 x15/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8216 GND x89/junc0 x89/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8217 x348/RWL1_junc RWL_11 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8218 x489/junc0 x489/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8219 WBL_13 WWL_22 x204/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8220 GND x675/junc1 x675/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8221 GND x17/junc1 x17/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8222 x917/RWL0_junc x917/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8223 GND x921/junc0 x921/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8224 x564/RWL0_junc x564/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8225 x829/RWL0_junc x829/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8226 x713/junc0 x713/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8227 GND x833/junc0 x833/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8228 x360/RWL1_junc RWL_1 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8229 VDD x975/junc0 x975/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8230 RBL0_29 RWL_29 x504/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8231 x783/junc1 WWL_23 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8232 WBL_28 WWL_20 x711/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8233 VDD x974/junc0 x974/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8234 VDD x300/junc0 x300/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8235 GND x199/junc0 x199/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8236 GND x200/junc0 x200/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8237 GND x208/junc0 x208/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8238 x985/RWL1_junc RWL_7 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8239 x368/RWL1_junc RWL_27 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8240 x96/junc0 x96/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8241 VDD x714/junc0 x714/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8242 x134/junc0 x134/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8243 x100/junc0 x100/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8244 GND x372/junc1 x372/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8245 GND x688/junc1 x688/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8246 x710/junc0 x710/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8247 x552/junc0 x552/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8248 x338/junc0 x338/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8249 x213/junc0 x213/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8250 GND x116/junc0 x116/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8251 x751/junc0 x751/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8252 VDD x314/junc0 x314/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8253 WBL_6 WWL_3 x226/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8254 GND x690/junc1 x690/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8255 x450/RWL0_junc x450/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8256 x20/RWL0_junc x20/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8257 x914/junc1 WWL_27 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8258 RBL0_30 RWL_20 x144/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8259 VDD x718/junc0 x718/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8260 x716/junc0 x716/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8261 WBL_17 WWL_5 x239/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8262 GND x930/junc0 x930/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8263 x909/junc1 WWL_0 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8264 x916/junc1 WWL_4 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8265 WBL_21 WWL_1 x721/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8266 GND x694/junc1 x694/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8267 RBL0_5 RWL_5 x153/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8268 x251/junc0 x251/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8269 x720/junc0 x720/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8270 RBL0_8 RWL_17 x232/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8271 GND x70/junc1 x70/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8272 x397/RWL1_junc RWL_4 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8273 x825/RWL1_junc RWL_12 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8274 WBL_13 WWL_23 x252/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8275 RBL0_12 RWL_13 x760/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8276 x928/RWL0_junc x928/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8277 x527/RWL0_junc x527/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8278 x762/junc0 x762/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8279 x72/RWL1_junc RWL_31 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8280 GND x246/junc0 x246/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8281 GND x934/junc0 x934/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8282 GND x150/junc0 x150/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8283 VDD x977/junc0 x977/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8284 x919/junc1 WWL_24 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8285 VDD x763/junc0 x763/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8286 x676/RWL0_junc x676/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8287 VDD x732/junc0 x732/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8288 x734/RWL0_junc x734/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8289 WBL_8 WWL_2 x293/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8290 RBL0_17 RWL_21 x788/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8291 x255/junc0 x255/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8292 x990/RWL1_junc RWL_8 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8293 RBL0_30 RWL_9 x183/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8294 x803/junc1 WWL_22 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8295 x148/junc0 x148/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8296 GND x416/junc1 x416/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8297 x146/junc0 x146/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8298 VDD x802/junc0 x802/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8299 x152/junc0 x152/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8300 GND x828/junc1 x828/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8301 x380/junc0 x380/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8302 x731/junc0 x731/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8303 WBL_15 WWL_10 x517/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8304 WBL_0 WWL_3 x272/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8305 x12/RWL1_junc RWL_24 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8306 x475/RWL0_junc x475/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8307 VDD x358/junc0 x358/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8308 WBL_6 WWL_4 x742/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8309 x361/junc0 x361/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8310 x78/RWL0_junc x78/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8311 x476/RWL0_junc x476/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8312 GND x171/junc0 x171/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8313 x737/junc0 x737/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8314 VDD x337/junc0 x337/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8315 WBL_25 WWL_2 x759/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8316 GND x113/junc1 x113/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8317 x915/junc1 WWL_1 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8318 GND x735/junc1 x735/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8319 x367/junc0 x367/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8320 x935/RWL0_junc x935/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8321 GND x1023/junc0 x1023/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8322 GND x124/junc1 x124/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8323 RBL0_8 RWL_18 x285/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8324 WBL_24 WWL_14 x699/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8325 GND x719/junc1 x719/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8326 x242/RWL1_junc RWL_5 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8327 WBL_13 WWL_24 x489/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8328 x561/RWL0_junc x561/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8329 GND x189/junc0 x189/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8330 WBL_18 WWL_28 x864/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8331 x524/junc0 x524/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8332 x943/junc1 WWL_5 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8333 x301/junc1 WWL_9 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8334 GND x850/junc1 x850/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8335 RBL0_2 RWL_24 x784/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8336 GND x356/junc0 x356/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8337 GND x291/junc0 x291/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8338 x292/junc0 x292/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8339 x500/RWL0_junc x500/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8340 x294/junc0 x294/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8341 VDD x393/junc0 x393/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8342 x931/junc1 WWL_21 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8343 RBL0_26 RWL_14 x219/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8344 VDD x395/junc0 x395/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8345 x1013/junc0 x1013/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8346 RBL0_17 RWL_22 x803/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8347 x823/junc1 WWL_23 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8348 x296/junc0 x296/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8349 WBL_15 WWL_11 x552/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8350 WBL_0 WWL_4 x710/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8351 x66/RWL1_junc RWL_17 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8352 WBL_2 WWL_9 x338/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8353 x68/RWL1_junc RWL_25 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8354 x901/RWL1_junc RWL_21 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8355 x125/RWL0_junc x125/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8356 VDD x404/junc0 x404/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8357 VDD x933/junc0 x933/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8358 x491/RWL0_junc x491/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8359 x324/junc0 x324/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8360 x406/junc0 x406/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8361 GND x215/junc0 x215/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8362 GND x860/junc0 x860/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8363 x634/junc1 WWL_2 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8364 x525/RWL1_junc RWL_6 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8365 WBL_9 WWL_17 x716/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8366 VDD x379/junc0 x379/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8367 GND x161/junc1 x161/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8368 GND x162/junc1 x162/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8369 x210/junc0 x210/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8370 GND x501/junc1 x501/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8371 x815/junc0 x815/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8372 x590/RWL0_junc x590/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8373 GND x1002/junc0 x1002/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8374 WBL_20 WWL_19 x1000/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8375 RBL0_8 RWL_19 x323/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8376 GND x169/junc1 x169/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8377 x149/RWL1_junc RWL_31 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8378 x428/RWL0_junc x428/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8379 x418/junc0 x418/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8380 GND x858/junc1 x858/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8381 x98/RWL1_junc RWL_2 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8382 GND x237/junc0 x237/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8383 x647/junc1 WWL_2 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8384 x325/junc0 x325/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8385 RBL0_11 RWL_17 x259/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8386 x52/junc0 x52/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8387 RBL0_2 RWL_25 x802/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8388 WBL_18 WWL_21 x762/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8389 GND x861/junc1 x861/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8390 x755/RWL0_junc x755/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8391 x329/junc0 x329/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8392 x863/RWL0_junc x863/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8393 x330/junc0 x330/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8394 x939/junc1 WWL_14 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8395 x236/junc0 x236/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8396 x768/junc0 x768/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8397 VDD x437/junc0 x437/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8398 x332/junc0 x332/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8399 VDD x983/junc0 x983/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8400 VDD x436/junc0 x436/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8401 RBL0_26 RWL_15 x267/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8402 RBL0_17 RWL_23 x823/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8403 x1016/junc1 WWL_24 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8404 WBL_11 WWL_2 x380/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8405 x119/RWL1_junc RWL_18 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8406 x556/RWL1_junc RWL_22 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8407 x172/RWL0_junc x172/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8408 x123/RWL1_junc RWL_26 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8409 VDD x188/junc0 x188/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8410 x442/junc0 x442/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8411 x534/junc0 x534/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8412 WBL_5 WWL_22 x361/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8413 GND x262/junc0 x262/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8414 x385/junc1 WWL_30 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8415 GND x872/junc0 x872/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8416 GND x206/junc1 x206/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8417 WBL_9 WWL_18 x737/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8418 x810/RWL0_junc x810/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8419 x184/RWL0_junc x184/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8420 GND x748/junc1 x748/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8421 x450/junc0 x450/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8422 WBL_29 WWL_12 x367/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8423 x621/RWL0_junc x621/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8424 x766/RWL0_junc x766/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8425 WBL_20 WWL_20 x276/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8426 GND x273/junc0 x273/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8427 VDD x578/junc0 x578/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8428 x623/junc1 WWL_9 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8429 x778/RWL0_junc x778/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8430 x812/junc0 x812/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8431 GND x870/junc1 x870/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8432 VDD x16/junc0 x16/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8433 GND x948/junc0 x948/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8434 x941/junc1 WWL_17 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8435 x147/RWL1_junc x61/RWL1 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8436 x366/junc0 x366/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8437 GND x676/junc0 x676/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8438 RBL0_11 RWL_18 x299/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8439 GND x797/junc1 x797/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8440 RBL0_2 RWL_26 x817/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8441 GND x880/junc0 x880/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8442 VDD x986/junc0 x986/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8443 x834/junc1 WWL_19 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8444 VDD x816/junc0 x816/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8445 GND x597/junc1 x597/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8446 x160/RWL1_junc RWL_21 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8447 RBL0_22 RWL_20 x1018/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8448 x373/junc0 x373/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8449 x286/junc0 x286/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8450 x244/junc0 x244/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8451 VDD x190/junc0 x190/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8452 VDD x673/junc0 x673/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8453 RBL0_26 RWL_16 x307/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8454 x837/junc1 WWL_25 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8455 WBL_5 WWL_29 x287/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8456 x589/RWL1_junc RWL_23 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8457 x166/RWL1_junc RWL_19 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8458 x1014/junc1 WWL_21 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8459 x916/RWL1_junc RWL_4 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8460 VDD x998/junc0 x998/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8461 WBL_14 WWL_15 x405/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8462 x580/RWL0_junc x580/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8463 x227/junc0 x227/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8464 WBL_5 WWL_23 x406/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8465 x428/junc1 WWL_31 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8466 x640/RWL0_junc x640/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8467 x950/RWL0_junc x950/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8468 x663/RWL0_junc x663/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8469 x476/junc0 x476/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8470 x417/junc1 WWL_9 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8471 x790/RWL0_junc x790/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8472 GND x884/junc1 x884/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8473 WBL_29 WWL_13 x815/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8474 x230/RWL0_junc x230/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8475 GND x885/junc1 x885/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8476 x284/RWL1_junc RWL_6 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8477 GND x952/junc0 x952/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8478 VDD x611/junc0 x611/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8479 x591/RWL0_junc x591/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8480 x192/RWL1_junc RWL_0 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8481 x841/junc1 WWL_22 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8482 RBL0_22 RWL_9 x937/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8483 GND x352/junc1 x352/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8484 WBL_23 WWL_19 x418/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8485 x410/junc0 x410/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8486 x946/junc1 WWL_18 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8487 x75/junc0 x75/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8488 x412/junc0 x412/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8489 x446/junc1 WWL_29 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8490 RBL0_11 RWL_19 x339/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8491 GND x415/junc0 x415/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8492 x163/junc0 x163/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8493 x34/junc0 x34/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8494 VDD x991/junc0 x991/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8495 x947/junc1 WWL_20 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8496 x685/junc0 x685/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8497 GND x279/junc1 x279/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8498 x204/RWL1_junc RWL_22 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8499 GND x891/junc0 x891/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8500 GND x244/junc0 x244/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8501 GND x782/junc1 x782/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8502 x792/RWL0_junc x792/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8503 x847/junc1 WWL_26 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8504 VDD x804/junc0 x804/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8505 x182/RWL0_junc x182/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8506 x180/RWL0_junc x180/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8507 x98/junc0 x98/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8508 x927/RWL1_junc RWL_5 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8509 x848/junc1 WWL_3 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8510 RBL0_13 RWL_6 x112/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8511 WBL_14 WWL_16 x442/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8512 x614/RWL0_junc x614/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8513 WBL_5 WWL_24 x534/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8514 x507/junc0 x507/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8515 x805/junc0 x805/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8516 GND x958/junc0 x958/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8517 GND x349/junc0 x349/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8518 x639/junc0 x639/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8519 GND x388/junc1 x388/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8520 GND x791/junc1 x791/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8521 GND x465/junc1 x465/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8522 GND x892/junc1 x892/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8523 x955/RWL0_junc x955/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8524 GND x959/junc0 x959/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8525 GND x428/junc0 x428/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8526 x893/RWL0_junc x893/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8527 x201/RWL0_junc x201/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8528 GND x497/junc0 x497/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8529 x833/junc0 x833/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8530 x235/RWL1_junc RWL_1 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8531 RBL0_31 RWL_2 x377/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8532 VDD x49/junc0 x49/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8533 x853/junc1 WWL_23 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8534 VDD x995/junc0 x995/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8535 WBL_23 WWL_20 x812/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8536 x448/junc0 x448/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8537 x249/RWL1_junc RWL_27 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8538 GND x454/junc0 x454/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8539 x90/junc0 x90/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8540 RBL0_0 RWL_21 x391/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8541 VDD x133/junc0 x133/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8542 x705/junc0 x705/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8543 GND x798/junc1 x798/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8544 x252/RWL1_junc RWL_23 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8545 GND x902/junc0 x902/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8546 GND x321/junc1 x321/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8547 x382/RWL1_junc RWL_30 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8548 GND x800/junc1 x800/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8549 x298/RWL0_junc x298/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8550 x679/RWL0_junc x679/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8551 x855/junc1 WWL_19 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8552 x65/junc1 WWL_27 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8553 RBL0_25 RWL_20 x403/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8554 VDD x824/junc0 x824/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8555 x681/RWL0_junc x681/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8556 x818/junc0 x818/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8557 GND x966/junc0 x966/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8558 x73/junc1 WWL_0 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8559 x954/junc1 WWL_4 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8560 RBL0_11 RWL_30 x174/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8561 GND x925/junc1 x925/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8562 x637/RWL0_junc x637/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8563 x466/junc0 x466/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8564 x839/junc0 x839/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8565 x229/junc0 x229/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8566 VDD x544/junc0 x544/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8567 RBL0_3 RWL_17 x1/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8568 x1005/RWL1_junc RWL_4 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8569 x118/junc0 x118/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8570 GND x430/junc1 x430/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8571 RBL0_7 RWL_13 x5/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8572 x641/RWL0_junc x641/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8573 GND x431/junc1 x431/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8574 x964/RWL0_junc x964/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8575 RBL0_27 RWL_7 x10/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8576 GND x531/junc0 x531/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8577 RBL0_31 x389/RWL1 x14/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8578 VDD x106/junc0 x106/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8579 x741/RWL1_junc RWL_28 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8580 x957/junc1 WWL_24 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8581 VDD x843/junc0 x843/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8582 WBL_3 WWL_2 x75/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8583 VDD x176/junc0 x176/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8584 x479/junc0 x479/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8585 RBL0_25 RWL_9 x26/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8586 x140/junc0 x140/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8587 x1010/junc0 x1010/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8588 RBL0_0 RWL_22 x27/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8589 x187/junc0 x187/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8590 WBL_10 WWL_10 x685/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8591 RBL0_21 RWL_28 x0/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8592 GND x362/junc1 x362/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8593 GND x365/junc1 x365/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8594 VDD x569/junc0 x569/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8595 x515/junc1 WWL_29 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8596 x489/junc0 x489/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8597 x340/RWL0_junc x340/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8598 x962/junc1 WWL_20 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8599 GND x485/junc0 x485/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8600 x702/RWL0_junc x702/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8601 x849/junc0 x849/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8602 x827/junc0 x827/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8603 GND x8/junc0 x8/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8604 RBL0_13 RWL_31 x776/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8605 x127/junc1 WWL_1 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8606 x577/junc0 x577/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8607 x496/junc0 x496/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8608 x969/RWL0_junc x969/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8609 GND x432/junc0 x432/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8610 WBL_28 WWL_6 x507/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8611 x851/junc0 x851/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8612 RBL0_12 RWL_10 x49/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8613 x704/junc0 x704/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8614 x965/junc1 WWL_17 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8615 WBL_19 WWL_14 x805/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8616 GND x376/junc1 x376/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8617 RBL0_3 RWL_18 x51/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8618 x472/RWL1_junc RWL_5 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8619 RBL0_16 RWL_6 x57/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8620 x665/RWL0_junc x665/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8621 x712/RWL0_junc x712/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8622 GND x438/junc0 x438/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8623 RBL0_27 RWL_8 x64/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8624 VDD x583/junc0 x583/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8625 GND x33/junc0 x33/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8626 GND x568/junc0 x568/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8627 x874/RWL1_junc RWL_13 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8628 x385/RWL1_junc RWL_30 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8629 WBL_1 WWL_21 x833/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8630 x515/RWL1_junc RWL_29 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8631 VDD x43/junc0 x43/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8632 x308/junc0 x308/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8633 VDD x592/junc0 x592/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8634 RBL0_21 RWL_14 x80/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8635 x223/junc0 x223/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8636 x221/junc0 x221/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8637 x511/junc0 x511/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8638 RBL0_0 RWL_23 x81/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8639 RBL0_17 RWL_30 x231/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8640 WBL_10 WWL_11 x705/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8641 GND x408/junc1 x408/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8642 RBL0_21 RWL_29 x54/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8643 WBL_14 WWL_30 x188/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8644 x333/RWL1_junc RWL_17 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8645 x1014/RWL1_junc RWL_21 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8646 x17/RWL0_junc x17/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8647 x378/RWL0_junc x378/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8648 VDD x601/junc0 x601/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8649 VDD x95/junc0 x95/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8650 x520/junc0 x520/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8651 x383/RWL0_junc x383/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8652 GND x458/junc0 x458/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8653 x859/junc0 x859/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8654 GND x145/junc0 x145/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8655 x753/junc1 WWL_2 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8656 VDD x212/junc0 x212/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8657 WBL_4 WWL_17 x818/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8658 GND x62/junc0 x62/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8659 GND x413/junc1 x413/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8660 x455/junc0 x455/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8661 x248/junc0 x248/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8662 x528/junc0 x528/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8663 x730/RWL0_junc x730/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8664 GND x976/junc0 x976/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8665 x179/junc1 WWL_10 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8666 WBL_28 WWL_7 x839/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8667 RBL0_12 RWL_11 x106/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8668 x970/junc1 WWL_18 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8669 GND x420/junc1 x420/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8670 RBL0_3 RWL_19 x110/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8671 x918/RWL0_junc x918/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8672 x615/junc0 x615/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8673 GND x922/junc0 x922/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8674 GND x917/junc1 x917/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8675 GND x767/junc0 x767/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8676 GND x469/junc0 x469/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8677 GND x923/junc0 x923/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8678 x359/RWL1_junc RWL_14 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8679 x539/junc0 x539/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8680 RBL0_6 RWL_17 x120/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8681 GND x829/junc1 x829/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8682 VDD x260/junc0 x260/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8683 GND x381/junc1 x381/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8684 x543/junc0 x543/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8685 WBL_24 WWL_28 x816/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8686 GND x443/junc1 x443/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8687 x547/junc0 x547/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8688 RBL0_30 RWL_7 x130/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8689 x694/RWL0_junc x694/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8690 VDD x100/junc0 x100/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8691 x198/junc1 WWL_14 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8692 x471/junc0 x471/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8693 x350/junc0 x350/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8694 VDD x624/junc0 x624/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8695 RBL0_21 RWL_15 x131/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8696 WBL_6 WWL_2 x187/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8697 WBL_14 WWL_31 x998/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8698 x107/junc1 WWL_25 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8699 x374/RWL1_junc RWL_18 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8700 x707/RWL1_junc RWL_22 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8701 x423/RWL0_junc x423/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8702 x628/junc0 x628/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8703 x557/junc0 x557/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8704 GND x488/junc0 x488/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8705 WBL_13 WWL_10 x849/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8706 GND x945/junc1 x945/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8707 GND x452/junc1 x452/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8708 WBL_4 WWL_18 x827/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8709 x874/RWL0_junc x874/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8710 x435/RWL0_junc x435/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8711 x593/junc1 WWL_28 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8712 GND x786/junc0 x786/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8713 WBL_24 WWL_12 x577/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8714 x746/RWL0_junc x746/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8715 x844/RWL0_junc x844/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8716 GND x126/junc0 x126/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8717 x220/junc1 WWL_11 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8718 WBL_28 WWL_8 x851/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8719 RBL0_12 RWL_12 x159/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8720 VDD x422/junc0 x422/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8721 x637/junc0 x637/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8722 WBL_11 WWL_29 x999/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8723 x877/junc0 x877/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8724 GND x928/junc1 x928/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8725 GND x132/junc0 x132/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8726 x405/RWL1_junc RWL_15 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8727 x495/junc0 x495/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8728 GND x978/junc0 x978/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8729 x232/junc1 WWL_17 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8730 x264/junc0 x264/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8731 x576/junc0 x576/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8732 RBL0_6 RWL_18 x167/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8733 WBL_20 WWL_30 x562/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8734 GND x933/junc0 x933/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8735 VDD x143/junc0 x143/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8736 x900/junc1 WWL_19 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8737 GND x734/junc1 x734/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8738 x411/RWL1_junc RWL_21 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8739 RBL0_17 RWL_20 x95/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8740 x579/junc0 x579/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8741 x503/junc0 x503/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8742 RBL0_30 RWL_8 x175/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8743 x653/RWL0_junc x653/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8744 VDD x784/junc0 x784/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8745 RBL0_21 RWL_16 x177/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8746 WBL_15 WWL_9 x223/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8747 WBL_0 WWL_2 x221/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8748 x158/junc1 WWL_26 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8749 x729/RWL1_junc RWL_23 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8750 x418/RWL1_junc RWL_19 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8751 x954/RWL1_junc RWL_4 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8752 WBL_9 WWL_15 x603/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8753 x850/RWL0_junc x850/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8754 VDD x651/junc0 x651/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8755 GND x951/junc1 x951/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8756 WBL_13 WWL_11 x859/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8757 x756/RWL0_junc x756/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8758 x980/RWL0_junc x980/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8759 GND x482/junc1 x482/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8760 GND x935/junc1 x935/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8761 WBL_24 WWL_13 x248/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8762 x467/RWL0_junc x467/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8763 GND x173/junc0 x173/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8764 VDD x459/junc0 x459/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8765 x194/junc0 x194/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8766 x440/RWL1_junc RWL_0 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8767 x632/RWL0_junc x632/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8768 GND x676/junc1 x676/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8769 x905/junc1 WWL_22 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8770 x336/junc0 x336/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8771 RBL0_17 RWL_9 x134/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8772 GND x561/junc1 x561/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8773 WBL_18 WWL_19 x615/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8774 GND x181/junc0 x181/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8775 x1019/junc1 WWL_10 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8776 x442/RWL1_junc RWL_16 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8777 x609/junc0 x609/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8778 x285/junc1 WWL_18 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8779 x610/junc0 x610/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8780 RBL0_6 RWL_19 x213/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8781 WBL_20 WWL_31 x842/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8782 GND x538/junc0 x538/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8783 x998/RWL0_junc x998/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8784 GND x612/junc0 x612/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8785 VDD x667/junc0 x667/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8786 x907/junc1 WWL_12 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8787 x415/junc0 x415/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8788 x534/junc0 x534/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8789 GND x1021/junc1 x1021/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8790 VDD x196/junc0 x196/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8791 GND x500/junc1 x500/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8792 x290/junc1 WWL_20 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8793 x865/junc0 x865/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8794 x450/RWL1_junc RWL_22 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8795 GND x940/junc0 x940/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8796 GND x19/junc1 x19/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8797 x962/RWL1_junc RWL_20 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8798 x319/junc0 x319/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8799 x799/junc0 x799/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8800 x434/RWL0_junc x434/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8801 WBL_20 WWL_6 x1010/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8802 x774/junc1 WWL_27 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8803 x963/RWL1_junc RWL_5 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8804 RBL0_8 RWL_6 x233/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8805 WBL_9 WWL_16 x628/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8806 x861/RWL0_junc x861/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8807 VDD x210/junc0 x210/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8808 x675/junc0 x675/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8809 WBL_17 WWL_29 x544/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8810 GND x513/junc1 x513/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8811 GND x590/junc1 x590/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8812 VDD x346/junc0 x346/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8813 GND x216/junc0 x216/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8814 GND x673/junc0 x673/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8815 x447/RWL0_junc x447/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8816 VDD x684/junc0 x684/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8817 x504/RWL0_junc x504/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8818 x912/junc1 WWL_15 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8819 x470/RWL1_junc RWL_1 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8820 RBL0_26 RWL_2 x255/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8821 VDD x325/junc0 x325/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8822 x913/junc1 WWL_23 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8823 VDD x225/junc0 x225/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8824 WBL_18 WWL_20 x877/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8825 x1020/junc1 WWL_11 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8826 x631/junc0 x631/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8827 x688/junc0 x688/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8828 x687/junc0 x687/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8829 GND x574/junc0 x574/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8830 x266/RWL1_junc RWL_9 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8831 GND x635/junc0 x635/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8832 x474/RWL1_junc RWL_27 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8833 GND x244/junc1 x244/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8834 x570/junc0 x570/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8835 x473/RWL1_junc RWL_13 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8836 VDD x236/junc0 x236/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8837 x572/junc0 x572/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8838 GND x1022/junc1 x1022/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8839 x819/junc1 WWL_13 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8840 x690/junc0 x690/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8841 x876/junc0 x876/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8842 GND x863/junc1 x863/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8843 x476/RWL1_junc RWL_23 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8844 GND x23/junc0 x23/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8845 GND x867/junc1 x867/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8846 x363/junc0 x363/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8847 x518/RWL0_junc x518/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8848 x247/junc1 WWL_19 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8849 x811/junc0 x811/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8850 WBL_20 WWL_7 x588/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8851 x984/RWL0_junc x984/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8852 x697/junc0 x697/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8853 x797/RWL0_junc x797/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8854 x648/junc0 x648/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8855 x903/junc0 x903/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8856 x104/RWL1_junc RWL_4 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8857 GND x428/junc1 x428/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8858 x757/RWL0_junc x757/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8859 GND x621/junc1 x621/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8860 GND x868/junc1 x868/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8861 RBL0_2 RWL_13 x292/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8862 VDD x394/junc0 x394/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8863 x920/junc1 WWL_6 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8864 RBL0_22 RWL_7 x294/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8865 GND x778/junc1 x778/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8866 GND x599/junc0 x599/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8867 GND x692/junc0 x692/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8868 VDD x523/junc0 x523/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8869 x921/junc1 WWL_16 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8870 RBL0_26 x389/RWL1 x296/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8871 VDD x366/junc0 x366/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8872 x58/RWL1_junc RWL_28 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8873 x982/junc1 WWL_24 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8874 VDD x275/junc0 x275/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8875 x887/junc0 x887/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8876 x708/junc0 x708/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8877 WBL_30 WWL_25 x662/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8878 VDD x427/junc0 x427/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8879 x507/RWL1_junc RWL_6 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8880 x508/RWL1_junc RWL_20 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8881 GND x949/junc0 x949/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8882 x602/junc0 x602/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8883 GND x73/junc0 x73/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8884 VDD x286/junc0 x286/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8885 x605/junc0 x605/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8886 x888/junc0 x888/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8887 GND x897/junc1 x897/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8888 WBL_5 WWL_10 x865/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8889 GND x573/junc1 x573/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8890 VDD x713/junc0 x713/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8891 x989/RWL0_junc x989/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8892 x683/junc1 WWL_29 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8893 x988/RWL0_junc x988/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8894 x639/junc0 x639/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8895 x554/RWL0_junc x554/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8896 x1018/junc1 WWL_20 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8897 x407/junc0 x407/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8898 WBL_29 WWL_0 x799/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8899 x793/junc0 x793/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8900 RBL0_13 RWL_4 x668/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8901 WBL_20 WWL_8 x617/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8902 GND x293/junc0 x293/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8903 x831/RWL0_junc x831/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8904 x719/junc0 x719/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8905 x672/junc0 x672/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8906 GND x622/junc0 x622/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8907 WBL_23 WWL_6 x675/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8908 x911/junc0 x911/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8909 GND x640/junc1 x640/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8910 RBL0_7 RWL_10 x325/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8911 GND x950/junc1 x950/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8912 GND x582/junc1 x582/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8913 x153/RWL1_junc RWL_5 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8914 RBL0_11 RWL_6 x329/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8915 x777/RWL0_junc x777/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8916 x809/junc0 x809/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8917 x722/junc0 x722/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8918 x724/junc0 x724/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8919 RBL0_31 RWL_0 x330/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8920 x985/junc1 WWL_7 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8921 VDD x725/junc0 x725/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8922 RBL0_22 RWL_8 x332/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8923 GND x591/junc1 x591/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8924 GND x994/junc0 x994/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8925 x536/RWL1_junc RWL_9 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8926 GND x709/junc0 x709/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8927 GND x715/junc0 x715/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8928 VDD x560/junc0 x560/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8929 x683/RWL1_junc RWL_29 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8930 x821/junc0 x821/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8931 WBL_31 WWL_22 x687/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8932 WBL_30 WWL_26 x688/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8933 x464/junc0 x464/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8934 x593/RWL1_junc RWL_28 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8935 x627/junc0 x627/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8936 GND x127/junc0 x127/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8937 WBL_14 WWL_3 x690/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8938 x514/junc0 x514/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8939 x733/junc0 x733/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8940 WBL_5 WWL_11 x876/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8941 GND x606/junc1 x606/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8942 x548/RWL1_junc RWL_17 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8943 x892/RWL0_junc x892/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8944 VDD x736/junc0 x736/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8945 x992/RWL0_junc x992/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8946 x993/RWL0_junc x993/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8947 RBL0_27 RWL_28 x265/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8948 x899/junc0 x899/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8949 x587/RWL0_junc x587/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8950 GND x638/junc0 x638/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8951 WBL_29 WWL_1 x811/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8952 GND x182/junc1 x182/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8953 x806/junc0 x806/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8954 x838/junc1 WWL_2 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8955 GND x180/junc1 x180/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8956 RBL0_13 RWL_5 x545/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8957 VDD x739/junc0 x739/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8958 GND x331/junc0 x331/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8959 GND x953/junc1 x953/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8960 x636/junc0 x636/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8961 x535/RWL0_junc x535/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8962 x473/junc0 x473/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8963 GND x864/junc0 x864/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8964 x691/junc0 x691/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8965 GND x996/junc0 x996/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8966 WBL_23 WWL_7 x903/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8967 x429/junc1 WWL_10 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8968 x453/junc0 x453/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8969 RBL0_7 RWL_11 x366/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8970 GND x616/junc1 x616/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8971 x155/RWL0_junc x155/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8972 x1019/RWL1_junc RWL_10 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8973 GND x960/junc0 x960/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8974 x981/junc0 x981/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8975 GND x955/junc1 x955/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8976 GND x845/junc0 x845/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8977 x822/junc0 x822/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8978 x922/junc0 x922/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8979 WBL_16 WWL_25 x85/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8980 x923/junc0 x923/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8981 x571/RWL1_junc RWL_14 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8982 RBL0_31 RWL_1 x373/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8983 x990/junc1 WWL_8 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8984 VDD x483/junc0 x483/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8985 GND x893/junc1 x893/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8986 x608/RWL0_junc x608/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8987 GND x201/junc1 x201/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8988 VDD x486/junc0 x486/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M8989 GND x586/junc1 x586/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8990 GND x997/junc0 x997/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8991 WBL_3 WWL_28 x53/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8992 GND x768/junc1 x768/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8993 x356/junc1 WWL_6 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8994 WBL_31 WWL_23 x708/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8995 x701/junc0 x701/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8996 RBL0_25 RWL_7 x384/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8997 x925/RWL0_junc x925/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8998 RBL0_15 RWL_27 x381/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M8999 WBL_30 WWL_27 x887/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9000 VDD x90/junc0 x90/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9001 x445/junc1 WWL_14 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9002 x371/junc0 x371/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9003 RBL0_0 RWL_20 x386/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9004 x71/RWL1_junc RWL_29 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9005 WBL_14 WWL_4 x888/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9006 x774/RWL1_junc RWL_27 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9007 x581/RWL1_junc RWL_18 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9008 x748/junc0 x748/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9009 GND x370/junc0 x370/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9010 RBL0_27 RWL_29 x302/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9011 x908/junc0 x908/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9012 GND x661/junc0 x661/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9013 GND x681/junc1 x681/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9014 WBL_26 WWL_30 x164/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9015 GND x961/junc1 x961/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9016 VDD x466/junc0 x466/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9017 x711/junc0 x711/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9018 WBL_19 WWL_12 x719/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9019 GND x663/junc0 x663/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9020 x860/junc1 WWL_15 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9021 GND x875/junc0 x875/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9022 RBL0_16 RWL_4 x410/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9023 x462/junc1 WWL_11 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9024 x480/junc0 x480/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9025 WBL_23 WWL_8 x911/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9026 RBL0_7 RWL_12 x412/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9027 GND x968/junc0 x968/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9028 GND x641/junc1 x641/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9029 GND x390/junc0 x390/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9030 x1020/RWL1_junc RWL_11 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9031 GND x964/junc1 x964/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9032 WBL_16 WWL_26 x722/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9033 x603/RWL1_junc RWL_15 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9034 RBL0_0 RWL_9 x417/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9035 WBL_1 WWL_19 x724/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9036 x1/junc1 WWL_17 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9037 x490/junc0 x490/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9038 x630/RWL0_junc x630/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9039 VDD x270/junc0 x270/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9040 x634/RWL0_junc x634/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9041 x10/junc1 WWL_7 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9042 x792/RWL1_junc RWL_21 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9043 x721/junc0 x721/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9044 WBL_31 WWL_24 x821/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9045 x1017/junc0 x1017/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9046 RBL0_25 RWL_8 x426/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9047 GND x537/junc1 x537/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9048 WBL_10 WWL_9 x464/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9049 x509/junc1 WWL_28 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9050 RBL0_20 RWL_24 x734/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9051 x317/junc0 x317/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9052 x615/RWL1_junc RWL_19 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9053 x536/junc0 x536/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9054 WBL_4 WWL_15 x162/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9055 GND x414/junc0 x414/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9056 x1019/RWL0_junc x1019/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9057 VDD x765/junc0 x765/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9058 WBL_26 WWL_31 x211/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9059 x228/RWL0_junc x228/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9060 x441/junc1 WWL_29 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9061 x1001/RWL0_junc x1001/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9062 x83/junc0 x83/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9063 WBL_28 WWL_5 x169/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9064 GND x659/junc1 x659/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9065 x872/junc1 WWL_16 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9066 GND x760/junc0 x760/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9067 GND x969/junc1 x969/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9068 WBL_19 WWL_13 x473/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9069 RBL0_16 RWL_5 x448/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9070 x553/junc0 x553/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9071 GND x972/junc0 x972/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9072 x517/junc0 x517/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9073 x752/RWL0_junc x752/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9074 WBL_27 WWL_17 x836/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9075 GND x665/junc1 x665/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9076 GND x712/junc1 x712/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9077 GND x433/junc0 x433/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9078 x862/RWL1_junc RWL_12 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9079 WBL_16 WWL_27 x922/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9080 x628/RWL1_junc RWL_16 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9081 x742/junc0 x742/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9082 WBL_1 WWL_20 x923/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9083 x51/junc1 WWL_18 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9084 x652/RWL0_junc x652/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9085 GND x696/junc0 x696/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9086 GND x788/junc0 x788/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9087 VDD x780/junc0 x780/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9088 x413/RWL0_junc x413/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9089 x948/junc1 WWL_12 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9090 x612/junc0 x612/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9091 VDD x781/junc0 x781/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9092 VDD x308/junc0 x308/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9093 x656/RWL0_junc x656/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9094 x64/junc1 WWL_8 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9095 x679/RWL1_junc RWL_22 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9096 x755/junc1 WWL_30 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9097 RBL0_28 RWL_21 x466/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9098 x1018/RWL1_junc RWL_20 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9099 RBL0_29 RWL_17 x1021/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9100 x699/junc0 x699/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9101 RBL0_20 RWL_25 x500/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9102 x121/junc0 x121/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9103 x924/RWL0_junc x924/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9104 x623/RWL0_junc x623/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9105 VDD x520/junc0 x520/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9106 RBL0_3 RWL_6 x118/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9107 x401/RWL1_junc RWL_24 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9108 WBL_4 WWL_16 x748/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9109 x1020/RWL0_junc x1020/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9110 VDD x455/junc0 x455/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9111 x791/junc0 x791/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9112 GND x975/junc0 x975/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9113 GND x974/junc0 x974/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9114 VDD x457/junc0 x457/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9115 x873/junc1 WWL_9 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9116 x243/junc0 x243/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9117 GND x682/junc1 x682/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9118 GND x657/junc1 x657/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9119 GND x730/junc1 x730/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9120 GND x749/junc0 x749/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9121 GND x784/junc0 x784/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9122 x710/junc0 x710/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9123 x552/junc0 x552/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9124 x764/RWL0_junc x764/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9125 WBL_27 WWL_18 x846/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9126 x952/junc1 WWL_15 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9127 RBL0_21 RWL_2 x479/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9128 VDD x539/junc0 x539/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9129 GND x918/junc1 x918/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9130 VDD x565/junc0 x565/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9131 VDD x59/junc0 x59/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9132 x751/junc0 x751/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9133 x766/junc1 WWL_28 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9134 x40/junc0 x40/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9135 x798/junc0 x798/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9136 GND x718/junc0 x718/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9137 x937/RWL1_junc RWL_9 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9138 GND x803/junc0 x803/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9139 VDD x471/junc0 x471/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9140 x452/RWL0_junc x452/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9141 x716/junc0 x716/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9142 x881/junc1 WWL_13 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9143 VDD x350/junc0 x350/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9144 x800/junc0 x800/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9145 x263/junc0 x263/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9146 x702/RWL1_junc RWL_23 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9147 x399/junc0 x399/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9148 VDD x801/junc0 x801/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9149 x858/junc1 WWL_17 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9150 x776/junc1 WWL_31 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9151 x546/junc1 WWL_21 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9152 RBL0_28 RWL_22 x496/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9153 RBL0_29 RWL_18 x1022/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9154 x720/junc0 x720/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9155 x686/RWL0_junc x686/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9156 RBL0_20 RWL_26 x863/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9157 x168/junc0 x168/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9158 WBL_13 WWL_9 x536/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9159 x662/RWL1_junc RWL_25 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9160 x1003/RWL0_junc x1003/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9161 x862/RWL0_junc x862/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9162 x762/junc0 x762/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9163 WBL_8 WWL_25 x899/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9164 x178/junc0 x178/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9165 x613/junc0 x613/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9166 x669/RWL1_junc RWL_2 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9167 GND x977/junc0 x977/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9168 GND x763/junc0 x763/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9169 VDD x38/junc0 x38/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9170 WBL_12 WWL_21 x83/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9171 GND x680/junc1 x680/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9172 x840/RWL0_junc x840/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9173 GND x746/junc1 x746/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9174 GND x926/junc1 x926/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9175 VDD x142/junc0 x142/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9176 x958/junc1 WWL_6 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9177 RBL0_17 RWL_7 x308/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9178 GND x802/junc0 x802/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9179 x731/junc0 x731/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9180 x585/junc0 x585/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9181 x959/junc1 WWL_16 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9182 RBL0_21 x61/RWL1 x511/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9183 VDD x576/junc0 x576/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9184 VDD x704/junc0 x704/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9185 x790/junc1 WWL_30 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9186 x15/RWL1_junc RWL_10 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9187 x649/RWL1_junc RWL_30 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9188 x197/junc0 x197/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9189 WBL_25 WWL_25 x279/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9190 x93/junc0 x93/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9191 VDD x619/junc0 x619/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9192 GND x979/junc0 x979/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9193 x675/RWL1_junc RWL_6 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9194 GND x823/junc0 x823/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9195 x17/RWL1_junc RWL_20 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9196 RBL0_14 RWL_21 x747/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9197 x737/junc0 x737/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9198 GND x337/junc0 x337/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9199 VDD x503/junc0 x503/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9200 RBL0_25 RWL_31 x676/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9201 x205/junc0 x205/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9202 x542/junc0 x542/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9203 GND x717/junc1 x717/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9204 x1004/RWL0_junc x1004/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9205 x870/junc1 WWL_18 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9206 RBL0_29 RWL_19 x897/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9207 x743/junc0 x743/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9208 x706/RWL0_junc x706/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9209 WBL_30 WWL_29 x739/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9210 RBL0_28 RWL_23 x528/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9211 WBL_24 WWL_0 x121/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9212 RBL0_8 RWL_4 x207/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9213 GND x75/junc0 x75/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9214 x688/RWL1_junc RWL_26 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9215 x895/RWL0_junc x895/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9216 x524/junc0 x524/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9217 x2/junc0 x2/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9218 x218/junc0 x218/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9219 WBL_18 WWL_6 x791/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9220 GND x756/junc1 x756/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9221 x222/junc0 x222/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9222 WBL_8 WWL_26 x908/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9223 x690/RWL1_junc x61/RWL1 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9224 RBL0_2 RWL_10 x539/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9225 GND x980/junc1 x980/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9226 x1021/RWL0_junc x1021/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9227 GND x787/junc0 x787/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9228 RBL0_6 RWL_6 x543/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9229 GND x703/junc1 x703/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9230 x852/RWL0_junc x852/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9231 VDD x194/junc0 x194/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9232 x137/junc0 x137/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9233 x1013/junc0 x1013/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9234 x391/RWL1_junc RWL_21 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9235 RBL0_26 RWL_0 x547/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9236 x596/junc1 WWL_7 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9237 VDD x825/junc0 x825/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9238 RBL0_17 RWL_8 x350/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9239 x694/RWL1_junc RWL_9 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9240 x134/junc1 WWL_9 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9241 GND x649/junc1 x649/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9242 GND x817/junc0 x817/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9243 VDD x1015/junc0 x1015/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9244 x324/junc1 WWL_31 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9245 x10/RWL1_junc RWL_7 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9246 x531/junc1 WWL_25 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9247 x70/RWL1_junc RWL_11 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9248 x880/junc0 x880/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9249 WBL_26 WWL_22 x40/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9250 VDD x643/junc0 x643/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9251 WBL_25 WWL_26 x798/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9252 x644/junc0 x644/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9253 x884/junc1 WWL_21 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9254 x885/junc1 WWL_14 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9255 RBL0_14 RWL_22 x761/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9256 x32/junc0 x32/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9257 GND x379/junc0 x379/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9258 WBL_9 WWL_3 x800/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9259 x253/junc0 x253/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9260 GND x738/junc1 x738/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9261 VDD x319/junc0 x319/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9262 x1007/RWL0_junc x1007/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9263 WBL_20 WWL_5 x1017/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9264 x728/RWL0_junc x728/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9265 WBL_24 WWL_1 x168/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9266 GND x434/junc1 x434/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9267 VDD x828/junc0 x828/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9268 RBL0_8 RWL_5 x256/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9269 x629/junc1 WWL_25 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9270 GND x129/junc0 x129/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9271 x52/junc0 x52/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9272 x55/junc0 x55/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9273 x269/junc0 x269/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9274 WBL_18 WWL_7 x178/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9275 x620/junc1 WWL_10 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9276 WBL_8 WWL_27 x882/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9277 RBL0_2 RWL_11 x576/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9278 x1022/RWL0_junc x1022/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9279 x509/RWL1_junc RWL_28 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9280 x154/junc0 x154/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9281 x409/RWL0_junc x409/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9282 x768/junc0 x768/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9283 GND x983/junc0 x983/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9284 x113/RWL1_junc RWL_14 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9285 GND x910/junc0 x910/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9286 x625/junc1 WWL_0 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9287 x883/junc0 x883/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9288 x1006/RWL0_junc x1006/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9289 x960/junc0 x960/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9290 WBL_11 WWL_25 x82/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9291 x27/RWL1_junc RWL_22 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9292 RBL0_26 RWL_1 x579/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9293 x626/junc1 WWL_8 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9294 VDD x76/junc0 x76/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9295 RBL0_29 RWL_30 x936/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9296 x740/RWL0_junc x740/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9297 GND x447/junc1 x447/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9298 VDD x660/junc0 x660/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9299 RBL0_21 RWL_31 x428/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9300 x647/junc0 x647/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9301 x124/RWL1_junc RWL_4 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9302 x64/RWL1_junc RWL_8 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9303 GND x188/junc0 x188/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9304 x33/junc1 WWL_6 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9305 x719/RWL1_junc RWL_12 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9306 x568/junc1 WWL_26 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9307 WBL_26 WWL_23 x93/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9308 VDD x570/junc0 x570/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9309 RBL0_10 RWL_27 x586/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9310 WBL_25 WWL_27 x197/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9311 VDD x572/junc0 x572/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9312 x669/junc0 x669/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9313 GND x13/junc1 x13/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9314 RBL0_14 RWL_23 x783/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9315 WBL_9 WWL_4 x205/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9316 VDD x363/junc0 x363/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9317 GND x578/junc0 x578/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9318 GND x30/junc1 x30/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9319 x341/RWL0_junc x341/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9320 x871/RWL0_junc x871/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9321 x747/RWL0_junc x747/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9322 x651/junc1 WWL_26 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9323 VDD x648/junc0 x648/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9324 x812/junc0 x812/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9325 GND x984/junc1 x984/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9326 x108/junc0 x108/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9327 x62/junc1 WWL_3 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9328 RBL0_11 RWL_4 x609/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9329 x645/junc1 WWL_11 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9330 WBL_18 WWL_8 x222/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9331 RBL0_2 RWL_12 x610/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9332 x821/junc0 x821/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9333 x897/RWL0_junc x897/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9334 GND x986/junc0 x986/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9335 x968/junc0 x968/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9336 GND x816/junc0 x816/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9337 x313/junc0 x313/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9338 x544/RWL1_junc RWL_29 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9339 x6/junc0 x6/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9340 x976/junc1 WWL_5 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9341 GND x987/junc0 x987/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9342 GND x757/junc1 x757/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9343 GND x190/junc0 x190/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9344 x161/RWL1_junc RWL_7 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9345 x650/junc1 WWL_1 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9346 WBL_11 WWL_26 x137/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9347 x81/RWL1_junc RWL_23 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9348 x162/RWL1_junc RWL_15 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9349 x519/junc0 x519/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9350 GND x956/junc1 x956/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9351 x750/RWL0_junc x750/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9352 GND x998/junc0 x998/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9353 VDD x97/junc0 x97/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9354 x753/RWL0_junc x753/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9355 x169/RWL1_junc RWL_5 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9356 x670/junc0 x670/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9357 x294/junc1 WWL_7 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9358 x1008/junc1 WWL_27 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9359 VDD x602/junc0 x602/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9360 WBL_26 WWL_24 x880/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9361 GND x67/junc1 x67/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9362 x227/junc0 x227/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9363 x858/RWL1_junc RWL_17 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9364 WBL_5 WWL_9 x644/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9365 GND x697/junc1 x697/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9366 x533/junc0 x533/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9367 GND x989/junc1 x989/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9368 x694/junc0 x694/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9369 GND x988/junc1 x988/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9370 GND x611/junc0 x611/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9371 VDD x123/junc0 x123/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9372 x392/RWL0_junc x392/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9373 x886/RWL0_junc x886/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9374 x761/RWL0_junc x761/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9375 x210/junc1 WWL_27 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9376 x258/junc0 x258/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9377 x343/junc0 x343/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9378 WBL_23 WWL_5 x420/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9379 GND x831/junc1 x831/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9380 GND x223/junc0 x223/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9381 GND x775/junc1 x775/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9382 GND x5/junc0 x5/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9383 x668/junc1 WWL_4 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9384 RBL0_11 RWL_5 x631/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9385 x163/junc0 x163/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9386 x972/junc0 x972/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9387 GND x991/junc0 x991/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9388 x685/junc0 x685/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9389 GND x234/junc0 x234/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9390 RBL0_17 RWL_31 x663/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9391 x357/junc0 x357/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9392 WBL_22 WWL_17 x154/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9393 GND x777/junc1 x777/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9394 GND x105/junc1 x105/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9395 x206/RWL1_junc RWL_8 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9396 x170/junc0 x170/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9397 WBL_11 WWL_27 x960/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9398 x748/RWL1_junc RWL_16 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9399 x769/RWL0_junc x769/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9400 GND x804/junc0 x804/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9401 x953/RWL0_junc x953/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9402 VDD x147/junc0 x147/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9403 x978/junc1 WWL_12 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9404 VDD x151/junc0 x151/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9405 WBL_0 WWL_29 x801/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9406 x771/RWL0_junc x771/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9407 x332/junc1 WWL_8 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9408 x973/junc0 x973/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9409 WBL_14 WWL_2 x669/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9410 x278/junc0 x278/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9411 x870/RWL1_junc RWL_18 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9412 RBL0_24 RWL_17 x814/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9413 RBL0_23 RWL_21 x648/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9414 x805/junc0 x805/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9415 x375/junc0 x375/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9416 x199/RWL0_junc x199/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9417 VDD x899/junc0 x899/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9418 GND x993/junc1 x993/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9419 GND x992/junc1 x992/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9420 x597/RWL1_junc RWL_24 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9421 VDD x166/junc0 x166/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9422 VDD x636/junc0 x636/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9423 x499/RWL0_junc x499/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9424 x99/junc0 x99/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9425 x783/RWL0_junc x783/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9426 x833/junc0 x833/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9427 x437/RWL0_junc x437/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9428 GND x49/junc0 x49/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9429 GND x995/junc0 x995/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9430 x974/junc0 x974/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9431 x975/junc0 x975/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9432 VDD x271/junc0 x271/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9433 x930/junc1 WWL_9 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9434 GND x535/junc1 x535/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9435 GND x796/junc1 x796/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9436 GND x772/junc1 x772/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9437 x208/junc0 x208/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9438 GND x835/junc0 x835/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9439 WBL_18 WWL_30 x704/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9440 WBL_31 WWL_10 x968/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9441 GND x1006/junc0 x1006/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9442 RBL0_15 RWL_14 x657/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9443 WBL_30 WWL_14 x313/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9444 RBL0_0 RWL_7 x658/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9445 x705/junc0 x705/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9446 WBL_22 WWL_18 x6/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9447 x173/junc1 WWL_15 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9448 GND x155/junc1 x155/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9449 GND x733/junc1 x733/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9450 x844/junc1 WWL_28 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9451 x314/junc0 x314/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9452 x863/junc0 x863/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9453 x884/RWL1_junc RWL_21 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9454 GND x824/junc0 x824/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9455 x885/RWL1_junc RWL_14 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9456 x794/RWL0_junc x794/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9457 x181/junc1 WWL_5 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9458 x842/junc0 x842/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9459 VDD x371/junc0 x371/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9460 x961/RWL0_junc x961/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9461 VDD x34/junc0 x34/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9462 x818/junc0 x818/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9463 x934/junc1 WWL_13 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9464 x867/junc0 x867/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9465 x487/junc0 x487/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9466 x594/junc0 x594/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9467 x352/RWL1_junc RWL_19 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9468 x917/junc1 WWL_17 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9469 x839/junc0 x839/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9470 VDD x204/junc0 x204/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9471 x700/junc1 WWL_21 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9472 RBL0_23 RWL_22 x672/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9473 RBL0_24 RWL_18 x826/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9474 x229/junc0 x229/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9475 x419/junc0 x419/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9476 x279/RWL1_junc RWL_25 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9477 x1009/RWL0_junc x1009/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9478 VDD x711/junc0 x711/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9479 x868/junc0 x868/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9480 x150/junc0 x150/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9481 WBL_3 WWL_25 x45/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9482 GND x106/junc0 x106/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9483 x246/junc0 x246/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9484 x782/RWL1_junc RWL_2 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9485 GND x843/junc0 x843/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9486 x763/junc0 x763/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9487 WBL_1 WWL_6 x258/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9488 x977/junc0 x977/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9489 VDD x309/junc0 x309/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9490 WBL_7 WWL_21 x343/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9491 GND x195/junc1 x195/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9492 GND x795/junc1 x795/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9493 VDD x311/junc0 x311/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9494 WBL_27 WWL_15 x52/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9495 x509/junc0 x509/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9496 WBL_18 WWL_31 x1015/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9497 WBL_31 WWL_11 x972/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9498 RBL0_15 RWL_15 x680/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9499 RBL0_0 RWL_8 x678/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9500 x726/junc0 x726/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9501 x216/junc1 WWL_16 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9502 x444/junc0 x444/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9503 x358/junc0 x358/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9504 x388/RWL1_junc RWL_22 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9505 GND x1000/junc0 x1000/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9506 x465/RWL1_junc RWL_15 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9507 x807/RWL0_junc x807/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9508 x791/RWL1_junc RWL_6 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9509 x849/junc0 x849/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9510 VDD x809/junc0 x809/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9511 RBL0_9 RWL_21 x832/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9512 x892/RWL1_junc RWL_20 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9513 x827/junc0 x827/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9514 VDD x1017/junc0 x1017/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9515 x451/junc0 x451/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9516 x149/junc0 x149/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9517 x1011/RWL0_junc x1011/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9518 x851/junc0 x851/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9519 VDD x252/junc0 x252/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9520 x928/junc1 WWL_18 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9521 WBL_9 WWL_29 x828/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9522 RBL0_24 RWL_19 x834/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9523 x282/junc0 x282/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9524 RBL0_23 RWL_23 x691/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9525 x23/junc1 WWL_3 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9526 WBL_19 WWL_0 x375/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9527 RBL0_3 RWL_4 x453/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9528 x798/RWL1_junc RWL_26 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9529 x943/RWL0_junc x943/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9530 x461/junc0 x461/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9531 GND x228/junc1 x228/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9532 GND x159/junc0 x159/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9533 WBL_3 WWL_26 x99/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9534 x291/junc0 x291/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9535 x800/RWL1_junc x61/RWL1 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9536 GND x1001/junc1 x1001/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9537 x814/RWL0_junc x814/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9538 GND x39/junc0 x39/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9539 WBL_1 WWL_7 x975/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9540 x297/RWL0_junc x297/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9541 WBL_16 WWL_14 x974/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9542 GND x808/junc1 x808/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9543 x819/RWL0_junc x819/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9544 x820/RWL0_junc x820/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9545 GND x43/junc0 x43/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9546 VDD x353/junc0 x353/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9547 x395/junc0 x395/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9548 VDD x272/junc0 x272/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9549 GND x919/junc1 x919/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9550 WBL_27 WWL_16 x108/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9551 RBL0_21 RWL_0 x701/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9552 x925/RWL1_junc RWL_9 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9553 RBL0_15 RWL_16 x703/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9554 x25/junc1 WWL_29 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9555 x294/RWL1_junc RWL_7 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9556 x1008/RWL1_junc RWL_27 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9557 x692/junc1 WWL_25 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9558 GND x95/junc0 x95/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9559 VDD x759/junc0 x759/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9560 x933/junc0 x933/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9561 WBL_21 WWL_22 x314/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9562 VDD x981/junc0 x981/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9563 x430/RWL1_junc RWL_23 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9564 x935/junc1 WWL_21 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9565 x431/RWL1_junc RWL_16 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9566 x859/junc0 x859/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9567 GND x212/junc0 x212/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9568 RBL0_9 RWL_22 x841/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9569 x306/junc0 x306/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9570 x477/junc0 x477/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9571 WBL_4 WWL_3 x867/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9572 x695/junc1 WWL_15 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9573 x949/junc1 WWL_19 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9574 RBL0_28 RWL_20 x711/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9575 VDD x699/junc0 x699/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9576 x1015/RWL0_junc x1015/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9577 x1012/RWL0_junc x1012/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9578 VDD x489/junc0 x489/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9579 x104/junc1 WWL_4 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9580 WBL_19 WWL_1 x419/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9581 GND x623/junc1 x623/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9582 RBL0_3 RWL_5 x480/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9583 x562/junc0 x562/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9584 x362/RWL1_junc RWL_0 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9585 WBL_12 WWL_19 x868/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9586 WBL_3 WWL_27 x150/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9587 x826/RWL0_junc x826/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9588 WBL_1 WWL_8 x977/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9589 x893/junc0 x893/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9590 x498/junc0 x498/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9591 GND x134/junc0 x134/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9592 GND x100/junc0 x100/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9593 x125/junc1 WWL_0 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9594 VDD x710/junc0 x710/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9595 x983/junc0 x983/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9596 GND x830/junc1 x830/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9597 WBL_6 WWL_25 x342/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9598 RBL0_21 RWL_1 x721/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9599 VDD x338/junc0 x338/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9600 x71/junc0 x71/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9601 x109/RWL0_junc x109/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9602 x666/junc0 x666/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9603 x376/RWL1_junc RWL_4 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9604 x332/RWL1_junc RWL_8 RBL1_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9605 x715/junc1 WWL_26 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9606 x994/junc1 WWL_22 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9607 VDD x716/junc0 x716/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9608 RBL0_28 RWL_9 x317/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9609 WBL_21 WWL_23 x358/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9610 RBL0_20 RWL_13 x447/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9611 RBL0_5 RWL_27 x727/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9612 x782/junc0 x782/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9613 VDD x604/junc0 x604/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9614 x345/junc0 x345/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9615 GND x441/junc0 x441/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9616 RBL0_9 RWL_23 x853/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9617 WBL_4 WWL_4 x451/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9618 x144/junc1 WWL_20 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9619 x37/junc1 WWL_16 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9620 VDD x720/junc0 x720/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9621 GND x128/junc0 x128/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9622 GND x422/junc0 x422/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9623 GND x646/junc1 x646/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9624 GND x304/junc1 x304/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9625 x929/RWL0_junc x929/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9626 x832/RWL0_junc x832/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9627 x842/junc0 x842/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9628 VDD x762/junc0 x762/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9629 x877/junc0 x877/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9630 GND x1003/junc1 x1003/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9631 x408/RWL1_junc RWL_1 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9632 x331/junc1 WWL_3 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9633 WBL_12 WWL_20 x461/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9634 RBL0_6 RWL_4 x742/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9635 x880/junc0 x880/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9636 x834/RWL0_junc x834/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9637 GND x143/junc0 x143/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9638 x986/junc0 x986/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9639 x530/junc0 x530/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9640 x529/junc0 x529/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9641 WBL_0 WWL_25 x591/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9642 x532/junc0 x532/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9643 x996/junc1 WWL_5 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9644 GND x148/junc0 x148/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9645 x413/RWL1_junc RWL_7 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9646 GND x840/junc1 x840/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9647 GND x152/junc0 x152/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9648 x172/junc1 WWL_1 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9649 VDD x731/junc0 x731/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9650 GND x327/junc1 x327/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9651 WBL_6 WWL_26 x395/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9652 x837/RWL0_junc x837/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9653 x632/RWL1_junc RWL_28 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9654 VDD x361/junc0 x361/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9655 x77/junc1 WWL_19 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9656 x838/RWL0_junc x838/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9657 x420/RWL1_junc RWL_5 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9658 RBL0_29 RWL_6 x956/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9659 x79/junc1 WWL_12 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9660 GND x1016/junc1 x1016/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9661 x997/junc1 WWL_23 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9662 x389/junc0 x389/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9663 x184/junc1 WWL_27 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9664 WBL_21 WWL_24 x933/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9665 RBL0_14 RWL_20 x866/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9666 VDD x737/junc0 x737/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9667 x917/RWL1_junc RWL_17 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9668 VDD x367/junc0 x367/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9669 RBL0_25 RWL_28 x741/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9670 x829/RWL1_junc RWL_13 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9671 x381/RWL1_junc RWL_27 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9672 x693/junc0 x693/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9673 x504/junc1 WWL_29 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9674 GND x61/junc0 x61/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9675 GND x1004/junc1 x1004/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9676 GND x459/junc0 x459/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9677 x844/RWL1_junc RWL_28 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9678 GND x344/junc1 x344/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9679 x938/RWL0_junc x938/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9680 x841/RWL0_junc x841/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9681 VDD x524/junc0 x524/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9682 x558/junc0 x558/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9683 WBL_18 WWL_5 x616/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9684 GND x895/junc1 x895/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9685 GND x292/junc0 x292/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9686 x207/junc1 WWL_4 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9687 RBL0_6 RWL_5 x751/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9688 x415/junc0 x415/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9689 x991/junc0 x991/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9690 GND x196/junc0 x196/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9691 x865/junc0 x865/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9692 WBL_0 WWL_26 x893/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9693 x386/RWL1_junc RWL_20 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9694 WBL_17 WWL_17 x498/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9695 x566/junc0 x566/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9696 RBL0_1 RWL_21 x833/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9697 GND x852/junc1 x852/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9698 x421/junc0 x421/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9699 x452/RWL1_junc RWL_8 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9700 RBL0_14 RWL_9 x873/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9701 GND x998/junc1 x998/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9702 WBL_6 WWL_27 x983/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9703 x653/RWL1_junc RWL_30 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9704 x504/RWL1_junc RWL_29 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9705 x847/RWL0_junc x847/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9706 x799/junc0 x799/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9707 VDD x406/junc0 x406/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9708 x41/junc1 WWL_24 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9709 x950/junc1 WWL_20 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9710 x502/junc1 WWL_13 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9711 x848/RWL0_junc x848/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9712 GND x564/junc1 x564/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9713 WBL_9 WWL_2 x782/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9714 GND x210/junc0 x210/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9715 x928/RWL1_junc RWL_18 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9716 RBL0_21 RWL_30 x385/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9717 RBL0_25 RWL_29 x515/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9718 RBL0_19 RWL_17 x879/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9719 VDD x815/junc0 x815/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9720 GND x854/junc1 x854/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9721 RBL0_18 RWL_21 x762/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9722 x714/junc0 x714/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9723 VDD x45/junc0 x45/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9724 GND x346/junc0 x346/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9725 WBL_8 WWL_14 x273/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9726 GND x856/junc1 x856/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9727 GND x1007/junc1 x1007/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9728 x734/RWL1_junc RWL_24 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9729 x467/RWL1_junc RWL_29 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9730 VDD x418/junc0 x418/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9731 x853/RWL0_junc x853/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9732 x674/RWL0_junc x674/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9733 VDD x52/junc0 x52/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9734 GND x325/junc0 x325/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9735 GND x225/junc0 x225/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9736 x417/RWL1_junc RWL_9 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9737 x995/junc0 x995/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9738 VDD x494/junc0 x494/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9739 x966/junc1 WWL_9 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9740 x918/junc0 x918/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9741 x369/junc0 x369/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9742 x454/junc0 x454/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9743 GND x236/junc0 x236/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9744 WBL_26 WWL_10 x986/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9745 GND x240/junc0 x240/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9746 x876/junc0 x876/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9747 WBL_0 WWL_27 x529/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9748 RBL0_10 RWL_14 x772/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9749 WBL_25 WWL_14 x530/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9750 GND x1023/junc1 x1023/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9751 RBL0_1 RWL_22 x246/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9752 WBL_17 WWL_18 x532/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9753 GND x409/junc1 x409/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9754 WBL_28 WWL_28 x809/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9755 x935/RWL1_junc RWL_21 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9756 x857/RWL0_junc x857/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9757 x811/junc0 x811/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9758 x433/junc1 WWL_5 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9759 VDD x442/junc0 x442/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9760 VDD x534/junc0 x534/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9761 GND x527/junc1 x527/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9762 x561/RWL1_junc RWL_19 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9763 x955/junc1 WWL_17 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9764 x903/junc0 x903/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9765 VDD x450/junc0 x450/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9766 x283/junc1 WWL_21 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9767 RBL0_18 RWL_22 x2/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9768 RBL0_19 RWL_18 x890/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9769 x468/junc0 x468/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9770 GND x869/junc1 x869/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9771 x956/RWL0_junc x956/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9772 VDD x506/junc0 x506/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9773 x1021/RWL1_junc RWL_17 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9774 x500/RWL1_junc RWL_25 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9775 x866/RWL0_junc x866/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9776 VDD x812/junc0 x812/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9777 x926/junc0 x926/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9778 GND x871/junc1 x871/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9779 GND x523/junc0 x523/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9780 GND x366/junc0 x366/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9781 x19/RWL1_junc RWL_2 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9782 GND x275/junc0 x275/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9783 x843/junc0 x843/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9784 x8/junc1 WWL_2 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9785 WBL_2 WWL_21 x558/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9786 VDD x526/junc0 x526/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9787 x485/RWL0_junc x485/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9788 x887/junc0 x887/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9789 x176/junc0 x176/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9790 WBL_22 WWL_15 x328/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9791 x829/junc0 x829/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9792 GND x286/junc0 x286/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9793 x888/junc0 x888/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9794 x298/junc1 WWL_14 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9795 WBL_26 WWL_11 x991/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9796 RBL0_10 RWL_15 x795/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9797 GND x1002/junc1 x1002/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9798 x484/junc0 x484/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9799 RBL0_1 RWL_23 x291/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9800 x629/junc0 x629/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9801 WBL_24 WWL_30 x981/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9802 GND x878/junc1 x878/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9803 x590/RWL1_junc RWL_22 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9804 x7/RWL0_junc x7/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9805 x793/junc0 x793/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9806 VDD x1013/junc0 x1013/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9807 RBL0_4 RWL_21 x896/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9808 x555/RWL1_junc RWL_31 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9809 x873/RWL0_junc x873/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9810 x964/junc1 WWL_18 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9811 x319/junc1 WWL_14 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9812 x911/junc0 x911/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9813 VDD x476/junc0 x476/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9814 RBL0_18 RWL_23 x55/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9815 RBL0_19 RWL_19 x900/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9816 VDD x607/junc0 x607/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9817 x1022/RWL1_junc RWL_18 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9818 x863/RWL1_junc RWL_26 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9819 x583/junc0 x583/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9820 x36/junc0 x36/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9821 GND x886/junc1 x886/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9822 GND x560/junc0 x560/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9823 GND x412/junc0 x412/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9824 x924/junc1 WWL_30 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9825 x867/RWL1_junc RWL_3 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9826 x516/RWL0_junc x516/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9827 x879/RWL0_junc x879/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9828 GND x312/junc0 x312/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9829 WBL_11 WWL_14 x995/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9830 x145/RWL0_junc x145/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9831 x881/RWL0_junc x881/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9832 x203/junc1 WWL_28 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9833 GND x34/junc0 x34/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9834 VDD x685/junc0 x685/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9835 WBL_30 WWL_12 x918/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9836 GND x957/junc1 x957/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9837 WBL_22 WWL_16 x369/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9838 x514/junc0 x514/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9839 RBL0_10 RWL_16 x808/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9840 x50/RWL0_junc x50/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9841 x184/RWL1_junc RWL_27 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9842 WBL_24 WWL_31 x604/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9843 x802/junc1 WWL_25 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9844 VDD x98/junc0 x98/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9845 GND x478/junc1 x478/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9846 x621/RWL1_junc RWL_23 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9847 x969/junc1 WWL_21 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9848 x806/junc0 x806/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9849 RBL0_4 RWL_22 x905/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9850 VDD x507/junc0 x507/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9851 x267/junc1 WWL_15 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9852 x979/junc1 WWL_19 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9853 VDD x805/junc0 x805/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9854 RBL0_23 RWL_20 x812/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9855 x684/RWL0_junc x684/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9856 VDD x639/junc0 x639/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9857 x671/RWL1_junc RWL_31 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9858 RBL0_31 RWL_24 x821/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9859 WBL_15 WWL_29 x250/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9860 x897/RWL1_junc RWL_19 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9861 x767/junc0 x767/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9862 x922/junc0 x922/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9863 x923/junc0 x923/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9864 WBL_21 WWL_29 x54/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9865 x573/RWL1_junc RWL_0 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9866 x260/junc0 x260/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9867 GND x499/junc1 x499/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9868 WBL_7 WWL_19 x926/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9869 x889/RWL0_junc x889/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9870 x117/junc0 x117/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9871 x932/junc1 WWL_31 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9872 x890/RWL0_junc x890/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9873 GND x90/junc0 x90/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9874 WBL_31 WWL_9 x176/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9875 VDD x705/junc0 x705/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9876 x936/RWL0_junc x936/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9877 WBL_30 WWL_13 x829/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9878 x378/junc1 WWL_0 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9879 GND x894/junc1 x894/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9880 x107/RWL0_junc x107/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9881 x640/RWL1_junc RWL_6 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9882 x211/RWL1_junc RWL_31 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9883 x391/junc1 WWL_21 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9884 x950/RWL1_junc RWL_20 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9885 x16/junc0 x16/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9886 x582/RWL1_junc RWL_4 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9887 RBL0_23 RWL_9 x533/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9888 x817/junc1 WWL_26 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9889 x97/junc1 WWL_22 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9890 VDD x818/junc0 x818/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9891 GND x510/junc1 x510/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9892 x19/junc0 x19/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9893 x22/junc0 x22/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9894 RBL0_4 RWL_23 x913/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9895 GND x466/junc0 x466/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9896 VDD x839/junc0 x839/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9897 GND x901/junc1 x901/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9898 x403/junc1 WWL_20 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9899 x307/junc1 WWL_16 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9900 x30/junc0 x30/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9901 VDD x229/junc0 x229/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9902 x126/junc0 x126/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9903 x786/junc0 x786/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9904 GND x380/junc0 x380/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9905 GND x891/junc1 x891/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9906 VDD x227/junc0 x227/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9907 GND x525/junc1 x525/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9908 RBL0_31 RWL_25 x163/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9909 x965/RWL0_junc x965/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9910 x896/RWL0_junc x896/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9911 GND x1009/junc1 x1009/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9912 x606/RWL1_junc RWL_1 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9913 RBL0_15 RWL_2 x646/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9914 x129/junc1 WWL_3 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9915 WBL_1 WWL_5 x584/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9916 WBL_16 WWL_12 x583/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9917 WBL_7 WWL_20 x36/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9918 x898/RWL0_junc x898/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9919 x933/junc0 x933/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9920 x900/RWL0_junc x900/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9921 x143/junc0 x143/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9922 x56/junc0 x56/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9923 x180/RWL1_junc RWL_2 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9924 x182/RWL1_junc RWL_9 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9925 GND x140/junc0 x140/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9926 GND x1010/junc0 x1010/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9927 x953/RWL1_junc RWL_7 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9928 x423/junc1 WWL_1 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9929 GND x541/junc1 x541/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9930 x752/RWL1_junc RWL_28 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9931 x158/RWL0_junc x158/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9932 RBL0_20 RWL_10 x840/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9933 GND x489/junc0 x489/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9934 VDD x849/junc0 x849/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9935 x339/junc1 WWL_19 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9936 x74/junc0 x74/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9937 x616/RWL1_junc RWL_5 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9938 RBL0_24 RWL_6 x920/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9939 x151/junc1 WWL_23 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9940 x435/junc1 WWL_27 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9941 RBL0_9 RWL_20 x89/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9942 VDD x827/junc0 x827/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9943 x955/RWL1_junc RWL_17 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9944 VDD x577/junc0 x577/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9945 RBL0_4 RWL_28 x58/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9946 x387/RWL1_junc RWL_31 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9947 GND x496/junc0 x496/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9948 x201/RWL1_junc RWL_13 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9949 x586/RWL1_junc RWL_27 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9950 x83/junc0 x83/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9951 VDD x851/junc0 x851/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9952 x87/junc0 x87/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9953 x764/junc1 WWL_29 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9954 GND x556/junc1 x556/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9955 x940/junc1 WWL_2 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9956 x173/junc0 x173/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9957 GND x424/junc0 x424/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9958 GND x1011/junc1 x1011/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9959 GND x902/junc1 x902/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9960 x970/RWL0_junc x970/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9961 x904/RWL0_junc x904/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9962 RBL0_31 RWL_26 x208/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9963 x905/RWL0_junc x905/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9964 VDD x642/junc0 x642/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9965 WBL_27 WWL_3 x468/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9966 GND x943/junc1 x943/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9967 RBL0_15 x61/RWL1 x344/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9968 WBL_16 WWL_13 x260/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9969 x453/junc1 WWL_4 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9970 x907/RWL0_junc x907/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9971 x612/junc0 x612/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9972 GND x308/junc0 x308/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9973 x298/RWL1_junc RWL_14 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9974 x196/junc0 x196/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9975 VDD x221/junc0 x221/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9976 x111/junc0 x111/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9977 x681/RWL1_junc RWL_3 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9978 x114/junc0 x114/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9979 x961/RWL1_junc RWL_8 RBL1_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9980 RBL0_9 RWL_9 x930/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9981 x402/RWL1_junc RWL_30 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9982 x987/junc1 WWL_6 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9983 x764/RWL1_junc RWL_29 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9984 x121/junc0 x121/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9985 RBL0_28 RWL_7 x839/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9986 RBL0_20 RWL_11 x852/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9987 GND x520/junc0 x520/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9988 VDD x859/junc0 x859/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9989 x34/junc1 WWL_24 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9990 x980/junc1 WWL_20 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9991 x641/RWL1_junc RWL_10 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9992 WBL_4 WWL_2 x19/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9993 GND x455/junc0 x455/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9994 x964/RWL1_junc RWL_18 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9995 x230/junc0 x230/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9996 RBL0_4 RWL_29 x683/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9997 VDD x248/junc0 x248/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M9998 GND x914/junc1 x914/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M9999 GND x528/junc0 x528/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10000 x135/junc0 x135/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10001 GND x457/junc0 x457/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10002 x243/junc0 x243/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10003 GND x589/junc1 x589/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10004 WBL_12 WWL_6 x30/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10005 x139/junc0 x139/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10006 GND x909/junc1 x909/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10007 RBL0_31 RWL_28 x593/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10008 WBL_3 WWL_14 x126/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10009 GND x916/junc1 x916/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10010 GND x1012/junc1 x1012/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10011 VDD x94/junc0 x94/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10012 GND x654/junc0 x654/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10013 VDD x615/junc0 x615/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10014 x785/RWL0_junc x785/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10015 x912/RWL0_junc x912/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10016 x913/RWL0_junc x913/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10017 VDD x328/junc0 x328/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10018 GND x539/junc0 x539/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10019 GND x565/junc0 x565/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10020 WBL_27 WWL_4 x132/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10021 x225/junc0 x225/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10022 GND x59/junc0 x59/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10023 x155/junc0 x155/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10024 x157/junc0 x157/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10025 x635/junc0 x635/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10026 GND x471/junc0 x471/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10027 GND x350/junc0 x350/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10028 x340/RWL1_junc RWL_15 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10029 WBL_21 WWL_10 x143/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10030 x263/junc0 x263/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10031 RBL0_5 RWL_14 x171/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10032 WBL_7 WWL_28 x1013/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10033 x14/junc1 WWL_3 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10034 x130/junc1 WWL_7 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10035 x969/RWL1_junc RWL_21 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10036 x60/RWL0_junc x60/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10037 RBL0_29 RWL_4 x1023/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10038 x168/junc0 x168/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10039 RBL0_28 RWL_8 x851/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10040 RBL0_20 RWL_12 x409/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10041 VDD x628/junc0 x628/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10042 GND x557/junc0 x557/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10043 x924/RWL1_junc RWL_30 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10044 x665/RWL1_junc RWL_11 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10045 x712/RWL1_junc RWL_19 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10046 VDD x29/junc0 x29/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10047 x178/junc0 x178/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10048 VDD x679/junc0 x679/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10049 GND x38/junc0 x38/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10050 x287/junc0 x287/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10051 x185/junc0 x185/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10052 x288/junc0 x288/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10053 RBL0_27 RWL_30 x84/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10054 WBL_12 WWL_7 x87/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10055 GND x915/junc1 x915/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10056 RBL0_31 RWL_29 x71/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10057 GND x927/junc1 x927/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10058 x920/RWL0_junc x920/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10059 x814/RWL1_junc RWL_17 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10060 VDD x637/junc0 x637/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10061 x89/RWL0_junc x89/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10062 x599/junc0 x599/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10063 VDD x877/junc0 x877/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10064 x191/junc0 x191/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10065 x195/junc0 x195/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10066 x921/RWL0_junc x921/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10067 GND x495/junc0 x495/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10068 GND x576/junc0 x576/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10069 GND x25/junc0 x25/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10070 GND x704/junc0 x704/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10071 x275/junc0 x275/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10072 x293/junc1 WWL_2 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10073 GND x115/junc0 x115/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10074 GND x63/junc1 x63/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10075 GND x973/junc1 x973/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10076 x197/junc0 x197/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10077 x427/junc0 x427/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10078 WBL_17 WWL_15 x779/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10079 x201/junc0 x201/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10080 GND x503/junc0 x503/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10081 x57/junc1 WWL_6 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10082 x517/junc1 WWL_10 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10083 x383/RWL1_junc RWL_16 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10084 x205/junc0 x205/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10085 RBL0_14 RWL_7 x215/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10086 x518/junc1 WWL_14 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10087 WBL_21 WWL_11 x196/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10088 RBL0_5 RWL_15 x860/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10089 WBL_3 WWL_30 x768/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10090 x209/junc0 x209/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10091 GND x931/junc1 x931/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10092 x657/RWL1_junc RWL_14 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10093 x984/junc1 WWL_4 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10094 x730/RWL1_junc RWL_22 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10095 RBL0_29 RWL_5 x1002/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10096 x175/junc1 WWL_8 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10097 x116/RWL0_junc x116/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10098 RBL0_14 RWL_31 x998/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10099 x930/RWL0_junc x930/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10100 x918/RWL1_junc RWL_12 RBL1_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10101 VDD x85/junc0 x85/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10102 x218/junc0 x218/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10103 VDD x86/junc0 x86/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10104 x222/junc0 x222/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10105 GND x1015/junc0 x1015/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10106 VDD x702/junc0 x702/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10107 WBL_8 WWL_12 x22/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10108 WBL_12 WWL_8 x139/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10109 GND x194/junc0 x194/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10110 x826/RWL1_junc RWL_18 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10111 VDD x336/junc0 x336/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10112 x658/RWL1_junc RWL_7 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10113 x725/junc0 x725/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10114 x238/junc0 x238/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10115 x241/junc0 x241/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10116 GND x610/junc0 x610/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10117 WBL_6 WWL_14 x225/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10118 GND x999/junc1 x999/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10119 x934/RWL0_junc x934/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10120 GND x534/junc0 x534/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10121 VDD x865/junc0 x865/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10122 WBL_25 WWL_12 x155/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10123 x689/RWL0_junc x689/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10124 GND x982/junc1 x982/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10125 RBL0_1 RWL_20 x923/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10126 WBL_17 WWL_16 x157/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10127 x988/junc1 WWL_0 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10128 x989/junc1 WWL_7 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10129 x552/junc1 WWL_11 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10130 RBL0_14 RWL_8 x262/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10131 x253/junc0 x253/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10132 x254/junc0 x254/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10133 RBL0_5 RWL_16 x872/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10134 GND x319/junc0 x319/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10135 VDD x799/junc0 x799/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10136 x435/RWL1_junc RWL_27 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10137 WBL_3 WWL_31 x244/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10138 GND x939/junc1 x939/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10139 GND x655/junc1 x655/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10140 x680/RWL1_junc RWL_15 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10141 x746/RWL1_junc RWL_23 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10142 VDD x675/junc0 x675/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10143 x131/junc1 WWL_15 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10144 x1000/junc1 WWL_19 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10145 x231/junc1 WWL_30 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10146 RBL0_18 RWL_20 x877/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10147 x102/RWL0_junc x102/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10148 x269/junc0 x269/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10149 VDD x723/junc0 x723/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10150 WBL_8 WWL_13 x594/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10151 x1023/RWL0_junc x1023/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10152 RBL0_26 RWL_24 x880/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10153 x154/junc0 x154/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10154 x186/junc0 x186/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10155 x834/RWL1_junc RWL_19 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10156 x845/junc0 x845/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10157 x960/junc0 x960/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10158 x717/RWL1_junc RWL_0 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10159 WBL_15 WWL_21 x599/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10160 WBL_0 WWL_14 x191/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10161 x486/junc0 x486/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10162 x678/RWL1_junc RWL_8 RBL1_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10163 RBL0_1 RWL_9 x786/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10164 WBL_2 WWL_19 x195/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10165 x372/junc0 x372/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10166 x189/RWL0_junc x189/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10167 VDD x688/junc0 x688/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10168 GND x570/junc0 x570/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10169 GND x572/junc0 x572/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10170 VDD x690/junc0 x690/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10171 x159/junc1 WWL_12 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10172 WBL_26 WWL_9 x427/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10173 VDD x876/junc0 x876/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10174 x709/RWL0_junc x709/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10175 GND x941/junc1 x941/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10176 WBL_25 WWL_13 x201/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10177 x446/RWL0_junc x446/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10178 GND x942/junc1 x942/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10179 x992/junc1 WWL_8 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10180 x993/junc1 WWL_1 WBLb_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10181 GND x874/junc1 x874/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10182 x295/junc0 x295/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10183 x265/junc1 WWL_28 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10184 GND x363/junc0 x363/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10185 x756/RWL1_junc RWL_6 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10186 x980/RWL1_junc RWL_20 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10187 VDD x811/junc0 x811/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10188 RBL0_10 RWL_31 x1006/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10189 RBL0_18 RWL_9 x693/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10190 GND x944/junc1 x944/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10191 GND x677/junc1 x677/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10192 x703/RWL1_junc RWL_16 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10193 GND x648/junc0 x648/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10194 x215/RWL0_junc x215/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10195 x91/junc0 x91/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10196 VDD x903/junc0 x903/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10197 x367/junc1 WWL_12 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10198 x177/junc1 WWL_16 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10199 GND x1014/junc1 x1014/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10200 x276/junc1 WWL_20 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10201 x304/junc0 x304/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10202 x663/junc1 WWL_31 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10203 GND x187/junc0 x187/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10204 x968/junc0 x968/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10205 x1002/RWL0_junc x1002/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10206 RBL0_26 RWL_25 x415/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10207 x6/junc0 x6/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10208 x313/junc0 x313/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10209 x316/junc0 x316/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10210 x390/junc0 x390/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10211 x738/RWL1_junc RWL_1 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10212 RBL0_10 RWL_2 x891/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10213 WBL_11 WWL_12 x725/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10214 x416/junc0 x416/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10215 WBL_2 WWL_20 x241/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10216 x237/RWL0_junc x237/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10217 VDD x887/junc0 x887/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10218 WBL_27 WWL_29 x302/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10219 x327/junc0 x327/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10220 GND x602/junc0 x602/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10221 x434/RWL1_junc RWL_9 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10222 GND x605/junc0 x605/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10223 VDD x888/junc0 x888/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10224 x760/junc1 WWL_13 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10225 GND x946/junc1 x946/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10226 VDD x744/junc0 x744/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10227 GND x698/junc1 x698/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10228 VDD x770/junc0 x770/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10229 x297/junc1 WWL_30 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10230 x334/junc0 x334/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10231 WBL_29 WWL_22 x254/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10232 GND x639/junc0 x639/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10233 GND x947/junc1 x947/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10234 GND x407/junc0 x407/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10235 VDD x793/junc0 x793/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10236 x213/junc1 WWL_19 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10237 RBL0_19 RWL_6 x958/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10238 GND x4/junc1 x4/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10239 x257/RWL0_junc x257/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10240 RBL0_4 RWL_20 x349/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10241 VDD x719/junc0 x719/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10242 GND x672/junc0 x672/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10243 x397/RWL0_junc x397/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10244 x262/RWL0_junc x262/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10245 x447/RWL1_junc RWL_13 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10246 x727/RWL1_junc RWL_27 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10247 x343/junc0 x343/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10248 x815/junc1 WWL_13 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10249 VDD x911/junc0 x911/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10250 x776/junc0 x776/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10251 x347/junc0 x347/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10252 GND x707/junc1 x707/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10253 GND x226/junc0 x226/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10254 x972/junc0 x972/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10255 x247/junc0 x247/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10256 x357/junc0 x357/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10257 RBL0_26 RWL_26 x454/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10258 x360/junc0 x360/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10259 WBL_22 WWL_3 x186/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10260 x433/junc0 x433/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10261 VDD x754/junc0 x754/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10262 RBL0_10 x61/RWL1 x902/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10263 x456/junc0 x456/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10264 WBL_11 WWL_13 x486/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10265 x948/RWL0_junc x948/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10266 x368/junc0 x368/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10267 WBL_14 WWL_25 x830/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10268 x518/RWL1_junc RWL_14 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10269 VDD x464/junc0 x464/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10270 GND x165/junc1 x165/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10271 x973/junc0 x973/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10272 GND x627/junc0 x627/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10273 VDD x514/junc0 x514/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10274 RBL0_4 RWL_9 x966/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10275 GND x48/junc1 x48/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10276 VDD x553/junc0 x553/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10277 x984/RWL1_junc RWL_4 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10278 VDD x654/junc0 x654/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10279 x148/junc1 WWL_6 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10280 x152/junc1 WWL_19 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10281 x375/junc0 x375/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10282 RBL0_23 RWL_7 x903/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10283 RBL0_13 RWL_27 x820/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10284 x251/junc1 WWL_31 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10285 GND x50/junc1 x50/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10286 WBL_29 WWL_23 x295/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10287 GND x899/junc0 x899/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10288 VDD x806/junc0 x806/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10289 x1001/junc1 WWL_20 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10290 x156/RWL1_junc RWL_28 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10291 x757/RWL1_junc RWL_10 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10292 GND x636/junc0 x636/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10293 x467/junc0 x467/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10294 x956/RWL1_junc RWL_6 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10295 VDD x473/junc0 x473/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10296 x242/RWL0_junc x242/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10297 x300/junc0 x300/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10298 GND x65/junc1 x65/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10299 GND x691/junc0 x691/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10300 x974/junc0 x974/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10301 x975/junc0 x975/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10302 x393/junc0 x393/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10303 x457/junc0 x457/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10304 GND x271/junc0 x271/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10305 x398/junc0 x398/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10306 GND x729/junc1 x729/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10307 WBL_7 WWL_6 x304/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10308 RBL0_10 RWL_28 x475/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10309 GND x73/junc1 x73/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10310 GND x954/junc1 x954/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10311 VDD x280/junc0 x280/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10312 VDD x697/junc0 x697/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10313 x200/junc1 WWL_29 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10314 x749/junc0 x749/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10315 x404/junc0 x404/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10316 RBL0_15 RWL_0 x909/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10317 WBL_30 WWL_0 x316/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10318 WBL_22 WWL_4 x390/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10319 x409/junc0 x409/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10320 x988/RWL1_junc RWL_0 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10321 GND x371/junc0 x371/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10322 x989/RWL1_junc RWL_7 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10323 WBL_14 WWL_26 x327/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10324 x554/RWL1_junc RWL_15 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10325 x487/junc0 x487/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10326 x901/RWL0_junc x901/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10327 x999/junc0 x999/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10328 x831/RWL1_junc RWL_5 RBL1_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10329 x296/junc1 WWL_3 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10330 x384/junc1 WWL_7 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10331 x419/junc0 x419/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10332 RBL0_24 RWL_4 x432/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10333 GND x107/junc1 x107/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10334 WBL_29 WWL_24 x334/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10335 x386/junc1 WWL_20 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10336 VDD x748/junc0 x748/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10337 RBL0_23 RWL_8 x911/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10338 GND x908/junc0 x908/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10339 x122/junc0 x122/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10340 x200/RWL1_junc RWL_29 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10341 GND x509/junc1 x509/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10342 GND x711/junc0 x711/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10343 x777/RWL1_junc RWL_11 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10344 x150/junc0 x150/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10345 GND x962/junc1 x962/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10346 x763/junc0 x763/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10347 x732/junc0 x732/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10348 x977/junc0 x977/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10349 x436/junc0 x436/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10350 GND x309/junc0 x309/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10351 x38/junc0 x38/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10352 x504/junc0 x504/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10353 GND x654/junc1 x654/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10354 WBL_7 WWL_7 x347/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10355 RBL0_10 RWL_29 x491/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10356 GND x127/junc1 x127/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10357 GND x963/junc1 x963/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10358 x958/RWL0_junc x958/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10359 VDD x797/junc0 x797/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10360 x349/RWL0_junc x349/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10361 x42/junc0 x42/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10362 x509/junc0 x509/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10363 x72/RWL0_junc x72/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10364 GND x965/junc1 x965/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10365 GND x490/junc0 x490/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10366 WBL_30 WWL_1 x360/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10367 RBL0_15 RWL_1 x915/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10368 GND x138/junc1 x138/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10369 x75/junc1 WWL_2 WBLb_3 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10370 x497/RWL0_junc x497/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10371 x444/junc0 x444/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10372 x619/junc0 x619/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10373 x231/RWL1_junc RWL_30 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10374 x502/RWL0_junc x502/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10375 x447/junc0 x447/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10376 GND x809/junc0 x809/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10377 x992/RWL1_junc RWL_8 RBL1_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10378 x993/RWL1_junc RWL_1 RBL1_1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10379 GND x1017/junc0 x1017/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10380 x329/junc1 WWL_6 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10381 x685/junc1 WWL_10 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10382 x587/RWL1_junc RWL_16 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10383 x451/junc0 x451/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10384 RBL0_9 RWL_7 x458/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10385 WBL_14 WWL_27 x368/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10386 x686/junc1 WWL_14 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10387 x556/RWL0_junc x556/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10388 x66/junc0 x66/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10389 x68/junc0 x68/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10390 GND x317/junc0 x317/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10391 x772/RWL1_junc RWL_14 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10392 x1003/junc1 WWL_4 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10393 RBL0_24 RWL_5 x976/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10394 x426/junc1 WWL_8 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10395 VDD x536/junc0 x536/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10396 GND x266/junc1 x266/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10397 GND x158/junc1 x158/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10398 x443/RWL0_junc x443/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10399 VDD x733/junc0 x733/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10400 GND x755/junc1 x755/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10401 RBL0_27 RWL_17 x836/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10402 GND x544/junc1 x544/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10403 x966/RWL0_junc x966/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10404 x155/RWL1_junc RWL_12 RBL1_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10405 RBL0_16 RWL_27 x922/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10406 VDD x82/junc0 x82/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10407 VDD x83/junc0 x83/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10408 x461/junc0 x461/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10409 RBL0_31 RWL_13 x767/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10410 WBL_3 WWL_12 x300/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10411 x787/junc0 x787/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10412 VDD x352/junc0 x352/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10413 WBL_16 WWL_0 x457/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10414 WBL_7 WWL_8 x398/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10415 GND x353/junc0 x353/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10416 x265/RWL1_junc RWL_28 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10417 VDD x810/junc0 x810/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10418 WBL_27 WWL_2 x714/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10419 GND x179/junc1 x179/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10420 x825/junc0 x825/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10421 x544/junc0 x544/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10422 GND x970/junc1 x970/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10423 x531/RWL0_junc x531/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10424 GND x425/junc0 x425/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10425 RBL0_23 RWL_28 x766/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10426 GND x981/junc0 x981/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10427 GND x822/junc0 x822/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10428 x1004/junc1 WWL_7 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10429 x705/junc1 WWL_11 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10430 RBL0_9 RWL_8 x488/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10431 GND x766/junc1 x766/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10432 x478/junc0 x478/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10433 x477/junc0 x477/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10434 x589/RWL0_junc x589/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10435 GND x699/junc0 x699/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10436 x286/junc1 WWL_5 WBLb_30 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10437 x456/junc0 x456/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10438 x119/junc0 x119/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10439 VDD x121/junc0 x121/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10440 GND x198/junc1 x198/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10441 x483/junc0 x483/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10442 x795/RWL1_junc RWL_15 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10443 x546/RWL0_junc x546/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10444 x562/junc0 x562/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10445 VDD x388/junc0 x388/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10446 VDD x791/junc0 x791/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10447 GND x1015/junc1 x1015/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10448 RBL0_27 RWL_18 x846/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10449 x8/RWL0_junc x8/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10450 x284/RWL0_junc x284/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10451 WBL_12 WWL_5 x869/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10452 x149/RWL0_junc x149/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10453 WBL_3 WWL_13 x732/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10454 x432/RWL0_junc x432/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10455 WBL_16 WWL_1 x38/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10456 RBL0_21 RWL_24 x933/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10457 VDD x141/junc0 x141/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10458 x498/junc0 x498/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10459 x437/junc0 x437/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10460 x501/junc0 x501/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10461 x499/junc0 x499/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10462 RBL0_18 RWL_31 x1015/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10463 x302/RWL1_junc RWL_29 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10464 x910/junc0 x910/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10465 x634/RWL1_junc RWL_2 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10466 GND x710/junc0 x710/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10467 x983/junc0 x983/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10468 GND x220/junc1 x220/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10469 WBL_10 WWL_21 x42/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10470 x660/junc0 x660/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10471 x438/RWL0_junc x438/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10472 x3/junc0 x3/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10473 GND x785/junc1 x785/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10474 VDD x798/junc0 x798/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10475 x568/RWL0_junc x568/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10476 RBL0_23 RWL_29 x230/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10477 GND x716/junc0 x716/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10478 x160/junc0 x160/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10479 VDD x800/junc0 x800/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10480 x412/junc1 WWL_12 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10481 WBL_21 WWL_9 x619/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10482 GND x232/junc1 x232/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10483 GND x399/junc0 x399/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10484 x1007/junc1 WWL_8 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10485 GND x790/junc1 x790/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10486 GND x230/junc1 x230/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10487 x510/junc0 x510/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10488 x485/junc1 WWL_28 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10489 GND x720/junc0 x720/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10490 x377/junc1 WWL_2 WBLb_31 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10491 x228/RWL1_junc RWL_6 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10492 x1001/RWL1_junc RWL_20 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10493 WBL_28 WWL_17 x66/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10494 VDD x168/junc0 x168/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10495 RBL0_12 RWL_21 x83/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10496 GND x245/junc1 x245/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10497 x808/RWL1_junc RWL_16 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10498 x174/junc0 x174/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10499 x310/RWL0_junc x310/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10500 x919/RWL1_junc RWL_24 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10501 GND x762/junc0 x762/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10502 x458/RWL0_junc x458/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10503 VDD x430/junc0 x430/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10504 VDD x178/junc0 x178/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10505 RBL0_27 RWL_19 x855/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10506 VDD x431/junc0 x431/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10507 x62/RWL0_junc x62/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10508 x525/junc0 x525/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10509 x986/junc0 x986/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10510 RBL0_30 RWL_17 x538/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10511 x530/junc0 x530/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10512 x976/RWL0_junc x976/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10513 x529/junc0 x529/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10514 RBL0_21 RWL_25 x612/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10515 x532/junc0 x532/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10516 x190/junc0 x190/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10517 x192/junc0 x192/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10518 x193/junc0 x193/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10519 x535/junc0 x535/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10520 GND x72/junc0 x72/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10521 x656/RWL1_junc x61/RWL1 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10522 GND x731/junc0 x731/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10523 RBL0_5 RWL_2 x940/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10524 WBL_6 WWL_12 x825/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10525 GND x9/junc1 x9/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10526 x469/RWL0_junc x469/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10527 VDD x197/junc0 x197/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10528 x541/junc0 x541/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10529 GND x737/junc0 x737/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10530 x448/junc1 WWL_5 WBLb_16 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10531 x223/junc1 WWL_9 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10532 x623/RWL1_junc RWL_9 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10533 x203/junc0 x203/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10534 VDD x205/junc0 x205/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10535 GND x1019/junc1 x1019/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10536 x5/junc1 WWL_13 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10537 x0/junc0 x0/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10538 GND x285/junc1 x285/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10539 x516/junc1 WWL_30 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10540 x549/junc0 x549/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10541 WBL_24 WWL_22 x478/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10542 GND x723/junc0 x723/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10543 GND x290/junc1 x290/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10544 GND x743/junc0 x743/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10545 x747/junc1 WWL_21 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10546 WBL_28 WWL_18 x119/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10547 VDD x214/junc0 x214/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10548 RBL0_12 RWL_22 x135/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10549 GND x35/junc1 x35/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10550 x481/RWL0_junc x481/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10551 x556/junc0 x556/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10552 x58/RWL0_junc x58/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10553 x72/junc0 x72/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10554 x351/RWL0_junc x351/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10555 GND x524/junc0 x524/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10556 x244/RWL0_junc x244/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10557 x830/RWL1_junc RWL_25 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10558 GND x2/junc0 x2/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10559 VDD x218/junc0 x218/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10560 x1005/RWL0_junc x1005/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10561 x488/RWL0_junc x488/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10562 VDD x463/junc0 x463/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10563 x558/junc0 x558/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10564 VDD x222/junc0 x222/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10565 x224/junc0 x224/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10566 WBL_13 WWL_29 x697/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10567 x991/junc0 x991/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10568 RBL0_30 RWL_18 x574/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10569 RBL0_21 RWL_26 x635/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10570 x569/junc0 x569/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10571 x566/junc0 x566/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10572 x235/junc0 x235/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10573 WBL_0 WWL_12 x499/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10574 WBL_15 WWL_19 x437/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10575 WBL_17 WWL_3 x501/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10576 x239/junc0 x239/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10577 RBL0_1 RWL_7 x975/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10578 VDD x243/junc0 x243/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10579 RBL0_5 RWL_3 x23/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10580 WBL_6 WWL_13 x660/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10581 x978/RWL0_junc x978/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10582 x249/junc0 x249/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10583 WBL_9 WWL_25 x894/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10584 x686/RWL1_junc RWL_14 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10585 VDD x644/junc0 x644/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10586 GND x315/junc1 x315/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10587 x646/RWL1_junc RWL_2 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10588 GND x32/junc0 x32/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10589 WBL_13 WWL_21 x160/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10590 VDD x253/junc0 x253/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10591 GND x1020/junc1 x1020/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10592 x231/junc0 x231/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10593 GND x323/junc1 x323/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10594 x1003/RWL1_junc RWL_4 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10595 x1010/junc1 WWL_6 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10596 x633/junc1 WWL_31 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10597 WBL_24 WWL_23 x510/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10598 RBL0_18 RWL_7 x178/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10599 RBL0_8 RWL_27 x882/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10600 GND x45/junc0 x45/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10601 VDD x261/junc0 x261/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10602 RBL0_12 RWL_23 x185/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10603 VDD x263/junc0 x263/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10604 WBL_8 WWL_0 x578/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10605 x840/RWL1_junc RWL_10 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10606 x589/junc0 x589/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10607 x683/RWL0_junc x683/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10608 GND x52/junc0 x52/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10609 x920/RWL1_junc RWL_6 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10610 x327/RWL1_junc RWL_26 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10611 x472/RWL0_junc x472/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10612 GND x55/junc0 x55/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10613 x995/junc0 x995/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10614 VDD x269/junc0 x269/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10615 x592/junc0 x592/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10616 x271/junc0 x271/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10617 GND x494/junc0 x494/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10618 x274/junc0 x274/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10619 WBL_2 WWL_6 x525/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10620 x496/junc1 WWL_22 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10621 VDD x277/junc0 x277/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10622 x133/junc0 x133/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10623 x835/junc0 x835/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10624 RBL0_30 RWL_19 x949/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10625 x601/junc0 x601/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10626 WBL_25 WWL_0 x192/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10627 RBL0_10 RWL_0 x73/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10628 WBL_15 WWL_20 x190/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10629 WBL_17 WWL_4 x193/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10630 WBL_0 WWL_13 x535/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10631 RBL0_1 RWL_8 x977/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10632 x334/junc0 x334/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10633 x289/junc0 x289/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10634 GND x647/junc0 x647/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10635 x1004/RWL1_junc RWL_7 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10636 VDD x669/junc0 x669/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10637 GND x355/junc1 x355/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10638 WBL_9 WWL_26 x541/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10639 x706/RWL1_junc RWL_15 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10640 x344/RWL1_junc x61/RWL1 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10641 x1014/RWL0_junc x1014/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10642 GND x862/junc1 x862/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10643 x663/junc0 x663/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10644 x895/RWL1_junc RWL_5 RBL1_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10645 x511/junc1 WWL_3 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10646 x588/junc1 WWL_7 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10647 RBL0_19 RWL_4 x622/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10648 WBL_24 WWL_24 x549/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10649 RBL0_18 RWL_8 x222/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10650 WBL_19 WWL_29 x733/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10651 GND x99/junc0 x99/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10652 GND x506/junc0 x506/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10653 VDD x542/junc0 x542/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10654 WBL_8 WWL_1 x611/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10655 GND x812/junc0 x812/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10656 x852/RWL1_junc RWL_11 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10657 x520/junc1 WWL_25 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10658 x618/junc0 x618/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10659 x788/junc1 WWL_21 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10660 GND x1018/junc1 x1018/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10661 GND x108/junc0 x108/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10662 x843/junc0 x843/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10663 x624/junc0 x624/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10664 x309/junc0 x309/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10665 GND x526/junc0 x526/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10666 WBL_2 WWL_7 x224/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10667 x528/junc1 WWL_23 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10668 VDD x313/junc0 x313/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10669 x318/junc0 x318/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10670 GND x519/junc0 x519/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10671 x794/junc1 WWL_0 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10672 WBL_25 WWL_1 x235/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10673 RBL0_10 RWL_1 x127/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10674 x854/RWL1_junc RWL_27 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10675 GND x396/junc1 x396/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10676 x629/junc0 x629/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10677 x673/RWL0_junc x673/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10678 x326/junc0 x326/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10679 x773/junc1 WWL_29 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10680 GND x670/junc0 x670/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10681 GND x985/junc1 x985/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10682 WBL_20 WWL_17 x804/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10683 GND x1013/junc0 x1013/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10684 x543/junc1 WWL_6 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10685 x1007/RWL1_junc RWL_8 RBL1_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10686 WBL_9 WWL_27 x249/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10687 x728/RWL1_junc RWL_16 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10688 GND x69/junc1 x69/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10689 RBL0_4 RWL_7 x638/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10690 x575/RWL0_junc x575/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10691 x707/RWL0_junc x707/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10692 x932/junc0 x932/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10693 x333/junc0 x333/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10694 GND x533/junc0 x533/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10695 x799/junc1 WWL_0 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10696 x171/RWL1_junc RWL_14 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10697 x1009/junc1 WWL_4 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10698 x617/junc1 WWL_8 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10699 VDD x694/junc0 x694/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10700 RBL0_19 RWL_5 x996/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10701 GND x937/junc1 x937/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10702 GND x257/junc1 x257/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10703 RBL0_22 RWL_17 x154/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10704 x1023/RWL1_junc RWL_4 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10705 x643/junc0 x643/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10706 x409/RWL1_junc RWL_12 RBL1_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10707 x557/junc1 WWL_26 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10708 VDD x341/junc0 x341/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10709 x33/junc0 x33/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10710 RBL0_11 RWL_27 x960/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10711 VDD x342/junc0 x342/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10712 VDD x343/junc0 x343/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10713 x36/junc0 x36/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10714 RBL0_26 RWL_13 x845/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10715 x39/junc0 x39/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10716 VDD x561/junc0 x561/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10717 WBL_11 WWL_0 x271/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10718 x212/RWL0_junc x212/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10719 WBL_2 WWL_8 x274/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10720 x485/RWL1_junc RWL_28 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10721 x608/junc1 WWL_24 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10722 VDD x357/junc0 x357/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10723 GND x685/junc0 x685/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10724 x359/junc0 x359/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10725 WBL_22 WWL_2 x133/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10726 GND x170/junc0 x170/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10727 GND x429/junc1 x429/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10728 x807/junc1 WWL_1 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10729 GND x112/junc1 x112/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10730 x598/RWL0_junc x598/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10731 x600/RWL0_junc x600/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10732 x651/junc0 x651/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10733 x692/RWL0_junc x692/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10734 x495/junc1 WWL_6 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10735 RBL0_2 RWL_28 x844/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10736 WBL_29 WWL_10 x289/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10737 RBL0_13 RWL_14 x904/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10738 WBL_20 WWL_18 x824/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10739 GND x990/junc1 x990/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10740 GND x883/junc0 x883/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10741 x1011/junc1 WWL_7 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10742 RBL0_4 RWL_8 x661/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10743 GND x844/junc1 x844/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10744 x655/junc0 x655/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10745 x695/RWL0_junc x695/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10746 x729/RWL0_junc x729/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10747 GND x805/junc0 x805/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10748 x503/junc1 WWL_5 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10749 x936/RWL1_junc RWL_30 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10750 x374/junc0 x374/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10751 VDD x375/junc0 x375/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10752 GND x445/junc1 x445/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10753 x76/junc0 x76/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10754 x860/RWL1_junc RWL_15 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10755 x811/junc1 WWL_1 WBLb_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10756 x700/RWL0_junc x700/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10757 x814/junc1 WWL_17 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10758 RBL0_31 RWL_10 x968/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10759 VDD x590/junc0 x590/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10760 RBL0_22 RWL_18 x6/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10761 x1002/RWL1_junc RWL_5 RBL1_29 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10762 RBL0_25 RWL_30 x653/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10763 x667/junc0 x667/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10764 x820/junc1 WWL_27 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10765 VDD x392/junc0 x392/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10766 x117/junc0 x117/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10767 WBL_7 WWL_5 x927/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10768 x622/RWL0_junc x622/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10769 VDD x400/junc0 x400/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10770 WBL_11 WWL_1 x309/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10771 x441/RWL0_junc x441/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10772 x516/RWL1_junc RWL_30 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10773 x674/junc0 x674/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10774 x145/RWL1_junc RWL_29 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10775 GND x705/junc0 x705/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10776 x753/RWL1_junc RWL_2 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10777 x405/junc0 x405/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10778 GND x462/junc1 x462/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10779 WBL_5 WWL_21 x318/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10780 GND x425/junc1 x425/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10781 VDD x863/junc0 x863/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10782 x18/RWL0_junc x18/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10783 x21/RWL0_junc x21/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10784 x715/RWL0_junc x715/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10785 GND x818/junc0 x818/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10786 RBL0_2 RWL_29 x467/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10787 x411/junc0 x411/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10788 x658/junc1 WWL_7 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10789 WBL_29 WWL_11 x326/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10790 RBL0_13 RWL_15 x912/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10791 VDD x867/junc0 x867/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10792 x610/junc1 WWL_12 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10793 x962/RWL0_junc x962/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10794 GND x1/junc1 x1/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10795 GND x594/junc0 x594/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10796 x1012/junc1 WWL_8 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10797 GND x467/junc1 x467/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10798 x37/RWL0_junc x37/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10799 x677/junc0 x677/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10800 GND x839/junc0 x839/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10801 GND x229/junc0 x229/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10802 x255/junc1 WWL_2 WBLb_26 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10803 WBL_23 WWL_17 x333/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10804 x126/junc0 x126/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10805 VDD x419/junc0 x419/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10806 GND x10/junc1 x10/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10807 RBL0_7 RWL_21 x343/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10808 x128/junc0 x128/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10809 GND x268/junc1 x268/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10810 x422/junc0 x422/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10811 x872/RWL1_junc RWL_16 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10812 GND x227/junc0 x227/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10813 x47/RWL0_junc x47/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10814 x957/RWL1_junc RWL_24 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10815 x638/RWL0_junc x638/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10816 RBL0_31 RWL_11 x972/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10817 VDD x621/junc0 x621/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10818 VDD x868/junc0 x868/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10819 x826/junc1 WWL_18 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10820 RBL0_22 RWL_19 x247/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10821 x739/junc0 x739/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10822 x996/RWL0_junc x996/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10823 x143/junc0 x143/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10824 RBL0_25 RWL_17 x696/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10825 x56/junc0 x56/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10826 WBL_5 WWL_28 x243/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10827 x439/junc0 x439/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10828 x440/junc0 x440/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10829 GND x726/junc0 x726/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10830 x771/RWL1_junc RWL_3 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10831 WBL_14 WWL_14 x359/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10832 x266/RWL0_junc x266/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10833 GND x202/junc1 x202/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10834 VDD x444/junc0 x444/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10835 x698/junc0 x698/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10836 x77/RWL0_junc x77/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10837 GND x849/junc0 x849/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10838 x79/RWL0_junc x79/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10839 GND x827/junc0 x827/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10840 x631/junc1 WWL_5 WBLb_11 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10841 x678/junc1 WWL_8 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10842 x464/junc1 WWL_9 WBLb_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10843 VDD x451/junc0 x451/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10844 RBL0_13 RWL_16 x921/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10845 GND x502/junc1 x502/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10846 x292/junc1 WWL_13 WBLb_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10847 GND x51/junc1 x51/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10848 x572/junc1 WWL_25 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10849 x4/junc0 x4/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10850 x12/junc0 x12/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10851 WBL_19 WWL_22 x655/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10852 GND x851/junc0 x851/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10853 x87/junc0 x87/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10854 WBL_28 WWL_30 x263/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10855 x832/junc1 WWL_21 WBLb_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10856 GND x282/junc0 x282/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10857 WBL_23 WWL_18 x374/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10858 RBL0_16 RWL_14 x974/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10859 GND x64/junc1 x64/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10860 RBL0_7 RWL_22 x393/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10861 x173/junc0 x173/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10862 GND x217/junc1 x217/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10863 x459/junc0 x459/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10864 x61/junc0 x61/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10865 x92/RWL0_junc x92/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10866 VDD x640/junc0 x640/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10867 x689/junc1 WWL_28 WBLb_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10868 GND x278/junc0 x278/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10869 x101/RWL0_junc x101/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10870 x894/RWL1_junc RWL_25 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10871 x788/RWL1_junc RWL_21 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10872 GND x642/junc0 x642/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10873 x370/RWL0_junc x370/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10874 VDD x460/junc0 x460/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10875 x104/RWL0_junc x104/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10876 x661/RWL0_junc x661/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10877 RBL0_31 RWL_12 x749/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10878 VDD x28/junc0 x28/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10879 VDD x461/junc0 x461/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10880 GND x72/junc1 x72/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10881 x836/junc1 WWL_17 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10882 x196/junc0 x196/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10883 RBL0_25 RWL_18 x718/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10884 x794/RWL1_junc RWL_0 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10885 x111/junc0 x111/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10886 x470/junc0 x470/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10887 WBL_10 WWL_19 x674/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10888 x346/RWL0_junc x346/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10889 x48/junc0 x48/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10890 x474/junc0 x474/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10891 WBL_4 WWL_25 x942/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10892 GND x859/junc0 x859/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10893 x891/RWL1_junc RWL_2 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10894 GND x306/junc0 x306/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10895 VDD x477/junc0 x477/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10896 GND x110/junc1 x110/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10897 x1009/RWL1_junc RWL_4 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10898 x605/junc1 WWL_26 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10899 WBL_28 WWL_15 x944/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10900 WBL_19 WWL_23 x677/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10901 RBL0_3 RWL_27 x150/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10902 WBL_28 WWL_31 x542/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10903 x139/junc0 x139/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10904 RBL0_16 RWL_15 x763/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10905 VDD x487/junc0 x487/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10906 RBL0_7 RWL_23 x436/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10907 x216/junc0 x216/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10908 GND x94/junc0 x94/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10909 x144/RWL0_junc x144/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10910 WBL_3 WWL_0 x422/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10911 VDD x492/junc0 x492/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10912 x684/junc0 x684/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10913 GND x546/junc1 x546/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10914 x803/RWL1_junc RWL_22 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10915 GND x328/junc0 x328/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10916 x414/RWL0_junc x414/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10917 x541/RWL1_junc RWL_26 RBL1_9 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10918 x153/RWL0_junc x153/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10919 x225/junc0 x225/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10920 VDD x493/junc0 x493/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10921 x494/junc0 x494/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10922 GND x284/junc1 x284/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10923 x232/RWL0_junc x232/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10924 VDD x893/junc0 x893/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10925 x672/junc1 WWL_22 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10926 VDD x498/junc0 x498/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10927 x760/RWL0_junc x760/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10928 x735/junc0 x735/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10929 x846/junc1 WWL_18 WBLb_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10930 x240/junc0 x240/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10931 RBL0_25 RWL_19 x979/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10932 x807/RWL1_junc RWL_1 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10933 x736/junc0 x736/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10934 RBL0_5 RWL_0 x337/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10935 WBL_10 WWL_20 x439/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10936 x549/junc0 x549/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10937 x505/junc0 x505/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10938 GND x666/junc0 x666/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10939 x1011/RWL1_junc RWL_7 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10940 x382/junc1 WWL_30 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10941 x508/junc0 x508/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10942 VDD x782/junc0 x782/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10943 GND x567/junc1 x567/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10944 VDD x509/junc0 x509/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10945 WBL_4 WWL_26 x698/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10946 GND x345/junc0 x345/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10947 x902/RWL1_junc x61/RWL1 RBL1_10 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10948 x788/RWL0_junc x788/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10949 x183/RWL0_junc x183/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10950 GND x463/junc0 x463/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10951 GND x29/junc0 x29/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10952 VDD x681/junc0 x681/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10953 x943/RWL1_junc RWL_5 RBL1_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10954 RBL0_27 RWL_6 x356/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10955 VDD x512/junc0 x512/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10956 GND x41/junc1 x41/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10957 x627/junc1 WWL_19 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10958 WBL_28 WWL_16 x4/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10959 x727/junc1 WWL_27 WBLb_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10960 RBL0_12 RWL_20 x461/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10961 WBL_19 WWL_24 x12/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10962 x288/junc0 x288/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10963 RBL0_16 RWL_16 x787/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10964 VDD x149/junc0 x149/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10965 GND x443/junc0 x443/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10966 GND x687/junc0 x687/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10967 WBL_3 WWL_1 x459/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10968 x599/junc0 x599/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10969 GND x877/junc0 x877/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10970 VDD x521/junc0 x521/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10971 x899/junc1 WWL_25 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10972 x191/junc0 x191/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10973 GND x310/junc1 x310/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10974 x522/junc0 x522/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10975 x523/junc0 x523/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10976 x823/RWL1_junc RWL_23 RBL1_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10977 GND x369/junc0 x369/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10978 x275/junc0 x275/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10979 x526/junc0 x526/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10980 x285/RWL0_junc x285/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10981 VDD x529/junc0 x529/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10982 x691/junc1 WWL_23 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10983 VDD x530/junc0 x530/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10984 VDD x532/junc0 x532/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10985 x741/junc1 WWL_28 WBLb_25 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10986 x857/junc1 WWL_0 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10987 RBL0_5 RWL_1 x379/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10988 x914/RWL1_junc RWL_27 RBL1_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10989 x209/junc0 x209/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10990 x784/RWL0_junc x784/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10991 x537/junc0 x537/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10992 x540/junc0 x540/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M10993 x136/RWL1_junc RWL_31 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10994 GND x389/junc0 x389/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10995 GND x596/junc1 x596/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10996 x909/RWL1_junc RWL_0 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10997 x1012/RWL1_junc RWL_8 RBL1_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10998 RBL0_12 RWL_9 x483/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M10999 x425/junc1 WWL_31 WBLb_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11000 WBL_13 WWL_19 x48/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11001 GND x335/junc1 x335/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11002 WBL_4 WWL_27 x474/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11003 x219/RWL0_junc x219/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11004 x803/RWL0_junc x803/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11005 x548/junc0 x548/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11006 GND x693/junc0 x693/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11007 GND x85/junc0 x85/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11008 GND x86/junc0 x86/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11009 VDD x550/junc0 x550/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11010 VDD x551/junc0 x551/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11011 x866/junc1 WWL_20 WBLb_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11012 VDD x925/junc0 x925/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11013 GND x96/junc1 x96/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11014 x801/junc0 x801/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11015 RBL0_17 RWL_17 x498/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11016 GND x481/junc1 x481/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11017 GND x708/junc0 x708/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11018 x432/RWL1_junc RWL_4 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11019 x994/junc0 x994/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11020 x759/junc0 x759/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11021 x270/junc0 x270/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11022 x908/junc1 WWL_26 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11023 VDD x558/junc0 x558/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11024 x238/junc0 x238/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11025 RBL0_6 RWL_27 x983/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11026 GND x351/junc1 x351/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11027 x241/junc0 x241/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11028 RBL0_21 RWL_13 x910/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11029 x559/junc0 x559/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11030 WBL_15 WWL_6 x684/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11031 x560/junc0 x560/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11032 x312/junc0 x312/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11033 GND x149/junc0 x149/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11034 VDD x712/junc0 x712/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11035 WBL_6 WWL_0 x494/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11036 VDD x562/junc0 x562/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11037 x740/junc1 WWL_24 WBLb_23 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11038 x323/RWL0_junc x323/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11039 VDD x566/junc0 x566/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11040 GND x865/junc0 x865/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11041 x571/junc0 x571/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11042 WBL_17 WWL_2 x735/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11043 GND x421/junc0 x421/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11044 GND x620/junc1 x620/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11045 x7/junc1 WWL_1 WBLb_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11046 GND x233/junc1 x233/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11047 x259/RWL0_junc x259/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11048 GND x799/junc0 x799/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11049 x765/junc0 x765/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11050 x802/RWL0_junc x802/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11051 x555/junc0 x555/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11052 GND x625/junc1 x625/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11053 WBL_24 WWL_10 x505/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11054 RBL0_8 RWL_14 x273/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11055 GND x626/junc1 x626/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11056 x915/RWL1_junc RWL_1 RBL1_15 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11057 WBL_13 WWL_20 x508/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11058 x618/junc0 x618/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11059 x267/RWL0_junc x267/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11060 x823/RWL0_junc x823/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11061 x580/junc0 x580/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11062 x456/RWL1_junc RWL_31 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11063 x709/RWL1_junc RWL_30 RBL1_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11064 x581/junc0 x581/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11065 x1017/junc1 WWL_5 WBLb_20 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11066 GND x714/junc0 x714/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11067 GND x722/junc0 x722/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11068 GND x724/junc0 x724/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11069 x63/RWL1_junc RWL_13 RBL1_14 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11070 x338/junc0 x338/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11071 VDD x584/junc0 x584/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11072 GND x146/junc1 x146/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11073 x283/RWL0_junc x283/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11074 RBL0_26 RWL_10 x986/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11075 x879/junc1 WWL_17 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11076 VDD x730/junc0 x730/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11077 x302/junc0 x302/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11078 RBL0_4 RWL_30 x402/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11079 RBL0_17 RWL_18 x532/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11080 x976/RWL1_junc RWL_5 RBL1_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11081 x569/junc1 WWL_19 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11082 x780/junc0 x780/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11083 RBL0_30 RWL_6 x987/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11084 x882/junc1 WWL_27 WBLb_8 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11085 x997/junc0 x997/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11086 x781/junc0 x781/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11087 WBL_15 WWL_7 x523/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11088 WBL_0 WWL_0 x522/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11089 x372/junc0 x372/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11090 WBL_2 WWL_5 x963/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11091 x931/RWL1_junc RWL_21 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11092 x836/RWL1_junc RWL_17 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11093 VDD x918/junc0 x918/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11094 VDD x595/junc0 x595/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11095 WBL_6 WWL_1 x526/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11096 VDD x842/junc0 x842/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11097 x785/junc0 x785/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11098 GND x876/junc0 x876/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11099 x838/RWL1_junc RWL_2 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11100 x603/junc0 x603/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11101 GND x645/junc1 x645/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11102 x689/RWL1_junc RWL_28 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11103 x789/junc0 x789/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11104 x864/RWL1_junc RWL_28 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11105 x299/RWL0_junc x299/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11106 GND x811/junc0 x811/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11107 x817/RWL0_junc x817/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11108 WBL_20 WWL_15 x111/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11109 WBL_24 WWL_11 x540/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11110 RBL0_8 RWL_15 x952/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11111 GND x650/junc1 x650/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11112 x1018/RWL0_junc x1018/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11113 GND x732/junc0 x732/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11114 RBL0_8 RWL_28 x752/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11115 x91/junc0 x91/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11116 x307/RWL0_junc x307/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11117 GND x903/junc0 x903/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11118 VDD x999/junc0 x999/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11119 x614/junc0 x614/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11120 WBL_11 WWL_28 x973/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11121 x479/junc1 WWL_2 WBLb_21 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11122 GND x1008/junc1 x1008/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11123 RBL0_2 RWL_21 x558/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11124 WBL_18 WWL_17 x548/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11125 GND x468/junc0 x468/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11126 GND x294/junc1 x294/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11127 x875/junc1 WWL_29 WBLb_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11128 x380/junc0 x380/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11129 x322/RWL0_junc x322/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11130 x889/junc1 WWL_10 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11131 x982/RWL1_junc RWL_24 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11132 x316/junc0 x316/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11133 x390/junc0 x390/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11134 RBL0_26 RWL_11 x991/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11135 VDD x746/junc0 x746/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11136 VDD x926/junc0 x926/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11137 x890/junc1 WWL_18 WBLb_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11138 RBL0_17 RWL_19 x569/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11139 x95/junc1 WWL_20 WBLb_17 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11140 x416/junc0 x416/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11141 WBL_15 WWL_8 x560/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11142 WBL_0 WWL_1 x559/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11143 GND x887/junc0 x887/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11144 x828/junc0 x828/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11145 x939/RWL1_junc RWL_14 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11146 RBL0_31 RWL_30 x924/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11147 x846/RWL1_junc RWL_18 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11148 x655/RWL1_junc RWL_22 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11149 VDD x829/junc0 x829/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11150 GND x210/junc1 x210/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11151 x9/junc0 x9/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11152 x11/junc0 x11/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11153 GND x888/junc0 x888/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11154 GND x484/junc0 x484/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11155 x848/RWL1_junc RWL_3 RBL1_2 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11156 GND x744/junc0 x744/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11157 GND x668/junc1 x668/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11158 WBL_9 WWL_14 x571/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11159 x937/RWL0_junc x937/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11160 GND x449/junc1 x449/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11161 GND x770/junc0 x770/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11162 VDD x629/junc0 x629/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11163 x446/RWL1_junc RWL_29 RBL1_12 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11164 GND x203/junc1 x203/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11165 x875/RWL1_junc RWL_29 RBL1_18 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11166 x339/RWL0_junc x339/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11167 GND x793/junc0 x793/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11168 WBL_20 WWL_16 x736/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11169 x751/junc1 WWL_5 WBLb_6 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11170 RBL0_8 RWL_16 x959/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11171 RBL0_8 RWL_29 x764/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11172 x35/junc0 x35/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11173 GND x575/junc1 x575/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11174 x142/junc0 x142/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11175 GND x911/junc0 x911/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11176 WBL_7 WWL_30 x487/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11177 x347/junc0 x347/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11178 x896/junc1 WWL_21 WBLb_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11179 WBL_18 WWL_18 x581/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11180 RBL0_11 RWL_14 x995/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11181 GND x332/junc1 x332/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11182 RBL0_2 RWL_22 x592/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11183 x424/junc0 x424/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11184 VDD x756/junc0 x756/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11185 x720/junc1 WWL_15 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11186 x364/RWL0_junc x364/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11187 x941/RWL1_junc RWL_17 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11188 x942/RWL1_junc RWL_25 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11189 x360/junc0 x360/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11190 x898/junc1 WWL_11 WBLb_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11191 VDD x703/junc0 x703/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11192 x433/junc0 x433/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11193 RBL0_26 RWL_12 x835/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11194 VDD x303/junc0 x303/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11195 VDD x36/junc0 x36/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11196 GND x754/junc0 x754/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11197 x649/junc0 x649/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11198 x855/RWL1_junc RWL_19 RBL1_27 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11199 x944/RWL1_junc RWL_15 RBL1_28 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11200 x815/junc0 x815/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11201 x368/junc0 x368/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11202 x677/RWL1_junc RWL_23 RBL1_19 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11203 x154/junc1 WWL_17 WBLb_22 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11204 x857/RWL1_junc RWL_0 RBL1_7 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11205 x63/junc0 x63/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11206 GND x514/junc0 x514/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11207 WBL_5 WWL_19 x785/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11208 x377/RWL0_junc x377/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11209 GND x545/junc1 x545/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11210 GND x174/junc1 x174/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11211 WBL_17 WWL_28 x509/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11212 GND x250/junc1 x250/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11213 x323/junc0 x323/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11214 x731/junc1 WWL_5 WBLb_0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11215 WBL_29 WWL_9 x789/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11216 GND x600/junc1 x600/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11217 GND x598/junc1 x598/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11218 x940/RWL1_junc RWL_2 RBL1_5 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11219 GND x806/junc0 x806/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11220 x565/RWL0_junc x565/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11221 x391/RWL0_junc x391/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11222 GND x695/junc1 x695/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11223 WBL_23 WWL_15 x245/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11224 x457/junc0 x457/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11225 WBL_7 WWL_31 x149/junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11226 x904/junc1 WWL_14 WBLb_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11227 x398/junc0 x398/junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11228 RBL0_11 RWL_15 x843/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11229 RBL0_2 RWL_23 x624/RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11230 GND x280/junc0 x280/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11231 x403/RWL0_junc x403/junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11232 x662/junc0 x662/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11233 x94/junc0 x94/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11234 VDD x664/junc0 x664/junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11235 GND x700/junc1 x700/RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11236 x743/junc1 WWL_16 WBLb_24 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11237 x102/junc0 x102/junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15

M11238 x946/RWL1_junc RWL_18 RBL1_13 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11239 x698/RWL1_junc RWL_26 RBL1_4 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

M11240 GND x773/junc0 x773/junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15

.ends

** hspice subcircuit dictionary
* x0	10T_1x8_magic_70/10T_toy_magic_2
* x1	10T_1x8_magic_29/10T_toy_magic_4
* x2	10T_1x8_magic_82/10T_toy_magic_5
* x3	10T_1x8_magic_16/10T_toy_magic_7
* x4	10T_1x8_magic_95/10T_toy_magic_3
* x5	10T_1x8_magic_10/10T_toy_magic_1
* x6	10T_1x8_magic_91/10T_toy_magic_0
* x7	10T_1x8_magic_3/10T_toy_magic_1
* x8	10T_1x8_magic_61/10T_toy_magic_2
* x9	10T_1x8_magic_51/10T_toy_magic_0
* x10	10T_1x8_magic_113/10T_toy_magic_4
* x11	10T_1x8_magic_28/10T_toy_magic_2
* x12	10T_1x8_magic_77/10T_toy_magic_4
* x13	10T_1x8_magic_34/10T_toy_magic_2
* x14	10T_1x8_magic_121/10T_toy_magic_1
* x15	10T_1x8_magic_105/10T_toy_magic_4
* x16	10T_1x8_magic_122/10T_toy_magic_4
* x17	10T_1x8_magic_43/10T_toy_magic_7
* x18	10T_1x8_magic_91/10T_toy_magic_7
* x19	10T_1x8_magic_0/10T_toy_magic_3
* x20	10T_1x8_magic_122/10T_toy_magic_5
* x21	10T_1x8_magic_12/10T_toy_magic_6
* x22	10T_1x8_magic_51/10T_toy_magic_7
* x23	10T_1x8_magic_1/10T_toy_magic_2
* x24	10T_1x8_magic_32/10T_toy_magic_3
* x25	10T_1x8_magic_68/10T_toy_magic_7
* x26	10T_1x8_magic_109/10T_toy_magic_6
* x27	10T_1x8_magic_26/10T_toy_magic_7
* x28	10T_1x8_magic_38/10T_toy_magic_4
* x29	10T_1x8_magic_29/10T_toy_magic_6
* x30	10T_1x8_magic_57/10T_toy_magic_3
* x31	10T_1x8_magic_53/10T_toy_magic_4
* x32	10T_1x8_magic_44/10T_toy_magic_6
* x33	10T_1x8_magic_114/10T_toy_magic_0
* x34	10T_1x8_magic_38/10T_toy_magic_5
* x35	10T_1x8_magic_94/10T_toy_magic_1
* x36	10T_1x8_magic_28/10T_toy_magic_1
* x37	10T_1x8_magic_95/10T_toy_magic_1
* x38	10T_1x8_magic_124/10T_toy_magic_7
* x39	10T_1x8_magic_47/10T_toy_magic_4
* x40	10T_1x8_magic_83/10T_toy_magic_5
* x41	10T_1x8_magic_38/10T_toy_magic_1
* x42	10T_1x8_magic_42/10T_toy_magic_5
* x43	10T_1x8_magic_29/10T_toy_magic_7
* x44	10T_1x8_magic_111/10T_toy_magic_5
* x45	10T_1x8_magic_21/10T_toy_magic_4
* x46	10T_1x8_magic_56/10T_toy_magic_5
* x47	10T_1x8_magic_83/10T_toy_magic_6
* x48	10T_1x8_magic_44/10T_toy_magic_2
* x49	10T_1x8_magic_53/10T_toy_magic_3
* x50	10T_1x8_magic_24/10T_toy_magic_6
* x51	10T_1x8_magic_30/10T_toy_magic_4
* x52	10T_1x8_magic_97/10T_toy_magic_4
* x53	10T_1x8_magic_20/10T_toy_magic_4
* x54	10T_1x8_magic_68/10T_toy_magic_2
* x55	10T_1x8_magic_80/10T_toy_magic_5
* x56	10T_1x8_magic_98/10T_toy_magic_3
* x57	10T_1x8_magic_114/10T_toy_magic_7
* x58	10T_1x8_magic_20/10T_toy_magic_3
* x59	10T_1x8_magic_70/10T_toy_magic_0
* x60	10T_1x8_magic_2/10T_toy_magic_5
* x61	10T_1x8_magic_120/10T_toy_magic_7
* x62	10T_1x8_magic_60/10T_toy_magic_2
* x63	10T_1x8_magic_50/10T_toy_magic_0
* x64	10T_1x8_magic_111/10T_toy_magic_4
* x65	10T_1x8_magic_72/10T_toy_magic_5
* x66	10T_1x8_magic_92/10T_toy_magic_3
* x67	10T_1x8_magic_32/10T_toy_magic_6
* x68	10T_1x8_magic_76/10T_toy_magic_4
* x69	10T_1x8_magic_121/10T_toy_magic_3
* x70	10T_1x8_magic_104/10T_toy_magic_4
* x71	10T_1x8_magic_69/10T_toy_magic_1
* x72	10T_1x8_magic_33/10T_toy_magic_4
* x73	10T_1x8_magic_63/10T_toy_magic_5
* x74	10T_1x8_magic_120/10T_toy_magic_4
* x75	10T_1x8_magic_0/10T_toy_magic_4
* x76	10T_1x8_magic_15/10T_toy_magic_1
* x77	10T_1x8_magic_88/10T_toy_magic_7
* x78	10T_1x8_magic_120/10T_toy_magic_5
* x79	10T_1x8_magic_11/10T_toy_magic_6
* x80	10T_1x8_magic_98/10T_toy_magic_2
* x81	10T_1x8_magic_23/10T_toy_magic_7
* x82	10T_1x8_magic_40/10T_toy_magic_4
* x83	10T_1x8_magic_42/10T_toy_magic_3
* x84	10T_1x8_magic_66/10T_toy_magic_4
* x85	10T_1x8_magic_76/10T_toy_magic_7
* x86	10T_1x8_magic_30/10T_toy_magic_6
* x87	10T_1x8_magic_56/10T_toy_magic_3
* x88	10T_1x8_magic_52/10T_toy_magic_4
* x89	10T_1x8_magic_43/10T_toy_magic_6
* x90	10T_1x8_magic_40/10T_toy_magic_5
* x91	10T_1x8_magic_79/10T_toy_magic_4
* x92	10T_1x8_magic_72/10T_toy_magic_2
* x93	10T_1x8_magic_81/10T_toy_magic_5
* x94	10T_1x8_magic_85/10T_toy_magic_1
* x95	10T_1x8_magic_86/10T_toy_magic_6
* x96	10T_1x8_magic_40/10T_toy_magic_1
* x97	10T_1x8_magic_41/10T_toy_magic_5
* x98	10T_1x8_magic_122/10T_toy_magic_3
* x99	10T_1x8_magic_22/10T_toy_magic_4
* x100	10T_1x8_magic_30/10T_toy_magic_7
* x101	10T_1x8_magic_81/10T_toy_magic_6
* x102	10T_1x8_magic_57/10T_toy_magic_5
* x103	10T_1x8_magic_55/10T_toy_magic_5
* x104	10T_1x8_magic_6/10T_toy_magic_2
* x105	10T_1x8_magic_70/10T_toy_magic_4
* x106	10T_1x8_magic_52/10T_toy_magic_3
* x107	10T_1x8_magic_21/10T_toy_magic_6
* x108	10T_1x8_magic_95/10T_toy_magic_4
* x109	10T_1x8_magic_77/10T_toy_magic_5
* x110	10T_1x8_magic_27/10T_toy_magic_4
* x111	10T_1x8_magic_96/10T_toy_magic_3
* x112	10T_1x8_magic_57/10T_toy_magic_2
* x113	10T_1x8_magic_8/10T_toy_magic_3
* x114	10T_1x8_magic_5/10T_toy_magic_3
* x115	10T_1x8_magic_68/10T_toy_magic_0
* x116	10T_1x8_magic_3/10T_toy_magic_5
* x117	10T_1x8_magic_71/10T_toy_magic_0
* x118	10T_1x8_magic_5/10T_toy_magic_4
* x119	10T_1x8_magic_93/10T_toy_magic_3
* x120	10T_1x8_magic_29/10T_toy_magic_0
* x121	10T_1x8_magic_127/10T_toy_magic_7
* x122	10T_1x8_magic_33/10T_toy_magic_6
* x123	10T_1x8_magic_74/10T_toy_magic_4
* x124	10T_1x8_magic_119/10T_toy_magic_3
* x125	10T_1x8_magic_126/10T_toy_magic_1
* x126	10T_1x8_magic_8/10T_toy_magic_4
* x127	10T_1x8_magic_62/10T_toy_magic_5
* x128	10T_1x8_magic_122/10T_toy_magic_7
* x129	10T_1x8_magic_1/10T_toy_magic_4
* x130	10T_1x8_magic_113/10T_toy_magic_0
* x131	10T_1x8_magic_96/10T_toy_magic_2
* x132	10T_1x8_magic_119/10T_toy_magic_4
* x133	10T_1x8_magic_122/10T_toy_magic_0
* x134	10T_1x8_magic_108/10T_toy_magic_6
* x135	10T_1x8_magic_41/10T_toy_magic_3
* x136	10T_1x8_magic_67/10T_toy_magic_4
* x137	10T_1x8_magic_36/10T_toy_magic_4
* x138	10T_1x8_magic_50/10T_toy_magic_6
* x139	10T_1x8_magic_55/10T_toy_magic_3
* x140	10T_1x8_magic_36/10T_toy_magic_5
* x141	10T_1x8_magic_87/10T_toy_magic_1
* x142	10T_1x8_magic_75/10T_toy_magic_4
* x143	10T_1x8_magic_105/10T_toy_magic_2
* x144	10T_1x8_magic_87/10T_toy_magic_0
* x145	10T_1x8_magic_17/10T_toy_magic_0
* x146	10T_1x8_magic_36/10T_toy_magic_1
* x147	10T_1x8_magic_120/10T_toy_magic_3
* x148	10T_1x8_magic_115/10T_toy_magic_6
* x149	10T_1x8_magic_16/10T_toy_magic_1
* x150	10T_1x8_magic_19/10T_toy_magic_4
* x151	10T_1x8_magic_39/10T_toy_magic_5
* x152	10T_1x8_magic_27/10T_toy_magic_7
* x153	10T_1x8_magic_7/10T_toy_magic_2
* x154	10T_1x8_magic_90/10T_toy_magic_0
* x155	10T_1x8_magic_103/10T_toy_magic_6
* x156	10T_1x8_magic_34/10T_toy_magic_0
* x157	10T_1x8_magic_94/10T_toy_magic_6
* x158	10T_1x8_magic_22/10T_toy_magic_6
* x159	10T_1x8_magic_51/10T_toy_magic_3
* x160	10T_1x8_magic_42/10T_toy_magic_2
* x161	10T_1x8_magic_56/10T_toy_magic_2
* x162	10T_1x8_magic_9/10T_toy_magic_3
* x163	10T_1x8_magic_79/10T_toy_magic_1
* x164	10T_1x8_magic_66/10T_toy_magic_5
* x165	10T_1x8_magic_109/10T_toy_magic_7
* x166	10T_1x8_magic_89/10T_toy_magic_3
* x167	10T_1x8_magic_30/10T_toy_magic_0
* x168	10T_1x8_magic_125/10T_toy_magic_7
* x169	10T_1x8_magic_118/10T_toy_magic_3
* x170	10T_1x8_magic_57/10T_toy_magic_0
* x171	10T_1x8_magic_8/10T_toy_magic_2
* x172	10T_1x8_magic_124/10T_toy_magic_1
* x173	10T_1x8_magic_9/10T_toy_magic_4
* x174	10T_1x8_magic_32/10T_toy_magic_4
* x175	10T_1x8_magic_111/10T_toy_magic_0
* x176	10T_1x8_magic_109/10T_toy_magic_1
* x177	10T_1x8_magic_94/10T_toy_magic_2
* x178	10T_1x8_magic_112/10T_toy_magic_5
* x179	10T_1x8_magic_53/10T_toy_magic_0
* x180	10T_1x8_magic_0/10T_toy_magic_6
* x181	10T_1x8_magic_118/10T_toy_magic_4
* x182	10T_1x8_magic_108/10T_toy_magic_7
* x183	10T_1x8_magic_109/10T_toy_magic_0
* x184	10T_1x8_magic_19/10T_toy_magic_1
* x185	10T_1x8_magic_39/10T_toy_magic_3
* x186	10T_1x8_magic_120/10T_toy_magic_0
* x187	10T_1x8_magic_0/10T_toy_magic_0
* x188	10T_1x8_magic_32/10T_toy_magic_0
* x189	10T_1x8_magic_105/10T_toy_magic_1
* x190	10T_1x8_magic_43/10T_toy_magic_1
* x191	10T_1x8_magic_8/10T_toy_magic_7
* x192	10T_1x8_magic_127/10T_toy_magic_6
* x193	10T_1x8_magic_116/10T_toy_magic_6
* x194	10T_1x8_magic_73/10T_toy_magic_4
* x195	10T_1x8_magic_27/10T_toy_magic_5
* x196	10T_1x8_magic_104/10T_toy_magic_2
* x197	10T_1x8_magic_73/10T_toy_magic_6
* x198	10T_1x8_magic_98/10T_toy_magic_1
* x199	10T_1x8_magic_32/10T_toy_magic_5
* x200	10T_1x8_magic_35/10T_toy_magic_0
* x201	10T_1x8_magic_101/10T_toy_magic_6
* x202	10T_1x8_magic_51/10T_toy_magic_6
* x203	10T_1x8_magic_34/10T_toy_magic_1
* x204	10T_1x8_magic_41/10T_toy_magic_2
* x205	10T_1x8_magic_59/10T_toy_magic_6
* x206	10T_1x8_magic_55/10T_toy_magic_2
* x207	10T_1x8_magic_59/10T_toy_magic_7
* x208	10T_1x8_magic_75/10T_toy_magic_1
* x209	10T_1x8_magic_79/10T_toy_magic_7
* x210	10T_1x8_magic_73/10T_toy_magic_2
* x211	10T_1x8_magic_67/10T_toy_magic_5
* x212	10T_1x8_magic_20/10T_toy_magic_6
* x213	10T_1x8_magic_27/10T_toy_magic_0
* x214	10T_1x8_magic_13/10T_toy_magic_4
* x215	10T_1x8_magic_56/10T_toy_magic_0
* x216	10T_1x8_magic_31/10T_toy_magic_4
* x217	10T_1x8_magic_94/10T_toy_magic_5
* x218	10T_1x8_magic_127/10T_toy_magic_4
* x219	10T_1x8_magic_99/10T_toy_magic_5
* x220	10T_1x8_magic_52/10T_toy_magic_0
* x221	10T_1x8_magic_0/10T_toy_magic_7
* x222	10T_1x8_magic_110/10T_toy_magic_5
* x223	10T_1x8_magic_54/10T_toy_magic_1
* x224	10T_1x8_magic_4/10T_toy_magic_5
* x225	10T_1x8_magic_8/10T_toy_magic_0
* x226	10T_1x8_magic_1/10T_toy_magic_0
* x227	10T_1x8_magic_70/10T_toy_magic_3
* x228	10T_1x8_magic_114/10T_toy_magic_2
* x229	10T_1x8_magic_96/10T_toy_magic_4
* x230	10T_1x8_magic_68/10T_toy_magic_1
* x231	10T_1x8_magic_65/10T_toy_magic_6
* x232	10T_1x8_magic_45/10T_toy_magic_7
* x233	10T_1x8_magic_57/10T_toy_magic_7
* x234	10T_1x8_magic_69/10T_toy_magic_7
* x235	10T_1x8_magic_125/10T_toy_magic_6
* x236	10T_1x8_magic_119/10T_toy_magic_0
* x237	10T_1x8_magic_104/10T_toy_magic_1
* x238	10T_1x8_magic_9/10T_toy_magic_7
* x239	10T_1x8_magic_117/10T_toy_magic_6
* x240	10T_1x8_magic_102/10T_toy_magic_2
* x241	10T_1x8_magic_28/10T_toy_magic_5
* x242	10T_1x8_magic_58/10T_toy_magic_1
* x243	10T_1x8_magic_20/10T_toy_magic_2
* x244	10T_1x8_magic_16/10T_toy_magic_4
* x245	10T_1x8_magic_96/10T_toy_magic_1
* x246	10T_1x8_magic_26/10T_toy_magic_6
* x247	10T_1x8_magic_88/10T_toy_magic_0
* x248	10T_1x8_magic_101/10T_toy_magic_7
* x249	10T_1x8_magic_37/10T_toy_magic_6
* x250	10T_1x8_magic_35/10T_toy_magic_1
* x251	10T_1x8_magic_64/10T_toy_magic_1
* x252	10T_1x8_magic_39/10T_toy_magic_2
* x253	10T_1x8_magic_58/10T_toy_magic_6
* x254	10T_1x8_magic_83/10T_toy_magic_2
* x255	10T_1x8_magic_123/10T_toy_magic_5
* x256	10T_1x8_magic_58/10T_toy_magic_7
* x257	10T_1x8_magic_73/10T_toy_magic_1
* x258	10T_1x8_magic_5/10T_toy_magic_6
* x259	10T_1x8_magic_45/10T_toy_magic_4
* x260	10T_1x8_magic_100/10T_toy_magic_7
* x261	10T_1x8_magic_12/10T_toy_magic_4
* x262	10T_1x8_magic_55/10T_toy_magic_0
* x263	10T_1x8_magic_66/10T_toy_magic_3
* x264	10T_1x8_magic_50/10T_toy_magic_1
* x265	10T_1x8_magic_71/10T_toy_magic_4
* x266	10T_1x8_magic_109/10T_toy_magic_4
* x267	10T_1x8_magic_97/10T_toy_magic_5
* x268	10T_1x8_magic_96/10T_toy_magic_5
* x269	10T_1x8_magic_125/10T_toy_magic_4
* x270	10T_1x8_magic_114/10T_toy_magic_6
* x271	10T_1x8_magic_63/10T_toy_magic_4
* x272	10T_1x8_magic_1/10T_toy_magic_7
* x273	10T_1x8_magic_49/10T_toy_magic_7
* x274	10T_1x8_magic_14/10T_toy_magic_5
* x275	10T_1x8_magic_9/10T_toy_magic_0
* x276	10T_1x8_magic_86/10T_toy_magic_3
* x277	10T_1x8_magic_84/10T_toy_magic_2
* x278	10T_1x8_magic_68/10T_toy_magic_3
* x279	10T_1x8_magic_79/10T_toy_magic_6
* x280	10T_1x8_magic_85/10T_toy_magic_5
* x281	10T_1x8_magic_112/10T_toy_magic_2
* x282	10T_1x8_magic_94/10T_toy_magic_4
* x283	10T_1x8_magic_84/10T_toy_magic_3
* x284	10T_1x8_magic_5/10T_toy_magic_2
* x285	10T_1x8_magic_46/10T_toy_magic_7
* x286	10T_1x8_magic_118/10T_toy_magic_0
* x287	10T_1x8_magic_17/10T_toy_magic_2
* x288	10T_1x8_magic_20/10T_toy_magic_7
* x289	10T_1x8_magic_107/10T_toy_magic_2
* x290	10T_1x8_magic_86/10T_toy_magic_4
* x291	10T_1x8_magic_23/10T_toy_magic_6
* x292	10T_1x8_magic_10/10T_toy_magic_5
* x293	10T_1x8_magic_61/10T_toy_magic_7
* x294	10T_1x8_magic_112/10T_toy_magic_0
* x295	10T_1x8_magic_81/10T_toy_magic_2
* x296	10T_1x8_magic_121/10T_toy_magic_5
* x297	10T_1x8_magic_65/10T_toy_magic_1
* x298	10T_1x8_magic_49/10T_toy_magic_3
* x299	10T_1x8_magic_46/10T_toy_magic_4
* x300	10T_1x8_magic_11/10T_toy_magic_4
* x301	10T_1x8_magic_108/10T_toy_magic_3
* x302	10T_1x8_magic_69/10T_toy_magic_4
* x303	10T_1x8_magic_24/10T_toy_magic_0
* x304	10T_1x8_magic_5/10T_toy_magic_1
* x305	10T_1x8_magic_13/10T_toy_magic_0
* x306	10T_1x8_magic_27/10T_toy_magic_3
* x307	10T_1x8_magic_95/10T_toy_magic_5
* x308	10T_1x8_magic_112/10T_toy_magic_6
* x309	10T_1x8_magic_62/10T_toy_magic_4
* x310	10T_1x8_magic_83/10T_toy_magic_0
* x311	10T_1x8_magic_74/10T_toy_magic_0
* x312	10T_1x8_magic_31/10T_toy_magic_0
* x313	10T_1x8_magic_99/10T_toy_magic_0
* x314	10T_1x8_magic_82/10T_toy_magic_2
* x315	10T_1x8_magic_108/10T_toy_magic_4
* x316	10T_1x8_magic_127/10T_toy_magic_0
* x317	10T_1x8_magic_109/10T_toy_magic_3
* x318	10T_1x8_magic_25/10T_toy_magic_2
* x319	10T_1x8_magic_99/10T_toy_magic_2
* x320	10T_1x8_magic_110/10T_toy_magic_2
* x321	10T_1x8_magic_4/10T_toy_magic_2
* x322	10T_1x8_magic_82/10T_toy_magic_3
* x323	10T_1x8_magic_44/10T_toy_magic_7
* x324	10T_1x8_magic_64/10T_toy_magic_4
* x325	10T_1x8_magic_13/10T_toy_magic_1
* x326	10T_1x8_magic_106/10T_toy_magic_2
* x327	10T_1x8_magic_36/10T_toy_magic_0
* x328	10T_1x8_magic_96/10T_toy_magic_0
* x329	10T_1x8_magic_57/10T_toy_magic_4
* x330	10T_1x8_magic_127/10T_toy_magic_1
* x331	10T_1x8_magic_60/10T_toy_magic_7
* x332	10T_1x8_magic_110/10T_toy_magic_0
* x333	10T_1x8_magic_90/10T_toy_magic_1
* x334	10T_1x8_magic_78/10T_toy_magic_2
* x335	10T_1x8_magic_120/10T_toy_magic_1
* x336	10T_1x8_magic_101/10T_toy_magic_4
* x337	10T_1x8_magic_2/10T_toy_magic_2
* x338	10T_1x8_magic_15/10T_toy_magic_5
* x339	10T_1x8_magic_44/10T_toy_magic_4
* x340	10T_1x8_magic_48/10T_toy_magic_3
* x341	10T_1x8_magic_45/10T_toy_magic_1
* x342	10T_1x8_magic_21/10T_toy_magic_0
* x343	10T_1x8_magic_25/10T_toy_magic_1
* x344	10T_1x8_magic_60/10T_toy_magic_1
* x345	10T_1x8_magic_51/10T_toy_magic_2
* x346	10T_1x8_magic_18/10T_toy_magic_0
* x347	10T_1x8_magic_4/10T_toy_magic_1
* x348	10T_1x8_magic_12/10T_toy_magic_0
* x349	10T_1x8_magic_28/10T_toy_magic_3
* x350	10T_1x8_magic_110/10T_toy_magic_6
* x351	10T_1x8_magic_81/10T_toy_magic_0
* x352	10T_1x8_magic_89/10T_toy_magic_1
* x353	10T_1x8_magic_72/10T_toy_magic_0
* x354	10T_1x8_magic_76/10T_toy_magic_0
* x355	10T_1x8_magic_123/10T_toy_magic_3
* x356	10T_1x8_magic_115/10T_toy_magic_4
* x357	10T_1x8_magic_97/10T_toy_magic_0
* x358	10T_1x8_magic_80/10T_toy_magic_2
* x359	10T_1x8_magic_49/10T_toy_magic_0
* x360	10T_1x8_magic_125/10T_toy_magic_0
* x361	10T_1x8_magic_26/10T_toy_magic_2
* x362	10T_1x8_magic_63/10T_toy_magic_0
* x363	10T_1x8_magic_97/10T_toy_magic_2
* x364	10T_1x8_magic_80/10T_toy_magic_3
* x365	10T_1x8_magic_14/10T_toy_magic_2
* x366	10T_1x8_magic_12/10T_toy_magic_1
* x367	10T_1x8_magic_103/10T_toy_magic_2
* x368	10T_1x8_magic_37/10T_toy_magic_0
* x369	10T_1x8_magic_94/10T_toy_magic_0
* x370	10T_1x8_magic_63/10T_toy_magic_2
* x371	10T_1x8_magic_116/10T_toy_magic_3
* x372	10T_1x8_magic_34/10T_toy_magic_6
* x373	10T_1x8_magic_125/10T_toy_magic_1
* x374	10T_1x8_magic_91/10T_toy_magic_1
* x375	10T_1x8_magic_126/10T_toy_magic_4
* x376	10T_1x8_magic_116/10T_toy_magic_1
* x377	10T_1x8_magic_123/10T_toy_magic_1
* x378	10T_1x8_magic_126/10T_toy_magic_5
* x379	10T_1x8_magic_3/10T_toy_magic_2
* x380	10T_1x8_magic_61/10T_toy_magic_4
* x381	10T_1x8_magic_37/10T_toy_magic_1
* x382	10T_1x8_magic_32/10T_toy_magic_1
* x383	10T_1x8_magic_47/10T_toy_magic_3
* x384	10T_1x8_magic_113/10T_toy_magic_6
* x385	10T_1x8_magic_65/10T_toy_magic_2
* x386	10T_1x8_magic_28/10T_toy_magic_7
* x387	10T_1x8_magic_16/10T_toy_magic_3
* x388	10T_1x8_magic_82/10T_toy_magic_7
* x389	10T_1x8_magic_121/10T_toy_magic_7
* x390	10T_1x8_magic_116/10T_toy_magic_0
* x391	10T_1x8_magic_25/10T_toy_magic_7
* x392	10T_1x8_magic_46/10T_toy_magic_1
* x393	10T_1x8_magic_26/10T_toy_magic_1
* x394	10T_1x8_magic_16/10T_toy_magic_0
* x395	10T_1x8_magic_22/10T_toy_magic_0
* x396	10T_1x8_magic_10/10T_toy_magic_3
* x397	10T_1x8_magic_59/10T_toy_magic_1
* x398	10T_1x8_magic_14/10T_toy_magic_1
* x399	10T_1x8_magic_50/10T_toy_magic_2
* x400	10T_1x8_magic_87/10T_toy_magic_5
* x401	10T_1x8_magic_78/10T_toy_magic_0
* x402	10T_1x8_magic_18/10T_toy_magic_3
* x403	10T_1x8_magic_87/10T_toy_magic_6
* x404	10T_1x8_magic_95/10T_toy_magic_0
* x405	10T_1x8_magic_48/10T_toy_magic_0
* x406	10T_1x8_magic_23/10T_toy_magic_2
* x407	10T_1x8_magic_95/10T_toy_magic_2
* x408	10T_1x8_magic_62/10T_toy_magic_0
* x409	10T_1x8_magic_102/10T_toy_magic_3
* x410	10T_1x8_magic_116/10T_toy_magic_7
* x411	10T_1x8_magic_42/10T_toy_magic_7
* x412	10T_1x8_magic_11/10T_toy_magic_1
* x413	10T_1x8_magic_56/10T_toy_magic_7
* x414	10T_1x8_magic_62/10T_toy_magic_2
* x415	10T_1x8_magic_79/10T_toy_magic_5
* x416	10T_1x8_magic_18/10T_toy_magic_2
* x417	10T_1x8_magic_15/10T_toy_magic_7
* x418	10T_1x8_magic_88/10T_toy_magic_1
* x419	10T_1x8_magic_124/10T_toy_magic_4
* x420	10T_1x8_magic_117/10T_toy_magic_1
* x421	10T_1x8_magic_57/10T_toy_magic_6
* x422	10T_1x8_magic_2/10T_toy_magic_4
* x423	10T_1x8_magic_124/10T_toy_magic_5
* x424	10T_1x8_magic_60/10T_toy_magic_4
* x425	10T_1x8_magic_33/10T_toy_magic_1
* x426	10T_1x8_magic_111/10T_toy_magic_6
* x427	10T_1x8_magic_109/10T_toy_magic_5
* x428	10T_1x8_magic_64/10T_toy_magic_2
* x429	10T_1x8_magic_53/10T_toy_magic_6
* x430	10T_1x8_magic_80/10T_toy_magic_7
* x431	10T_1x8_magic_31/10T_toy_magic_6
* x432	10T_1x8_magic_119/10T_toy_magic_7
* x433	10T_1x8_magic_117/10T_toy_magic_0
* x434	10T_1x8_magic_54/10T_toy_magic_4
* x435	10T_1x8_magic_19/10T_toy_magic_5
* x436	10T_1x8_magic_23/10T_toy_magic_1
* x437	10T_1x8_magic_44/10T_toy_magic_1
* x438	10T_1x8_magic_105/10T_toy_magic_5
* x439	10T_1x8_magic_43/10T_toy_magic_5
* x440	10T_1x8_magic_126/10T_toy_magic_3
* x441	10T_1x8_magic_17/10T_toy_magic_6
* x442	10T_1x8_magic_47/10T_toy_magic_0
* x443	10T_1x8_magic_67/10T_toy_magic_2
* x444	10T_1x8_magic_72/10T_toy_magic_3
* x445	10T_1x8_magic_98/10T_toy_magic_5
* x446	10T_1x8_magic_35/10T_toy_magic_3
* x447	10T_1x8_magic_100/10T_toy_magic_3
* x448	10T_1x8_magic_117/10T_toy_magic_7
* x449	10T_1x8_magic_11/10T_toy_magic_3
* x450	10T_1x8_magic_41/10T_toy_magic_7
* x451	10T_1x8_magic_6/10T_toy_magic_3
* x452	10T_1x8_magic_55/10T_toy_magic_7
* x453	10T_1x8_magic_6/10T_toy_magic_4
* x454	10T_1x8_magic_75/10T_toy_magic_5
* x455	10T_1x8_magic_73/10T_toy_magic_7
* x456	10T_1x8_magic_16/10T_toy_magic_2
* x457	10T_1x8_magic_126/10T_toy_magic_7
* x458	10T_1x8_magic_56/10T_toy_magic_6
* x459	10T_1x8_magic_3/10T_toy_magic_4
* x460	10T_1x8_magic_126/10T_toy_magic_0
* x461	10T_1x8_magic_43/10T_toy_magic_3
* x462	10T_1x8_magic_52/10T_toy_magic_6
* x463	10T_1x8_magic_77/10T_toy_magic_7
* x464	10T_1x8_magic_54/10T_toy_magic_5
* x465	10T_1x8_magic_9/10T_toy_magic_6
* x466	10T_1x8_magic_85/10T_toy_magic_3
* x467	10T_1x8_magic_17/10T_toy_magic_5
* x468	10T_1x8_magic_121/10T_toy_magic_4
* x469	10T_1x8_magic_104/10T_toy_magic_5
* x470	10T_1x8_magic_124/10T_toy_magic_3
* x471	10T_1x8_magic_119/10T_toy_magic_6
* x472	10T_1x8_magic_58/10T_toy_magic_5
* x473	10T_1x8_magic_100/10T_toy_magic_4
* x474	10T_1x8_magic_19/10T_toy_magic_3
* x475	10T_1x8_magic_34/10T_toy_magic_5
* x476	10T_1x8_magic_39/10T_toy_magic_7
* x477	10T_1x8_magic_7/10T_toy_magic_3
* x478	10T_1x8_magic_83/10T_toy_magic_7
* x479	10T_1x8_magic_122/10T_toy_magic_2
* x480	10T_1x8_magic_7/10T_toy_magic_4
* x481	10T_1x8_magic_73/10T_toy_magic_5
* x482	10T_1x8_magic_45/10T_toy_magic_3
* x483	10T_1x8_magic_54/10T_toy_magic_3
* x484	10T_1x8_magic_11/10T_toy_magic_2
* x485	10T_1x8_magic_20/10T_toy_magic_0
* x486	10T_1x8_magic_50/10T_toy_magic_4
* x487	10T_1x8_magic_18/10T_toy_magic_1
* x488	10T_1x8_magic_55/10T_toy_magic_6
* x489	10T_1x8_magic_38/10T_toy_magic_2
* x490	10T_1x8_magic_50/10T_toy_magic_5
* x491	10T_1x8_magic_35/10T_toy_magic_5
* x492	10T_1x8_magic_113/10T_toy_magic_1
* x493	10T_1x8_magic_124/10T_toy_magic_0
* x494	10T_1x8_magic_2/10T_toy_magic_0
* x495	10T_1x8_magic_5/10T_toy_magic_7
* x496	10T_1x8_magic_83/10T_toy_magic_3
* x497	10T_1x8_magic_38/10T_toy_magic_3
* x498	10T_1x8_magic_90/10T_toy_magic_6
* x499	10T_1x8_magic_11/10T_toy_magic_7
* x500	10T_1x8_magic_76/10T_toy_magic_3
* x501	10T_1x8_magic_120/10T_toy_magic_6
* x502	10T_1x8_magic_10/10T_toy_magic_6
* x503	10T_1x8_magic_118/10T_toy_magic_6
* x504	10T_1x8_magic_69/10T_toy_magic_2
* x505	10T_1x8_magic_107/10T_toy_magic_7
* x506	10T_1x8_magic_18/10T_toy_magic_6
* x507	10T_1x8_magic_115/10T_toy_magic_3
* x508	10T_1x8_magic_43/10T_toy_magic_2
* x509	10T_1x8_magic_70/10T_toy_magic_6
* x510	10T_1x8_magic_81/10T_toy_magic_7
* x511	10T_1x8_magic_120/10T_toy_magic_2
* x512	10T_1x8_magic_105/10T_toy_magic_7
* x513	10T_1x8_magic_46/10T_toy_magic_3
* x514	10T_1x8_magic_58/10T_toy_magic_0
* x515	10T_1x8_magic_69/10T_toy_magic_6
* x516	10T_1x8_magic_18/10T_toy_magic_5
* x517	10T_1x8_magic_53/10T_toy_magic_1
* x518	10T_1x8_magic_8/10T_toy_magic_1
* x519	10T_1x8_magic_10/10T_toy_magic_2
* x520	10T_1x8_magic_40/10T_toy_magic_2
* x521	10T_1x8_magic_111/10T_toy_magic_1
* x522	10T_1x8_magic_2/10T_toy_magic_7
* x523	10T_1x8_magic_56/10T_toy_magic_1
* x524	10T_1x8_magic_99/10T_toy_magic_4
* x525	10T_1x8_magic_5/10T_toy_magic_5
* x526	10T_1x8_magic_3/10T_toy_magic_0
* x527	10T_1x8_magic_74/10T_toy_magic_6
* x528	10T_1x8_magic_81/10T_toy_magic_3
* x529	10T_1x8_magic_19/10T_toy_magic_7
* x530	10T_1x8_magic_99/10T_toy_magic_6
* x531	10T_1x8_magic_40/10T_toy_magic_3
* x532	10T_1x8_magic_91/10T_toy_magic_6
* x533	10T_1x8_magic_108/10T_toy_magic_1
* x534	10T_1x8_magic_24/10T_toy_magic_2
* x535	10T_1x8_magic_10/10T_toy_magic_7
* x536	10T_1x8_magic_54/10T_toy_magic_2
* x537	10T_1x8_magic_66/10T_toy_magic_0
* x538	10T_1x8_magic_92/10T_toy_magic_0
* x539	10T_1x8_magic_13/10T_toy_magic_5
* x540	10T_1x8_magic_106/10T_toy_magic_7
* x541	10T_1x8_magic_36/10T_toy_magic_6
* x542	10T_1x8_magic_67/10T_toy_magic_3
* x543	10T_1x8_magic_5/10T_toy_magic_0
* x544	10T_1x8_magic_68/10T_toy_magic_6
* x545	10T_1x8_magic_58/10T_toy_magic_2
* x546	10T_1x8_magic_85/10T_toy_magic_0
* x547	10T_1x8_magic_127/10T_toy_magic_5
* x548	10T_1x8_magic_90/10T_toy_magic_5
* x549	10T_1x8_magic_78/10T_toy_magic_7
* x550	10T_1x8_magic_6/10T_toy_magic_6
* x551	10T_1x8_magic_104/10T_toy_magic_7
* x552	10T_1x8_magic_52/10T_toy_magic_1
* x553	10T_1x8_magic_64/10T_toy_magic_7
* x554	10T_1x8_magic_9/10T_toy_magic_1
* x555	10T_1x8_magic_67/10T_toy_magic_0
* x556	10T_1x8_magic_83/10T_toy_magic_4
* x557	10T_1x8_magic_36/10T_toy_magic_2
* x558	10T_1x8_magic_25/10T_toy_magic_5
* x559	10T_1x8_magic_3/10T_toy_magic_7
* x560	10T_1x8_magic_55/10T_toy_magic_1
* x561	10T_1x8_magic_89/10T_toy_magic_5
* x562	10T_1x8_magic_65/10T_toy_magic_3
* x563	10T_1x8_magic_72/10T_toy_magic_6
* x564	10T_1x8_magic_76/10T_toy_magic_6
* x565	10T_1x8_magic_70/10T_toy_magic_7
* x566	10T_1x8_magic_97/10T_toy_magic_6
* x567	10T_1x8_magic_122/10T_toy_magic_1
* x568	10T_1x8_magic_36/10T_toy_magic_3
* x569	10T_1x8_magic_88/10T_toy_magic_6
* x570	10T_1x8_magic_45/10T_toy_magic_0
* x571	10T_1x8_magic_49/10T_toy_magic_6
* x572	10T_1x8_magic_21/10T_toy_magic_2
* x573	10T_1x8_magic_63/10T_toy_magic_6
* x574	10T_1x8_magic_93/10T_toy_magic_0
* x575	10T_1x8_magic_99/10T_toy_magic_1
* x576	10T_1x8_magic_12/10T_toy_magic_5
* x577	10T_1x8_magic_103/10T_toy_magic_7
* x578	10T_1x8_magic_63/10T_toy_magic_7
* x579	10T_1x8_magic_125/10T_toy_magic_5
* x580	10T_1x8_magic_107/10T_toy_magic_4
* x581	10T_1x8_magic_91/10T_toy_magic_5
* x582	10T_1x8_magic_116/10T_toy_magic_5
* x583	10T_1x8_magic_102/10T_toy_magic_7
* x584	10T_1x8_magic_7/10T_toy_magic_6
* x585	10T_1x8_magic_51/10T_toy_magic_1
* x586	10T_1x8_magic_37/10T_toy_magic_5
* x587	10T_1x8_magic_31/10T_toy_magic_1
* x588	10T_1x8_magic_112/10T_toy_magic_3
* x589	10T_1x8_magic_81/10T_toy_magic_4
* x590	10T_1x8_magic_41/10T_toy_magic_4
* x591	10T_1x8_magic_21/10T_toy_magic_7
* x592	10T_1x8_magic_26/10T_toy_magic_5
* x593	10T_1x8_magic_71/10T_toy_magic_1
* x594	10T_1x8_magic_50/10T_toy_magic_7
* x595	10T_1x8_magic_86/10T_toy_magic_2
* x596	10T_1x8_magic_112/10T_toy_magic_4
* x597	10T_1x8_magic_78/10T_toy_magic_6
* x598	10T_1x8_magic_13/10T_toy_magic_6
* x599	10T_1x8_magic_42/10T_toy_magic_1
* x600	10T_1x8_magic_90/10T_toy_magic_7
* x601	10T_1x8_magic_95/10T_toy_magic_6
* x602	10T_1x8_magic_46/10T_toy_magic_0
* x603	10T_1x8_magic_48/10T_toy_magic_6
* x604	10T_1x8_magic_67/10T_toy_magic_7
* x605	10T_1x8_magic_22/10T_toy_magic_2
* x606	10T_1x8_magic_62/10T_toy_magic_6
* x607	10T_1x8_magic_16/10T_toy_magic_6
* x608	10T_1x8_magic_78/10T_toy_magic_3
* x609	10T_1x8_magic_59/10T_toy_magic_4
* x610	10T_1x8_magic_11/10T_toy_magic_5
* x611	10T_1x8_magic_62/10T_toy_magic_7
* x612	10T_1x8_magic_76/10T_toy_magic_2
* x613	10T_1x8_magic_33/10T_toy_magic_3
* x614	10T_1x8_magic_106/10T_toy_magic_4
* x615	10T_1x8_magic_88/10T_toy_magic_5
* x616	10T_1x8_magic_117/10T_toy_magic_5
* x617	10T_1x8_magic_110/10T_toy_magic_3
* x618	10T_1x8_magic_78/10T_toy_magic_4
* x619	10T_1x8_magic_108/10T_toy_magic_2
* x620	10T_1x8_magic_13/10T_toy_magic_3
* x621	10T_1x8_magic_39/10T_toy_magic_4
* x622	10T_1x8_magic_116/10T_toy_magic_4
* x623	10T_1x8_magic_15/10T_toy_magic_0
* x624	10T_1x8_magic_23/10T_toy_magic_5
* x625	10T_1x8_magic_127/10T_toy_magic_3
* x626	10T_1x8_magic_110/10T_toy_magic_4
* x627	10T_1x8_magic_44/10T_toy_magic_0
* x628	10T_1x8_magic_47/10T_toy_magic_6
* x629	10T_1x8_magic_79/10T_toy_magic_2
* x630	10T_1x8_magic_79/10T_toy_magic_3
* x631	10T_1x8_magic_58/10T_toy_magic_4
* x632	10T_1x8_magic_71/10T_toy_magic_2
* x633	10T_1x8_magic_16/10T_toy_magic_5
* x634	10T_1x8_magic_61/10T_toy_magic_3
* x635	10T_1x8_magic_74/10T_toy_magic_2
* x636	10T_1x8_magic_72/10T_toy_magic_4
* x637	10T_1x8_magic_103/10T_toy_magic_4
* x638	10T_1x8_magic_4/10T_toy_magic_3
* x639	10T_1x8_magic_38/10T_toy_magic_7
* x640	10T_1x8_magic_115/10T_toy_magic_1
* x641	10T_1x8_magic_107/10T_toy_magic_0
* x642	10T_1x8_magic_98/10T_toy_magic_0
* x643	10T_1x8_magic_123/10T_toy_magic_0
* x644	10T_1x8_magic_15/10T_toy_magic_2
* x645	10T_1x8_magic_12/10T_toy_magic_3
* x646	10T_1x8_magic_61/10T_toy_magic_1
* x647	10T_1x8_magic_123/10T_toy_magic_2
* x648	10T_1x8_magic_84/10T_toy_magic_1
* x649	10T_1x8_magic_18/10T_toy_magic_7
* x650	10T_1x8_magic_125/10T_toy_magic_3
* x651	10T_1x8_magic_75/10T_toy_magic_2
* x652	10T_1x8_magic_75/10T_toy_magic_3
* x653	10T_1x8_magic_66/10T_toy_magic_6
* x654	10T_1x8_magic_64/10T_toy_magic_0
* x655	10T_1x8_magic_82/10T_toy_magic_4
* x656	10T_1x8_magic_60/10T_toy_magic_3
* x657	10T_1x8_magic_49/10T_toy_magic_1
* x658	10T_1x8_magic_4/10T_toy_magic_7
* x659	10T_1x8_magic_29/10T_toy_magic_1
* x660	10T_1x8_magic_10/10T_toy_magic_0
* x661	10T_1x8_magic_14/10T_toy_magic_3
* x662	10T_1x8_magic_79/10T_toy_magic_0
* x663	10T_1x8_magic_64/10T_toy_magic_6
* x664	10T_1x8_magic_113/10T_toy_magic_5
* x665	10T_1x8_magic_106/10T_toy_magic_0
* x666	10T_1x8_magic_123/10T_toy_magic_7
* x667	10T_1x8_magic_121/10T_toy_magic_0
* x668	10T_1x8_magic_59/10T_toy_magic_2
* x669	10T_1x8_magic_61/10T_toy_magic_0
* x670	10T_1x8_magic_121/10T_toy_magic_2
* x671	10T_1x8_magic_33/10T_toy_magic_7
* x672	10T_1x8_magic_82/10T_toy_magic_1
* x673	10T_1x8_magic_24/10T_toy_magic_1
* x674	10T_1x8_magic_44/10T_toy_magic_5
* x675	10T_1x8_magic_114/10T_toy_magic_1
* x676	10T_1x8_magic_67/10T_toy_magic_6
* x677	10T_1x8_magic_80/10T_toy_magic_4
* x678	10T_1x8_magic_14/10T_toy_magic_7
* x679	10T_1x8_magic_26/10T_toy_magic_4
* x680	10T_1x8_magic_48/10T_toy_magic_1
* x681	10T_1x8_magic_1/10T_toy_magic_6
* x682	10T_1x8_magic_30/10T_toy_magic_1
* x683	10T_1x8_magic_17/10T_toy_magic_3
* x684	10T_1x8_magic_57/10T_toy_magic_1
* x685	10T_1x8_magic_53/10T_toy_magic_5
* x686	10T_1x8_magic_8/10T_toy_magic_5
* x687	10T_1x8_magic_83/10T_toy_magic_1
* x688	10T_1x8_magic_75/10T_toy_magic_0
* x689	10T_1x8_magic_34/10T_toy_magic_3
* x690	10T_1x8_magic_60/10T_toy_magic_0
* x691	10T_1x8_magic_80/10T_toy_magic_1
* x692	10T_1x8_magic_21/10T_toy_magic_1
* x693	10T_1x8_magic_108/10T_toy_magic_5
* x694	10T_1x8_magic_54/10T_toy_magic_7
* x695	10T_1x8_magic_97/10T_toy_magic_1
* x696	10T_1x8_magic_92/10T_toy_magic_6
* x697	10T_1x8_magic_35/10T_toy_magic_2
* x698	10T_1x8_magic_22/10T_toy_magic_3
* x699	10T_1x8_magic_99/10T_toy_magic_7
* x700	10T_1x8_magic_85/10T_toy_magic_6
* x701	10T_1x8_magic_126/10T_toy_magic_2
* x702	10T_1x8_magic_23/10T_toy_magic_4
* x703	10T_1x8_magic_47/10T_toy_magic_1
* x704	10T_1x8_magic_65/10T_toy_magic_5
* x705	10T_1x8_magic_52/10T_toy_magic_5
* x706	10T_1x8_magic_9/10T_toy_magic_5
* x707	10T_1x8_magic_82/10T_toy_magic_0
* x708	10T_1x8_magic_81/10T_toy_magic_1
* x709	10T_1x8_magic_32/10T_toy_magic_7
* x710	10T_1x8_magic_6/10T_toy_magic_7
* x711	10T_1x8_magic_87/10T_toy_magic_3
* x712	10T_1x8_magic_88/10T_toy_magic_2
* x713	10T_1x8_magic_17/10T_toy_magic_4
* x714	10T_1x8_magic_123/10T_toy_magic_4
* x715	10T_1x8_magic_22/10T_toy_magic_1
* x716	10T_1x8_magic_45/10T_toy_magic_6
* x717	10T_1x8_magic_2/10T_toy_magic_3
* x718	10T_1x8_magic_93/10T_toy_magic_6
* x719	10T_1x8_magic_102/10T_toy_magic_4
* x720	10T_1x8_magic_97/10T_toy_magic_7
* x721	10T_1x8_magic_124/10T_toy_magic_2
* x722	10T_1x8_magic_74/10T_toy_magic_7
* x723	10T_1x8_magic_24/10T_toy_magic_4
* x724	10T_1x8_magic_27/10T_toy_magic_6
* x725	10T_1x8_magic_51/10T_toy_magic_4
* x726	10T_1x8_magic_51/10T_toy_magic_5
* x727	10T_1x8_magic_19/10T_toy_magic_2
* x728	10T_1x8_magic_31/10T_toy_magic_5
* x729	10T_1x8_magic_80/10T_toy_magic_0
* x730	10T_1x8_magic_26/10T_toy_magic_0
* x731	10T_1x8_magic_7/10T_toy_magic_7
* x732	10T_1x8_magic_10/10T_toy_magic_4
* x733	10T_1x8_magic_68/10T_toy_magic_4
* x734	10T_1x8_magic_77/10T_toy_magic_3
* x735	10T_1x8_magic_122/10T_toy_magic_6
* x736	10T_1x8_magic_94/10T_toy_magic_3
* x737	10T_1x8_magic_46/10T_toy_magic_6
* x738	10T_1x8_magic_3/10T_toy_magic_3
* x739	10T_1x8_magic_69/10T_toy_magic_0
* x740	10T_1x8_magic_77/10T_toy_magic_1
* x741	10T_1x8_magic_71/10T_toy_magic_6
* x742	10T_1x8_magic_6/10T_toy_magic_0
* x743	10T_1x8_magic_95/10T_toy_magic_7
* x744	10T_1x8_magic_65/10T_toy_magic_7
* x745	10T_1x8_magic_77/10T_toy_magic_0
* x746	10T_1x8_magic_23/10T_toy_magic_0
* x747	10T_1x8_magic_42/10T_toy_magic_0
* x748	10T_1x8_magic_31/10T_toy_magic_3
* x749	10T_1x8_magic_103/10T_toy_magic_1
* x750	10T_1x8_magic_76/10T_toy_magic_1
* x751	10T_1x8_magic_7/10T_toy_magic_0
* x752	10T_1x8_magic_34/10T_toy_magic_7
* x753	10T_1x8_magic_0/10T_toy_magic_1
* x754	10T_1x8_magic_71/10T_toy_magic_5
* x755	10T_1x8_magic_32/10T_toy_magic_2
* x756	10T_1x8_magic_115/10T_toy_magic_5
* x757	10T_1x8_magic_107/10T_toy_magic_6
* x758	10T_1x8_magic_98/10T_toy_magic_6
* x759	10T_1x8_magic_123/10T_toy_magic_6
* x760	10T_1x8_magic_50/10T_toy_magic_3
* x761	10T_1x8_magic_41/10T_toy_magic_0
* x762	10T_1x8_magic_84/10T_toy_magic_5
* x763	10T_1x8_magic_96/10T_toy_magic_7
* x764	10T_1x8_magic_35/10T_toy_magic_7
* x765	10T_1x8_magic_75/10T_toy_magic_7
* x766	10T_1x8_magic_70/10T_toy_magic_1
* x767	10T_1x8_magic_101/10T_toy_magic_1
* x768	10T_1x8_magic_18/10T_toy_magic_4
* x769	10T_1x8_magic_74/10T_toy_magic_1
* x770	10T_1x8_magic_65/10T_toy_magic_0
* x771	10T_1x8_magic_1/10T_toy_magic_1
* x772	10T_1x8_magic_49/10T_toy_magic_5
* x773	10T_1x8_magic_69/10T_toy_magic_5
* x774	10T_1x8_magic_19/10T_toy_magic_6
* x775	10T_1x8_magic_29/10T_toy_magic_5
* x776	10T_1x8_magic_33/10T_toy_magic_2
* x777	10T_1x8_magic_106/10T_toy_magic_6
* x778	10T_1x8_magic_24/10T_toy_magic_7
* x779	10T_1x8_magic_96/10T_toy_magic_6
* x780	10T_1x8_magic_121/10T_toy_magic_6
* x781	10T_1x8_magic_31/10T_toy_magic_7
* x782	10T_1x8_magic_61/10T_toy_magic_6
* x783	10T_1x8_magic_39/10T_toy_magic_0
* x784	10T_1x8_magic_24/10T_toy_magic_5
* x785	10T_1x8_magic_27/10T_toy_magic_2
* x786	10T_1x8_magic_15/10T_toy_magic_6
* x787	10T_1x8_magic_94/10T_toy_magic_7
* x788	10T_1x8_magic_84/10T_toy_magic_6
* x789	10T_1x8_magic_109/10T_toy_magic_2
* x790	10T_1x8_magic_65/10T_toy_magic_4
* x791	10T_1x8_magic_114/10T_toy_magic_5
* x792	10T_1x8_magic_25/10T_toy_magic_4
* x793	10T_1x8_magic_53/10T_toy_magic_7
* x794	10T_1x8_magic_63/10T_toy_magic_3
* x795	10T_1x8_magic_48/10T_toy_magic_5
* x796	10T_1x8_magic_30/10T_toy_magic_5
* x797	10T_1x8_magic_102/10T_toy_magic_0
* x798	10T_1x8_magic_75/10T_toy_magic_6
* x799	10T_1x8_magic_127/10T_toy_magic_2
* x800	10T_1x8_magic_60/10T_toy_magic_6
* x801	10T_1x8_magic_17/10T_toy_magic_7
* x802	10T_1x8_magic_21/10T_toy_magic_5
* x803	10T_1x8_magic_82/10T_toy_magic_6
* x804	10T_1x8_magic_90/10T_toy_magic_3
* x805	10T_1x8_magic_98/10T_toy_magic_4
* x806	10T_1x8_magic_52/10T_toy_magic_7
* x807	10T_1x8_magic_62/10T_toy_magic_3
* x808	10T_1x8_magic_47/10T_toy_magic_5
* x809	10T_1x8_magic_71/10T_toy_magic_3
* x810	10T_1x8_magic_100/10T_toy_magic_0
* x811	10T_1x8_magic_125/10T_toy_magic_2
* x812	10T_1x8_magic_86/10T_toy_magic_1
* x813	10T_1x8_magic_85/10T_toy_magic_2
* x814	10T_1x8_magic_92/10T_toy_magic_7
* x815	10T_1x8_magic_101/10T_toy_magic_2
* x816	10T_1x8_magic_71/10T_toy_magic_7
* x817	10T_1x8_magic_22/10T_toy_magic_5
* x818	10T_1x8_magic_29/10T_toy_magic_3
* x819	10T_1x8_magic_101/10T_toy_magic_3
* x820	10T_1x8_magic_37/10T_toy_magic_2
* x821	10T_1x8_magic_78/10T_toy_magic_1
* x822	10T_1x8_magic_69/10T_toy_magic_3
* x823	10T_1x8_magic_80/10T_toy_magic_6
* x824	10T_1x8_magic_91/10T_toy_magic_3
* x825	10T_1x8_magic_11/10T_toy_magic_0
* x826	10T_1x8_magic_93/10T_toy_magic_7
* x827	10T_1x8_magic_30/10T_toy_magic_3
* x828	10T_1x8_magic_35/10T_toy_magic_6
* x829	10T_1x8_magic_101/10T_toy_magic_0
* x830	10T_1x8_magic_40/10T_toy_magic_0
* x831	10T_1x8_magic_118/10T_toy_magic_1
* x832	10T_1x8_magic_42/10T_toy_magic_6
* x833	10T_1x8_magic_25/10T_toy_magic_6
* x834	10T_1x8_magic_89/10T_toy_magic_7
* x835	10T_1x8_magic_103/10T_toy_magic_5
* x836	10T_1x8_magic_92/10T_toy_magic_4
* x837	10T_1x8_magic_76/10T_toy_magic_5
* x838	10T_1x8_magic_0/10T_toy_magic_5
* x839	10T_1x8_magic_113/10T_toy_magic_3
* x840	10T_1x8_magic_105/10T_toy_magic_3
* x841	10T_1x8_magic_41/10T_toy_magic_6
* x842	10T_1x8_magic_64/10T_toy_magic_3
* x843	10T_1x8_magic_48/10T_toy_magic_4
* x844	10T_1x8_magic_20/10T_toy_magic_5
* x845	10T_1x8_magic_101/10T_toy_magic_5
* x846	10T_1x8_magic_93/10T_toy_magic_4
* x847	10T_1x8_magic_74/10T_toy_magic_5
* x848	10T_1x8_magic_1/10T_toy_magic_5
* x849	10T_1x8_magic_53/10T_toy_magic_2
* x850	10T_1x8_magic_105/10T_toy_magic_0
* x851	10T_1x8_magic_111/10T_toy_magic_3
* x852	10T_1x8_magic_104/10T_toy_magic_3
* x853	10T_1x8_magic_39/10T_toy_magic_6
* x854	10T_1x8_magic_73/10T_toy_magic_3
* x855	10T_1x8_magic_89/10T_toy_magic_4
* x856	10T_1x8_magic_59/10T_toy_magic_3
* x857	10T_1x8_magic_2/10T_toy_magic_1
* x858	10T_1x8_magic_92/10T_toy_magic_1
* x859	10T_1x8_magic_52/10T_toy_magic_2
* x860	10T_1x8_magic_9/10T_toy_magic_2
* x861	10T_1x8_magic_104/10T_toy_magic_0
* x862	10T_1x8_magic_102/10T_toy_magic_6
* x863	10T_1x8_magic_74/10T_toy_magic_3
* x864	10T_1x8_magic_70/10T_toy_magic_5
* x865	10T_1x8_magic_13/10T_toy_magic_2
* x866	10T_1x8_magic_43/10T_toy_magic_0
* x867	10T_1x8_magic_1/10T_toy_magic_3
* x868	10T_1x8_magic_44/10T_toy_magic_3
* x869	10T_1x8_magic_58/10T_toy_magic_3
* x870	10T_1x8_magic_93/10T_toy_magic_1
* x871	10T_1x8_magic_13/10T_toy_magic_7
* x872	10T_1x8_magic_31/10T_toy_magic_2
* x873	10T_1x8_magic_54/10T_toy_magic_0
* x874	10T_1x8_magic_100/10T_toy_magic_6
* x875	10T_1x8_magic_68/10T_toy_magic_5
* x876	10T_1x8_magic_12/10T_toy_magic_2
* x877	10T_1x8_magic_86/10T_toy_magic_5
* x878	10T_1x8_magic_85/10T_toy_magic_7
* x879	10T_1x8_magic_90/10T_toy_magic_4
* x880	10T_1x8_magic_78/10T_toy_magic_5
* x881	10T_1x8_magic_100/10T_toy_magic_1
* x882	10T_1x8_magic_37/10T_toy_magic_7
* x883	10T_1x8_magic_17/10T_toy_magic_1
* x884	10T_1x8_magic_84/10T_toy_magic_7
* x885	10T_1x8_magic_8/10T_toy_magic_6
* x886	10T_1x8_magic_12/10T_toy_magic_7
* x887	10T_1x8_magic_73/10T_toy_magic_0
* x888	10T_1x8_magic_59/10T_toy_magic_0
* x889	10T_1x8_magic_107/10T_toy_magic_3
* x890	10T_1x8_magic_91/10T_toy_magic_4
* x891	10T_1x8_magic_61/10T_toy_magic_5
* x892	10T_1x8_magic_28/10T_toy_magic_4
* x893	10T_1x8_magic_22/10T_toy_magic_7
* x894	10T_1x8_magic_40/10T_toy_magic_6
* x895	10T_1x8_magic_118/10T_toy_magic_5
* x896	10T_1x8_magic_25/10T_toy_magic_3
* x897	10T_1x8_magic_89/10T_toy_magic_2
* x898	10T_1x8_magic_106/10T_toy_magic_3
* x899	10T_1x8_magic_40/10T_toy_magic_7
* x900	10T_1x8_magic_88/10T_toy_magic_4
* x901	10T_1x8_magic_85/10T_toy_magic_4
* x902	10T_1x8_magic_60/10T_toy_magic_5
* x903	10T_1x8_magic_112/10T_toy_magic_1
* x904	10T_1x8_magic_49/10T_toy_magic_2
* x905	10T_1x8_magic_26/10T_toy_magic_3
* x906	10T_1x8_magic_87/10T_toy_magic_2
* x907	10T_1x8_magic_103/10T_toy_magic_3
* x908	10T_1x8_magic_36/10T_toy_magic_7
* x909	10T_1x8_magic_63/10T_toy_magic_1
* x910	10T_1x8_magic_100/10T_toy_magic_2
* x911	10T_1x8_magic_110/10T_toy_magic_1
* x912	10T_1x8_magic_48/10T_toy_magic_2
* x913	10T_1x8_magic_23/10T_toy_magic_3
* x914	10T_1x8_magic_72/10T_toy_magic_1
* x915	10T_1x8_magic_62/10T_toy_magic_1
* x916	10T_1x8_magic_6/10T_toy_magic_1
* x917	10T_1x8_magic_92/10T_toy_magic_5
* x918	10T_1x8_magic_103/10T_toy_magic_0
* x919	10T_1x8_magic_38/10T_toy_magic_0
* x920	10T_1x8_magic_115/10T_toy_magic_7
* x921	10T_1x8_magic_47/10T_toy_magic_2
* x922	10T_1x8_magic_72/10T_toy_magic_7
* x923	10T_1x8_magic_28/10T_toy_magic_6
* x924	10T_1x8_magic_66/10T_toy_magic_1
* x925	10T_1x8_magic_15/10T_toy_magic_4
* x926	10T_1x8_magic_27/10T_toy_magic_1
* x927	10T_1x8_magic_7/10T_toy_magic_1
* x928	10T_1x8_magic_93/10T_toy_magic_5
* x929	10T_1x8_magic_45/10T_toy_magic_5
* x930	10T_1x8_magic_54/10T_toy_magic_6
* x931	10T_1x8_magic_84/10T_toy_magic_4
* x932	10T_1x8_magic_67/10T_toy_magic_1
* x933	10T_1x8_magic_77/10T_toy_magic_2
* x934	10T_1x8_magic_100/10T_toy_magic_5
* x935	10T_1x8_magic_42/10T_toy_magic_4
* x936	10T_1x8_magic_66/10T_toy_magic_2
* x937	10T_1x8_magic_108/10T_toy_magic_0
* x938	10T_1x8_magic_46/10T_toy_magic_5
* x939	10T_1x8_magic_99/10T_toy_magic_3
* x940	10T_1x8_magic_0/10T_toy_magic_2
* x941	10T_1x8_magic_45/10T_toy_magic_2
* x942	10T_1x8_magic_21/10T_toy_magic_3
* x943	10T_1x8_magic_117/10T_toy_magic_2
* x944	10T_1x8_magic_97/10T_toy_magic_3
* x945	10T_1x8_magic_126/10T_toy_magic_6
* x946	10T_1x8_magic_46/10T_toy_magic_2
* x947	10T_1x8_magic_87/10T_toy_magic_7
* x948	10T_1x8_magic_102/10T_toy_magic_1
* x949	10T_1x8_magic_89/10T_toy_magic_0
* x950	10T_1x8_magic_86/10T_toy_magic_7
* x951	10T_1x8_magic_124/10T_toy_magic_6
* x952	10T_1x8_magic_48/10T_toy_magic_7
* x953	10T_1x8_magic_4/10T_toy_magic_4
* x954	10T_1x8_magic_6/10T_toy_magic_5
* x955	10T_1x8_magic_90/10T_toy_magic_2
* x956	10T_1x8_magic_115/10T_toy_magic_2
* x957	10T_1x8_magic_38/10T_toy_magic_6
* x958	10T_1x8_magic_114/10T_toy_magic_4
* x959	10T_1x8_magic_47/10T_toy_magic_7
* x960	10T_1x8_magic_37/10T_toy_magic_4
* x961	10T_1x8_magic_14/10T_toy_magic_4
* x962	10T_1x8_magic_87/10T_toy_magic_4
* x963	10T_1x8_magic_7/10T_toy_magic_5
* x964	10T_1x8_magic_91/10T_toy_magic_2
* x965	10T_1x8_magic_29/10T_toy_magic_2
* x966	10T_1x8_magic_15/10T_toy_magic_3
* x967	10T_1x8_magic_113/10T_toy_magic_2
* x968	10T_1x8_magic_107/10T_toy_magic_1
* x969	10T_1x8_magic_25/10T_toy_magic_0
* x970	10T_1x8_magic_30/10T_toy_magic_2
* x971	10T_1x8_magic_111/10T_toy_magic_2
* x972	10T_1x8_magic_106/10T_toy_magic_1
* x973	10T_1x8_magic_34/10T_toy_magic_4
* x974	10T_1x8_magic_98/10T_toy_magic_7
* x975	10T_1x8_magic_4/10T_toy_magic_6
* x976	10T_1x8_magic_118/10T_toy_magic_7
* x977	10T_1x8_magic_14/10T_toy_magic_6
* x978	10T_1x8_magic_102/10T_toy_magic_5
* x979	10T_1x8_magic_89/10T_toy_magic_6
* x980	10T_1x8_magic_43/10T_toy_magic_4
* x981	10T_1x8_magic_66/10T_toy_magic_7
* x982	10T_1x8_magic_24/10T_toy_magic_3
* x983	10T_1x8_magic_19/10T_toy_magic_0
* x984	10T_1x8_magic_119/10T_toy_magic_1
* x985	10T_1x8_magic_113/10T_toy_magic_7
* x986	10T_1x8_magic_107/10T_toy_magic_5
* x987	10T_1x8_magic_115/10T_toy_magic_0
* x988	10T_1x8_magic_2/10T_toy_magic_6
* x989	10T_1x8_magic_112/10T_toy_magic_7
* x990	10T_1x8_magic_111/10T_toy_magic_7
* x991	10T_1x8_magic_106/10T_toy_magic_5
* x992	10T_1x8_magic_110/10T_toy_magic_7
* x993	10T_1x8_magic_3/10T_toy_magic_6
* x994	10T_1x8_magic_41/10T_toy_magic_1
* x995	10T_1x8_magic_49/10T_toy_magic_4
* x996	10T_1x8_magic_117/10T_toy_magic_4
* x997	10T_1x8_magic_39/10T_toy_magic_1
* x998	10T_1x8_magic_33/10T_toy_magic_0
* x999	10T_1x8_magic_35/10T_toy_magic_4
* x1000	10T_1x8_magic_88/10T_toy_magic_3
* x1001	10T_1x8_magic_28/10T_toy_magic_0
* x1002	10T_1x8_magic_118/10T_toy_magic_2
* x1003	10T_1x8_magic_119/10T_toy_magic_5
* x1004	10T_1x8_magic_56/10T_toy_magic_4
* x1005	10T_1x8_magic_59/10T_toy_magic_5
* x1006	10T_1x8_magic_33/10T_toy_magic_5
* x1007	10T_1x8_magic_55/10T_toy_magic_4
* x1008	10T_1x8_magic_37/10T_toy_magic_3
* x1009	10T_1x8_magic_116/10T_toy_magic_2
* x1010	10T_1x8_magic_114/10T_toy_magic_3
* x1011	10T_1x8_magic_4/10T_toy_magic_0
* x1012	10T_1x8_magic_14/10T_toy_magic_0
* x1013	10T_1x8_magic_20/10T_toy_magic_1
* x1014	10T_1x8_magic_84/10T_toy_magic_0
* x1015	10T_1x8_magic_64/10T_toy_magic_5
* x1016	10T_1x8_magic_77/10T_toy_magic_6
* x1017	10T_1x8_magic_117/10T_toy_magic_3
* x1018	10T_1x8_magic_86/10T_toy_magic_0
* x1019	10T_1x8_magic_105/10T_toy_magic_6
* x1020	10T_1x8_magic_104/10T_toy_magic_6
* x1021	10T_1x8_magic_92/10T_toy_magic_2
* x1022	10T_1x8_magic_93/10T_toy_magic_2
* x1023	10T_1x8_magic_119/10T_toy_magic_2
