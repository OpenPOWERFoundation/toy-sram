** sch_path: /home/rjridle/osu-toy-sram/xschem/10T_toy_xschem.sch
.subckt 10T_toy_xschem WWL RWL0 RWL1 WBL WBLb RBL0 RBL1
*.PININFO WWL:I RWL0:I RWL1:I WBL:I WBLb:I RBL0:O RBL1:O
x1 net1 net2 VDD GND INVX1
x2 net2 net1 VDD GND INVX1
XM1 net2 WWL WBL GND sky130_fd_pr__nfet_01v8 L=0.15 W=1
XM2 WBLb WWL net1 GND sky130_fd_pr__nfet_01v8 L=0.15 W=1
XM3 net3 net2 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1
XM4 RBL0 RWL0 net3 GND sky130_fd_pr__nfet_01v8 L=0.15 W=1
XM5 net4 net1 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1
XM6 RBL1 RWL1 net4 GND sky130_fd_pr__nfet_01v8 L=0.15 W=1
.ends

* expanding   symbol:  INVX1.sym # of pins=2
** sym_path: /home/rjridle/osu-toy-sram/xschem/INVX1.sym
** sch_path: /home/rjridle/osu-toy-sram/xschem/INVX1.sch
.subckt INVX1  Y A  VDD  GND
*.PININFO A:I Y:O
XM1 Y A GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1
XM2 Y A VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1
.ends

.end
