module local_eval (
   inout VDD,
   inout GND,
   //input PRE_L_b,
   input RBL_L_b,
   input PRE_R_b,
   input RBL_R_b,
   output RBL_O
);
endmodule