magic
tech sky130A
magscale 1 2
timestamp 1639519430
<< error_s >>
rect 49 453 79 485
rect 167 481 199 487
rect 150 471 216 481
rect 34 451 79 453
rect 34 445 53 451
rect 24 437 53 445
rect 17 431 53 437
rect 68 431 74 451
rect 116 445 122 453
rect 129 451 237 471
rect 87 435 122 445
rect 167 437 183 451
rect 87 431 138 435
rect 17 429 138 431
rect 167 429 174 437
rect 192 429 199 451
rect 244 445 250 453
rect 287 451 317 485
rect 244 435 279 445
rect 228 431 279 435
rect 292 431 298 451
rect 326 445 332 453
rect 341 445 354 453
rect 325 431 354 445
rect 228 429 354 431
rect -1 421 59 429
rect -1 409 33 421
rect 34 409 59 421
rect -1 401 59 409
rect 68 417 74 429
rect 87 425 138 429
rect 87 421 199 425
rect 87 417 104 421
rect 116 419 199 421
rect 228 421 298 429
rect 68 409 104 417
rect 68 401 112 409
rect 24 385 53 401
rect 34 329 53 385
rect 68 329 74 401
rect 79 399 112 401
rect 121 399 138 419
rect 228 409 272 421
rect 279 415 298 421
rect 325 421 367 429
rect 325 417 332 421
rect 274 409 298 415
rect 228 401 298 409
rect 310 409 332 417
rect 333 409 367 421
rect 310 401 367 409
rect 79 398 200 399
rect 239 398 287 401
rect 79 387 287 398
rect 87 385 103 387
rect 90 329 96 385
rect 104 381 120 387
rect 129 365 159 376
rect 174 371 200 387
rect 250 384 262 387
rect 220 382 221 383
rect 221 381 230 382
rect 221 376 231 381
rect 236 376 242 381
rect 124 360 166 365
rect 207 360 242 376
rect 124 342 175 360
rect 207 342 253 360
rect 113 329 175 342
rect 191 329 253 342
rect 270 329 276 369
rect 292 329 298 401
rect 325 385 354 401
rect 326 329 332 385
rect 34 323 332 329
rect 341 323 354 385
rect 25 241 354 323
rect 25 227 341 241
rect 26 225 123 227
rect 26 219 54 225
rect 25 211 54 219
rect 18 205 54 211
rect 69 209 123 225
rect 129 225 160 227
rect 129 209 130 225
rect 69 207 139 209
rect 69 205 75 207
rect 88 205 139 207
rect 18 203 139 205
rect 168 203 175 227
rect 183 225 238 227
rect 245 225 318 227
rect 188 215 235 225
rect 193 209 235 215
rect 245 209 299 225
rect 327 219 355 227
rect 193 207 299 209
rect 193 205 280 207
rect 293 205 299 207
rect 326 205 355 219
rect 193 203 200 205
rect 229 203 355 205
rect 0 195 60 203
rect 0 183 34 195
rect 35 183 60 195
rect 0 175 60 183
rect 69 191 75 203
rect 88 199 139 203
rect 88 195 167 199
rect 88 191 105 195
rect 116 193 167 195
rect 229 195 299 203
rect 69 183 105 191
rect 69 175 113 183
rect 25 169 54 175
rect 69 169 75 175
rect 80 173 113 175
rect 122 173 139 193
rect 229 183 273 195
rect 280 189 299 195
rect 326 195 368 203
rect 326 191 333 195
rect 275 183 299 189
rect 229 175 299 183
rect 311 183 333 191
rect 334 183 368 195
rect 311 175 368 183
rect 80 172 201 173
rect 240 172 288 175
rect 80 169 288 172
rect 293 169 299 175
rect 326 169 355 175
rect 25 159 355 169
rect 26 97 355 159
rect 35 15 54 97
rect 69 69 75 97
rect 91 91 97 97
rect 125 84 146 97
rect 87 73 109 83
rect 125 79 131 84
rect 133 79 145 84
rect 167 81 175 89
rect 208 84 224 97
rect 271 83 277 97
rect 145 77 147 79
rect 87 69 121 73
rect 167 71 185 81
rect 247 71 281 83
rect 167 69 281 71
rect 293 69 299 97
rect 69 61 299 69
rect 69 55 75 61
rect 80 55 130 61
rect 238 55 299 61
rect 69 39 137 55
rect 231 52 299 55
rect 145 43 299 52
rect 231 39 299 43
rect 69 15 75 39
rect 85 31 103 39
rect 87 23 103 31
rect 117 15 123 39
rect 168 37 175 39
rect 193 37 200 39
rect 168 35 200 37
rect 167 29 201 35
rect 151 17 217 29
rect 245 23 263 39
rect 49 13 50 15
rect 75 -17 80 1
rect 130 -1 238 17
rect 245 15 251 23
rect 293 15 299 39
rect 318 13 319 93
rect 327 15 333 97
rect 342 15 355 97
rect 130 -17 160 -1
rect 168 -15 238 -1
rect 200 -17 238 -15
rect 288 -17 293 1
rect 200 -35 236 -17
use sram_sp  sram_sp_1
timestamp 1639519430
transform 0 1 25 -1 0 467
box -26 -26 312 342
use sram_sp  sram_sp_0
timestamp 1639519430
transform 0 1 26 -1 0 241
box -26 -26 312 342
<< end >>
