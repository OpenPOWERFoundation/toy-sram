VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO 10T_16x8_magic
  CLASS BLOCK ;
  FOREIGN 10T_16x8_magic ;
  ORIGIN 0.035 0.020 ;
  SIZE 23.190 BY 21.830 ;
  PIN RBL1_0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 0.000 20.440 0.075 20.650 ;
        RECT 0.000 19.090 0.075 19.300 ;
        RECT 0.000 17.740 0.075 17.950 ;
        RECT 0.000 16.390 0.075 16.600 ;
        RECT 0.000 15.040 0.075 15.250 ;
        RECT 0.000 13.690 0.075 13.900 ;
        RECT 0.000 12.340 0.075 12.550 ;
        RECT 0.000 10.990 0.075 11.200 ;
        RECT 0.000 9.640 0.075 9.850 ;
        RECT 0.000 8.290 0.075 8.500 ;
        RECT 0.000 6.940 0.075 7.150 ;
        RECT 0.000 5.590 0.075 5.800 ;
        RECT 0.000 4.240 0.075 4.450 ;
        RECT 0.000 2.890 0.075 3.100 ;
        RECT 0.000 1.540 0.075 1.750 ;
        RECT 0.000 0.190 0.075 0.400 ;
    END
  END RBL1_0
  PIN RBL0_0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 2.685 20.440 2.760 20.650 ;
        RECT 2.685 19.090 2.760 19.300 ;
        RECT 2.685 17.740 2.760 17.950 ;
        RECT 2.685 16.390 2.760 16.600 ;
        RECT 2.685 15.040 2.760 15.250 ;
        RECT 2.685 13.690 2.760 13.900 ;
        RECT 2.685 12.340 2.760 12.550 ;
        RECT 2.685 10.990 2.760 11.200 ;
        RECT 2.685 9.640 2.760 9.850 ;
        RECT 2.685 8.290 2.760 8.500 ;
        RECT 2.685 6.940 2.760 7.150 ;
        RECT 2.685 5.590 2.760 5.800 ;
        RECT 2.685 4.240 2.760 4.450 ;
        RECT 2.685 2.890 2.760 3.100 ;
        RECT 2.685 1.540 2.760 1.750 ;
        RECT 2.685 0.190 2.760 0.400 ;
    END
  END RBL0_0
  PIN RBL1_1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 2.900 20.440 2.975 20.650 ;
        RECT 2.900 19.090 2.975 19.300 ;
        RECT 2.900 17.740 2.975 17.950 ;
        RECT 2.900 16.390 2.975 16.600 ;
        RECT 2.900 15.040 2.975 15.250 ;
        RECT 2.900 13.690 2.975 13.900 ;
        RECT 2.900 12.340 2.975 12.550 ;
        RECT 2.900 10.990 2.975 11.200 ;
        RECT 2.900 9.640 2.975 9.850 ;
        RECT 2.900 8.290 2.975 8.500 ;
        RECT 2.900 6.940 2.975 7.150 ;
        RECT 2.900 5.590 2.975 5.800 ;
        RECT 2.900 4.240 2.975 4.450 ;
        RECT 2.900 2.890 2.975 3.100 ;
        RECT 2.900 1.540 2.975 1.750 ;
        RECT 2.900 0.190 2.975 0.400 ;
    END
  END RBL1_1
  PIN RBL0_1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 5.585 20.440 5.660 20.650 ;
        RECT 5.585 19.090 5.660 19.300 ;
        RECT 5.585 17.740 5.660 17.950 ;
        RECT 5.585 16.390 5.660 16.600 ;
        RECT 5.585 15.040 5.660 15.250 ;
        RECT 5.585 13.690 5.660 13.900 ;
        RECT 5.585 12.340 5.660 12.550 ;
        RECT 5.585 10.990 5.660 11.200 ;
        RECT 5.585 9.640 5.660 9.850 ;
        RECT 5.585 8.290 5.660 8.500 ;
        RECT 5.585 6.940 5.660 7.150 ;
        RECT 5.585 5.590 5.660 5.800 ;
        RECT 5.585 4.240 5.660 4.450 ;
        RECT 5.585 2.890 5.660 3.100 ;
        RECT 5.585 1.540 5.660 1.750 ;
        RECT 5.585 0.190 5.660 0.400 ;
    END
  END RBL0_1
  PIN RBL1_2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 5.800 20.440 5.875 20.650 ;
        RECT 5.800 19.090 5.875 19.300 ;
        RECT 5.800 17.740 5.875 17.950 ;
        RECT 5.800 16.390 5.875 16.600 ;
        RECT 5.800 15.040 5.875 15.250 ;
        RECT 5.800 13.690 5.875 13.900 ;
        RECT 5.800 12.340 5.875 12.550 ;
        RECT 5.800 10.990 5.875 11.200 ;
        RECT 5.800 9.640 5.875 9.850 ;
        RECT 5.800 8.290 5.875 8.500 ;
        RECT 5.800 6.940 5.875 7.150 ;
        RECT 5.800 5.590 5.875 5.800 ;
        RECT 5.800 4.240 5.875 4.450 ;
        RECT 5.800 2.890 5.875 3.100 ;
        RECT 5.800 1.540 5.875 1.750 ;
        RECT 5.800 0.190 5.875 0.400 ;
    END
  END RBL1_2
  PIN RBL0_2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 8.485 20.440 8.560 20.650 ;
        RECT 8.485 19.090 8.560 19.300 ;
        RECT 8.485 17.740 8.560 17.950 ;
        RECT 8.485 16.390 8.560 16.600 ;
        RECT 8.485 15.040 8.560 15.250 ;
        RECT 8.485 13.690 8.560 13.900 ;
        RECT 8.485 12.340 8.560 12.550 ;
        RECT 8.485 10.990 8.560 11.200 ;
        RECT 8.485 9.640 8.560 9.850 ;
        RECT 8.485 8.290 8.560 8.500 ;
        RECT 8.485 6.940 8.560 7.150 ;
        RECT 8.485 5.590 8.560 5.800 ;
        RECT 8.485 4.240 8.560 4.450 ;
        RECT 8.485 2.890 8.560 3.100 ;
        RECT 8.485 1.540 8.560 1.750 ;
        RECT 8.485 0.190 8.560 0.400 ;
    END
  END RBL0_2
  PIN RBL1_3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 8.700 20.440 8.775 20.650 ;
        RECT 8.700 19.090 8.775 19.300 ;
        RECT 8.700 17.740 8.775 17.950 ;
        RECT 8.700 16.390 8.775 16.600 ;
        RECT 8.700 15.040 8.775 15.250 ;
        RECT 8.700 13.690 8.775 13.900 ;
        RECT 8.700 12.340 8.775 12.550 ;
        RECT 8.700 10.990 8.775 11.200 ;
        RECT 8.700 9.640 8.775 9.850 ;
        RECT 8.700 8.290 8.775 8.500 ;
        RECT 8.700 6.940 8.775 7.150 ;
        RECT 8.700 5.590 8.775 5.800 ;
        RECT 8.700 4.240 8.775 4.450 ;
        RECT 8.700 2.890 8.775 3.100 ;
        RECT 8.700 1.540 8.775 1.750 ;
        RECT 8.700 0.190 8.775 0.400 ;
    END
  END RBL1_3
  PIN RBL0_3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 11.385 20.440 11.460 20.650 ;
        RECT 11.385 19.090 11.460 19.300 ;
        RECT 11.385 17.740 11.460 17.950 ;
        RECT 11.385 16.390 11.460 16.600 ;
        RECT 11.385 15.040 11.460 15.250 ;
        RECT 11.385 13.690 11.460 13.900 ;
        RECT 11.385 12.340 11.460 12.550 ;
        RECT 11.385 10.990 11.460 11.200 ;
        RECT 11.385 9.640 11.460 9.850 ;
        RECT 11.385 8.290 11.460 8.500 ;
        RECT 11.385 6.940 11.460 7.150 ;
        RECT 11.385 5.590 11.460 5.800 ;
        RECT 11.385 4.240 11.460 4.450 ;
        RECT 11.385 2.890 11.460 3.100 ;
        RECT 11.385 1.540 11.460 1.750 ;
        RECT 11.385 0.190 11.460 0.400 ;
    END
  END RBL0_3
  PIN RBL1_4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 11.600 20.440 11.675 20.650 ;
        RECT 11.600 19.090 11.675 19.300 ;
        RECT 11.600 17.740 11.675 17.950 ;
        RECT 11.600 16.390 11.675 16.600 ;
        RECT 11.600 15.040 11.675 15.250 ;
        RECT 11.600 13.690 11.675 13.900 ;
        RECT 11.600 12.340 11.675 12.550 ;
        RECT 11.600 10.990 11.675 11.200 ;
        RECT 11.600 9.640 11.675 9.850 ;
        RECT 11.600 8.290 11.675 8.500 ;
        RECT 11.600 6.940 11.675 7.150 ;
        RECT 11.600 5.590 11.675 5.800 ;
        RECT 11.600 4.240 11.675 4.450 ;
        RECT 11.600 2.890 11.675 3.100 ;
        RECT 11.600 1.540 11.675 1.750 ;
        RECT 11.600 0.190 11.675 0.400 ;
    END
  END RBL1_4
  PIN RBL0_4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 14.285 20.440 14.360 20.650 ;
        RECT 14.285 19.090 14.360 19.300 ;
        RECT 14.285 17.740 14.360 17.950 ;
        RECT 14.285 16.390 14.360 16.600 ;
        RECT 14.285 15.040 14.360 15.250 ;
        RECT 14.285 13.690 14.360 13.900 ;
        RECT 14.285 12.340 14.360 12.550 ;
        RECT 14.285 10.990 14.360 11.200 ;
        RECT 14.285 9.640 14.360 9.850 ;
        RECT 14.285 8.290 14.360 8.500 ;
        RECT 14.285 6.940 14.360 7.150 ;
        RECT 14.285 5.590 14.360 5.800 ;
        RECT 14.285 4.240 14.360 4.450 ;
        RECT 14.285 2.890 14.360 3.100 ;
        RECT 14.285 1.540 14.360 1.750 ;
        RECT 14.285 0.190 14.360 0.400 ;
    END
  END RBL0_4
  PIN RBL1_5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 14.500 20.440 14.575 20.650 ;
        RECT 14.500 19.090 14.575 19.300 ;
        RECT 14.500 17.740 14.575 17.950 ;
        RECT 14.500 16.390 14.575 16.600 ;
        RECT 14.500 15.040 14.575 15.250 ;
        RECT 14.500 13.690 14.575 13.900 ;
        RECT 14.500 12.340 14.575 12.550 ;
        RECT 14.500 10.990 14.575 11.200 ;
        RECT 14.500 9.640 14.575 9.850 ;
        RECT 14.500 8.290 14.575 8.500 ;
        RECT 14.500 6.940 14.575 7.150 ;
        RECT 14.500 5.590 14.575 5.800 ;
        RECT 14.500 4.240 14.575 4.450 ;
        RECT 14.500 2.890 14.575 3.100 ;
        RECT 14.500 1.540 14.575 1.750 ;
        RECT 14.500 0.190 14.575 0.400 ;
    END
  END RBL1_5
  PIN RBL0_5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 17.185 20.440 17.260 20.650 ;
        RECT 17.185 19.090 17.260 19.300 ;
        RECT 17.185 17.740 17.260 17.950 ;
        RECT 17.185 16.390 17.260 16.600 ;
        RECT 17.185 15.040 17.260 15.250 ;
        RECT 17.185 13.690 17.260 13.900 ;
        RECT 17.185 12.340 17.260 12.550 ;
        RECT 17.185 10.990 17.260 11.200 ;
        RECT 17.185 9.640 17.260 9.850 ;
        RECT 17.185 8.290 17.260 8.500 ;
        RECT 17.185 6.940 17.260 7.150 ;
        RECT 17.185 5.590 17.260 5.800 ;
        RECT 17.185 4.240 17.260 4.450 ;
        RECT 17.185 2.890 17.260 3.100 ;
        RECT 17.185 1.540 17.260 1.750 ;
        RECT 17.185 0.190 17.260 0.400 ;
    END
  END RBL0_5
  PIN RBL1_6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 17.400 20.440 17.475 20.650 ;
        RECT 17.400 19.090 17.475 19.300 ;
        RECT 17.400 17.740 17.475 17.950 ;
        RECT 17.400 16.390 17.475 16.600 ;
        RECT 17.400 15.040 17.475 15.250 ;
        RECT 17.400 13.690 17.475 13.900 ;
        RECT 17.400 12.340 17.475 12.550 ;
        RECT 17.400 10.990 17.475 11.200 ;
        RECT 17.400 9.640 17.475 9.850 ;
        RECT 17.400 8.290 17.475 8.500 ;
        RECT 17.400 6.940 17.475 7.150 ;
        RECT 17.400 5.590 17.475 5.800 ;
        RECT 17.400 4.240 17.475 4.450 ;
        RECT 17.400 2.890 17.475 3.100 ;
        RECT 17.400 1.540 17.475 1.750 ;
        RECT 17.400 0.190 17.475 0.400 ;
    END
  END RBL1_6
  PIN RBL0_6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 20.085 20.440 20.160 20.650 ;
        RECT 20.085 19.090 20.160 19.300 ;
        RECT 20.085 17.740 20.160 17.950 ;
        RECT 20.085 16.390 20.160 16.600 ;
        RECT 20.085 15.040 20.160 15.250 ;
        RECT 20.085 13.690 20.160 13.900 ;
        RECT 20.085 12.340 20.160 12.550 ;
        RECT 20.085 10.990 20.160 11.200 ;
        RECT 20.085 9.640 20.160 9.850 ;
        RECT 20.085 8.290 20.160 8.500 ;
        RECT 20.085 6.940 20.160 7.150 ;
        RECT 20.085 5.590 20.160 5.800 ;
        RECT 20.085 4.240 20.160 4.450 ;
        RECT 20.085 2.890 20.160 3.100 ;
        RECT 20.085 1.540 20.160 1.750 ;
        RECT 20.085 0.190 20.160 0.400 ;
    END
  END RBL0_6
  PIN RBL1_7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 20.300 20.440 20.375 20.650 ;
        RECT 20.300 19.090 20.375 19.300 ;
        RECT 20.300 17.740 20.375 17.950 ;
        RECT 20.300 16.390 20.375 16.600 ;
        RECT 20.300 15.040 20.375 15.250 ;
        RECT 20.300 13.690 20.375 13.900 ;
        RECT 20.300 12.340 20.375 12.550 ;
        RECT 20.300 10.990 20.375 11.200 ;
        RECT 20.300 9.640 20.375 9.850 ;
        RECT 20.300 8.290 20.375 8.500 ;
        RECT 20.300 6.940 20.375 7.150 ;
        RECT 20.300 5.590 20.375 5.800 ;
        RECT 20.300 4.240 20.375 4.450 ;
        RECT 20.300 2.890 20.375 3.100 ;
        RECT 20.300 1.540 20.375 1.750 ;
        RECT 20.300 0.190 20.375 0.400 ;
    END
  END RBL1_7
  PIN RBL0_7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 22.985 20.440 23.060 20.650 ;
        RECT 22.985 19.090 23.060 19.300 ;
        RECT 22.985 17.740 23.060 17.950 ;
        RECT 22.985 16.390 23.060 16.600 ;
        RECT 22.985 15.040 23.060 15.250 ;
        RECT 22.985 13.690 23.060 13.900 ;
        RECT 22.985 12.340 23.060 12.550 ;
        RECT 22.985 10.990 23.060 11.200 ;
        RECT 22.985 9.640 23.060 9.850 ;
        RECT 22.985 8.290 23.060 8.500 ;
        RECT 22.985 6.940 23.060 7.150 ;
        RECT 22.985 5.590 23.060 5.800 ;
        RECT 22.985 4.240 23.060 4.450 ;
        RECT 22.985 2.890 23.060 3.100 ;
        RECT 22.985 1.540 23.060 1.750 ;
        RECT 22.985 0.190 23.060 0.400 ;
    END
  END RBL0_7
  PIN WBL_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.386800 ;
    PORT
      LAYER li1 ;
        RECT 2.320 21.170 2.395 21.315 ;
        RECT 2.320 19.820 2.395 19.965 ;
        RECT 2.320 18.470 2.395 18.615 ;
        RECT 2.320 17.120 2.395 17.265 ;
        RECT 2.320 15.770 2.395 15.915 ;
        RECT 2.320 14.420 2.395 14.565 ;
        RECT 2.320 13.070 2.395 13.215 ;
        RECT 2.320 11.720 2.395 11.865 ;
        RECT 2.320 10.370 2.395 10.515 ;
        RECT 2.320 9.020 2.395 9.165 ;
        RECT 2.320 7.670 2.395 7.815 ;
        RECT 2.320 6.320 2.395 6.465 ;
        RECT 2.320 4.970 2.395 5.115 ;
        RECT 2.320 3.620 2.395 3.765 ;
        RECT 2.320 2.270 2.395 2.415 ;
        RECT 2.320 0.920 2.395 1.065 ;
    END
  END WBL_0
  PIN WBLb_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.369600 ;
    PORT
      LAYER li1 ;
        RECT 0.370 21.170 0.445 21.310 ;
        RECT 0.370 19.820 0.445 19.960 ;
        RECT 0.370 18.470 0.445 18.610 ;
        RECT 0.370 17.120 0.445 17.260 ;
        RECT 0.370 15.770 0.445 15.910 ;
        RECT 0.370 14.420 0.445 14.560 ;
        RECT 0.370 13.070 0.445 13.210 ;
        RECT 0.370 11.720 0.445 11.860 ;
        RECT 0.370 10.370 0.445 10.510 ;
        RECT 0.370 9.020 0.445 9.160 ;
        RECT 0.370 7.670 0.445 7.810 ;
        RECT 0.370 6.320 0.445 6.460 ;
        RECT 0.370 4.970 0.445 5.110 ;
        RECT 0.370 3.620 0.445 3.760 ;
        RECT 0.370 2.270 0.445 2.410 ;
        RECT 0.370 0.920 0.445 1.060 ;
    END
  END WBLb_0
  PIN WBL_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.386800 ;
    PORT
      LAYER li1 ;
        RECT 5.220 21.170 5.295 21.315 ;
        RECT 5.220 19.820 5.295 19.965 ;
        RECT 5.220 18.470 5.295 18.615 ;
        RECT 5.220 17.120 5.295 17.265 ;
        RECT 5.220 15.770 5.295 15.915 ;
        RECT 5.220 14.420 5.295 14.565 ;
        RECT 5.220 13.070 5.295 13.215 ;
        RECT 5.220 11.720 5.295 11.865 ;
        RECT 5.220 10.370 5.295 10.515 ;
        RECT 5.220 9.020 5.295 9.165 ;
        RECT 5.220 7.670 5.295 7.815 ;
        RECT 5.220 6.320 5.295 6.465 ;
        RECT 5.220 4.970 5.295 5.115 ;
        RECT 5.220 3.620 5.295 3.765 ;
        RECT 5.220 2.270 5.295 2.415 ;
        RECT 5.220 0.920 5.295 1.065 ;
    END
  END WBL_1
  PIN WBLb_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.369600 ;
    PORT
      LAYER li1 ;
        RECT 3.270 21.170 3.345 21.310 ;
        RECT 3.270 19.820 3.345 19.960 ;
        RECT 3.270 18.470 3.345 18.610 ;
        RECT 3.270 17.120 3.345 17.260 ;
        RECT 3.270 15.770 3.345 15.910 ;
        RECT 3.270 14.420 3.345 14.560 ;
        RECT 3.270 13.070 3.345 13.210 ;
        RECT 3.270 11.720 3.345 11.860 ;
        RECT 3.270 10.370 3.345 10.510 ;
        RECT 3.270 9.020 3.345 9.160 ;
        RECT 3.270 7.670 3.345 7.810 ;
        RECT 3.270 6.320 3.345 6.460 ;
        RECT 3.270 4.970 3.345 5.110 ;
        RECT 3.270 3.620 3.345 3.760 ;
        RECT 3.270 2.270 3.345 2.410 ;
        RECT 3.270 0.920 3.345 1.060 ;
    END
  END WBLb_1
  PIN WBL_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.386800 ;
    PORT
      LAYER li1 ;
        RECT 8.120 21.170 8.195 21.315 ;
        RECT 8.120 19.820 8.195 19.965 ;
        RECT 8.120 18.470 8.195 18.615 ;
        RECT 8.120 17.120 8.195 17.265 ;
        RECT 8.120 15.770 8.195 15.915 ;
        RECT 8.120 14.420 8.195 14.565 ;
        RECT 8.120 13.070 8.195 13.215 ;
        RECT 8.120 11.720 8.195 11.865 ;
        RECT 8.120 10.370 8.195 10.515 ;
        RECT 8.120 9.020 8.195 9.165 ;
        RECT 8.120 7.670 8.195 7.815 ;
        RECT 8.120 6.320 8.195 6.465 ;
        RECT 8.120 4.970 8.195 5.115 ;
        RECT 8.120 3.620 8.195 3.765 ;
        RECT 8.120 2.270 8.195 2.415 ;
        RECT 8.120 0.920 8.195 1.065 ;
    END
  END WBL_2
  PIN WBLb_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.369600 ;
    PORT
      LAYER li1 ;
        RECT 6.170 21.170 6.245 21.310 ;
        RECT 6.170 19.820 6.245 19.960 ;
        RECT 6.170 18.470 6.245 18.610 ;
        RECT 6.170 17.120 6.245 17.260 ;
        RECT 6.170 15.770 6.245 15.910 ;
        RECT 6.170 14.420 6.245 14.560 ;
        RECT 6.170 13.070 6.245 13.210 ;
        RECT 6.170 11.720 6.245 11.860 ;
        RECT 6.170 10.370 6.245 10.510 ;
        RECT 6.170 9.020 6.245 9.160 ;
        RECT 6.170 7.670 6.245 7.810 ;
        RECT 6.170 6.320 6.245 6.460 ;
        RECT 6.170 4.970 6.245 5.110 ;
        RECT 6.170 3.620 6.245 3.760 ;
        RECT 6.170 2.270 6.245 2.410 ;
        RECT 6.170 0.920 6.245 1.060 ;
    END
  END WBLb_2
  PIN WBL_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.386800 ;
    PORT
      LAYER li1 ;
        RECT 11.020 21.170 11.095 21.315 ;
        RECT 11.020 19.820 11.095 19.965 ;
        RECT 11.020 18.470 11.095 18.615 ;
        RECT 11.020 17.120 11.095 17.265 ;
        RECT 11.020 15.770 11.095 15.915 ;
        RECT 11.020 14.420 11.095 14.565 ;
        RECT 11.020 13.070 11.095 13.215 ;
        RECT 11.020 11.720 11.095 11.865 ;
        RECT 11.020 10.370 11.095 10.515 ;
        RECT 11.020 9.020 11.095 9.165 ;
        RECT 11.020 7.670 11.095 7.815 ;
        RECT 11.020 6.320 11.095 6.465 ;
        RECT 11.020 4.970 11.095 5.115 ;
        RECT 11.020 3.620 11.095 3.765 ;
        RECT 11.020 2.270 11.095 2.415 ;
        RECT 11.020 0.920 11.095 1.065 ;
    END
  END WBL_3
  PIN WBLb_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.369600 ;
    PORT
      LAYER li1 ;
        RECT 9.070 21.170 9.145 21.310 ;
        RECT 9.070 19.820 9.145 19.960 ;
        RECT 9.070 18.470 9.145 18.610 ;
        RECT 9.070 17.120 9.145 17.260 ;
        RECT 9.070 15.770 9.145 15.910 ;
        RECT 9.070 14.420 9.145 14.560 ;
        RECT 9.070 13.070 9.145 13.210 ;
        RECT 9.070 11.720 9.145 11.860 ;
        RECT 9.070 10.370 9.145 10.510 ;
        RECT 9.070 9.020 9.145 9.160 ;
        RECT 9.070 7.670 9.145 7.810 ;
        RECT 9.070 6.320 9.145 6.460 ;
        RECT 9.070 4.970 9.145 5.110 ;
        RECT 9.070 3.620 9.145 3.760 ;
        RECT 9.070 2.270 9.145 2.410 ;
        RECT 9.070 0.920 9.145 1.060 ;
    END
  END WBLb_3
  PIN WBL_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.386800 ;
    PORT
      LAYER li1 ;
        RECT 13.920 21.170 13.995 21.315 ;
        RECT 13.920 19.820 13.995 19.965 ;
        RECT 13.920 18.470 13.995 18.615 ;
        RECT 13.920 17.120 13.995 17.265 ;
        RECT 13.920 15.770 13.995 15.915 ;
        RECT 13.920 14.420 13.995 14.565 ;
        RECT 13.920 13.070 13.995 13.215 ;
        RECT 13.920 11.720 13.995 11.865 ;
        RECT 13.920 10.370 13.995 10.515 ;
        RECT 13.920 9.020 13.995 9.165 ;
        RECT 13.920 7.670 13.995 7.815 ;
        RECT 13.920 6.320 13.995 6.465 ;
        RECT 13.920 4.970 13.995 5.115 ;
        RECT 13.920 3.620 13.995 3.765 ;
        RECT 13.920 2.270 13.995 2.415 ;
        RECT 13.920 0.920 13.995 1.065 ;
    END
  END WBL_4
  PIN WBLb_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.369600 ;
    PORT
      LAYER li1 ;
        RECT 11.970 21.170 12.045 21.310 ;
        RECT 11.970 19.820 12.045 19.960 ;
        RECT 11.970 18.470 12.045 18.610 ;
        RECT 11.970 17.120 12.045 17.260 ;
        RECT 11.970 15.770 12.045 15.910 ;
        RECT 11.970 14.420 12.045 14.560 ;
        RECT 11.970 13.070 12.045 13.210 ;
        RECT 11.970 11.720 12.045 11.860 ;
        RECT 11.970 10.370 12.045 10.510 ;
        RECT 11.970 9.020 12.045 9.160 ;
        RECT 11.970 7.670 12.045 7.810 ;
        RECT 11.970 6.320 12.045 6.460 ;
        RECT 11.970 4.970 12.045 5.110 ;
        RECT 11.970 3.620 12.045 3.760 ;
        RECT 11.970 2.270 12.045 2.410 ;
        RECT 11.970 0.920 12.045 1.060 ;
    END
  END WBLb_4
  PIN WBL_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.386800 ;
    PORT
      LAYER li1 ;
        RECT 16.820 21.170 16.895 21.315 ;
        RECT 16.820 19.820 16.895 19.965 ;
        RECT 16.820 18.470 16.895 18.615 ;
        RECT 16.820 17.120 16.895 17.265 ;
        RECT 16.820 15.770 16.895 15.915 ;
        RECT 16.820 14.420 16.895 14.565 ;
        RECT 16.820 13.070 16.895 13.215 ;
        RECT 16.820 11.720 16.895 11.865 ;
        RECT 16.820 10.370 16.895 10.515 ;
        RECT 16.820 9.020 16.895 9.165 ;
        RECT 16.820 7.670 16.895 7.815 ;
        RECT 16.820 6.320 16.895 6.465 ;
        RECT 16.820 4.970 16.895 5.115 ;
        RECT 16.820 3.620 16.895 3.765 ;
        RECT 16.820 2.270 16.895 2.415 ;
        RECT 16.820 0.920 16.895 1.065 ;
    END
  END WBL_5
  PIN WBLb_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.369600 ;
    PORT
      LAYER li1 ;
        RECT 14.870 21.170 14.945 21.310 ;
        RECT 14.870 19.820 14.945 19.960 ;
        RECT 14.870 18.470 14.945 18.610 ;
        RECT 14.870 17.120 14.945 17.260 ;
        RECT 14.870 15.770 14.945 15.910 ;
        RECT 14.870 14.420 14.945 14.560 ;
        RECT 14.870 13.070 14.945 13.210 ;
        RECT 14.870 11.720 14.945 11.860 ;
        RECT 14.870 10.370 14.945 10.510 ;
        RECT 14.870 9.020 14.945 9.160 ;
        RECT 14.870 7.670 14.945 7.810 ;
        RECT 14.870 6.320 14.945 6.460 ;
        RECT 14.870 4.970 14.945 5.110 ;
        RECT 14.870 3.620 14.945 3.760 ;
        RECT 14.870 2.270 14.945 2.410 ;
        RECT 14.870 0.920 14.945 1.060 ;
    END
  END WBLb_5
  PIN WBL_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.386800 ;
    PORT
      LAYER li1 ;
        RECT 19.720 21.170 19.795 21.315 ;
        RECT 19.720 19.820 19.795 19.965 ;
        RECT 19.720 18.470 19.795 18.615 ;
        RECT 19.720 17.120 19.795 17.265 ;
        RECT 19.720 15.770 19.795 15.915 ;
        RECT 19.720 14.420 19.795 14.565 ;
        RECT 19.720 13.070 19.795 13.215 ;
        RECT 19.720 11.720 19.795 11.865 ;
        RECT 19.720 10.370 19.795 10.515 ;
        RECT 19.720 9.020 19.795 9.165 ;
        RECT 19.720 7.670 19.795 7.815 ;
        RECT 19.720 6.320 19.795 6.465 ;
        RECT 19.720 4.970 19.795 5.115 ;
        RECT 19.720 3.620 19.795 3.765 ;
        RECT 19.720 2.270 19.795 2.415 ;
        RECT 19.720 0.920 19.795 1.065 ;
    END
  END WBL_6
  PIN WBLb_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.369600 ;
    PORT
      LAYER li1 ;
        RECT 17.770 21.170 17.845 21.310 ;
        RECT 17.770 19.820 17.845 19.960 ;
        RECT 17.770 18.470 17.845 18.610 ;
        RECT 17.770 17.120 17.845 17.260 ;
        RECT 17.770 15.770 17.845 15.910 ;
        RECT 17.770 14.420 17.845 14.560 ;
        RECT 17.770 13.070 17.845 13.210 ;
        RECT 17.770 11.720 17.845 11.860 ;
        RECT 17.770 10.370 17.845 10.510 ;
        RECT 17.770 9.020 17.845 9.160 ;
        RECT 17.770 7.670 17.845 7.810 ;
        RECT 17.770 6.320 17.845 6.460 ;
        RECT 17.770 4.970 17.845 5.110 ;
        RECT 17.770 3.620 17.845 3.760 ;
        RECT 17.770 2.270 17.845 2.410 ;
        RECT 17.770 0.920 17.845 1.060 ;
    END
  END WBLb_6
  PIN WBL_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.386800 ;
    PORT
      LAYER li1 ;
        RECT 22.620 21.170 22.695 21.315 ;
        RECT 22.620 19.820 22.695 19.965 ;
        RECT 22.620 18.470 22.695 18.615 ;
        RECT 22.620 17.120 22.695 17.265 ;
        RECT 22.620 15.770 22.695 15.915 ;
        RECT 22.620 14.420 22.695 14.565 ;
        RECT 22.620 13.070 22.695 13.215 ;
        RECT 22.620 11.720 22.695 11.865 ;
        RECT 22.620 10.370 22.695 10.515 ;
        RECT 22.620 9.020 22.695 9.165 ;
        RECT 22.620 7.670 22.695 7.815 ;
        RECT 22.620 6.320 22.695 6.465 ;
        RECT 22.620 4.970 22.695 5.115 ;
        RECT 22.620 3.620 22.695 3.765 ;
        RECT 22.620 2.270 22.695 2.415 ;
        RECT 22.620 0.920 22.695 1.065 ;
    END
  END WBL_7
  PIN WBLb_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.369600 ;
    PORT
      LAYER li1 ;
        RECT 20.670 21.170 20.745 21.310 ;
        RECT 20.670 19.820 20.745 19.960 ;
        RECT 20.670 18.470 20.745 18.610 ;
        RECT 20.670 17.120 20.745 17.260 ;
        RECT 20.670 15.770 20.745 15.910 ;
        RECT 20.670 14.420 20.745 14.560 ;
        RECT 20.670 13.070 20.745 13.210 ;
        RECT 20.670 11.720 20.745 11.860 ;
        RECT 20.670 10.370 20.745 10.510 ;
        RECT 20.670 9.020 20.745 9.160 ;
        RECT 20.670 7.670 20.745 7.810 ;
        RECT 20.670 6.320 20.745 6.460 ;
        RECT 20.670 4.970 20.745 5.110 ;
        RECT 20.670 3.620 20.745 3.760 ;
        RECT 20.670 2.270 20.745 2.410 ;
        RECT 20.670 0.920 20.745 1.060 ;
    END
  END WBLb_7
  PIN RWL_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.504000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 20.760 0.365 20.930 ;
        RECT 2.395 20.760 2.545 20.930 ;
        RECT 3.115 20.760 3.265 20.930 ;
        RECT 5.295 20.760 5.445 20.930 ;
        RECT 6.015 20.760 6.165 20.930 ;
        RECT 8.195 20.760 8.345 20.930 ;
        RECT 8.915 20.760 9.065 20.930 ;
        RECT 11.095 20.760 11.245 20.930 ;
        RECT 11.815 20.760 11.965 20.930 ;
        RECT 13.995 20.760 14.145 20.930 ;
        RECT 14.715 20.760 14.865 20.930 ;
        RECT 16.895 20.760 17.045 20.930 ;
        RECT 17.615 20.760 17.765 20.930 ;
        RECT 19.795 20.760 19.945 20.930 ;
        RECT 20.515 20.760 20.665 20.930 ;
        RECT 22.695 20.760 22.845 20.930 ;
      LAYER met1 ;
        RECT 0.000 20.760 22.845 20.930 ;
    END
  END RWL_0
  PIN RWL_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.504000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 19.410 0.365 19.580 ;
        RECT 2.395 19.410 2.545 19.580 ;
        RECT 3.115 19.410 3.265 19.580 ;
        RECT 5.295 19.410 5.445 19.580 ;
        RECT 6.015 19.410 6.165 19.580 ;
        RECT 8.195 19.410 8.345 19.580 ;
        RECT 8.915 19.410 9.065 19.580 ;
        RECT 11.095 19.410 11.245 19.580 ;
        RECT 11.815 19.410 11.965 19.580 ;
        RECT 13.995 19.410 14.145 19.580 ;
        RECT 14.715 19.410 14.865 19.580 ;
        RECT 16.895 19.410 17.045 19.580 ;
        RECT 17.615 19.410 17.765 19.580 ;
        RECT 19.795 19.410 19.945 19.580 ;
        RECT 20.515 19.410 20.665 19.580 ;
        RECT 22.695 19.410 22.845 19.580 ;
      LAYER met1 ;
        RECT 0.000 19.410 22.845 19.580 ;
    END
  END RWL_1
  PIN RWL_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.504000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 18.060 0.365 18.230 ;
        RECT 2.395 18.060 2.545 18.230 ;
        RECT 3.115 18.060 3.265 18.230 ;
        RECT 5.295 18.060 5.445 18.230 ;
        RECT 6.015 18.060 6.165 18.230 ;
        RECT 8.195 18.060 8.345 18.230 ;
        RECT 8.915 18.060 9.065 18.230 ;
        RECT 11.095 18.060 11.245 18.230 ;
        RECT 11.815 18.060 11.965 18.230 ;
        RECT 13.995 18.060 14.145 18.230 ;
        RECT 14.715 18.060 14.865 18.230 ;
        RECT 16.895 18.060 17.045 18.230 ;
        RECT 17.615 18.060 17.765 18.230 ;
        RECT 19.795 18.060 19.945 18.230 ;
        RECT 20.515 18.060 20.665 18.230 ;
        RECT 22.695 18.060 22.845 18.230 ;
      LAYER met1 ;
        RECT 0.000 18.060 22.845 18.230 ;
    END
  END RWL_2
  PIN RWL_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.504000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 16.710 0.365 16.880 ;
        RECT 2.395 16.710 2.545 16.880 ;
        RECT 3.115 16.710 3.265 16.880 ;
        RECT 5.295 16.710 5.445 16.880 ;
        RECT 6.015 16.710 6.165 16.880 ;
        RECT 8.195 16.710 8.345 16.880 ;
        RECT 8.915 16.710 9.065 16.880 ;
        RECT 11.095 16.710 11.245 16.880 ;
        RECT 11.815 16.710 11.965 16.880 ;
        RECT 13.995 16.710 14.145 16.880 ;
        RECT 14.715 16.710 14.865 16.880 ;
        RECT 16.895 16.710 17.045 16.880 ;
        RECT 17.615 16.710 17.765 16.880 ;
        RECT 19.795 16.710 19.945 16.880 ;
        RECT 20.515 16.710 20.665 16.880 ;
        RECT 22.695 16.710 22.845 16.880 ;
      LAYER met1 ;
        RECT 0.000 16.710 22.845 16.880 ;
    END
  END RWL_3
  PIN RWL_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.504000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 15.360 0.365 15.530 ;
        RECT 2.395 15.360 2.545 15.530 ;
        RECT 3.115 15.360 3.265 15.530 ;
        RECT 5.295 15.360 5.445 15.530 ;
        RECT 6.015 15.360 6.165 15.530 ;
        RECT 8.195 15.360 8.345 15.530 ;
        RECT 8.915 15.360 9.065 15.530 ;
        RECT 11.095 15.360 11.245 15.530 ;
        RECT 11.815 15.360 11.965 15.530 ;
        RECT 13.995 15.360 14.145 15.530 ;
        RECT 14.715 15.360 14.865 15.530 ;
        RECT 16.895 15.360 17.045 15.530 ;
        RECT 17.615 15.360 17.765 15.530 ;
        RECT 19.795 15.360 19.945 15.530 ;
        RECT 20.515 15.360 20.665 15.530 ;
        RECT 22.695 15.360 22.845 15.530 ;
      LAYER met1 ;
        RECT 0.000 15.360 22.845 15.530 ;
    END
  END RWL_4
  PIN RWL_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.504000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 14.010 0.365 14.180 ;
        RECT 2.395 14.010 2.545 14.180 ;
        RECT 3.115 14.010 3.265 14.180 ;
        RECT 5.295 14.010 5.445 14.180 ;
        RECT 6.015 14.010 6.165 14.180 ;
        RECT 8.195 14.010 8.345 14.180 ;
        RECT 8.915 14.010 9.065 14.180 ;
        RECT 11.095 14.010 11.245 14.180 ;
        RECT 11.815 14.010 11.965 14.180 ;
        RECT 13.995 14.010 14.145 14.180 ;
        RECT 14.715 14.010 14.865 14.180 ;
        RECT 16.895 14.010 17.045 14.180 ;
        RECT 17.615 14.010 17.765 14.180 ;
        RECT 19.795 14.010 19.945 14.180 ;
        RECT 20.515 14.010 20.665 14.180 ;
        RECT 22.695 14.010 22.845 14.180 ;
      LAYER met1 ;
        RECT 0.000 14.010 22.845 14.180 ;
    END
  END RWL_5
  PIN RWL_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.504000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 12.660 0.365 12.830 ;
        RECT 2.395 12.660 2.545 12.830 ;
        RECT 3.115 12.660 3.265 12.830 ;
        RECT 5.295 12.660 5.445 12.830 ;
        RECT 6.015 12.660 6.165 12.830 ;
        RECT 8.195 12.660 8.345 12.830 ;
        RECT 8.915 12.660 9.065 12.830 ;
        RECT 11.095 12.660 11.245 12.830 ;
        RECT 11.815 12.660 11.965 12.830 ;
        RECT 13.995 12.660 14.145 12.830 ;
        RECT 14.715 12.660 14.865 12.830 ;
        RECT 16.895 12.660 17.045 12.830 ;
        RECT 17.615 12.660 17.765 12.830 ;
        RECT 19.795 12.660 19.945 12.830 ;
        RECT 20.515 12.660 20.665 12.830 ;
        RECT 22.695 12.660 22.845 12.830 ;
      LAYER met1 ;
        RECT 0.000 12.660 22.845 12.830 ;
    END
  END RWL_6
  PIN RWL_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.504000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 11.310 0.365 11.480 ;
        RECT 2.395 11.310 2.545 11.480 ;
        RECT 3.115 11.310 3.265 11.480 ;
        RECT 5.295 11.310 5.445 11.480 ;
        RECT 6.015 11.310 6.165 11.480 ;
        RECT 8.195 11.310 8.345 11.480 ;
        RECT 8.915 11.310 9.065 11.480 ;
        RECT 11.095 11.310 11.245 11.480 ;
        RECT 11.815 11.310 11.965 11.480 ;
        RECT 13.995 11.310 14.145 11.480 ;
        RECT 14.715 11.310 14.865 11.480 ;
        RECT 16.895 11.310 17.045 11.480 ;
        RECT 17.615 11.310 17.765 11.480 ;
        RECT 19.795 11.310 19.945 11.480 ;
        RECT 20.515 11.310 20.665 11.480 ;
        RECT 22.695 11.310 22.845 11.480 ;
      LAYER met1 ;
        RECT 0.000 11.310 22.845 11.480 ;
    END
  END RWL_7
  PIN RWL_8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.504000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 9.960 0.365 10.130 ;
        RECT 2.395 9.960 2.545 10.130 ;
        RECT 3.115 9.960 3.265 10.130 ;
        RECT 5.295 9.960 5.445 10.130 ;
        RECT 6.015 9.960 6.165 10.130 ;
        RECT 8.195 9.960 8.345 10.130 ;
        RECT 8.915 9.960 9.065 10.130 ;
        RECT 11.095 9.960 11.245 10.130 ;
        RECT 11.815 9.960 11.965 10.130 ;
        RECT 13.995 9.960 14.145 10.130 ;
        RECT 14.715 9.960 14.865 10.130 ;
        RECT 16.895 9.960 17.045 10.130 ;
        RECT 17.615 9.960 17.765 10.130 ;
        RECT 19.795 9.960 19.945 10.130 ;
        RECT 20.515 9.960 20.665 10.130 ;
        RECT 22.695 9.960 22.845 10.130 ;
      LAYER met1 ;
        RECT 0.000 9.960 22.845 10.130 ;
    END
  END RWL_8
  PIN RWL_9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.504000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 8.610 0.365 8.780 ;
        RECT 2.395 8.610 2.545 8.780 ;
        RECT 3.115 8.610 3.265 8.780 ;
        RECT 5.295 8.610 5.445 8.780 ;
        RECT 6.015 8.610 6.165 8.780 ;
        RECT 8.195 8.610 8.345 8.780 ;
        RECT 8.915 8.610 9.065 8.780 ;
        RECT 11.095 8.610 11.245 8.780 ;
        RECT 11.815 8.610 11.965 8.780 ;
        RECT 13.995 8.610 14.145 8.780 ;
        RECT 14.715 8.610 14.865 8.780 ;
        RECT 16.895 8.610 17.045 8.780 ;
        RECT 17.615 8.610 17.765 8.780 ;
        RECT 19.795 8.610 19.945 8.780 ;
        RECT 20.515 8.610 20.665 8.780 ;
        RECT 22.695 8.610 22.845 8.780 ;
      LAYER met1 ;
        RECT 0.000 8.610 22.845 8.780 ;
    END
  END RWL_9
  PIN RWL_10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.504000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 7.260 0.365 7.430 ;
        RECT 2.395 7.260 2.545 7.430 ;
        RECT 3.115 7.260 3.265 7.430 ;
        RECT 5.295 7.260 5.445 7.430 ;
        RECT 6.015 7.260 6.165 7.430 ;
        RECT 8.195 7.260 8.345 7.430 ;
        RECT 8.915 7.260 9.065 7.430 ;
        RECT 11.095 7.260 11.245 7.430 ;
        RECT 11.815 7.260 11.965 7.430 ;
        RECT 13.995 7.260 14.145 7.430 ;
        RECT 14.715 7.260 14.865 7.430 ;
        RECT 16.895 7.260 17.045 7.430 ;
        RECT 17.615 7.260 17.765 7.430 ;
        RECT 19.795 7.260 19.945 7.430 ;
        RECT 20.515 7.260 20.665 7.430 ;
        RECT 22.695 7.260 22.845 7.430 ;
      LAYER met1 ;
        RECT 0.000 7.260 22.845 7.430 ;
    END
  END RWL_10
  PIN RWL_11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.504000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 5.910 0.365 6.080 ;
        RECT 2.395 5.910 2.545 6.080 ;
        RECT 3.115 5.910 3.265 6.080 ;
        RECT 5.295 5.910 5.445 6.080 ;
        RECT 6.015 5.910 6.165 6.080 ;
        RECT 8.195 5.910 8.345 6.080 ;
        RECT 8.915 5.910 9.065 6.080 ;
        RECT 11.095 5.910 11.245 6.080 ;
        RECT 11.815 5.910 11.965 6.080 ;
        RECT 13.995 5.910 14.145 6.080 ;
        RECT 14.715 5.910 14.865 6.080 ;
        RECT 16.895 5.910 17.045 6.080 ;
        RECT 17.615 5.910 17.765 6.080 ;
        RECT 19.795 5.910 19.945 6.080 ;
        RECT 20.515 5.910 20.665 6.080 ;
        RECT 22.695 5.910 22.845 6.080 ;
      LAYER met1 ;
        RECT 0.000 5.910 22.845 6.080 ;
    END
  END RWL_11
  PIN RWL_12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.504000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 4.560 0.365 4.730 ;
        RECT 2.395 4.560 2.545 4.730 ;
        RECT 3.115 4.560 3.265 4.730 ;
        RECT 5.295 4.560 5.445 4.730 ;
        RECT 6.015 4.560 6.165 4.730 ;
        RECT 8.195 4.560 8.345 4.730 ;
        RECT 8.915 4.560 9.065 4.730 ;
        RECT 11.095 4.560 11.245 4.730 ;
        RECT 11.815 4.560 11.965 4.730 ;
        RECT 13.995 4.560 14.145 4.730 ;
        RECT 14.715 4.560 14.865 4.730 ;
        RECT 16.895 4.560 17.045 4.730 ;
        RECT 17.615 4.560 17.765 4.730 ;
        RECT 19.795 4.560 19.945 4.730 ;
        RECT 20.515 4.560 20.665 4.730 ;
        RECT 22.695 4.560 22.845 4.730 ;
      LAYER met1 ;
        RECT 0.000 4.560 22.845 4.730 ;
    END
  END RWL_12
  PIN RWL_13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.504000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 3.210 0.365 3.380 ;
        RECT 2.395 3.210 2.545 3.380 ;
        RECT 3.115 3.210 3.265 3.380 ;
        RECT 5.295 3.210 5.445 3.380 ;
        RECT 6.015 3.210 6.165 3.380 ;
        RECT 8.195 3.210 8.345 3.380 ;
        RECT 8.915 3.210 9.065 3.380 ;
        RECT 11.095 3.210 11.245 3.380 ;
        RECT 11.815 3.210 11.965 3.380 ;
        RECT 13.995 3.210 14.145 3.380 ;
        RECT 14.715 3.210 14.865 3.380 ;
        RECT 16.895 3.210 17.045 3.380 ;
        RECT 17.615 3.210 17.765 3.380 ;
        RECT 19.795 3.210 19.945 3.380 ;
        RECT 20.515 3.210 20.665 3.380 ;
        RECT 22.695 3.210 22.845 3.380 ;
      LAYER met1 ;
        RECT 0.000 3.210 22.845 3.380 ;
    END
  END RWL_13
  PIN RWL_14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.504000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 1.860 0.365 2.030 ;
        RECT 2.395 1.860 2.545 2.030 ;
        RECT 3.115 1.860 3.265 2.030 ;
        RECT 5.295 1.860 5.445 2.030 ;
        RECT 6.015 1.860 6.165 2.030 ;
        RECT 8.195 1.860 8.345 2.030 ;
        RECT 8.915 1.860 9.065 2.030 ;
        RECT 11.095 1.860 11.245 2.030 ;
        RECT 11.815 1.860 11.965 2.030 ;
        RECT 13.995 1.860 14.145 2.030 ;
        RECT 14.715 1.860 14.865 2.030 ;
        RECT 16.895 1.860 17.045 2.030 ;
        RECT 17.615 1.860 17.765 2.030 ;
        RECT 19.795 1.860 19.945 2.030 ;
        RECT 20.515 1.860 20.665 2.030 ;
        RECT 22.695 1.860 22.845 2.030 ;
      LAYER met1 ;
        RECT 0.000 1.860 22.845 2.030 ;
    END
  END RWL_14
  PIN RWL_15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.504000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 0.510 0.365 0.680 ;
        RECT 2.395 0.510 2.545 0.680 ;
        RECT 3.115 0.510 3.265 0.680 ;
        RECT 5.295 0.510 5.445 0.680 ;
        RECT 6.015 0.510 6.165 0.680 ;
        RECT 8.195 0.510 8.345 0.680 ;
        RECT 8.915 0.510 9.065 0.680 ;
        RECT 11.095 0.510 11.245 0.680 ;
        RECT 11.815 0.510 11.965 0.680 ;
        RECT 13.995 0.510 14.145 0.680 ;
        RECT 14.715 0.510 14.865 0.680 ;
        RECT 16.895 0.510 17.045 0.680 ;
        RECT 17.615 0.510 17.765 0.680 ;
        RECT 19.795 0.510 19.945 0.680 ;
        RECT 20.515 0.510 20.665 0.680 ;
        RECT 22.695 0.510 22.845 0.680 ;
      LAYER met1 ;
        RECT 0.000 0.510 22.845 0.680 ;
    END
  END RWL_15
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER nwell ;
        RECT 0.990 20.970 1.755 21.450 ;
        RECT 3.890 20.970 4.655 21.450 ;
        RECT 6.790 20.970 7.555 21.450 ;
        RECT 9.690 20.970 10.455 21.450 ;
        RECT 12.590 20.970 13.355 21.450 ;
        RECT 15.490 20.970 16.255 21.450 ;
        RECT 18.390 20.970 19.155 21.450 ;
        RECT 21.290 20.970 22.055 21.450 ;
      LAYER li1 ;
        RECT 1.300 21.380 1.460 21.450 ;
        RECT 4.200 21.380 4.360 21.450 ;
        RECT 7.100 21.380 7.260 21.450 ;
        RECT 10.000 21.380 10.160 21.450 ;
        RECT 12.900 21.380 13.060 21.450 ;
        RECT 15.800 21.380 15.960 21.450 ;
        RECT 18.700 21.380 18.860 21.450 ;
        RECT 21.600 21.380 21.760 21.450 ;
        RECT 1.310 21.370 1.450 21.380 ;
        RECT 4.210 21.370 4.350 21.380 ;
        RECT 7.110 21.370 7.250 21.380 ;
        RECT 10.010 21.370 10.150 21.380 ;
        RECT 12.910 21.370 13.050 21.380 ;
        RECT 15.810 21.370 15.950 21.380 ;
        RECT 18.710 21.370 18.850 21.380 ;
        RECT 21.610 21.370 21.750 21.380 ;
      LAYER met1 ;
        RECT 0.000 21.380 23.060 21.450 ;
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER pwell ;
        RECT 0.000 20.740 0.850 21.600 ;
        RECT 1.910 20.740 3.750 21.600 ;
        RECT 4.810 20.740 6.650 21.600 ;
        RECT 7.710 20.740 9.550 21.600 ;
        RECT 10.610 20.740 12.450 21.600 ;
        RECT 13.510 20.740 15.350 21.600 ;
        RECT 16.410 20.740 18.250 21.600 ;
        RECT 19.310 20.740 21.150 21.600 ;
        RECT 22.210 20.740 23.060 21.600 ;
        RECT 0.000 20.250 23.060 20.740 ;
        RECT 0.000 19.390 0.850 20.250 ;
        RECT 1.910 19.390 3.750 20.250 ;
        RECT 4.810 19.390 6.650 20.250 ;
        RECT 7.710 19.390 9.550 20.250 ;
        RECT 10.610 19.390 12.450 20.250 ;
        RECT 13.510 19.390 15.350 20.250 ;
        RECT 16.410 19.390 18.250 20.250 ;
        RECT 19.310 19.390 21.150 20.250 ;
        RECT 22.210 19.390 23.060 20.250 ;
        RECT 0.000 18.900 23.060 19.390 ;
        RECT 0.000 18.040 0.850 18.900 ;
        RECT 1.910 18.040 3.750 18.900 ;
        RECT 4.810 18.040 6.650 18.900 ;
        RECT 7.710 18.040 9.550 18.900 ;
        RECT 10.610 18.040 12.450 18.900 ;
        RECT 13.510 18.040 15.350 18.900 ;
        RECT 16.410 18.040 18.250 18.900 ;
        RECT 19.310 18.040 21.150 18.900 ;
        RECT 22.210 18.040 23.060 18.900 ;
        RECT 0.000 17.550 23.060 18.040 ;
        RECT 0.000 16.690 0.850 17.550 ;
        RECT 1.910 16.690 3.750 17.550 ;
        RECT 4.810 16.690 6.650 17.550 ;
        RECT 7.710 16.690 9.550 17.550 ;
        RECT 10.610 16.690 12.450 17.550 ;
        RECT 13.510 16.690 15.350 17.550 ;
        RECT 16.410 16.690 18.250 17.550 ;
        RECT 19.310 16.690 21.150 17.550 ;
        RECT 22.210 16.690 23.060 17.550 ;
        RECT 0.000 16.200 23.060 16.690 ;
        RECT 0.000 15.340 0.850 16.200 ;
        RECT 1.910 15.340 3.750 16.200 ;
        RECT 4.810 15.340 6.650 16.200 ;
        RECT 7.710 15.340 9.550 16.200 ;
        RECT 10.610 15.340 12.450 16.200 ;
        RECT 13.510 15.340 15.350 16.200 ;
        RECT 16.410 15.340 18.250 16.200 ;
        RECT 19.310 15.340 21.150 16.200 ;
        RECT 22.210 15.340 23.060 16.200 ;
        RECT 0.000 14.850 23.060 15.340 ;
        RECT 0.000 13.990 0.850 14.850 ;
        RECT 1.910 13.990 3.750 14.850 ;
        RECT 4.810 13.990 6.650 14.850 ;
        RECT 7.710 13.990 9.550 14.850 ;
        RECT 10.610 13.990 12.450 14.850 ;
        RECT 13.510 13.990 15.350 14.850 ;
        RECT 16.410 13.990 18.250 14.850 ;
        RECT 19.310 13.990 21.150 14.850 ;
        RECT 22.210 13.990 23.060 14.850 ;
        RECT 0.000 13.500 23.060 13.990 ;
        RECT 0.000 12.640 0.850 13.500 ;
        RECT 1.910 12.640 3.750 13.500 ;
        RECT 4.810 12.640 6.650 13.500 ;
        RECT 7.710 12.640 9.550 13.500 ;
        RECT 10.610 12.640 12.450 13.500 ;
        RECT 13.510 12.640 15.350 13.500 ;
        RECT 16.410 12.640 18.250 13.500 ;
        RECT 19.310 12.640 21.150 13.500 ;
        RECT 22.210 12.640 23.060 13.500 ;
        RECT 0.000 12.150 23.060 12.640 ;
        RECT 0.000 11.290 0.850 12.150 ;
        RECT 1.910 11.290 3.750 12.150 ;
        RECT 4.810 11.290 6.650 12.150 ;
        RECT 7.710 11.290 9.550 12.150 ;
        RECT 10.610 11.290 12.450 12.150 ;
        RECT 13.510 11.290 15.350 12.150 ;
        RECT 16.410 11.290 18.250 12.150 ;
        RECT 19.310 11.290 21.150 12.150 ;
        RECT 22.210 11.290 23.060 12.150 ;
        RECT 0.000 10.800 23.060 11.290 ;
        RECT 0.000 9.940 0.850 10.800 ;
        RECT 1.910 9.940 3.750 10.800 ;
        RECT 4.810 9.940 6.650 10.800 ;
        RECT 7.710 9.940 9.550 10.800 ;
        RECT 10.610 9.940 12.450 10.800 ;
        RECT 13.510 9.940 15.350 10.800 ;
        RECT 16.410 9.940 18.250 10.800 ;
        RECT 19.310 9.940 21.150 10.800 ;
        RECT 22.210 9.940 23.060 10.800 ;
        RECT 0.000 9.450 23.060 9.940 ;
        RECT 0.000 8.590 0.850 9.450 ;
        RECT 1.910 8.590 3.750 9.450 ;
        RECT 4.810 8.590 6.650 9.450 ;
        RECT 7.710 8.590 9.550 9.450 ;
        RECT 10.610 8.590 12.450 9.450 ;
        RECT 13.510 8.590 15.350 9.450 ;
        RECT 16.410 8.590 18.250 9.450 ;
        RECT 19.310 8.590 21.150 9.450 ;
        RECT 22.210 8.590 23.060 9.450 ;
        RECT 0.000 8.100 23.060 8.590 ;
        RECT 0.000 7.240 0.850 8.100 ;
        RECT 1.910 7.240 3.750 8.100 ;
        RECT 4.810 7.240 6.650 8.100 ;
        RECT 7.710 7.240 9.550 8.100 ;
        RECT 10.610 7.240 12.450 8.100 ;
        RECT 13.510 7.240 15.350 8.100 ;
        RECT 16.410 7.240 18.250 8.100 ;
        RECT 19.310 7.240 21.150 8.100 ;
        RECT 22.210 7.240 23.060 8.100 ;
        RECT 0.000 6.750 23.060 7.240 ;
        RECT 0.000 5.890 0.850 6.750 ;
        RECT 1.910 5.890 3.750 6.750 ;
        RECT 4.810 5.890 6.650 6.750 ;
        RECT 7.710 5.890 9.550 6.750 ;
        RECT 10.610 5.890 12.450 6.750 ;
        RECT 13.510 5.890 15.350 6.750 ;
        RECT 16.410 5.890 18.250 6.750 ;
        RECT 19.310 5.890 21.150 6.750 ;
        RECT 22.210 5.890 23.060 6.750 ;
        RECT 0.000 5.400 23.060 5.890 ;
        RECT 0.000 4.540 0.850 5.400 ;
        RECT 1.910 4.540 3.750 5.400 ;
        RECT 4.810 4.540 6.650 5.400 ;
        RECT 7.710 4.540 9.550 5.400 ;
        RECT 10.610 4.540 12.450 5.400 ;
        RECT 13.510 4.540 15.350 5.400 ;
        RECT 16.410 4.540 18.250 5.400 ;
        RECT 19.310 4.540 21.150 5.400 ;
        RECT 22.210 4.540 23.060 5.400 ;
        RECT 0.000 4.050 23.060 4.540 ;
        RECT 0.000 3.190 0.850 4.050 ;
        RECT 1.910 3.190 3.750 4.050 ;
        RECT 4.810 3.190 6.650 4.050 ;
        RECT 7.710 3.190 9.550 4.050 ;
        RECT 10.610 3.190 12.450 4.050 ;
        RECT 13.510 3.190 15.350 4.050 ;
        RECT 16.410 3.190 18.250 4.050 ;
        RECT 19.310 3.190 21.150 4.050 ;
        RECT 22.210 3.190 23.060 4.050 ;
        RECT 0.000 2.700 23.060 3.190 ;
        RECT 0.000 1.840 0.850 2.700 ;
        RECT 1.910 1.840 3.750 2.700 ;
        RECT 4.810 1.840 6.650 2.700 ;
        RECT 7.710 1.840 9.550 2.700 ;
        RECT 10.610 1.840 12.450 2.700 ;
        RECT 13.510 1.840 15.350 2.700 ;
        RECT 16.410 1.840 18.250 2.700 ;
        RECT 19.310 1.840 21.150 2.700 ;
        RECT 22.210 1.840 23.060 2.700 ;
        RECT 0.000 1.350 23.060 1.840 ;
        RECT 0.000 0.490 0.850 1.350 ;
        RECT 1.910 0.490 3.750 1.350 ;
        RECT 4.810 0.490 6.650 1.350 ;
        RECT 7.710 0.490 9.550 1.350 ;
        RECT 10.610 0.490 12.450 1.350 ;
        RECT 13.510 0.490 15.350 1.350 ;
        RECT 16.410 0.490 18.250 1.350 ;
        RECT 19.310 0.490 21.150 1.350 ;
        RECT 22.210 0.490 23.060 1.350 ;
        RECT 0.000 0.000 23.060 0.490 ;
      LAYER li1 ;
        RECT 1.310 20.320 1.450 20.330 ;
        RECT 4.210 20.320 4.350 20.330 ;
        RECT 7.110 20.320 7.250 20.330 ;
        RECT 10.010 20.320 10.150 20.330 ;
        RECT 12.910 20.320 13.050 20.330 ;
        RECT 15.810 20.320 15.950 20.330 ;
        RECT 18.710 20.320 18.850 20.330 ;
        RECT 21.610 20.320 21.750 20.330 ;
        RECT 1.300 20.250 1.460 20.320 ;
        RECT 4.200 20.250 4.360 20.320 ;
        RECT 7.100 20.250 7.260 20.320 ;
        RECT 10.000 20.250 10.160 20.320 ;
        RECT 12.900 20.250 13.060 20.320 ;
        RECT 15.800 20.250 15.960 20.320 ;
        RECT 18.700 20.250 18.860 20.320 ;
        RECT 21.600 20.250 21.760 20.320 ;
        RECT 1.310 18.970 1.450 18.980 ;
        RECT 4.210 18.970 4.350 18.980 ;
        RECT 7.110 18.970 7.250 18.980 ;
        RECT 10.010 18.970 10.150 18.980 ;
        RECT 12.910 18.970 13.050 18.980 ;
        RECT 15.810 18.970 15.950 18.980 ;
        RECT 18.710 18.970 18.850 18.980 ;
        RECT 21.610 18.970 21.750 18.980 ;
        RECT 1.300 18.900 1.460 18.970 ;
        RECT 4.200 18.900 4.360 18.970 ;
        RECT 7.100 18.900 7.260 18.970 ;
        RECT 10.000 18.900 10.160 18.970 ;
        RECT 12.900 18.900 13.060 18.970 ;
        RECT 15.800 18.900 15.960 18.970 ;
        RECT 18.700 18.900 18.860 18.970 ;
        RECT 21.600 18.900 21.760 18.970 ;
        RECT 1.310 17.620 1.450 17.630 ;
        RECT 4.210 17.620 4.350 17.630 ;
        RECT 7.110 17.620 7.250 17.630 ;
        RECT 10.010 17.620 10.150 17.630 ;
        RECT 12.910 17.620 13.050 17.630 ;
        RECT 15.810 17.620 15.950 17.630 ;
        RECT 18.710 17.620 18.850 17.630 ;
        RECT 21.610 17.620 21.750 17.630 ;
        RECT 1.300 17.550 1.460 17.620 ;
        RECT 4.200 17.550 4.360 17.620 ;
        RECT 7.100 17.550 7.260 17.620 ;
        RECT 10.000 17.550 10.160 17.620 ;
        RECT 12.900 17.550 13.060 17.620 ;
        RECT 15.800 17.550 15.960 17.620 ;
        RECT 18.700 17.550 18.860 17.620 ;
        RECT 21.600 17.550 21.760 17.620 ;
        RECT 1.310 16.270 1.450 16.280 ;
        RECT 4.210 16.270 4.350 16.280 ;
        RECT 7.110 16.270 7.250 16.280 ;
        RECT 10.010 16.270 10.150 16.280 ;
        RECT 12.910 16.270 13.050 16.280 ;
        RECT 15.810 16.270 15.950 16.280 ;
        RECT 18.710 16.270 18.850 16.280 ;
        RECT 21.610 16.270 21.750 16.280 ;
        RECT 1.300 16.200 1.460 16.270 ;
        RECT 4.200 16.200 4.360 16.270 ;
        RECT 7.100 16.200 7.260 16.270 ;
        RECT 10.000 16.200 10.160 16.270 ;
        RECT 12.900 16.200 13.060 16.270 ;
        RECT 15.800 16.200 15.960 16.270 ;
        RECT 18.700 16.200 18.860 16.270 ;
        RECT 21.600 16.200 21.760 16.270 ;
        RECT 1.310 14.920 1.450 14.930 ;
        RECT 4.210 14.920 4.350 14.930 ;
        RECT 7.110 14.920 7.250 14.930 ;
        RECT 10.010 14.920 10.150 14.930 ;
        RECT 12.910 14.920 13.050 14.930 ;
        RECT 15.810 14.920 15.950 14.930 ;
        RECT 18.710 14.920 18.850 14.930 ;
        RECT 21.610 14.920 21.750 14.930 ;
        RECT 1.300 14.850 1.460 14.920 ;
        RECT 4.200 14.850 4.360 14.920 ;
        RECT 7.100 14.850 7.260 14.920 ;
        RECT 10.000 14.850 10.160 14.920 ;
        RECT 12.900 14.850 13.060 14.920 ;
        RECT 15.800 14.850 15.960 14.920 ;
        RECT 18.700 14.850 18.860 14.920 ;
        RECT 21.600 14.850 21.760 14.920 ;
        RECT 1.310 13.570 1.450 13.580 ;
        RECT 4.210 13.570 4.350 13.580 ;
        RECT 7.110 13.570 7.250 13.580 ;
        RECT 10.010 13.570 10.150 13.580 ;
        RECT 12.910 13.570 13.050 13.580 ;
        RECT 15.810 13.570 15.950 13.580 ;
        RECT 18.710 13.570 18.850 13.580 ;
        RECT 21.610 13.570 21.750 13.580 ;
        RECT 1.300 13.500 1.460 13.570 ;
        RECT 4.200 13.500 4.360 13.570 ;
        RECT 7.100 13.500 7.260 13.570 ;
        RECT 10.000 13.500 10.160 13.570 ;
        RECT 12.900 13.500 13.060 13.570 ;
        RECT 15.800 13.500 15.960 13.570 ;
        RECT 18.700 13.500 18.860 13.570 ;
        RECT 21.600 13.500 21.760 13.570 ;
        RECT 1.310 12.220 1.450 12.230 ;
        RECT 4.210 12.220 4.350 12.230 ;
        RECT 7.110 12.220 7.250 12.230 ;
        RECT 10.010 12.220 10.150 12.230 ;
        RECT 12.910 12.220 13.050 12.230 ;
        RECT 15.810 12.220 15.950 12.230 ;
        RECT 18.710 12.220 18.850 12.230 ;
        RECT 21.610 12.220 21.750 12.230 ;
        RECT 1.300 12.150 1.460 12.220 ;
        RECT 4.200 12.150 4.360 12.220 ;
        RECT 7.100 12.150 7.260 12.220 ;
        RECT 10.000 12.150 10.160 12.220 ;
        RECT 12.900 12.150 13.060 12.220 ;
        RECT 15.800 12.150 15.960 12.220 ;
        RECT 18.700 12.150 18.860 12.220 ;
        RECT 21.600 12.150 21.760 12.220 ;
        RECT 1.310 10.870 1.450 10.880 ;
        RECT 4.210 10.870 4.350 10.880 ;
        RECT 7.110 10.870 7.250 10.880 ;
        RECT 10.010 10.870 10.150 10.880 ;
        RECT 12.910 10.870 13.050 10.880 ;
        RECT 15.810 10.870 15.950 10.880 ;
        RECT 18.710 10.870 18.850 10.880 ;
        RECT 21.610 10.870 21.750 10.880 ;
        RECT 1.300 10.800 1.460 10.870 ;
        RECT 4.200 10.800 4.360 10.870 ;
        RECT 7.100 10.800 7.260 10.870 ;
        RECT 10.000 10.800 10.160 10.870 ;
        RECT 12.900 10.800 13.060 10.870 ;
        RECT 15.800 10.800 15.960 10.870 ;
        RECT 18.700 10.800 18.860 10.870 ;
        RECT 21.600 10.800 21.760 10.870 ;
        RECT 1.310 9.520 1.450 9.530 ;
        RECT 4.210 9.520 4.350 9.530 ;
        RECT 7.110 9.520 7.250 9.530 ;
        RECT 10.010 9.520 10.150 9.530 ;
        RECT 12.910 9.520 13.050 9.530 ;
        RECT 15.810 9.520 15.950 9.530 ;
        RECT 18.710 9.520 18.850 9.530 ;
        RECT 21.610 9.520 21.750 9.530 ;
        RECT 1.300 9.450 1.460 9.520 ;
        RECT 4.200 9.450 4.360 9.520 ;
        RECT 7.100 9.450 7.260 9.520 ;
        RECT 10.000 9.450 10.160 9.520 ;
        RECT 12.900 9.450 13.060 9.520 ;
        RECT 15.800 9.450 15.960 9.520 ;
        RECT 18.700 9.450 18.860 9.520 ;
        RECT 21.600 9.450 21.760 9.520 ;
        RECT 1.310 8.170 1.450 8.180 ;
        RECT 4.210 8.170 4.350 8.180 ;
        RECT 7.110 8.170 7.250 8.180 ;
        RECT 10.010 8.170 10.150 8.180 ;
        RECT 12.910 8.170 13.050 8.180 ;
        RECT 15.810 8.170 15.950 8.180 ;
        RECT 18.710 8.170 18.850 8.180 ;
        RECT 21.610 8.170 21.750 8.180 ;
        RECT 1.300 8.100 1.460 8.170 ;
        RECT 4.200 8.100 4.360 8.170 ;
        RECT 7.100 8.100 7.260 8.170 ;
        RECT 10.000 8.100 10.160 8.170 ;
        RECT 12.900 8.100 13.060 8.170 ;
        RECT 15.800 8.100 15.960 8.170 ;
        RECT 18.700 8.100 18.860 8.170 ;
        RECT 21.600 8.100 21.760 8.170 ;
        RECT 1.310 6.820 1.450 6.830 ;
        RECT 4.210 6.820 4.350 6.830 ;
        RECT 7.110 6.820 7.250 6.830 ;
        RECT 10.010 6.820 10.150 6.830 ;
        RECT 12.910 6.820 13.050 6.830 ;
        RECT 15.810 6.820 15.950 6.830 ;
        RECT 18.710 6.820 18.850 6.830 ;
        RECT 21.610 6.820 21.750 6.830 ;
        RECT 1.300 6.750 1.460 6.820 ;
        RECT 4.200 6.750 4.360 6.820 ;
        RECT 7.100 6.750 7.260 6.820 ;
        RECT 10.000 6.750 10.160 6.820 ;
        RECT 12.900 6.750 13.060 6.820 ;
        RECT 15.800 6.750 15.960 6.820 ;
        RECT 18.700 6.750 18.860 6.820 ;
        RECT 21.600 6.750 21.760 6.820 ;
        RECT 1.310 5.470 1.450 5.480 ;
        RECT 4.210 5.470 4.350 5.480 ;
        RECT 7.110 5.470 7.250 5.480 ;
        RECT 10.010 5.470 10.150 5.480 ;
        RECT 12.910 5.470 13.050 5.480 ;
        RECT 15.810 5.470 15.950 5.480 ;
        RECT 18.710 5.470 18.850 5.480 ;
        RECT 21.610 5.470 21.750 5.480 ;
        RECT 1.300 5.400 1.460 5.470 ;
        RECT 4.200 5.400 4.360 5.470 ;
        RECT 7.100 5.400 7.260 5.470 ;
        RECT 10.000 5.400 10.160 5.470 ;
        RECT 12.900 5.400 13.060 5.470 ;
        RECT 15.800 5.400 15.960 5.470 ;
        RECT 18.700 5.400 18.860 5.470 ;
        RECT 21.600 5.400 21.760 5.470 ;
        RECT 1.310 4.120 1.450 4.130 ;
        RECT 4.210 4.120 4.350 4.130 ;
        RECT 7.110 4.120 7.250 4.130 ;
        RECT 10.010 4.120 10.150 4.130 ;
        RECT 12.910 4.120 13.050 4.130 ;
        RECT 15.810 4.120 15.950 4.130 ;
        RECT 18.710 4.120 18.850 4.130 ;
        RECT 21.610 4.120 21.750 4.130 ;
        RECT 1.300 4.050 1.460 4.120 ;
        RECT 4.200 4.050 4.360 4.120 ;
        RECT 7.100 4.050 7.260 4.120 ;
        RECT 10.000 4.050 10.160 4.120 ;
        RECT 12.900 4.050 13.060 4.120 ;
        RECT 15.800 4.050 15.960 4.120 ;
        RECT 18.700 4.050 18.860 4.120 ;
        RECT 21.600 4.050 21.760 4.120 ;
        RECT 1.310 2.770 1.450 2.780 ;
        RECT 4.210 2.770 4.350 2.780 ;
        RECT 7.110 2.770 7.250 2.780 ;
        RECT 10.010 2.770 10.150 2.780 ;
        RECT 12.910 2.770 13.050 2.780 ;
        RECT 15.810 2.770 15.950 2.780 ;
        RECT 18.710 2.770 18.850 2.780 ;
        RECT 21.610 2.770 21.750 2.780 ;
        RECT 1.300 2.700 1.460 2.770 ;
        RECT 4.200 2.700 4.360 2.770 ;
        RECT 7.100 2.700 7.260 2.770 ;
        RECT 10.000 2.700 10.160 2.770 ;
        RECT 12.900 2.700 13.060 2.770 ;
        RECT 15.800 2.700 15.960 2.770 ;
        RECT 18.700 2.700 18.860 2.770 ;
        RECT 21.600 2.700 21.760 2.770 ;
        RECT 1.310 1.420 1.450 1.430 ;
        RECT 4.210 1.420 4.350 1.430 ;
        RECT 7.110 1.420 7.250 1.430 ;
        RECT 10.010 1.420 10.150 1.430 ;
        RECT 12.910 1.420 13.050 1.430 ;
        RECT 15.810 1.420 15.950 1.430 ;
        RECT 18.710 1.420 18.850 1.430 ;
        RECT 21.610 1.420 21.750 1.430 ;
        RECT 1.300 1.350 1.460 1.420 ;
        RECT 4.200 1.350 4.360 1.420 ;
        RECT 7.100 1.350 7.260 1.420 ;
        RECT 10.000 1.350 10.160 1.420 ;
        RECT 12.900 1.350 13.060 1.420 ;
        RECT 15.800 1.350 15.960 1.420 ;
        RECT 18.700 1.350 18.860 1.420 ;
        RECT 21.600 1.350 21.760 1.420 ;
        RECT 1.310 0.070 1.450 0.080 ;
        RECT 4.210 0.070 4.350 0.080 ;
        RECT 7.110 0.070 7.250 0.080 ;
        RECT 10.010 0.070 10.150 0.080 ;
        RECT 12.910 0.070 13.050 0.080 ;
        RECT 15.810 0.070 15.950 0.080 ;
        RECT 18.710 0.070 18.850 0.080 ;
        RECT 21.610 0.070 21.750 0.080 ;
        RECT 1.300 0.000 1.460 0.070 ;
        RECT 4.200 0.000 4.360 0.070 ;
        RECT 7.100 0.000 7.260 0.070 ;
        RECT 10.000 0.000 10.160 0.070 ;
        RECT 12.900 0.000 13.060 0.070 ;
        RECT 15.800 0.000 15.960 0.070 ;
        RECT 18.700 0.000 18.860 0.070 ;
        RECT 21.600 0.000 21.760 0.070 ;
      LAYER met1 ;
        RECT 0.000 20.250 23.060 20.320 ;
        RECT 0.000 18.900 23.060 18.970 ;
        RECT 0.000 17.550 23.060 17.620 ;
        RECT 0.000 16.200 23.060 16.270 ;
        RECT 0.000 14.850 23.060 14.920 ;
        RECT 0.000 13.500 23.060 13.570 ;
        RECT 0.000 12.150 23.060 12.220 ;
        RECT 0.000 10.800 23.060 10.870 ;
        RECT 0.000 9.450 23.060 9.520 ;
        RECT 0.000 8.100 23.060 8.170 ;
        RECT 0.000 6.750 23.060 6.820 ;
        RECT 0.000 5.400 23.060 5.470 ;
        RECT 0.000 4.050 23.060 4.120 ;
        RECT 0.000 2.700 23.060 2.770 ;
        RECT 0.000 1.350 23.060 1.420 ;
        RECT 0.000 0.000 23.060 0.070 ;
    END
  END GND
  OBS
      LAYER nwell ;
        RECT 0.990 19.620 1.755 20.100 ;
        RECT 3.890 19.620 4.655 20.100 ;
        RECT 6.790 19.620 7.555 20.100 ;
        RECT 9.690 19.620 10.455 20.100 ;
        RECT 12.590 19.620 13.355 20.100 ;
        RECT 15.490 19.620 16.255 20.100 ;
        RECT 18.390 19.620 19.155 20.100 ;
        RECT 21.290 19.620 22.055 20.100 ;
        RECT 0.990 18.270 1.755 18.750 ;
        RECT 3.890 18.270 4.655 18.750 ;
        RECT 6.790 18.270 7.555 18.750 ;
        RECT 9.690 18.270 10.455 18.750 ;
        RECT 12.590 18.270 13.355 18.750 ;
        RECT 15.490 18.270 16.255 18.750 ;
        RECT 18.390 18.270 19.155 18.750 ;
        RECT 21.290 18.270 22.055 18.750 ;
        RECT 0.990 16.920 1.755 17.400 ;
        RECT 3.890 16.920 4.655 17.400 ;
        RECT 6.790 16.920 7.555 17.400 ;
        RECT 9.690 16.920 10.455 17.400 ;
        RECT 12.590 16.920 13.355 17.400 ;
        RECT 15.490 16.920 16.255 17.400 ;
        RECT 18.390 16.920 19.155 17.400 ;
        RECT 21.290 16.920 22.055 17.400 ;
        RECT 0.990 15.570 1.755 16.050 ;
        RECT 3.890 15.570 4.655 16.050 ;
        RECT 6.790 15.570 7.555 16.050 ;
        RECT 9.690 15.570 10.455 16.050 ;
        RECT 12.590 15.570 13.355 16.050 ;
        RECT 15.490 15.570 16.255 16.050 ;
        RECT 18.390 15.570 19.155 16.050 ;
        RECT 21.290 15.570 22.055 16.050 ;
        RECT 0.990 14.220 1.755 14.700 ;
        RECT 3.890 14.220 4.655 14.700 ;
        RECT 6.790 14.220 7.555 14.700 ;
        RECT 9.690 14.220 10.455 14.700 ;
        RECT 12.590 14.220 13.355 14.700 ;
        RECT 15.490 14.220 16.255 14.700 ;
        RECT 18.390 14.220 19.155 14.700 ;
        RECT 21.290 14.220 22.055 14.700 ;
        RECT 0.990 12.870 1.755 13.350 ;
        RECT 3.890 12.870 4.655 13.350 ;
        RECT 6.790 12.870 7.555 13.350 ;
        RECT 9.690 12.870 10.455 13.350 ;
        RECT 12.590 12.870 13.355 13.350 ;
        RECT 15.490 12.870 16.255 13.350 ;
        RECT 18.390 12.870 19.155 13.350 ;
        RECT 21.290 12.870 22.055 13.350 ;
        RECT 0.990 11.520 1.755 12.000 ;
        RECT 3.890 11.520 4.655 12.000 ;
        RECT 6.790 11.520 7.555 12.000 ;
        RECT 9.690 11.520 10.455 12.000 ;
        RECT 12.590 11.520 13.355 12.000 ;
        RECT 15.490 11.520 16.255 12.000 ;
        RECT 18.390 11.520 19.155 12.000 ;
        RECT 21.290 11.520 22.055 12.000 ;
        RECT 0.990 10.170 1.755 10.650 ;
        RECT 3.890 10.170 4.655 10.650 ;
        RECT 6.790 10.170 7.555 10.650 ;
        RECT 9.690 10.170 10.455 10.650 ;
        RECT 12.590 10.170 13.355 10.650 ;
        RECT 15.490 10.170 16.255 10.650 ;
        RECT 18.390 10.170 19.155 10.650 ;
        RECT 21.290 10.170 22.055 10.650 ;
        RECT 0.990 8.820 1.755 9.300 ;
        RECT 3.890 8.820 4.655 9.300 ;
        RECT 6.790 8.820 7.555 9.300 ;
        RECT 9.690 8.820 10.455 9.300 ;
        RECT 12.590 8.820 13.355 9.300 ;
        RECT 15.490 8.820 16.255 9.300 ;
        RECT 18.390 8.820 19.155 9.300 ;
        RECT 21.290 8.820 22.055 9.300 ;
        RECT 0.990 7.470 1.755 7.950 ;
        RECT 3.890 7.470 4.655 7.950 ;
        RECT 6.790 7.470 7.555 7.950 ;
        RECT 9.690 7.470 10.455 7.950 ;
        RECT 12.590 7.470 13.355 7.950 ;
        RECT 15.490 7.470 16.255 7.950 ;
        RECT 18.390 7.470 19.155 7.950 ;
        RECT 21.290 7.470 22.055 7.950 ;
        RECT 0.990 6.120 1.755 6.600 ;
        RECT 3.890 6.120 4.655 6.600 ;
        RECT 6.790 6.120 7.555 6.600 ;
        RECT 9.690 6.120 10.455 6.600 ;
        RECT 12.590 6.120 13.355 6.600 ;
        RECT 15.490 6.120 16.255 6.600 ;
        RECT 18.390 6.120 19.155 6.600 ;
        RECT 21.290 6.120 22.055 6.600 ;
        RECT 0.990 4.770 1.755 5.250 ;
        RECT 3.890 4.770 4.655 5.250 ;
        RECT 6.790 4.770 7.555 5.250 ;
        RECT 9.690 4.770 10.455 5.250 ;
        RECT 12.590 4.770 13.355 5.250 ;
        RECT 15.490 4.770 16.255 5.250 ;
        RECT 18.390 4.770 19.155 5.250 ;
        RECT 21.290 4.770 22.055 5.250 ;
        RECT 0.990 3.420 1.755 3.900 ;
        RECT 3.890 3.420 4.655 3.900 ;
        RECT 6.790 3.420 7.555 3.900 ;
        RECT 9.690 3.420 10.455 3.900 ;
        RECT 12.590 3.420 13.355 3.900 ;
        RECT 15.490 3.420 16.255 3.900 ;
        RECT 18.390 3.420 19.155 3.900 ;
        RECT 21.290 3.420 22.055 3.900 ;
        RECT 0.990 2.070 1.755 2.550 ;
        RECT 3.890 2.070 4.655 2.550 ;
        RECT 6.790 2.070 7.555 2.550 ;
        RECT 9.690 2.070 10.455 2.550 ;
        RECT 12.590 2.070 13.355 2.550 ;
        RECT 15.490 2.070 16.255 2.550 ;
        RECT 18.390 2.070 19.155 2.550 ;
        RECT 21.290 2.070 22.055 2.550 ;
        RECT 0.990 0.720 1.755 1.200 ;
        RECT 3.890 0.720 4.655 1.200 ;
        RECT 6.790 0.720 7.555 1.200 ;
        RECT 9.690 0.720 10.455 1.200 ;
        RECT 12.590 0.720 13.355 1.200 ;
        RECT 15.490 0.720 16.255 1.200 ;
        RECT 18.390 0.720 19.155 1.200 ;
        RECT 21.290 0.720 22.055 1.200 ;
      LAYER li1 ;
        RECT 0.775 21.170 0.850 21.310 ;
        RECT 0.990 21.120 1.065 21.260 ;
        RECT 1.695 21.180 1.755 21.260 ;
        POLYGON 1.695 21.180 1.755 21.180 1.755 21.120 ;
        RECT 1.910 21.170 1.985 21.310 ;
        RECT 3.675 21.170 3.750 21.310 ;
        RECT 3.890 21.120 3.965 21.260 ;
        RECT 4.595 21.180 4.655 21.260 ;
        POLYGON 4.595 21.180 4.655 21.180 4.655 21.120 ;
        RECT 4.810 21.170 4.885 21.310 ;
        RECT 6.575 21.170 6.650 21.310 ;
        RECT 6.790 21.120 6.865 21.260 ;
        RECT 7.495 21.180 7.555 21.260 ;
        POLYGON 7.495 21.180 7.555 21.180 7.555 21.120 ;
        RECT 7.710 21.170 7.785 21.310 ;
        RECT 9.475 21.170 9.550 21.310 ;
        RECT 9.690 21.120 9.765 21.260 ;
        RECT 10.395 21.180 10.455 21.260 ;
        POLYGON 10.395 21.180 10.455 21.180 10.455 21.120 ;
        RECT 10.610 21.170 10.685 21.310 ;
        RECT 12.375 21.170 12.450 21.310 ;
        RECT 12.590 21.120 12.665 21.260 ;
        RECT 13.295 21.180 13.355 21.260 ;
        POLYGON 13.295 21.180 13.355 21.180 13.355 21.120 ;
        RECT 13.510 21.170 13.585 21.310 ;
        RECT 15.275 21.170 15.350 21.310 ;
        RECT 15.490 21.120 15.565 21.260 ;
        RECT 16.195 21.180 16.255 21.260 ;
        POLYGON 16.195 21.180 16.255 21.180 16.255 21.120 ;
        RECT 16.410 21.170 16.485 21.310 ;
        RECT 18.175 21.170 18.250 21.310 ;
        RECT 18.390 21.120 18.465 21.260 ;
        RECT 19.095 21.180 19.155 21.260 ;
        POLYGON 19.095 21.180 19.155 21.180 19.155 21.120 ;
        RECT 19.310 21.170 19.385 21.310 ;
        RECT 21.075 21.170 21.150 21.310 ;
        RECT 21.290 21.120 21.365 21.260 ;
        RECT 21.995 21.180 22.055 21.260 ;
        POLYGON 21.995 21.180 22.055 21.180 22.055 21.120 ;
        RECT 22.210 21.170 22.285 21.310 ;
        RECT 0.720 20.650 0.870 20.820 ;
        RECT 1.110 20.785 1.260 20.955 ;
        RECT 1.500 20.785 1.650 20.955 ;
        RECT 1.890 20.650 2.040 20.820 ;
        RECT 3.620 20.650 3.770 20.820 ;
        RECT 4.010 20.785 4.160 20.955 ;
        RECT 4.400 20.785 4.550 20.955 ;
        RECT 4.790 20.650 4.940 20.820 ;
        RECT 6.520 20.650 6.670 20.820 ;
        RECT 6.910 20.785 7.060 20.955 ;
        RECT 7.300 20.785 7.450 20.955 ;
        RECT 7.690 20.650 7.840 20.820 ;
        RECT 9.420 20.650 9.570 20.820 ;
        RECT 9.810 20.785 9.960 20.955 ;
        RECT 10.200 20.785 10.350 20.955 ;
        RECT 10.590 20.650 10.740 20.820 ;
        RECT 12.320 20.650 12.470 20.820 ;
        RECT 12.710 20.785 12.860 20.955 ;
        RECT 13.100 20.785 13.250 20.955 ;
        RECT 13.490 20.650 13.640 20.820 ;
        RECT 15.220 20.650 15.370 20.820 ;
        RECT 15.610 20.785 15.760 20.955 ;
        RECT 16.000 20.785 16.150 20.955 ;
        RECT 16.390 20.650 16.540 20.820 ;
        RECT 18.120 20.650 18.270 20.820 ;
        RECT 18.510 20.785 18.660 20.955 ;
        RECT 18.900 20.785 19.050 20.955 ;
        RECT 19.290 20.650 19.440 20.820 ;
        RECT 21.020 20.650 21.170 20.820 ;
        RECT 21.410 20.785 21.560 20.955 ;
        RECT 21.800 20.785 21.950 20.955 ;
        RECT 22.190 20.650 22.340 20.820 ;
        RECT 0.985 20.565 1.035 20.600 ;
        POLYGON 1.035 20.600 1.070 20.565 1.035 20.565 ;
        RECT 0.985 20.440 1.070 20.565 ;
        RECT 1.690 20.440 1.775 20.600 ;
        RECT 3.885 20.565 3.935 20.600 ;
        POLYGON 3.935 20.600 3.970 20.565 3.935 20.565 ;
        RECT 3.885 20.440 3.970 20.565 ;
        RECT 4.590 20.440 4.675 20.600 ;
        RECT 6.785 20.565 6.835 20.600 ;
        POLYGON 6.835 20.600 6.870 20.565 6.835 20.565 ;
        RECT 6.785 20.440 6.870 20.565 ;
        RECT 7.490 20.440 7.575 20.600 ;
        RECT 9.685 20.565 9.735 20.600 ;
        POLYGON 9.735 20.600 9.770 20.565 9.735 20.565 ;
        RECT 9.685 20.440 9.770 20.565 ;
        RECT 10.390 20.440 10.475 20.600 ;
        RECT 12.585 20.565 12.635 20.600 ;
        POLYGON 12.635 20.600 12.670 20.565 12.635 20.565 ;
        RECT 12.585 20.440 12.670 20.565 ;
        RECT 13.290 20.440 13.375 20.600 ;
        RECT 15.485 20.565 15.535 20.600 ;
        POLYGON 15.535 20.600 15.570 20.565 15.535 20.565 ;
        RECT 15.485 20.440 15.570 20.565 ;
        RECT 16.190 20.440 16.275 20.600 ;
        RECT 18.385 20.565 18.435 20.600 ;
        POLYGON 18.435 20.600 18.470 20.565 18.435 20.565 ;
        RECT 18.385 20.440 18.470 20.565 ;
        RECT 19.090 20.440 19.175 20.600 ;
        RECT 21.285 20.565 21.335 20.600 ;
        POLYGON 21.335 20.600 21.370 20.565 21.335 20.565 ;
        RECT 21.285 20.440 21.370 20.565 ;
        RECT 21.990 20.440 22.075 20.600 ;
        RECT 1.300 20.030 1.460 20.100 ;
        RECT 4.200 20.030 4.360 20.100 ;
        RECT 7.100 20.030 7.260 20.100 ;
        RECT 10.000 20.030 10.160 20.100 ;
        RECT 12.900 20.030 13.060 20.100 ;
        RECT 15.800 20.030 15.960 20.100 ;
        RECT 18.700 20.030 18.860 20.100 ;
        RECT 21.600 20.030 21.760 20.100 ;
        RECT 1.310 20.020 1.450 20.030 ;
        RECT 4.210 20.020 4.350 20.030 ;
        RECT 7.110 20.020 7.250 20.030 ;
        RECT 10.010 20.020 10.150 20.030 ;
        RECT 12.910 20.020 13.050 20.030 ;
        RECT 15.810 20.020 15.950 20.030 ;
        RECT 18.710 20.020 18.850 20.030 ;
        RECT 21.610 20.020 21.750 20.030 ;
        RECT 0.775 19.820 0.850 19.960 ;
        RECT 0.990 19.770 1.065 19.910 ;
        RECT 1.695 19.830 1.755 19.910 ;
        POLYGON 1.695 19.830 1.755 19.830 1.755 19.770 ;
        RECT 1.910 19.820 1.985 19.960 ;
        RECT 3.675 19.820 3.750 19.960 ;
        RECT 3.890 19.770 3.965 19.910 ;
        RECT 4.595 19.830 4.655 19.910 ;
        POLYGON 4.595 19.830 4.655 19.830 4.655 19.770 ;
        RECT 4.810 19.820 4.885 19.960 ;
        RECT 6.575 19.820 6.650 19.960 ;
        RECT 6.790 19.770 6.865 19.910 ;
        RECT 7.495 19.830 7.555 19.910 ;
        POLYGON 7.495 19.830 7.555 19.830 7.555 19.770 ;
        RECT 7.710 19.820 7.785 19.960 ;
        RECT 9.475 19.820 9.550 19.960 ;
        RECT 9.690 19.770 9.765 19.910 ;
        RECT 10.395 19.830 10.455 19.910 ;
        POLYGON 10.395 19.830 10.455 19.830 10.455 19.770 ;
        RECT 10.610 19.820 10.685 19.960 ;
        RECT 12.375 19.820 12.450 19.960 ;
        RECT 12.590 19.770 12.665 19.910 ;
        RECT 13.295 19.830 13.355 19.910 ;
        POLYGON 13.295 19.830 13.355 19.830 13.355 19.770 ;
        RECT 13.510 19.820 13.585 19.960 ;
        RECT 15.275 19.820 15.350 19.960 ;
        RECT 15.490 19.770 15.565 19.910 ;
        RECT 16.195 19.830 16.255 19.910 ;
        POLYGON 16.195 19.830 16.255 19.830 16.255 19.770 ;
        RECT 16.410 19.820 16.485 19.960 ;
        RECT 18.175 19.820 18.250 19.960 ;
        RECT 18.390 19.770 18.465 19.910 ;
        RECT 19.095 19.830 19.155 19.910 ;
        POLYGON 19.095 19.830 19.155 19.830 19.155 19.770 ;
        RECT 19.310 19.820 19.385 19.960 ;
        RECT 21.075 19.820 21.150 19.960 ;
        RECT 21.290 19.770 21.365 19.910 ;
        RECT 21.995 19.830 22.055 19.910 ;
        POLYGON 21.995 19.830 22.055 19.830 22.055 19.770 ;
        RECT 22.210 19.820 22.285 19.960 ;
        RECT 0.720 19.300 0.870 19.470 ;
        RECT 1.110 19.435 1.260 19.605 ;
        RECT 1.500 19.435 1.650 19.605 ;
        RECT 1.890 19.300 2.040 19.470 ;
        RECT 3.620 19.300 3.770 19.470 ;
        RECT 4.010 19.435 4.160 19.605 ;
        RECT 4.400 19.435 4.550 19.605 ;
        RECT 4.790 19.300 4.940 19.470 ;
        RECT 6.520 19.300 6.670 19.470 ;
        RECT 6.910 19.435 7.060 19.605 ;
        RECT 7.300 19.435 7.450 19.605 ;
        RECT 7.690 19.300 7.840 19.470 ;
        RECT 9.420 19.300 9.570 19.470 ;
        RECT 9.810 19.435 9.960 19.605 ;
        RECT 10.200 19.435 10.350 19.605 ;
        RECT 10.590 19.300 10.740 19.470 ;
        RECT 12.320 19.300 12.470 19.470 ;
        RECT 12.710 19.435 12.860 19.605 ;
        RECT 13.100 19.435 13.250 19.605 ;
        RECT 13.490 19.300 13.640 19.470 ;
        RECT 15.220 19.300 15.370 19.470 ;
        RECT 15.610 19.435 15.760 19.605 ;
        RECT 16.000 19.435 16.150 19.605 ;
        RECT 16.390 19.300 16.540 19.470 ;
        RECT 18.120 19.300 18.270 19.470 ;
        RECT 18.510 19.435 18.660 19.605 ;
        RECT 18.900 19.435 19.050 19.605 ;
        RECT 19.290 19.300 19.440 19.470 ;
        RECT 21.020 19.300 21.170 19.470 ;
        RECT 21.410 19.435 21.560 19.605 ;
        RECT 21.800 19.435 21.950 19.605 ;
        RECT 22.190 19.300 22.340 19.470 ;
        RECT 0.985 19.215 1.035 19.250 ;
        POLYGON 1.035 19.250 1.070 19.215 1.035 19.215 ;
        RECT 0.985 19.090 1.070 19.215 ;
        RECT 1.690 19.090 1.775 19.250 ;
        RECT 3.885 19.215 3.935 19.250 ;
        POLYGON 3.935 19.250 3.970 19.215 3.935 19.215 ;
        RECT 3.885 19.090 3.970 19.215 ;
        RECT 4.590 19.090 4.675 19.250 ;
        RECT 6.785 19.215 6.835 19.250 ;
        POLYGON 6.835 19.250 6.870 19.215 6.835 19.215 ;
        RECT 6.785 19.090 6.870 19.215 ;
        RECT 7.490 19.090 7.575 19.250 ;
        RECT 9.685 19.215 9.735 19.250 ;
        POLYGON 9.735 19.250 9.770 19.215 9.735 19.215 ;
        RECT 9.685 19.090 9.770 19.215 ;
        RECT 10.390 19.090 10.475 19.250 ;
        RECT 12.585 19.215 12.635 19.250 ;
        POLYGON 12.635 19.250 12.670 19.215 12.635 19.215 ;
        RECT 12.585 19.090 12.670 19.215 ;
        RECT 13.290 19.090 13.375 19.250 ;
        RECT 15.485 19.215 15.535 19.250 ;
        POLYGON 15.535 19.250 15.570 19.215 15.535 19.215 ;
        RECT 15.485 19.090 15.570 19.215 ;
        RECT 16.190 19.090 16.275 19.250 ;
        RECT 18.385 19.215 18.435 19.250 ;
        POLYGON 18.435 19.250 18.470 19.215 18.435 19.215 ;
        RECT 18.385 19.090 18.470 19.215 ;
        RECT 19.090 19.090 19.175 19.250 ;
        RECT 21.285 19.215 21.335 19.250 ;
        POLYGON 21.335 19.250 21.370 19.215 21.335 19.215 ;
        RECT 21.285 19.090 21.370 19.215 ;
        RECT 21.990 19.090 22.075 19.250 ;
        RECT 1.300 18.680 1.460 18.750 ;
        RECT 4.200 18.680 4.360 18.750 ;
        RECT 7.100 18.680 7.260 18.750 ;
        RECT 10.000 18.680 10.160 18.750 ;
        RECT 12.900 18.680 13.060 18.750 ;
        RECT 15.800 18.680 15.960 18.750 ;
        RECT 18.700 18.680 18.860 18.750 ;
        RECT 21.600 18.680 21.760 18.750 ;
        RECT 1.310 18.670 1.450 18.680 ;
        RECT 4.210 18.670 4.350 18.680 ;
        RECT 7.110 18.670 7.250 18.680 ;
        RECT 10.010 18.670 10.150 18.680 ;
        RECT 12.910 18.670 13.050 18.680 ;
        RECT 15.810 18.670 15.950 18.680 ;
        RECT 18.710 18.670 18.850 18.680 ;
        RECT 21.610 18.670 21.750 18.680 ;
        RECT 0.775 18.470 0.850 18.610 ;
        RECT 0.990 18.420 1.065 18.560 ;
        RECT 1.695 18.480 1.755 18.560 ;
        POLYGON 1.695 18.480 1.755 18.480 1.755 18.420 ;
        RECT 1.910 18.470 1.985 18.610 ;
        RECT 3.675 18.470 3.750 18.610 ;
        RECT 3.890 18.420 3.965 18.560 ;
        RECT 4.595 18.480 4.655 18.560 ;
        POLYGON 4.595 18.480 4.655 18.480 4.655 18.420 ;
        RECT 4.810 18.470 4.885 18.610 ;
        RECT 6.575 18.470 6.650 18.610 ;
        RECT 6.790 18.420 6.865 18.560 ;
        RECT 7.495 18.480 7.555 18.560 ;
        POLYGON 7.495 18.480 7.555 18.480 7.555 18.420 ;
        RECT 7.710 18.470 7.785 18.610 ;
        RECT 9.475 18.470 9.550 18.610 ;
        RECT 9.690 18.420 9.765 18.560 ;
        RECT 10.395 18.480 10.455 18.560 ;
        POLYGON 10.395 18.480 10.455 18.480 10.455 18.420 ;
        RECT 10.610 18.470 10.685 18.610 ;
        RECT 12.375 18.470 12.450 18.610 ;
        RECT 12.590 18.420 12.665 18.560 ;
        RECT 13.295 18.480 13.355 18.560 ;
        POLYGON 13.295 18.480 13.355 18.480 13.355 18.420 ;
        RECT 13.510 18.470 13.585 18.610 ;
        RECT 15.275 18.470 15.350 18.610 ;
        RECT 15.490 18.420 15.565 18.560 ;
        RECT 16.195 18.480 16.255 18.560 ;
        POLYGON 16.195 18.480 16.255 18.480 16.255 18.420 ;
        RECT 16.410 18.470 16.485 18.610 ;
        RECT 18.175 18.470 18.250 18.610 ;
        RECT 18.390 18.420 18.465 18.560 ;
        RECT 19.095 18.480 19.155 18.560 ;
        POLYGON 19.095 18.480 19.155 18.480 19.155 18.420 ;
        RECT 19.310 18.470 19.385 18.610 ;
        RECT 21.075 18.470 21.150 18.610 ;
        RECT 21.290 18.420 21.365 18.560 ;
        RECT 21.995 18.480 22.055 18.560 ;
        POLYGON 21.995 18.480 22.055 18.480 22.055 18.420 ;
        RECT 22.210 18.470 22.285 18.610 ;
        RECT 0.720 17.950 0.870 18.120 ;
        RECT 1.110 18.085 1.260 18.255 ;
        RECT 1.500 18.085 1.650 18.255 ;
        RECT 1.890 17.950 2.040 18.120 ;
        RECT 3.620 17.950 3.770 18.120 ;
        RECT 4.010 18.085 4.160 18.255 ;
        RECT 4.400 18.085 4.550 18.255 ;
        RECT 4.790 17.950 4.940 18.120 ;
        RECT 6.520 17.950 6.670 18.120 ;
        RECT 6.910 18.085 7.060 18.255 ;
        RECT 7.300 18.085 7.450 18.255 ;
        RECT 7.690 17.950 7.840 18.120 ;
        RECT 9.420 17.950 9.570 18.120 ;
        RECT 9.810 18.085 9.960 18.255 ;
        RECT 10.200 18.085 10.350 18.255 ;
        RECT 10.590 17.950 10.740 18.120 ;
        RECT 12.320 17.950 12.470 18.120 ;
        RECT 12.710 18.085 12.860 18.255 ;
        RECT 13.100 18.085 13.250 18.255 ;
        RECT 13.490 17.950 13.640 18.120 ;
        RECT 15.220 17.950 15.370 18.120 ;
        RECT 15.610 18.085 15.760 18.255 ;
        RECT 16.000 18.085 16.150 18.255 ;
        RECT 16.390 17.950 16.540 18.120 ;
        RECT 18.120 17.950 18.270 18.120 ;
        RECT 18.510 18.085 18.660 18.255 ;
        RECT 18.900 18.085 19.050 18.255 ;
        RECT 19.290 17.950 19.440 18.120 ;
        RECT 21.020 17.950 21.170 18.120 ;
        RECT 21.410 18.085 21.560 18.255 ;
        RECT 21.800 18.085 21.950 18.255 ;
        RECT 22.190 17.950 22.340 18.120 ;
        RECT 0.985 17.865 1.035 17.900 ;
        POLYGON 1.035 17.900 1.070 17.865 1.035 17.865 ;
        RECT 0.985 17.740 1.070 17.865 ;
        RECT 1.690 17.740 1.775 17.900 ;
        RECT 3.885 17.865 3.935 17.900 ;
        POLYGON 3.935 17.900 3.970 17.865 3.935 17.865 ;
        RECT 3.885 17.740 3.970 17.865 ;
        RECT 4.590 17.740 4.675 17.900 ;
        RECT 6.785 17.865 6.835 17.900 ;
        POLYGON 6.835 17.900 6.870 17.865 6.835 17.865 ;
        RECT 6.785 17.740 6.870 17.865 ;
        RECT 7.490 17.740 7.575 17.900 ;
        RECT 9.685 17.865 9.735 17.900 ;
        POLYGON 9.735 17.900 9.770 17.865 9.735 17.865 ;
        RECT 9.685 17.740 9.770 17.865 ;
        RECT 10.390 17.740 10.475 17.900 ;
        RECT 12.585 17.865 12.635 17.900 ;
        POLYGON 12.635 17.900 12.670 17.865 12.635 17.865 ;
        RECT 12.585 17.740 12.670 17.865 ;
        RECT 13.290 17.740 13.375 17.900 ;
        RECT 15.485 17.865 15.535 17.900 ;
        POLYGON 15.535 17.900 15.570 17.865 15.535 17.865 ;
        RECT 15.485 17.740 15.570 17.865 ;
        RECT 16.190 17.740 16.275 17.900 ;
        RECT 18.385 17.865 18.435 17.900 ;
        POLYGON 18.435 17.900 18.470 17.865 18.435 17.865 ;
        RECT 18.385 17.740 18.470 17.865 ;
        RECT 19.090 17.740 19.175 17.900 ;
        RECT 21.285 17.865 21.335 17.900 ;
        POLYGON 21.335 17.900 21.370 17.865 21.335 17.865 ;
        RECT 21.285 17.740 21.370 17.865 ;
        RECT 21.990 17.740 22.075 17.900 ;
        RECT 1.300 17.330 1.460 17.400 ;
        RECT 4.200 17.330 4.360 17.400 ;
        RECT 7.100 17.330 7.260 17.400 ;
        RECT 10.000 17.330 10.160 17.400 ;
        RECT 12.900 17.330 13.060 17.400 ;
        RECT 15.800 17.330 15.960 17.400 ;
        RECT 18.700 17.330 18.860 17.400 ;
        RECT 21.600 17.330 21.760 17.400 ;
        RECT 1.310 17.320 1.450 17.330 ;
        RECT 4.210 17.320 4.350 17.330 ;
        RECT 7.110 17.320 7.250 17.330 ;
        RECT 10.010 17.320 10.150 17.330 ;
        RECT 12.910 17.320 13.050 17.330 ;
        RECT 15.810 17.320 15.950 17.330 ;
        RECT 18.710 17.320 18.850 17.330 ;
        RECT 21.610 17.320 21.750 17.330 ;
        RECT 0.775 17.120 0.850 17.260 ;
        RECT 0.990 17.070 1.065 17.210 ;
        RECT 1.695 17.130 1.755 17.210 ;
        POLYGON 1.695 17.130 1.755 17.130 1.755 17.070 ;
        RECT 1.910 17.120 1.985 17.260 ;
        RECT 3.675 17.120 3.750 17.260 ;
        RECT 3.890 17.070 3.965 17.210 ;
        RECT 4.595 17.130 4.655 17.210 ;
        POLYGON 4.595 17.130 4.655 17.130 4.655 17.070 ;
        RECT 4.810 17.120 4.885 17.260 ;
        RECT 6.575 17.120 6.650 17.260 ;
        RECT 6.790 17.070 6.865 17.210 ;
        RECT 7.495 17.130 7.555 17.210 ;
        POLYGON 7.495 17.130 7.555 17.130 7.555 17.070 ;
        RECT 7.710 17.120 7.785 17.260 ;
        RECT 9.475 17.120 9.550 17.260 ;
        RECT 9.690 17.070 9.765 17.210 ;
        RECT 10.395 17.130 10.455 17.210 ;
        POLYGON 10.395 17.130 10.455 17.130 10.455 17.070 ;
        RECT 10.610 17.120 10.685 17.260 ;
        RECT 12.375 17.120 12.450 17.260 ;
        RECT 12.590 17.070 12.665 17.210 ;
        RECT 13.295 17.130 13.355 17.210 ;
        POLYGON 13.295 17.130 13.355 17.130 13.355 17.070 ;
        RECT 13.510 17.120 13.585 17.260 ;
        RECT 15.275 17.120 15.350 17.260 ;
        RECT 15.490 17.070 15.565 17.210 ;
        RECT 16.195 17.130 16.255 17.210 ;
        POLYGON 16.195 17.130 16.255 17.130 16.255 17.070 ;
        RECT 16.410 17.120 16.485 17.260 ;
        RECT 18.175 17.120 18.250 17.260 ;
        RECT 18.390 17.070 18.465 17.210 ;
        RECT 19.095 17.130 19.155 17.210 ;
        POLYGON 19.095 17.130 19.155 17.130 19.155 17.070 ;
        RECT 19.310 17.120 19.385 17.260 ;
        RECT 21.075 17.120 21.150 17.260 ;
        RECT 21.290 17.070 21.365 17.210 ;
        RECT 21.995 17.130 22.055 17.210 ;
        POLYGON 21.995 17.130 22.055 17.130 22.055 17.070 ;
        RECT 22.210 17.120 22.285 17.260 ;
        RECT 0.720 16.600 0.870 16.770 ;
        RECT 1.110 16.735 1.260 16.905 ;
        RECT 1.500 16.735 1.650 16.905 ;
        RECT 1.890 16.600 2.040 16.770 ;
        RECT 3.620 16.600 3.770 16.770 ;
        RECT 4.010 16.735 4.160 16.905 ;
        RECT 4.400 16.735 4.550 16.905 ;
        RECT 4.790 16.600 4.940 16.770 ;
        RECT 6.520 16.600 6.670 16.770 ;
        RECT 6.910 16.735 7.060 16.905 ;
        RECT 7.300 16.735 7.450 16.905 ;
        RECT 7.690 16.600 7.840 16.770 ;
        RECT 9.420 16.600 9.570 16.770 ;
        RECT 9.810 16.735 9.960 16.905 ;
        RECT 10.200 16.735 10.350 16.905 ;
        RECT 10.590 16.600 10.740 16.770 ;
        RECT 12.320 16.600 12.470 16.770 ;
        RECT 12.710 16.735 12.860 16.905 ;
        RECT 13.100 16.735 13.250 16.905 ;
        RECT 13.490 16.600 13.640 16.770 ;
        RECT 15.220 16.600 15.370 16.770 ;
        RECT 15.610 16.735 15.760 16.905 ;
        RECT 16.000 16.735 16.150 16.905 ;
        RECT 16.390 16.600 16.540 16.770 ;
        RECT 18.120 16.600 18.270 16.770 ;
        RECT 18.510 16.735 18.660 16.905 ;
        RECT 18.900 16.735 19.050 16.905 ;
        RECT 19.290 16.600 19.440 16.770 ;
        RECT 21.020 16.600 21.170 16.770 ;
        RECT 21.410 16.735 21.560 16.905 ;
        RECT 21.800 16.735 21.950 16.905 ;
        RECT 22.190 16.600 22.340 16.770 ;
        RECT 0.985 16.515 1.035 16.550 ;
        POLYGON 1.035 16.550 1.070 16.515 1.035 16.515 ;
        RECT 0.985 16.390 1.070 16.515 ;
        RECT 1.690 16.390 1.775 16.550 ;
        RECT 3.885 16.515 3.935 16.550 ;
        POLYGON 3.935 16.550 3.970 16.515 3.935 16.515 ;
        RECT 3.885 16.390 3.970 16.515 ;
        RECT 4.590 16.390 4.675 16.550 ;
        RECT 6.785 16.515 6.835 16.550 ;
        POLYGON 6.835 16.550 6.870 16.515 6.835 16.515 ;
        RECT 6.785 16.390 6.870 16.515 ;
        RECT 7.490 16.390 7.575 16.550 ;
        RECT 9.685 16.515 9.735 16.550 ;
        POLYGON 9.735 16.550 9.770 16.515 9.735 16.515 ;
        RECT 9.685 16.390 9.770 16.515 ;
        RECT 10.390 16.390 10.475 16.550 ;
        RECT 12.585 16.515 12.635 16.550 ;
        POLYGON 12.635 16.550 12.670 16.515 12.635 16.515 ;
        RECT 12.585 16.390 12.670 16.515 ;
        RECT 13.290 16.390 13.375 16.550 ;
        RECT 15.485 16.515 15.535 16.550 ;
        POLYGON 15.535 16.550 15.570 16.515 15.535 16.515 ;
        RECT 15.485 16.390 15.570 16.515 ;
        RECT 16.190 16.390 16.275 16.550 ;
        RECT 18.385 16.515 18.435 16.550 ;
        POLYGON 18.435 16.550 18.470 16.515 18.435 16.515 ;
        RECT 18.385 16.390 18.470 16.515 ;
        RECT 19.090 16.390 19.175 16.550 ;
        RECT 21.285 16.515 21.335 16.550 ;
        POLYGON 21.335 16.550 21.370 16.515 21.335 16.515 ;
        RECT 21.285 16.390 21.370 16.515 ;
        RECT 21.990 16.390 22.075 16.550 ;
        RECT 1.300 15.980 1.460 16.050 ;
        RECT 4.200 15.980 4.360 16.050 ;
        RECT 7.100 15.980 7.260 16.050 ;
        RECT 10.000 15.980 10.160 16.050 ;
        RECT 12.900 15.980 13.060 16.050 ;
        RECT 15.800 15.980 15.960 16.050 ;
        RECT 18.700 15.980 18.860 16.050 ;
        RECT 21.600 15.980 21.760 16.050 ;
        RECT 1.310 15.970 1.450 15.980 ;
        RECT 4.210 15.970 4.350 15.980 ;
        RECT 7.110 15.970 7.250 15.980 ;
        RECT 10.010 15.970 10.150 15.980 ;
        RECT 12.910 15.970 13.050 15.980 ;
        RECT 15.810 15.970 15.950 15.980 ;
        RECT 18.710 15.970 18.850 15.980 ;
        RECT 21.610 15.970 21.750 15.980 ;
        RECT 0.775 15.770 0.850 15.910 ;
        RECT 0.990 15.720 1.065 15.860 ;
        RECT 1.695 15.780 1.755 15.860 ;
        POLYGON 1.695 15.780 1.755 15.780 1.755 15.720 ;
        RECT 1.910 15.770 1.985 15.910 ;
        RECT 3.675 15.770 3.750 15.910 ;
        RECT 3.890 15.720 3.965 15.860 ;
        RECT 4.595 15.780 4.655 15.860 ;
        POLYGON 4.595 15.780 4.655 15.780 4.655 15.720 ;
        RECT 4.810 15.770 4.885 15.910 ;
        RECT 6.575 15.770 6.650 15.910 ;
        RECT 6.790 15.720 6.865 15.860 ;
        RECT 7.495 15.780 7.555 15.860 ;
        POLYGON 7.495 15.780 7.555 15.780 7.555 15.720 ;
        RECT 7.710 15.770 7.785 15.910 ;
        RECT 9.475 15.770 9.550 15.910 ;
        RECT 9.690 15.720 9.765 15.860 ;
        RECT 10.395 15.780 10.455 15.860 ;
        POLYGON 10.395 15.780 10.455 15.780 10.455 15.720 ;
        RECT 10.610 15.770 10.685 15.910 ;
        RECT 12.375 15.770 12.450 15.910 ;
        RECT 12.590 15.720 12.665 15.860 ;
        RECT 13.295 15.780 13.355 15.860 ;
        POLYGON 13.295 15.780 13.355 15.780 13.355 15.720 ;
        RECT 13.510 15.770 13.585 15.910 ;
        RECT 15.275 15.770 15.350 15.910 ;
        RECT 15.490 15.720 15.565 15.860 ;
        RECT 16.195 15.780 16.255 15.860 ;
        POLYGON 16.195 15.780 16.255 15.780 16.255 15.720 ;
        RECT 16.410 15.770 16.485 15.910 ;
        RECT 18.175 15.770 18.250 15.910 ;
        RECT 18.390 15.720 18.465 15.860 ;
        RECT 19.095 15.780 19.155 15.860 ;
        POLYGON 19.095 15.780 19.155 15.780 19.155 15.720 ;
        RECT 19.310 15.770 19.385 15.910 ;
        RECT 21.075 15.770 21.150 15.910 ;
        RECT 21.290 15.720 21.365 15.860 ;
        RECT 21.995 15.780 22.055 15.860 ;
        POLYGON 21.995 15.780 22.055 15.780 22.055 15.720 ;
        RECT 22.210 15.770 22.285 15.910 ;
        RECT 0.720 15.250 0.870 15.420 ;
        RECT 1.110 15.385 1.260 15.555 ;
        RECT 1.500 15.385 1.650 15.555 ;
        RECT 1.890 15.250 2.040 15.420 ;
        RECT 3.620 15.250 3.770 15.420 ;
        RECT 4.010 15.385 4.160 15.555 ;
        RECT 4.400 15.385 4.550 15.555 ;
        RECT 4.790 15.250 4.940 15.420 ;
        RECT 6.520 15.250 6.670 15.420 ;
        RECT 6.910 15.385 7.060 15.555 ;
        RECT 7.300 15.385 7.450 15.555 ;
        RECT 7.690 15.250 7.840 15.420 ;
        RECT 9.420 15.250 9.570 15.420 ;
        RECT 9.810 15.385 9.960 15.555 ;
        RECT 10.200 15.385 10.350 15.555 ;
        RECT 10.590 15.250 10.740 15.420 ;
        RECT 12.320 15.250 12.470 15.420 ;
        RECT 12.710 15.385 12.860 15.555 ;
        RECT 13.100 15.385 13.250 15.555 ;
        RECT 13.490 15.250 13.640 15.420 ;
        RECT 15.220 15.250 15.370 15.420 ;
        RECT 15.610 15.385 15.760 15.555 ;
        RECT 16.000 15.385 16.150 15.555 ;
        RECT 16.390 15.250 16.540 15.420 ;
        RECT 18.120 15.250 18.270 15.420 ;
        RECT 18.510 15.385 18.660 15.555 ;
        RECT 18.900 15.385 19.050 15.555 ;
        RECT 19.290 15.250 19.440 15.420 ;
        RECT 21.020 15.250 21.170 15.420 ;
        RECT 21.410 15.385 21.560 15.555 ;
        RECT 21.800 15.385 21.950 15.555 ;
        RECT 22.190 15.250 22.340 15.420 ;
        RECT 0.985 15.165 1.035 15.200 ;
        POLYGON 1.035 15.200 1.070 15.165 1.035 15.165 ;
        RECT 0.985 15.040 1.070 15.165 ;
        RECT 1.690 15.040 1.775 15.200 ;
        RECT 3.885 15.165 3.935 15.200 ;
        POLYGON 3.935 15.200 3.970 15.165 3.935 15.165 ;
        RECT 3.885 15.040 3.970 15.165 ;
        RECT 4.590 15.040 4.675 15.200 ;
        RECT 6.785 15.165 6.835 15.200 ;
        POLYGON 6.835 15.200 6.870 15.165 6.835 15.165 ;
        RECT 6.785 15.040 6.870 15.165 ;
        RECT 7.490 15.040 7.575 15.200 ;
        RECT 9.685 15.165 9.735 15.200 ;
        POLYGON 9.735 15.200 9.770 15.165 9.735 15.165 ;
        RECT 9.685 15.040 9.770 15.165 ;
        RECT 10.390 15.040 10.475 15.200 ;
        RECT 12.585 15.165 12.635 15.200 ;
        POLYGON 12.635 15.200 12.670 15.165 12.635 15.165 ;
        RECT 12.585 15.040 12.670 15.165 ;
        RECT 13.290 15.040 13.375 15.200 ;
        RECT 15.485 15.165 15.535 15.200 ;
        POLYGON 15.535 15.200 15.570 15.165 15.535 15.165 ;
        RECT 15.485 15.040 15.570 15.165 ;
        RECT 16.190 15.040 16.275 15.200 ;
        RECT 18.385 15.165 18.435 15.200 ;
        POLYGON 18.435 15.200 18.470 15.165 18.435 15.165 ;
        RECT 18.385 15.040 18.470 15.165 ;
        RECT 19.090 15.040 19.175 15.200 ;
        RECT 21.285 15.165 21.335 15.200 ;
        POLYGON 21.335 15.200 21.370 15.165 21.335 15.165 ;
        RECT 21.285 15.040 21.370 15.165 ;
        RECT 21.990 15.040 22.075 15.200 ;
        RECT 1.300 14.630 1.460 14.700 ;
        RECT 4.200 14.630 4.360 14.700 ;
        RECT 7.100 14.630 7.260 14.700 ;
        RECT 10.000 14.630 10.160 14.700 ;
        RECT 12.900 14.630 13.060 14.700 ;
        RECT 15.800 14.630 15.960 14.700 ;
        RECT 18.700 14.630 18.860 14.700 ;
        RECT 21.600 14.630 21.760 14.700 ;
        RECT 1.310 14.620 1.450 14.630 ;
        RECT 4.210 14.620 4.350 14.630 ;
        RECT 7.110 14.620 7.250 14.630 ;
        RECT 10.010 14.620 10.150 14.630 ;
        RECT 12.910 14.620 13.050 14.630 ;
        RECT 15.810 14.620 15.950 14.630 ;
        RECT 18.710 14.620 18.850 14.630 ;
        RECT 21.610 14.620 21.750 14.630 ;
        RECT 0.775 14.420 0.850 14.560 ;
        RECT 0.990 14.370 1.065 14.510 ;
        RECT 1.695 14.430 1.755 14.510 ;
        POLYGON 1.695 14.430 1.755 14.430 1.755 14.370 ;
        RECT 1.910 14.420 1.985 14.560 ;
        RECT 3.675 14.420 3.750 14.560 ;
        RECT 3.890 14.370 3.965 14.510 ;
        RECT 4.595 14.430 4.655 14.510 ;
        POLYGON 4.595 14.430 4.655 14.430 4.655 14.370 ;
        RECT 4.810 14.420 4.885 14.560 ;
        RECT 6.575 14.420 6.650 14.560 ;
        RECT 6.790 14.370 6.865 14.510 ;
        RECT 7.495 14.430 7.555 14.510 ;
        POLYGON 7.495 14.430 7.555 14.430 7.555 14.370 ;
        RECT 7.710 14.420 7.785 14.560 ;
        RECT 9.475 14.420 9.550 14.560 ;
        RECT 9.690 14.370 9.765 14.510 ;
        RECT 10.395 14.430 10.455 14.510 ;
        POLYGON 10.395 14.430 10.455 14.430 10.455 14.370 ;
        RECT 10.610 14.420 10.685 14.560 ;
        RECT 12.375 14.420 12.450 14.560 ;
        RECT 12.590 14.370 12.665 14.510 ;
        RECT 13.295 14.430 13.355 14.510 ;
        POLYGON 13.295 14.430 13.355 14.430 13.355 14.370 ;
        RECT 13.510 14.420 13.585 14.560 ;
        RECT 15.275 14.420 15.350 14.560 ;
        RECT 15.490 14.370 15.565 14.510 ;
        RECT 16.195 14.430 16.255 14.510 ;
        POLYGON 16.195 14.430 16.255 14.430 16.255 14.370 ;
        RECT 16.410 14.420 16.485 14.560 ;
        RECT 18.175 14.420 18.250 14.560 ;
        RECT 18.390 14.370 18.465 14.510 ;
        RECT 19.095 14.430 19.155 14.510 ;
        POLYGON 19.095 14.430 19.155 14.430 19.155 14.370 ;
        RECT 19.310 14.420 19.385 14.560 ;
        RECT 21.075 14.420 21.150 14.560 ;
        RECT 21.290 14.370 21.365 14.510 ;
        RECT 21.995 14.430 22.055 14.510 ;
        POLYGON 21.995 14.430 22.055 14.430 22.055 14.370 ;
        RECT 22.210 14.420 22.285 14.560 ;
        RECT 0.720 13.900 0.870 14.070 ;
        RECT 1.110 14.035 1.260 14.205 ;
        RECT 1.500 14.035 1.650 14.205 ;
        RECT 1.890 13.900 2.040 14.070 ;
        RECT 3.620 13.900 3.770 14.070 ;
        RECT 4.010 14.035 4.160 14.205 ;
        RECT 4.400 14.035 4.550 14.205 ;
        RECT 4.790 13.900 4.940 14.070 ;
        RECT 6.520 13.900 6.670 14.070 ;
        RECT 6.910 14.035 7.060 14.205 ;
        RECT 7.300 14.035 7.450 14.205 ;
        RECT 7.690 13.900 7.840 14.070 ;
        RECT 9.420 13.900 9.570 14.070 ;
        RECT 9.810 14.035 9.960 14.205 ;
        RECT 10.200 14.035 10.350 14.205 ;
        RECT 10.590 13.900 10.740 14.070 ;
        RECT 12.320 13.900 12.470 14.070 ;
        RECT 12.710 14.035 12.860 14.205 ;
        RECT 13.100 14.035 13.250 14.205 ;
        RECT 13.490 13.900 13.640 14.070 ;
        RECT 15.220 13.900 15.370 14.070 ;
        RECT 15.610 14.035 15.760 14.205 ;
        RECT 16.000 14.035 16.150 14.205 ;
        RECT 16.390 13.900 16.540 14.070 ;
        RECT 18.120 13.900 18.270 14.070 ;
        RECT 18.510 14.035 18.660 14.205 ;
        RECT 18.900 14.035 19.050 14.205 ;
        RECT 19.290 13.900 19.440 14.070 ;
        RECT 21.020 13.900 21.170 14.070 ;
        RECT 21.410 14.035 21.560 14.205 ;
        RECT 21.800 14.035 21.950 14.205 ;
        RECT 22.190 13.900 22.340 14.070 ;
        RECT 0.985 13.815 1.035 13.850 ;
        POLYGON 1.035 13.850 1.070 13.815 1.035 13.815 ;
        RECT 0.985 13.690 1.070 13.815 ;
        RECT 1.690 13.690 1.775 13.850 ;
        RECT 3.885 13.815 3.935 13.850 ;
        POLYGON 3.935 13.850 3.970 13.815 3.935 13.815 ;
        RECT 3.885 13.690 3.970 13.815 ;
        RECT 4.590 13.690 4.675 13.850 ;
        RECT 6.785 13.815 6.835 13.850 ;
        POLYGON 6.835 13.850 6.870 13.815 6.835 13.815 ;
        RECT 6.785 13.690 6.870 13.815 ;
        RECT 7.490 13.690 7.575 13.850 ;
        RECT 9.685 13.815 9.735 13.850 ;
        POLYGON 9.735 13.850 9.770 13.815 9.735 13.815 ;
        RECT 9.685 13.690 9.770 13.815 ;
        RECT 10.390 13.690 10.475 13.850 ;
        RECT 12.585 13.815 12.635 13.850 ;
        POLYGON 12.635 13.850 12.670 13.815 12.635 13.815 ;
        RECT 12.585 13.690 12.670 13.815 ;
        RECT 13.290 13.690 13.375 13.850 ;
        RECT 15.485 13.815 15.535 13.850 ;
        POLYGON 15.535 13.850 15.570 13.815 15.535 13.815 ;
        RECT 15.485 13.690 15.570 13.815 ;
        RECT 16.190 13.690 16.275 13.850 ;
        RECT 18.385 13.815 18.435 13.850 ;
        POLYGON 18.435 13.850 18.470 13.815 18.435 13.815 ;
        RECT 18.385 13.690 18.470 13.815 ;
        RECT 19.090 13.690 19.175 13.850 ;
        RECT 21.285 13.815 21.335 13.850 ;
        POLYGON 21.335 13.850 21.370 13.815 21.335 13.815 ;
        RECT 21.285 13.690 21.370 13.815 ;
        RECT 21.990 13.690 22.075 13.850 ;
        RECT 1.300 13.280 1.460 13.350 ;
        RECT 4.200 13.280 4.360 13.350 ;
        RECT 7.100 13.280 7.260 13.350 ;
        RECT 10.000 13.280 10.160 13.350 ;
        RECT 12.900 13.280 13.060 13.350 ;
        RECT 15.800 13.280 15.960 13.350 ;
        RECT 18.700 13.280 18.860 13.350 ;
        RECT 21.600 13.280 21.760 13.350 ;
        RECT 1.310 13.270 1.450 13.280 ;
        RECT 4.210 13.270 4.350 13.280 ;
        RECT 7.110 13.270 7.250 13.280 ;
        RECT 10.010 13.270 10.150 13.280 ;
        RECT 12.910 13.270 13.050 13.280 ;
        RECT 15.810 13.270 15.950 13.280 ;
        RECT 18.710 13.270 18.850 13.280 ;
        RECT 21.610 13.270 21.750 13.280 ;
        RECT 0.775 13.070 0.850 13.210 ;
        RECT 0.990 13.020 1.065 13.160 ;
        RECT 1.695 13.080 1.755 13.160 ;
        POLYGON 1.695 13.080 1.755 13.080 1.755 13.020 ;
        RECT 1.910 13.070 1.985 13.210 ;
        RECT 3.675 13.070 3.750 13.210 ;
        RECT 3.890 13.020 3.965 13.160 ;
        RECT 4.595 13.080 4.655 13.160 ;
        POLYGON 4.595 13.080 4.655 13.080 4.655 13.020 ;
        RECT 4.810 13.070 4.885 13.210 ;
        RECT 6.575 13.070 6.650 13.210 ;
        RECT 6.790 13.020 6.865 13.160 ;
        RECT 7.495 13.080 7.555 13.160 ;
        POLYGON 7.495 13.080 7.555 13.080 7.555 13.020 ;
        RECT 7.710 13.070 7.785 13.210 ;
        RECT 9.475 13.070 9.550 13.210 ;
        RECT 9.690 13.020 9.765 13.160 ;
        RECT 10.395 13.080 10.455 13.160 ;
        POLYGON 10.395 13.080 10.455 13.080 10.455 13.020 ;
        RECT 10.610 13.070 10.685 13.210 ;
        RECT 12.375 13.070 12.450 13.210 ;
        RECT 12.590 13.020 12.665 13.160 ;
        RECT 13.295 13.080 13.355 13.160 ;
        POLYGON 13.295 13.080 13.355 13.080 13.355 13.020 ;
        RECT 13.510 13.070 13.585 13.210 ;
        RECT 15.275 13.070 15.350 13.210 ;
        RECT 15.490 13.020 15.565 13.160 ;
        RECT 16.195 13.080 16.255 13.160 ;
        POLYGON 16.195 13.080 16.255 13.080 16.255 13.020 ;
        RECT 16.410 13.070 16.485 13.210 ;
        RECT 18.175 13.070 18.250 13.210 ;
        RECT 18.390 13.020 18.465 13.160 ;
        RECT 19.095 13.080 19.155 13.160 ;
        POLYGON 19.095 13.080 19.155 13.080 19.155 13.020 ;
        RECT 19.310 13.070 19.385 13.210 ;
        RECT 21.075 13.070 21.150 13.210 ;
        RECT 21.290 13.020 21.365 13.160 ;
        RECT 21.995 13.080 22.055 13.160 ;
        POLYGON 21.995 13.080 22.055 13.080 22.055 13.020 ;
        RECT 22.210 13.070 22.285 13.210 ;
        RECT 0.720 12.550 0.870 12.720 ;
        RECT 1.110 12.685 1.260 12.855 ;
        RECT 1.500 12.685 1.650 12.855 ;
        RECT 1.890 12.550 2.040 12.720 ;
        RECT 3.620 12.550 3.770 12.720 ;
        RECT 4.010 12.685 4.160 12.855 ;
        RECT 4.400 12.685 4.550 12.855 ;
        RECT 4.790 12.550 4.940 12.720 ;
        RECT 6.520 12.550 6.670 12.720 ;
        RECT 6.910 12.685 7.060 12.855 ;
        RECT 7.300 12.685 7.450 12.855 ;
        RECT 7.690 12.550 7.840 12.720 ;
        RECT 9.420 12.550 9.570 12.720 ;
        RECT 9.810 12.685 9.960 12.855 ;
        RECT 10.200 12.685 10.350 12.855 ;
        RECT 10.590 12.550 10.740 12.720 ;
        RECT 12.320 12.550 12.470 12.720 ;
        RECT 12.710 12.685 12.860 12.855 ;
        RECT 13.100 12.685 13.250 12.855 ;
        RECT 13.490 12.550 13.640 12.720 ;
        RECT 15.220 12.550 15.370 12.720 ;
        RECT 15.610 12.685 15.760 12.855 ;
        RECT 16.000 12.685 16.150 12.855 ;
        RECT 16.390 12.550 16.540 12.720 ;
        RECT 18.120 12.550 18.270 12.720 ;
        RECT 18.510 12.685 18.660 12.855 ;
        RECT 18.900 12.685 19.050 12.855 ;
        RECT 19.290 12.550 19.440 12.720 ;
        RECT 21.020 12.550 21.170 12.720 ;
        RECT 21.410 12.685 21.560 12.855 ;
        RECT 21.800 12.685 21.950 12.855 ;
        RECT 22.190 12.550 22.340 12.720 ;
        RECT 0.985 12.465 1.035 12.500 ;
        POLYGON 1.035 12.500 1.070 12.465 1.035 12.465 ;
        RECT 0.985 12.340 1.070 12.465 ;
        RECT 1.690 12.340 1.775 12.500 ;
        RECT 3.885 12.465 3.935 12.500 ;
        POLYGON 3.935 12.500 3.970 12.465 3.935 12.465 ;
        RECT 3.885 12.340 3.970 12.465 ;
        RECT 4.590 12.340 4.675 12.500 ;
        RECT 6.785 12.465 6.835 12.500 ;
        POLYGON 6.835 12.500 6.870 12.465 6.835 12.465 ;
        RECT 6.785 12.340 6.870 12.465 ;
        RECT 7.490 12.340 7.575 12.500 ;
        RECT 9.685 12.465 9.735 12.500 ;
        POLYGON 9.735 12.500 9.770 12.465 9.735 12.465 ;
        RECT 9.685 12.340 9.770 12.465 ;
        RECT 10.390 12.340 10.475 12.500 ;
        RECT 12.585 12.465 12.635 12.500 ;
        POLYGON 12.635 12.500 12.670 12.465 12.635 12.465 ;
        RECT 12.585 12.340 12.670 12.465 ;
        RECT 13.290 12.340 13.375 12.500 ;
        RECT 15.485 12.465 15.535 12.500 ;
        POLYGON 15.535 12.500 15.570 12.465 15.535 12.465 ;
        RECT 15.485 12.340 15.570 12.465 ;
        RECT 16.190 12.340 16.275 12.500 ;
        RECT 18.385 12.465 18.435 12.500 ;
        POLYGON 18.435 12.500 18.470 12.465 18.435 12.465 ;
        RECT 18.385 12.340 18.470 12.465 ;
        RECT 19.090 12.340 19.175 12.500 ;
        RECT 21.285 12.465 21.335 12.500 ;
        POLYGON 21.335 12.500 21.370 12.465 21.335 12.465 ;
        RECT 21.285 12.340 21.370 12.465 ;
        RECT 21.990 12.340 22.075 12.500 ;
        RECT 1.300 11.930 1.460 12.000 ;
        RECT 4.200 11.930 4.360 12.000 ;
        RECT 7.100 11.930 7.260 12.000 ;
        RECT 10.000 11.930 10.160 12.000 ;
        RECT 12.900 11.930 13.060 12.000 ;
        RECT 15.800 11.930 15.960 12.000 ;
        RECT 18.700 11.930 18.860 12.000 ;
        RECT 21.600 11.930 21.760 12.000 ;
        RECT 1.310 11.920 1.450 11.930 ;
        RECT 4.210 11.920 4.350 11.930 ;
        RECT 7.110 11.920 7.250 11.930 ;
        RECT 10.010 11.920 10.150 11.930 ;
        RECT 12.910 11.920 13.050 11.930 ;
        RECT 15.810 11.920 15.950 11.930 ;
        RECT 18.710 11.920 18.850 11.930 ;
        RECT 21.610 11.920 21.750 11.930 ;
        RECT 0.775 11.720 0.850 11.860 ;
        RECT 0.990 11.670 1.065 11.810 ;
        RECT 1.695 11.730 1.755 11.810 ;
        POLYGON 1.695 11.730 1.755 11.730 1.755 11.670 ;
        RECT 1.910 11.720 1.985 11.860 ;
        RECT 3.675 11.720 3.750 11.860 ;
        RECT 3.890 11.670 3.965 11.810 ;
        RECT 4.595 11.730 4.655 11.810 ;
        POLYGON 4.595 11.730 4.655 11.730 4.655 11.670 ;
        RECT 4.810 11.720 4.885 11.860 ;
        RECT 6.575 11.720 6.650 11.860 ;
        RECT 6.790 11.670 6.865 11.810 ;
        RECT 7.495 11.730 7.555 11.810 ;
        POLYGON 7.495 11.730 7.555 11.730 7.555 11.670 ;
        RECT 7.710 11.720 7.785 11.860 ;
        RECT 9.475 11.720 9.550 11.860 ;
        RECT 9.690 11.670 9.765 11.810 ;
        RECT 10.395 11.730 10.455 11.810 ;
        POLYGON 10.395 11.730 10.455 11.730 10.455 11.670 ;
        RECT 10.610 11.720 10.685 11.860 ;
        RECT 12.375 11.720 12.450 11.860 ;
        RECT 12.590 11.670 12.665 11.810 ;
        RECT 13.295 11.730 13.355 11.810 ;
        POLYGON 13.295 11.730 13.355 11.730 13.355 11.670 ;
        RECT 13.510 11.720 13.585 11.860 ;
        RECT 15.275 11.720 15.350 11.860 ;
        RECT 15.490 11.670 15.565 11.810 ;
        RECT 16.195 11.730 16.255 11.810 ;
        POLYGON 16.195 11.730 16.255 11.730 16.255 11.670 ;
        RECT 16.410 11.720 16.485 11.860 ;
        RECT 18.175 11.720 18.250 11.860 ;
        RECT 18.390 11.670 18.465 11.810 ;
        RECT 19.095 11.730 19.155 11.810 ;
        POLYGON 19.095 11.730 19.155 11.730 19.155 11.670 ;
        RECT 19.310 11.720 19.385 11.860 ;
        RECT 21.075 11.720 21.150 11.860 ;
        RECT 21.290 11.670 21.365 11.810 ;
        RECT 21.995 11.730 22.055 11.810 ;
        POLYGON 21.995 11.730 22.055 11.730 22.055 11.670 ;
        RECT 22.210 11.720 22.285 11.860 ;
        RECT 0.720 11.200 0.870 11.370 ;
        RECT 1.110 11.335 1.260 11.505 ;
        RECT 1.500 11.335 1.650 11.505 ;
        RECT 1.890 11.200 2.040 11.370 ;
        RECT 3.620 11.200 3.770 11.370 ;
        RECT 4.010 11.335 4.160 11.505 ;
        RECT 4.400 11.335 4.550 11.505 ;
        RECT 4.790 11.200 4.940 11.370 ;
        RECT 6.520 11.200 6.670 11.370 ;
        RECT 6.910 11.335 7.060 11.505 ;
        RECT 7.300 11.335 7.450 11.505 ;
        RECT 7.690 11.200 7.840 11.370 ;
        RECT 9.420 11.200 9.570 11.370 ;
        RECT 9.810 11.335 9.960 11.505 ;
        RECT 10.200 11.335 10.350 11.505 ;
        RECT 10.590 11.200 10.740 11.370 ;
        RECT 12.320 11.200 12.470 11.370 ;
        RECT 12.710 11.335 12.860 11.505 ;
        RECT 13.100 11.335 13.250 11.505 ;
        RECT 13.490 11.200 13.640 11.370 ;
        RECT 15.220 11.200 15.370 11.370 ;
        RECT 15.610 11.335 15.760 11.505 ;
        RECT 16.000 11.335 16.150 11.505 ;
        RECT 16.390 11.200 16.540 11.370 ;
        RECT 18.120 11.200 18.270 11.370 ;
        RECT 18.510 11.335 18.660 11.505 ;
        RECT 18.900 11.335 19.050 11.505 ;
        RECT 19.290 11.200 19.440 11.370 ;
        RECT 21.020 11.200 21.170 11.370 ;
        RECT 21.410 11.335 21.560 11.505 ;
        RECT 21.800 11.335 21.950 11.505 ;
        RECT 22.190 11.200 22.340 11.370 ;
        RECT 0.985 11.115 1.035 11.150 ;
        POLYGON 1.035 11.150 1.070 11.115 1.035 11.115 ;
        RECT 0.985 10.990 1.070 11.115 ;
        RECT 1.690 10.990 1.775 11.150 ;
        RECT 3.885 11.115 3.935 11.150 ;
        POLYGON 3.935 11.150 3.970 11.115 3.935 11.115 ;
        RECT 3.885 10.990 3.970 11.115 ;
        RECT 4.590 10.990 4.675 11.150 ;
        RECT 6.785 11.115 6.835 11.150 ;
        POLYGON 6.835 11.150 6.870 11.115 6.835 11.115 ;
        RECT 6.785 10.990 6.870 11.115 ;
        RECT 7.490 10.990 7.575 11.150 ;
        RECT 9.685 11.115 9.735 11.150 ;
        POLYGON 9.735 11.150 9.770 11.115 9.735 11.115 ;
        RECT 9.685 10.990 9.770 11.115 ;
        RECT 10.390 10.990 10.475 11.150 ;
        RECT 12.585 11.115 12.635 11.150 ;
        POLYGON 12.635 11.150 12.670 11.115 12.635 11.115 ;
        RECT 12.585 10.990 12.670 11.115 ;
        RECT 13.290 10.990 13.375 11.150 ;
        RECT 15.485 11.115 15.535 11.150 ;
        POLYGON 15.535 11.150 15.570 11.115 15.535 11.115 ;
        RECT 15.485 10.990 15.570 11.115 ;
        RECT 16.190 10.990 16.275 11.150 ;
        RECT 18.385 11.115 18.435 11.150 ;
        POLYGON 18.435 11.150 18.470 11.115 18.435 11.115 ;
        RECT 18.385 10.990 18.470 11.115 ;
        RECT 19.090 10.990 19.175 11.150 ;
        RECT 21.285 11.115 21.335 11.150 ;
        POLYGON 21.335 11.150 21.370 11.115 21.335 11.115 ;
        RECT 21.285 10.990 21.370 11.115 ;
        RECT 21.990 10.990 22.075 11.150 ;
        RECT 1.300 10.580 1.460 10.650 ;
        RECT 4.200 10.580 4.360 10.650 ;
        RECT 7.100 10.580 7.260 10.650 ;
        RECT 10.000 10.580 10.160 10.650 ;
        RECT 12.900 10.580 13.060 10.650 ;
        RECT 15.800 10.580 15.960 10.650 ;
        RECT 18.700 10.580 18.860 10.650 ;
        RECT 21.600 10.580 21.760 10.650 ;
        RECT 1.310 10.570 1.450 10.580 ;
        RECT 4.210 10.570 4.350 10.580 ;
        RECT 7.110 10.570 7.250 10.580 ;
        RECT 10.010 10.570 10.150 10.580 ;
        RECT 12.910 10.570 13.050 10.580 ;
        RECT 15.810 10.570 15.950 10.580 ;
        RECT 18.710 10.570 18.850 10.580 ;
        RECT 21.610 10.570 21.750 10.580 ;
        RECT 0.775 10.370 0.850 10.510 ;
        RECT 0.990 10.320 1.065 10.460 ;
        RECT 1.695 10.380 1.755 10.460 ;
        POLYGON 1.695 10.380 1.755 10.380 1.755 10.320 ;
        RECT 1.910 10.370 1.985 10.510 ;
        RECT 3.675 10.370 3.750 10.510 ;
        RECT 3.890 10.320 3.965 10.460 ;
        RECT 4.595 10.380 4.655 10.460 ;
        POLYGON 4.595 10.380 4.655 10.380 4.655 10.320 ;
        RECT 4.810 10.370 4.885 10.510 ;
        RECT 6.575 10.370 6.650 10.510 ;
        RECT 6.790 10.320 6.865 10.460 ;
        RECT 7.495 10.380 7.555 10.460 ;
        POLYGON 7.495 10.380 7.555 10.380 7.555 10.320 ;
        RECT 7.710 10.370 7.785 10.510 ;
        RECT 9.475 10.370 9.550 10.510 ;
        RECT 9.690 10.320 9.765 10.460 ;
        RECT 10.395 10.380 10.455 10.460 ;
        POLYGON 10.395 10.380 10.455 10.380 10.455 10.320 ;
        RECT 10.610 10.370 10.685 10.510 ;
        RECT 12.375 10.370 12.450 10.510 ;
        RECT 12.590 10.320 12.665 10.460 ;
        RECT 13.295 10.380 13.355 10.460 ;
        POLYGON 13.295 10.380 13.355 10.380 13.355 10.320 ;
        RECT 13.510 10.370 13.585 10.510 ;
        RECT 15.275 10.370 15.350 10.510 ;
        RECT 15.490 10.320 15.565 10.460 ;
        RECT 16.195 10.380 16.255 10.460 ;
        POLYGON 16.195 10.380 16.255 10.380 16.255 10.320 ;
        RECT 16.410 10.370 16.485 10.510 ;
        RECT 18.175 10.370 18.250 10.510 ;
        RECT 18.390 10.320 18.465 10.460 ;
        RECT 19.095 10.380 19.155 10.460 ;
        POLYGON 19.095 10.380 19.155 10.380 19.155 10.320 ;
        RECT 19.310 10.370 19.385 10.510 ;
        RECT 21.075 10.370 21.150 10.510 ;
        RECT 21.290 10.320 21.365 10.460 ;
        RECT 21.995 10.380 22.055 10.460 ;
        POLYGON 21.995 10.380 22.055 10.380 22.055 10.320 ;
        RECT 22.210 10.370 22.285 10.510 ;
        RECT 0.720 9.850 0.870 10.020 ;
        RECT 1.110 9.985 1.260 10.155 ;
        RECT 1.500 9.985 1.650 10.155 ;
        RECT 1.890 9.850 2.040 10.020 ;
        RECT 3.620 9.850 3.770 10.020 ;
        RECT 4.010 9.985 4.160 10.155 ;
        RECT 4.400 9.985 4.550 10.155 ;
        RECT 4.790 9.850 4.940 10.020 ;
        RECT 6.520 9.850 6.670 10.020 ;
        RECT 6.910 9.985 7.060 10.155 ;
        RECT 7.300 9.985 7.450 10.155 ;
        RECT 7.690 9.850 7.840 10.020 ;
        RECT 9.420 9.850 9.570 10.020 ;
        RECT 9.810 9.985 9.960 10.155 ;
        RECT 10.200 9.985 10.350 10.155 ;
        RECT 10.590 9.850 10.740 10.020 ;
        RECT 12.320 9.850 12.470 10.020 ;
        RECT 12.710 9.985 12.860 10.155 ;
        RECT 13.100 9.985 13.250 10.155 ;
        RECT 13.490 9.850 13.640 10.020 ;
        RECT 15.220 9.850 15.370 10.020 ;
        RECT 15.610 9.985 15.760 10.155 ;
        RECT 16.000 9.985 16.150 10.155 ;
        RECT 16.390 9.850 16.540 10.020 ;
        RECT 18.120 9.850 18.270 10.020 ;
        RECT 18.510 9.985 18.660 10.155 ;
        RECT 18.900 9.985 19.050 10.155 ;
        RECT 19.290 9.850 19.440 10.020 ;
        RECT 21.020 9.850 21.170 10.020 ;
        RECT 21.410 9.985 21.560 10.155 ;
        RECT 21.800 9.985 21.950 10.155 ;
        RECT 22.190 9.850 22.340 10.020 ;
        RECT 0.985 9.765 1.035 9.800 ;
        POLYGON 1.035 9.800 1.070 9.765 1.035 9.765 ;
        RECT 0.985 9.640 1.070 9.765 ;
        RECT 1.690 9.640 1.775 9.800 ;
        RECT 3.885 9.765 3.935 9.800 ;
        POLYGON 3.935 9.800 3.970 9.765 3.935 9.765 ;
        RECT 3.885 9.640 3.970 9.765 ;
        RECT 4.590 9.640 4.675 9.800 ;
        RECT 6.785 9.765 6.835 9.800 ;
        POLYGON 6.835 9.800 6.870 9.765 6.835 9.765 ;
        RECT 6.785 9.640 6.870 9.765 ;
        RECT 7.490 9.640 7.575 9.800 ;
        RECT 9.685 9.765 9.735 9.800 ;
        POLYGON 9.735 9.800 9.770 9.765 9.735 9.765 ;
        RECT 9.685 9.640 9.770 9.765 ;
        RECT 10.390 9.640 10.475 9.800 ;
        RECT 12.585 9.765 12.635 9.800 ;
        POLYGON 12.635 9.800 12.670 9.765 12.635 9.765 ;
        RECT 12.585 9.640 12.670 9.765 ;
        RECT 13.290 9.640 13.375 9.800 ;
        RECT 15.485 9.765 15.535 9.800 ;
        POLYGON 15.535 9.800 15.570 9.765 15.535 9.765 ;
        RECT 15.485 9.640 15.570 9.765 ;
        RECT 16.190 9.640 16.275 9.800 ;
        RECT 18.385 9.765 18.435 9.800 ;
        POLYGON 18.435 9.800 18.470 9.765 18.435 9.765 ;
        RECT 18.385 9.640 18.470 9.765 ;
        RECT 19.090 9.640 19.175 9.800 ;
        RECT 21.285 9.765 21.335 9.800 ;
        POLYGON 21.335 9.800 21.370 9.765 21.335 9.765 ;
        RECT 21.285 9.640 21.370 9.765 ;
        RECT 21.990 9.640 22.075 9.800 ;
        RECT 1.300 9.230 1.460 9.300 ;
        RECT 4.200 9.230 4.360 9.300 ;
        RECT 7.100 9.230 7.260 9.300 ;
        RECT 10.000 9.230 10.160 9.300 ;
        RECT 12.900 9.230 13.060 9.300 ;
        RECT 15.800 9.230 15.960 9.300 ;
        RECT 18.700 9.230 18.860 9.300 ;
        RECT 21.600 9.230 21.760 9.300 ;
        RECT 1.310 9.220 1.450 9.230 ;
        RECT 4.210 9.220 4.350 9.230 ;
        RECT 7.110 9.220 7.250 9.230 ;
        RECT 10.010 9.220 10.150 9.230 ;
        RECT 12.910 9.220 13.050 9.230 ;
        RECT 15.810 9.220 15.950 9.230 ;
        RECT 18.710 9.220 18.850 9.230 ;
        RECT 21.610 9.220 21.750 9.230 ;
        RECT 0.775 9.020 0.850 9.160 ;
        RECT 0.990 8.970 1.065 9.110 ;
        RECT 1.695 9.030 1.755 9.110 ;
        POLYGON 1.695 9.030 1.755 9.030 1.755 8.970 ;
        RECT 1.910 9.020 1.985 9.160 ;
        RECT 3.675 9.020 3.750 9.160 ;
        RECT 3.890 8.970 3.965 9.110 ;
        RECT 4.595 9.030 4.655 9.110 ;
        POLYGON 4.595 9.030 4.655 9.030 4.655 8.970 ;
        RECT 4.810 9.020 4.885 9.160 ;
        RECT 6.575 9.020 6.650 9.160 ;
        RECT 6.790 8.970 6.865 9.110 ;
        RECT 7.495 9.030 7.555 9.110 ;
        POLYGON 7.495 9.030 7.555 9.030 7.555 8.970 ;
        RECT 7.710 9.020 7.785 9.160 ;
        RECT 9.475 9.020 9.550 9.160 ;
        RECT 9.690 8.970 9.765 9.110 ;
        RECT 10.395 9.030 10.455 9.110 ;
        POLYGON 10.395 9.030 10.455 9.030 10.455 8.970 ;
        RECT 10.610 9.020 10.685 9.160 ;
        RECT 12.375 9.020 12.450 9.160 ;
        RECT 12.590 8.970 12.665 9.110 ;
        RECT 13.295 9.030 13.355 9.110 ;
        POLYGON 13.295 9.030 13.355 9.030 13.355 8.970 ;
        RECT 13.510 9.020 13.585 9.160 ;
        RECT 15.275 9.020 15.350 9.160 ;
        RECT 15.490 8.970 15.565 9.110 ;
        RECT 16.195 9.030 16.255 9.110 ;
        POLYGON 16.195 9.030 16.255 9.030 16.255 8.970 ;
        RECT 16.410 9.020 16.485 9.160 ;
        RECT 18.175 9.020 18.250 9.160 ;
        RECT 18.390 8.970 18.465 9.110 ;
        RECT 19.095 9.030 19.155 9.110 ;
        POLYGON 19.095 9.030 19.155 9.030 19.155 8.970 ;
        RECT 19.310 9.020 19.385 9.160 ;
        RECT 21.075 9.020 21.150 9.160 ;
        RECT 21.290 8.970 21.365 9.110 ;
        RECT 21.995 9.030 22.055 9.110 ;
        POLYGON 21.995 9.030 22.055 9.030 22.055 8.970 ;
        RECT 22.210 9.020 22.285 9.160 ;
        RECT 0.720 8.500 0.870 8.670 ;
        RECT 1.110 8.635 1.260 8.805 ;
        RECT 1.500 8.635 1.650 8.805 ;
        RECT 1.890 8.500 2.040 8.670 ;
        RECT 3.620 8.500 3.770 8.670 ;
        RECT 4.010 8.635 4.160 8.805 ;
        RECT 4.400 8.635 4.550 8.805 ;
        RECT 4.790 8.500 4.940 8.670 ;
        RECT 6.520 8.500 6.670 8.670 ;
        RECT 6.910 8.635 7.060 8.805 ;
        RECT 7.300 8.635 7.450 8.805 ;
        RECT 7.690 8.500 7.840 8.670 ;
        RECT 9.420 8.500 9.570 8.670 ;
        RECT 9.810 8.635 9.960 8.805 ;
        RECT 10.200 8.635 10.350 8.805 ;
        RECT 10.590 8.500 10.740 8.670 ;
        RECT 12.320 8.500 12.470 8.670 ;
        RECT 12.710 8.635 12.860 8.805 ;
        RECT 13.100 8.635 13.250 8.805 ;
        RECT 13.490 8.500 13.640 8.670 ;
        RECT 15.220 8.500 15.370 8.670 ;
        RECT 15.610 8.635 15.760 8.805 ;
        RECT 16.000 8.635 16.150 8.805 ;
        RECT 16.390 8.500 16.540 8.670 ;
        RECT 18.120 8.500 18.270 8.670 ;
        RECT 18.510 8.635 18.660 8.805 ;
        RECT 18.900 8.635 19.050 8.805 ;
        RECT 19.290 8.500 19.440 8.670 ;
        RECT 21.020 8.500 21.170 8.670 ;
        RECT 21.410 8.635 21.560 8.805 ;
        RECT 21.800 8.635 21.950 8.805 ;
        RECT 22.190 8.500 22.340 8.670 ;
        RECT 0.985 8.415 1.035 8.450 ;
        POLYGON 1.035 8.450 1.070 8.415 1.035 8.415 ;
        RECT 0.985 8.290 1.070 8.415 ;
        RECT 1.690 8.290 1.775 8.450 ;
        RECT 3.885 8.415 3.935 8.450 ;
        POLYGON 3.935 8.450 3.970 8.415 3.935 8.415 ;
        RECT 3.885 8.290 3.970 8.415 ;
        RECT 4.590 8.290 4.675 8.450 ;
        RECT 6.785 8.415 6.835 8.450 ;
        POLYGON 6.835 8.450 6.870 8.415 6.835 8.415 ;
        RECT 6.785 8.290 6.870 8.415 ;
        RECT 7.490 8.290 7.575 8.450 ;
        RECT 9.685 8.415 9.735 8.450 ;
        POLYGON 9.735 8.450 9.770 8.415 9.735 8.415 ;
        RECT 9.685 8.290 9.770 8.415 ;
        RECT 10.390 8.290 10.475 8.450 ;
        RECT 12.585 8.415 12.635 8.450 ;
        POLYGON 12.635 8.450 12.670 8.415 12.635 8.415 ;
        RECT 12.585 8.290 12.670 8.415 ;
        RECT 13.290 8.290 13.375 8.450 ;
        RECT 15.485 8.415 15.535 8.450 ;
        POLYGON 15.535 8.450 15.570 8.415 15.535 8.415 ;
        RECT 15.485 8.290 15.570 8.415 ;
        RECT 16.190 8.290 16.275 8.450 ;
        RECT 18.385 8.415 18.435 8.450 ;
        POLYGON 18.435 8.450 18.470 8.415 18.435 8.415 ;
        RECT 18.385 8.290 18.470 8.415 ;
        RECT 19.090 8.290 19.175 8.450 ;
        RECT 21.285 8.415 21.335 8.450 ;
        POLYGON 21.335 8.450 21.370 8.415 21.335 8.415 ;
        RECT 21.285 8.290 21.370 8.415 ;
        RECT 21.990 8.290 22.075 8.450 ;
        RECT 1.300 7.880 1.460 7.950 ;
        RECT 4.200 7.880 4.360 7.950 ;
        RECT 7.100 7.880 7.260 7.950 ;
        RECT 10.000 7.880 10.160 7.950 ;
        RECT 12.900 7.880 13.060 7.950 ;
        RECT 15.800 7.880 15.960 7.950 ;
        RECT 18.700 7.880 18.860 7.950 ;
        RECT 21.600 7.880 21.760 7.950 ;
        RECT 1.310 7.870 1.450 7.880 ;
        RECT 4.210 7.870 4.350 7.880 ;
        RECT 7.110 7.870 7.250 7.880 ;
        RECT 10.010 7.870 10.150 7.880 ;
        RECT 12.910 7.870 13.050 7.880 ;
        RECT 15.810 7.870 15.950 7.880 ;
        RECT 18.710 7.870 18.850 7.880 ;
        RECT 21.610 7.870 21.750 7.880 ;
        RECT 0.775 7.670 0.850 7.810 ;
        RECT 0.990 7.620 1.065 7.760 ;
        RECT 1.695 7.680 1.755 7.760 ;
        POLYGON 1.695 7.680 1.755 7.680 1.755 7.620 ;
        RECT 1.910 7.670 1.985 7.810 ;
        RECT 3.675 7.670 3.750 7.810 ;
        RECT 3.890 7.620 3.965 7.760 ;
        RECT 4.595 7.680 4.655 7.760 ;
        POLYGON 4.595 7.680 4.655 7.680 4.655 7.620 ;
        RECT 4.810 7.670 4.885 7.810 ;
        RECT 6.575 7.670 6.650 7.810 ;
        RECT 6.790 7.620 6.865 7.760 ;
        RECT 7.495 7.680 7.555 7.760 ;
        POLYGON 7.495 7.680 7.555 7.680 7.555 7.620 ;
        RECT 7.710 7.670 7.785 7.810 ;
        RECT 9.475 7.670 9.550 7.810 ;
        RECT 9.690 7.620 9.765 7.760 ;
        RECT 10.395 7.680 10.455 7.760 ;
        POLYGON 10.395 7.680 10.455 7.680 10.455 7.620 ;
        RECT 10.610 7.670 10.685 7.810 ;
        RECT 12.375 7.670 12.450 7.810 ;
        RECT 12.590 7.620 12.665 7.760 ;
        RECT 13.295 7.680 13.355 7.760 ;
        POLYGON 13.295 7.680 13.355 7.680 13.355 7.620 ;
        RECT 13.510 7.670 13.585 7.810 ;
        RECT 15.275 7.670 15.350 7.810 ;
        RECT 15.490 7.620 15.565 7.760 ;
        RECT 16.195 7.680 16.255 7.760 ;
        POLYGON 16.195 7.680 16.255 7.680 16.255 7.620 ;
        RECT 16.410 7.670 16.485 7.810 ;
        RECT 18.175 7.670 18.250 7.810 ;
        RECT 18.390 7.620 18.465 7.760 ;
        RECT 19.095 7.680 19.155 7.760 ;
        POLYGON 19.095 7.680 19.155 7.680 19.155 7.620 ;
        RECT 19.310 7.670 19.385 7.810 ;
        RECT 21.075 7.670 21.150 7.810 ;
        RECT 21.290 7.620 21.365 7.760 ;
        RECT 21.995 7.680 22.055 7.760 ;
        POLYGON 21.995 7.680 22.055 7.680 22.055 7.620 ;
        RECT 22.210 7.670 22.285 7.810 ;
        RECT 0.720 7.150 0.870 7.320 ;
        RECT 1.110 7.285 1.260 7.455 ;
        RECT 1.500 7.285 1.650 7.455 ;
        RECT 1.890 7.150 2.040 7.320 ;
        RECT 3.620 7.150 3.770 7.320 ;
        RECT 4.010 7.285 4.160 7.455 ;
        RECT 4.400 7.285 4.550 7.455 ;
        RECT 4.790 7.150 4.940 7.320 ;
        RECT 6.520 7.150 6.670 7.320 ;
        RECT 6.910 7.285 7.060 7.455 ;
        RECT 7.300 7.285 7.450 7.455 ;
        RECT 7.690 7.150 7.840 7.320 ;
        RECT 9.420 7.150 9.570 7.320 ;
        RECT 9.810 7.285 9.960 7.455 ;
        RECT 10.200 7.285 10.350 7.455 ;
        RECT 10.590 7.150 10.740 7.320 ;
        RECT 12.320 7.150 12.470 7.320 ;
        RECT 12.710 7.285 12.860 7.455 ;
        RECT 13.100 7.285 13.250 7.455 ;
        RECT 13.490 7.150 13.640 7.320 ;
        RECT 15.220 7.150 15.370 7.320 ;
        RECT 15.610 7.285 15.760 7.455 ;
        RECT 16.000 7.285 16.150 7.455 ;
        RECT 16.390 7.150 16.540 7.320 ;
        RECT 18.120 7.150 18.270 7.320 ;
        RECT 18.510 7.285 18.660 7.455 ;
        RECT 18.900 7.285 19.050 7.455 ;
        RECT 19.290 7.150 19.440 7.320 ;
        RECT 21.020 7.150 21.170 7.320 ;
        RECT 21.410 7.285 21.560 7.455 ;
        RECT 21.800 7.285 21.950 7.455 ;
        RECT 22.190 7.150 22.340 7.320 ;
        RECT 0.985 7.065 1.035 7.100 ;
        POLYGON 1.035 7.100 1.070 7.065 1.035 7.065 ;
        RECT 0.985 6.940 1.070 7.065 ;
        RECT 1.690 6.940 1.775 7.100 ;
        RECT 3.885 7.065 3.935 7.100 ;
        POLYGON 3.935 7.100 3.970 7.065 3.935 7.065 ;
        RECT 3.885 6.940 3.970 7.065 ;
        RECT 4.590 6.940 4.675 7.100 ;
        RECT 6.785 7.065 6.835 7.100 ;
        POLYGON 6.835 7.100 6.870 7.065 6.835 7.065 ;
        RECT 6.785 6.940 6.870 7.065 ;
        RECT 7.490 6.940 7.575 7.100 ;
        RECT 9.685 7.065 9.735 7.100 ;
        POLYGON 9.735 7.100 9.770 7.065 9.735 7.065 ;
        RECT 9.685 6.940 9.770 7.065 ;
        RECT 10.390 6.940 10.475 7.100 ;
        RECT 12.585 7.065 12.635 7.100 ;
        POLYGON 12.635 7.100 12.670 7.065 12.635 7.065 ;
        RECT 12.585 6.940 12.670 7.065 ;
        RECT 13.290 6.940 13.375 7.100 ;
        RECT 15.485 7.065 15.535 7.100 ;
        POLYGON 15.535 7.100 15.570 7.065 15.535 7.065 ;
        RECT 15.485 6.940 15.570 7.065 ;
        RECT 16.190 6.940 16.275 7.100 ;
        RECT 18.385 7.065 18.435 7.100 ;
        POLYGON 18.435 7.100 18.470 7.065 18.435 7.065 ;
        RECT 18.385 6.940 18.470 7.065 ;
        RECT 19.090 6.940 19.175 7.100 ;
        RECT 21.285 7.065 21.335 7.100 ;
        POLYGON 21.335 7.100 21.370 7.065 21.335 7.065 ;
        RECT 21.285 6.940 21.370 7.065 ;
        RECT 21.990 6.940 22.075 7.100 ;
        RECT 1.300 6.530 1.460 6.600 ;
        RECT 4.200 6.530 4.360 6.600 ;
        RECT 7.100 6.530 7.260 6.600 ;
        RECT 10.000 6.530 10.160 6.600 ;
        RECT 12.900 6.530 13.060 6.600 ;
        RECT 15.800 6.530 15.960 6.600 ;
        RECT 18.700 6.530 18.860 6.600 ;
        RECT 21.600 6.530 21.760 6.600 ;
        RECT 1.310 6.520 1.450 6.530 ;
        RECT 4.210 6.520 4.350 6.530 ;
        RECT 7.110 6.520 7.250 6.530 ;
        RECT 10.010 6.520 10.150 6.530 ;
        RECT 12.910 6.520 13.050 6.530 ;
        RECT 15.810 6.520 15.950 6.530 ;
        RECT 18.710 6.520 18.850 6.530 ;
        RECT 21.610 6.520 21.750 6.530 ;
        RECT 0.775 6.320 0.850 6.460 ;
        RECT 0.990 6.270 1.065 6.410 ;
        RECT 1.695 6.330 1.755 6.410 ;
        POLYGON 1.695 6.330 1.755 6.330 1.755 6.270 ;
        RECT 1.910 6.320 1.985 6.460 ;
        RECT 3.675 6.320 3.750 6.460 ;
        RECT 3.890 6.270 3.965 6.410 ;
        RECT 4.595 6.330 4.655 6.410 ;
        POLYGON 4.595 6.330 4.655 6.330 4.655 6.270 ;
        RECT 4.810 6.320 4.885 6.460 ;
        RECT 6.575 6.320 6.650 6.460 ;
        RECT 6.790 6.270 6.865 6.410 ;
        RECT 7.495 6.330 7.555 6.410 ;
        POLYGON 7.495 6.330 7.555 6.330 7.555 6.270 ;
        RECT 7.710 6.320 7.785 6.460 ;
        RECT 9.475 6.320 9.550 6.460 ;
        RECT 9.690 6.270 9.765 6.410 ;
        RECT 10.395 6.330 10.455 6.410 ;
        POLYGON 10.395 6.330 10.455 6.330 10.455 6.270 ;
        RECT 10.610 6.320 10.685 6.460 ;
        RECT 12.375 6.320 12.450 6.460 ;
        RECT 12.590 6.270 12.665 6.410 ;
        RECT 13.295 6.330 13.355 6.410 ;
        POLYGON 13.295 6.330 13.355 6.330 13.355 6.270 ;
        RECT 13.510 6.320 13.585 6.460 ;
        RECT 15.275 6.320 15.350 6.460 ;
        RECT 15.490 6.270 15.565 6.410 ;
        RECT 16.195 6.330 16.255 6.410 ;
        POLYGON 16.195 6.330 16.255 6.330 16.255 6.270 ;
        RECT 16.410 6.320 16.485 6.460 ;
        RECT 18.175 6.320 18.250 6.460 ;
        RECT 18.390 6.270 18.465 6.410 ;
        RECT 19.095 6.330 19.155 6.410 ;
        POLYGON 19.095 6.330 19.155 6.330 19.155 6.270 ;
        RECT 19.310 6.320 19.385 6.460 ;
        RECT 21.075 6.320 21.150 6.460 ;
        RECT 21.290 6.270 21.365 6.410 ;
        RECT 21.995 6.330 22.055 6.410 ;
        POLYGON 21.995 6.330 22.055 6.330 22.055 6.270 ;
        RECT 22.210 6.320 22.285 6.460 ;
        RECT 0.720 5.800 0.870 5.970 ;
        RECT 1.110 5.935 1.260 6.105 ;
        RECT 1.500 5.935 1.650 6.105 ;
        RECT 1.890 5.800 2.040 5.970 ;
        RECT 3.620 5.800 3.770 5.970 ;
        RECT 4.010 5.935 4.160 6.105 ;
        RECT 4.400 5.935 4.550 6.105 ;
        RECT 4.790 5.800 4.940 5.970 ;
        RECT 6.520 5.800 6.670 5.970 ;
        RECT 6.910 5.935 7.060 6.105 ;
        RECT 7.300 5.935 7.450 6.105 ;
        RECT 7.690 5.800 7.840 5.970 ;
        RECT 9.420 5.800 9.570 5.970 ;
        RECT 9.810 5.935 9.960 6.105 ;
        RECT 10.200 5.935 10.350 6.105 ;
        RECT 10.590 5.800 10.740 5.970 ;
        RECT 12.320 5.800 12.470 5.970 ;
        RECT 12.710 5.935 12.860 6.105 ;
        RECT 13.100 5.935 13.250 6.105 ;
        RECT 13.490 5.800 13.640 5.970 ;
        RECT 15.220 5.800 15.370 5.970 ;
        RECT 15.610 5.935 15.760 6.105 ;
        RECT 16.000 5.935 16.150 6.105 ;
        RECT 16.390 5.800 16.540 5.970 ;
        RECT 18.120 5.800 18.270 5.970 ;
        RECT 18.510 5.935 18.660 6.105 ;
        RECT 18.900 5.935 19.050 6.105 ;
        RECT 19.290 5.800 19.440 5.970 ;
        RECT 21.020 5.800 21.170 5.970 ;
        RECT 21.410 5.935 21.560 6.105 ;
        RECT 21.800 5.935 21.950 6.105 ;
        RECT 22.190 5.800 22.340 5.970 ;
        RECT 0.985 5.715 1.035 5.750 ;
        POLYGON 1.035 5.750 1.070 5.715 1.035 5.715 ;
        RECT 0.985 5.590 1.070 5.715 ;
        RECT 1.690 5.590 1.775 5.750 ;
        RECT 3.885 5.715 3.935 5.750 ;
        POLYGON 3.935 5.750 3.970 5.715 3.935 5.715 ;
        RECT 3.885 5.590 3.970 5.715 ;
        RECT 4.590 5.590 4.675 5.750 ;
        RECT 6.785 5.715 6.835 5.750 ;
        POLYGON 6.835 5.750 6.870 5.715 6.835 5.715 ;
        RECT 6.785 5.590 6.870 5.715 ;
        RECT 7.490 5.590 7.575 5.750 ;
        RECT 9.685 5.715 9.735 5.750 ;
        POLYGON 9.735 5.750 9.770 5.715 9.735 5.715 ;
        RECT 9.685 5.590 9.770 5.715 ;
        RECT 10.390 5.590 10.475 5.750 ;
        RECT 12.585 5.715 12.635 5.750 ;
        POLYGON 12.635 5.750 12.670 5.715 12.635 5.715 ;
        RECT 12.585 5.590 12.670 5.715 ;
        RECT 13.290 5.590 13.375 5.750 ;
        RECT 15.485 5.715 15.535 5.750 ;
        POLYGON 15.535 5.750 15.570 5.715 15.535 5.715 ;
        RECT 15.485 5.590 15.570 5.715 ;
        RECT 16.190 5.590 16.275 5.750 ;
        RECT 18.385 5.715 18.435 5.750 ;
        POLYGON 18.435 5.750 18.470 5.715 18.435 5.715 ;
        RECT 18.385 5.590 18.470 5.715 ;
        RECT 19.090 5.590 19.175 5.750 ;
        RECT 21.285 5.715 21.335 5.750 ;
        POLYGON 21.335 5.750 21.370 5.715 21.335 5.715 ;
        RECT 21.285 5.590 21.370 5.715 ;
        RECT 21.990 5.590 22.075 5.750 ;
        RECT 1.300 5.180 1.460 5.250 ;
        RECT 4.200 5.180 4.360 5.250 ;
        RECT 7.100 5.180 7.260 5.250 ;
        RECT 10.000 5.180 10.160 5.250 ;
        RECT 12.900 5.180 13.060 5.250 ;
        RECT 15.800 5.180 15.960 5.250 ;
        RECT 18.700 5.180 18.860 5.250 ;
        RECT 21.600 5.180 21.760 5.250 ;
        RECT 1.310 5.170 1.450 5.180 ;
        RECT 4.210 5.170 4.350 5.180 ;
        RECT 7.110 5.170 7.250 5.180 ;
        RECT 10.010 5.170 10.150 5.180 ;
        RECT 12.910 5.170 13.050 5.180 ;
        RECT 15.810 5.170 15.950 5.180 ;
        RECT 18.710 5.170 18.850 5.180 ;
        RECT 21.610 5.170 21.750 5.180 ;
        RECT 0.775 4.970 0.850 5.110 ;
        RECT 0.990 4.920 1.065 5.060 ;
        RECT 1.695 4.980 1.755 5.060 ;
        POLYGON 1.695 4.980 1.755 4.980 1.755 4.920 ;
        RECT 1.910 4.970 1.985 5.110 ;
        RECT 3.675 4.970 3.750 5.110 ;
        RECT 3.890 4.920 3.965 5.060 ;
        RECT 4.595 4.980 4.655 5.060 ;
        POLYGON 4.595 4.980 4.655 4.980 4.655 4.920 ;
        RECT 4.810 4.970 4.885 5.110 ;
        RECT 6.575 4.970 6.650 5.110 ;
        RECT 6.790 4.920 6.865 5.060 ;
        RECT 7.495 4.980 7.555 5.060 ;
        POLYGON 7.495 4.980 7.555 4.980 7.555 4.920 ;
        RECT 7.710 4.970 7.785 5.110 ;
        RECT 9.475 4.970 9.550 5.110 ;
        RECT 9.690 4.920 9.765 5.060 ;
        RECT 10.395 4.980 10.455 5.060 ;
        POLYGON 10.395 4.980 10.455 4.980 10.455 4.920 ;
        RECT 10.610 4.970 10.685 5.110 ;
        RECT 12.375 4.970 12.450 5.110 ;
        RECT 12.590 4.920 12.665 5.060 ;
        RECT 13.295 4.980 13.355 5.060 ;
        POLYGON 13.295 4.980 13.355 4.980 13.355 4.920 ;
        RECT 13.510 4.970 13.585 5.110 ;
        RECT 15.275 4.970 15.350 5.110 ;
        RECT 15.490 4.920 15.565 5.060 ;
        RECT 16.195 4.980 16.255 5.060 ;
        POLYGON 16.195 4.980 16.255 4.980 16.255 4.920 ;
        RECT 16.410 4.970 16.485 5.110 ;
        RECT 18.175 4.970 18.250 5.110 ;
        RECT 18.390 4.920 18.465 5.060 ;
        RECT 19.095 4.980 19.155 5.060 ;
        POLYGON 19.095 4.980 19.155 4.980 19.155 4.920 ;
        RECT 19.310 4.970 19.385 5.110 ;
        RECT 21.075 4.970 21.150 5.110 ;
        RECT 21.290 4.920 21.365 5.060 ;
        RECT 21.995 4.980 22.055 5.060 ;
        POLYGON 21.995 4.980 22.055 4.980 22.055 4.920 ;
        RECT 22.210 4.970 22.285 5.110 ;
        RECT 0.720 4.450 0.870 4.620 ;
        RECT 1.110 4.585 1.260 4.755 ;
        RECT 1.500 4.585 1.650 4.755 ;
        RECT 1.890 4.450 2.040 4.620 ;
        RECT 3.620 4.450 3.770 4.620 ;
        RECT 4.010 4.585 4.160 4.755 ;
        RECT 4.400 4.585 4.550 4.755 ;
        RECT 4.790 4.450 4.940 4.620 ;
        RECT 6.520 4.450 6.670 4.620 ;
        RECT 6.910 4.585 7.060 4.755 ;
        RECT 7.300 4.585 7.450 4.755 ;
        RECT 7.690 4.450 7.840 4.620 ;
        RECT 9.420 4.450 9.570 4.620 ;
        RECT 9.810 4.585 9.960 4.755 ;
        RECT 10.200 4.585 10.350 4.755 ;
        RECT 10.590 4.450 10.740 4.620 ;
        RECT 12.320 4.450 12.470 4.620 ;
        RECT 12.710 4.585 12.860 4.755 ;
        RECT 13.100 4.585 13.250 4.755 ;
        RECT 13.490 4.450 13.640 4.620 ;
        RECT 15.220 4.450 15.370 4.620 ;
        RECT 15.610 4.585 15.760 4.755 ;
        RECT 16.000 4.585 16.150 4.755 ;
        RECT 16.390 4.450 16.540 4.620 ;
        RECT 18.120 4.450 18.270 4.620 ;
        RECT 18.510 4.585 18.660 4.755 ;
        RECT 18.900 4.585 19.050 4.755 ;
        RECT 19.290 4.450 19.440 4.620 ;
        RECT 21.020 4.450 21.170 4.620 ;
        RECT 21.410 4.585 21.560 4.755 ;
        RECT 21.800 4.585 21.950 4.755 ;
        RECT 22.190 4.450 22.340 4.620 ;
        RECT 0.985 4.365 1.035 4.400 ;
        POLYGON 1.035 4.400 1.070 4.365 1.035 4.365 ;
        RECT 0.985 4.240 1.070 4.365 ;
        RECT 1.690 4.240 1.775 4.400 ;
        RECT 3.885 4.365 3.935 4.400 ;
        POLYGON 3.935 4.400 3.970 4.365 3.935 4.365 ;
        RECT 3.885 4.240 3.970 4.365 ;
        RECT 4.590 4.240 4.675 4.400 ;
        RECT 6.785 4.365 6.835 4.400 ;
        POLYGON 6.835 4.400 6.870 4.365 6.835 4.365 ;
        RECT 6.785 4.240 6.870 4.365 ;
        RECT 7.490 4.240 7.575 4.400 ;
        RECT 9.685 4.365 9.735 4.400 ;
        POLYGON 9.735 4.400 9.770 4.365 9.735 4.365 ;
        RECT 9.685 4.240 9.770 4.365 ;
        RECT 10.390 4.240 10.475 4.400 ;
        RECT 12.585 4.365 12.635 4.400 ;
        POLYGON 12.635 4.400 12.670 4.365 12.635 4.365 ;
        RECT 12.585 4.240 12.670 4.365 ;
        RECT 13.290 4.240 13.375 4.400 ;
        RECT 15.485 4.365 15.535 4.400 ;
        POLYGON 15.535 4.400 15.570 4.365 15.535 4.365 ;
        RECT 15.485 4.240 15.570 4.365 ;
        RECT 16.190 4.240 16.275 4.400 ;
        RECT 18.385 4.365 18.435 4.400 ;
        POLYGON 18.435 4.400 18.470 4.365 18.435 4.365 ;
        RECT 18.385 4.240 18.470 4.365 ;
        RECT 19.090 4.240 19.175 4.400 ;
        RECT 21.285 4.365 21.335 4.400 ;
        POLYGON 21.335 4.400 21.370 4.365 21.335 4.365 ;
        RECT 21.285 4.240 21.370 4.365 ;
        RECT 21.990 4.240 22.075 4.400 ;
        RECT 1.300 3.830 1.460 3.900 ;
        RECT 4.200 3.830 4.360 3.900 ;
        RECT 7.100 3.830 7.260 3.900 ;
        RECT 10.000 3.830 10.160 3.900 ;
        RECT 12.900 3.830 13.060 3.900 ;
        RECT 15.800 3.830 15.960 3.900 ;
        RECT 18.700 3.830 18.860 3.900 ;
        RECT 21.600 3.830 21.760 3.900 ;
        RECT 1.310 3.820 1.450 3.830 ;
        RECT 4.210 3.820 4.350 3.830 ;
        RECT 7.110 3.820 7.250 3.830 ;
        RECT 10.010 3.820 10.150 3.830 ;
        RECT 12.910 3.820 13.050 3.830 ;
        RECT 15.810 3.820 15.950 3.830 ;
        RECT 18.710 3.820 18.850 3.830 ;
        RECT 21.610 3.820 21.750 3.830 ;
        RECT 0.775 3.620 0.850 3.760 ;
        RECT 0.990 3.570 1.065 3.710 ;
        RECT 1.695 3.630 1.755 3.710 ;
        POLYGON 1.695 3.630 1.755 3.630 1.755 3.570 ;
        RECT 1.910 3.620 1.985 3.760 ;
        RECT 3.675 3.620 3.750 3.760 ;
        RECT 3.890 3.570 3.965 3.710 ;
        RECT 4.595 3.630 4.655 3.710 ;
        POLYGON 4.595 3.630 4.655 3.630 4.655 3.570 ;
        RECT 4.810 3.620 4.885 3.760 ;
        RECT 6.575 3.620 6.650 3.760 ;
        RECT 6.790 3.570 6.865 3.710 ;
        RECT 7.495 3.630 7.555 3.710 ;
        POLYGON 7.495 3.630 7.555 3.630 7.555 3.570 ;
        RECT 7.710 3.620 7.785 3.760 ;
        RECT 9.475 3.620 9.550 3.760 ;
        RECT 9.690 3.570 9.765 3.710 ;
        RECT 10.395 3.630 10.455 3.710 ;
        POLYGON 10.395 3.630 10.455 3.630 10.455 3.570 ;
        RECT 10.610 3.620 10.685 3.760 ;
        RECT 12.375 3.620 12.450 3.760 ;
        RECT 12.590 3.570 12.665 3.710 ;
        RECT 13.295 3.630 13.355 3.710 ;
        POLYGON 13.295 3.630 13.355 3.630 13.355 3.570 ;
        RECT 13.510 3.620 13.585 3.760 ;
        RECT 15.275 3.620 15.350 3.760 ;
        RECT 15.490 3.570 15.565 3.710 ;
        RECT 16.195 3.630 16.255 3.710 ;
        POLYGON 16.195 3.630 16.255 3.630 16.255 3.570 ;
        RECT 16.410 3.620 16.485 3.760 ;
        RECT 18.175 3.620 18.250 3.760 ;
        RECT 18.390 3.570 18.465 3.710 ;
        RECT 19.095 3.630 19.155 3.710 ;
        POLYGON 19.095 3.630 19.155 3.630 19.155 3.570 ;
        RECT 19.310 3.620 19.385 3.760 ;
        RECT 21.075 3.620 21.150 3.760 ;
        RECT 21.290 3.570 21.365 3.710 ;
        RECT 21.995 3.630 22.055 3.710 ;
        POLYGON 21.995 3.630 22.055 3.630 22.055 3.570 ;
        RECT 22.210 3.620 22.285 3.760 ;
        RECT 0.720 3.100 0.870 3.270 ;
        RECT 1.110 3.235 1.260 3.405 ;
        RECT 1.500 3.235 1.650 3.405 ;
        RECT 1.890 3.100 2.040 3.270 ;
        RECT 3.620 3.100 3.770 3.270 ;
        RECT 4.010 3.235 4.160 3.405 ;
        RECT 4.400 3.235 4.550 3.405 ;
        RECT 4.790 3.100 4.940 3.270 ;
        RECT 6.520 3.100 6.670 3.270 ;
        RECT 6.910 3.235 7.060 3.405 ;
        RECT 7.300 3.235 7.450 3.405 ;
        RECT 7.690 3.100 7.840 3.270 ;
        RECT 9.420 3.100 9.570 3.270 ;
        RECT 9.810 3.235 9.960 3.405 ;
        RECT 10.200 3.235 10.350 3.405 ;
        RECT 10.590 3.100 10.740 3.270 ;
        RECT 12.320 3.100 12.470 3.270 ;
        RECT 12.710 3.235 12.860 3.405 ;
        RECT 13.100 3.235 13.250 3.405 ;
        RECT 13.490 3.100 13.640 3.270 ;
        RECT 15.220 3.100 15.370 3.270 ;
        RECT 15.610 3.235 15.760 3.405 ;
        RECT 16.000 3.235 16.150 3.405 ;
        RECT 16.390 3.100 16.540 3.270 ;
        RECT 18.120 3.100 18.270 3.270 ;
        RECT 18.510 3.235 18.660 3.405 ;
        RECT 18.900 3.235 19.050 3.405 ;
        RECT 19.290 3.100 19.440 3.270 ;
        RECT 21.020 3.100 21.170 3.270 ;
        RECT 21.410 3.235 21.560 3.405 ;
        RECT 21.800 3.235 21.950 3.405 ;
        RECT 22.190 3.100 22.340 3.270 ;
        RECT 0.985 3.015 1.035 3.050 ;
        POLYGON 1.035 3.050 1.070 3.015 1.035 3.015 ;
        RECT 0.985 2.890 1.070 3.015 ;
        RECT 1.690 2.890 1.775 3.050 ;
        RECT 3.885 3.015 3.935 3.050 ;
        POLYGON 3.935 3.050 3.970 3.015 3.935 3.015 ;
        RECT 3.885 2.890 3.970 3.015 ;
        RECT 4.590 2.890 4.675 3.050 ;
        RECT 6.785 3.015 6.835 3.050 ;
        POLYGON 6.835 3.050 6.870 3.015 6.835 3.015 ;
        RECT 6.785 2.890 6.870 3.015 ;
        RECT 7.490 2.890 7.575 3.050 ;
        RECT 9.685 3.015 9.735 3.050 ;
        POLYGON 9.735 3.050 9.770 3.015 9.735 3.015 ;
        RECT 9.685 2.890 9.770 3.015 ;
        RECT 10.390 2.890 10.475 3.050 ;
        RECT 12.585 3.015 12.635 3.050 ;
        POLYGON 12.635 3.050 12.670 3.015 12.635 3.015 ;
        RECT 12.585 2.890 12.670 3.015 ;
        RECT 13.290 2.890 13.375 3.050 ;
        RECT 15.485 3.015 15.535 3.050 ;
        POLYGON 15.535 3.050 15.570 3.015 15.535 3.015 ;
        RECT 15.485 2.890 15.570 3.015 ;
        RECT 16.190 2.890 16.275 3.050 ;
        RECT 18.385 3.015 18.435 3.050 ;
        POLYGON 18.435 3.050 18.470 3.015 18.435 3.015 ;
        RECT 18.385 2.890 18.470 3.015 ;
        RECT 19.090 2.890 19.175 3.050 ;
        RECT 21.285 3.015 21.335 3.050 ;
        POLYGON 21.335 3.050 21.370 3.015 21.335 3.015 ;
        RECT 21.285 2.890 21.370 3.015 ;
        RECT 21.990 2.890 22.075 3.050 ;
        RECT 1.300 2.480 1.460 2.550 ;
        RECT 4.200 2.480 4.360 2.550 ;
        RECT 7.100 2.480 7.260 2.550 ;
        RECT 10.000 2.480 10.160 2.550 ;
        RECT 12.900 2.480 13.060 2.550 ;
        RECT 15.800 2.480 15.960 2.550 ;
        RECT 18.700 2.480 18.860 2.550 ;
        RECT 21.600 2.480 21.760 2.550 ;
        RECT 1.310 2.470 1.450 2.480 ;
        RECT 4.210 2.470 4.350 2.480 ;
        RECT 7.110 2.470 7.250 2.480 ;
        RECT 10.010 2.470 10.150 2.480 ;
        RECT 12.910 2.470 13.050 2.480 ;
        RECT 15.810 2.470 15.950 2.480 ;
        RECT 18.710 2.470 18.850 2.480 ;
        RECT 21.610 2.470 21.750 2.480 ;
        RECT 0.775 2.270 0.850 2.410 ;
        RECT 0.990 2.220 1.065 2.360 ;
        RECT 1.695 2.280 1.755 2.360 ;
        POLYGON 1.695 2.280 1.755 2.280 1.755 2.220 ;
        RECT 1.910 2.270 1.985 2.410 ;
        RECT 3.675 2.270 3.750 2.410 ;
        RECT 3.890 2.220 3.965 2.360 ;
        RECT 4.595 2.280 4.655 2.360 ;
        POLYGON 4.595 2.280 4.655 2.280 4.655 2.220 ;
        RECT 4.810 2.270 4.885 2.410 ;
        RECT 6.575 2.270 6.650 2.410 ;
        RECT 6.790 2.220 6.865 2.360 ;
        RECT 7.495 2.280 7.555 2.360 ;
        POLYGON 7.495 2.280 7.555 2.280 7.555 2.220 ;
        RECT 7.710 2.270 7.785 2.410 ;
        RECT 9.475 2.270 9.550 2.410 ;
        RECT 9.690 2.220 9.765 2.360 ;
        RECT 10.395 2.280 10.455 2.360 ;
        POLYGON 10.395 2.280 10.455 2.280 10.455 2.220 ;
        RECT 10.610 2.270 10.685 2.410 ;
        RECT 12.375 2.270 12.450 2.410 ;
        RECT 12.590 2.220 12.665 2.360 ;
        RECT 13.295 2.280 13.355 2.360 ;
        POLYGON 13.295 2.280 13.355 2.280 13.355 2.220 ;
        RECT 13.510 2.270 13.585 2.410 ;
        RECT 15.275 2.270 15.350 2.410 ;
        RECT 15.490 2.220 15.565 2.360 ;
        RECT 16.195 2.280 16.255 2.360 ;
        POLYGON 16.195 2.280 16.255 2.280 16.255 2.220 ;
        RECT 16.410 2.270 16.485 2.410 ;
        RECT 18.175 2.270 18.250 2.410 ;
        RECT 18.390 2.220 18.465 2.360 ;
        RECT 19.095 2.280 19.155 2.360 ;
        POLYGON 19.095 2.280 19.155 2.280 19.155 2.220 ;
        RECT 19.310 2.270 19.385 2.410 ;
        RECT 21.075 2.270 21.150 2.410 ;
        RECT 21.290 2.220 21.365 2.360 ;
        RECT 21.995 2.280 22.055 2.360 ;
        POLYGON 21.995 2.280 22.055 2.280 22.055 2.220 ;
        RECT 22.210 2.270 22.285 2.410 ;
        RECT 0.720 1.750 0.870 1.920 ;
        RECT 1.110 1.885 1.260 2.055 ;
        RECT 1.500 1.885 1.650 2.055 ;
        RECT 1.890 1.750 2.040 1.920 ;
        RECT 3.620 1.750 3.770 1.920 ;
        RECT 4.010 1.885 4.160 2.055 ;
        RECT 4.400 1.885 4.550 2.055 ;
        RECT 4.790 1.750 4.940 1.920 ;
        RECT 6.520 1.750 6.670 1.920 ;
        RECT 6.910 1.885 7.060 2.055 ;
        RECT 7.300 1.885 7.450 2.055 ;
        RECT 7.690 1.750 7.840 1.920 ;
        RECT 9.420 1.750 9.570 1.920 ;
        RECT 9.810 1.885 9.960 2.055 ;
        RECT 10.200 1.885 10.350 2.055 ;
        RECT 10.590 1.750 10.740 1.920 ;
        RECT 12.320 1.750 12.470 1.920 ;
        RECT 12.710 1.885 12.860 2.055 ;
        RECT 13.100 1.885 13.250 2.055 ;
        RECT 13.490 1.750 13.640 1.920 ;
        RECT 15.220 1.750 15.370 1.920 ;
        RECT 15.610 1.885 15.760 2.055 ;
        RECT 16.000 1.885 16.150 2.055 ;
        RECT 16.390 1.750 16.540 1.920 ;
        RECT 18.120 1.750 18.270 1.920 ;
        RECT 18.510 1.885 18.660 2.055 ;
        RECT 18.900 1.885 19.050 2.055 ;
        RECT 19.290 1.750 19.440 1.920 ;
        RECT 21.020 1.750 21.170 1.920 ;
        RECT 21.410 1.885 21.560 2.055 ;
        RECT 21.800 1.885 21.950 2.055 ;
        RECT 22.190 1.750 22.340 1.920 ;
        RECT 0.985 1.665 1.035 1.700 ;
        POLYGON 1.035 1.700 1.070 1.665 1.035 1.665 ;
        RECT 0.985 1.540 1.070 1.665 ;
        RECT 1.690 1.540 1.775 1.700 ;
        RECT 3.885 1.665 3.935 1.700 ;
        POLYGON 3.935 1.700 3.970 1.665 3.935 1.665 ;
        RECT 3.885 1.540 3.970 1.665 ;
        RECT 4.590 1.540 4.675 1.700 ;
        RECT 6.785 1.665 6.835 1.700 ;
        POLYGON 6.835 1.700 6.870 1.665 6.835 1.665 ;
        RECT 6.785 1.540 6.870 1.665 ;
        RECT 7.490 1.540 7.575 1.700 ;
        RECT 9.685 1.665 9.735 1.700 ;
        POLYGON 9.735 1.700 9.770 1.665 9.735 1.665 ;
        RECT 9.685 1.540 9.770 1.665 ;
        RECT 10.390 1.540 10.475 1.700 ;
        RECT 12.585 1.665 12.635 1.700 ;
        POLYGON 12.635 1.700 12.670 1.665 12.635 1.665 ;
        RECT 12.585 1.540 12.670 1.665 ;
        RECT 13.290 1.540 13.375 1.700 ;
        RECT 15.485 1.665 15.535 1.700 ;
        POLYGON 15.535 1.700 15.570 1.665 15.535 1.665 ;
        RECT 15.485 1.540 15.570 1.665 ;
        RECT 16.190 1.540 16.275 1.700 ;
        RECT 18.385 1.665 18.435 1.700 ;
        POLYGON 18.435 1.700 18.470 1.665 18.435 1.665 ;
        RECT 18.385 1.540 18.470 1.665 ;
        RECT 19.090 1.540 19.175 1.700 ;
        RECT 21.285 1.665 21.335 1.700 ;
        POLYGON 21.335 1.700 21.370 1.665 21.335 1.665 ;
        RECT 21.285 1.540 21.370 1.665 ;
        RECT 21.990 1.540 22.075 1.700 ;
        RECT 1.300 1.130 1.460 1.200 ;
        RECT 4.200 1.130 4.360 1.200 ;
        RECT 7.100 1.130 7.260 1.200 ;
        RECT 10.000 1.130 10.160 1.200 ;
        RECT 12.900 1.130 13.060 1.200 ;
        RECT 15.800 1.130 15.960 1.200 ;
        RECT 18.700 1.130 18.860 1.200 ;
        RECT 21.600 1.130 21.760 1.200 ;
        RECT 1.310 1.120 1.450 1.130 ;
        RECT 4.210 1.120 4.350 1.130 ;
        RECT 7.110 1.120 7.250 1.130 ;
        RECT 10.010 1.120 10.150 1.130 ;
        RECT 12.910 1.120 13.050 1.130 ;
        RECT 15.810 1.120 15.950 1.130 ;
        RECT 18.710 1.120 18.850 1.130 ;
        RECT 21.610 1.120 21.750 1.130 ;
        RECT 0.775 0.920 0.850 1.060 ;
        RECT 0.990 0.870 1.065 1.010 ;
        RECT 1.695 0.930 1.755 1.010 ;
        POLYGON 1.695 0.930 1.755 0.930 1.755 0.870 ;
        RECT 1.910 0.920 1.985 1.060 ;
        RECT 3.675 0.920 3.750 1.060 ;
        RECT 3.890 0.870 3.965 1.010 ;
        RECT 4.595 0.930 4.655 1.010 ;
        POLYGON 4.595 0.930 4.655 0.930 4.655 0.870 ;
        RECT 4.810 0.920 4.885 1.060 ;
        RECT 6.575 0.920 6.650 1.060 ;
        RECT 6.790 0.870 6.865 1.010 ;
        RECT 7.495 0.930 7.555 1.010 ;
        POLYGON 7.495 0.930 7.555 0.930 7.555 0.870 ;
        RECT 7.710 0.920 7.785 1.060 ;
        RECT 9.475 0.920 9.550 1.060 ;
        RECT 9.690 0.870 9.765 1.010 ;
        RECT 10.395 0.930 10.455 1.010 ;
        POLYGON 10.395 0.930 10.455 0.930 10.455 0.870 ;
        RECT 10.610 0.920 10.685 1.060 ;
        RECT 12.375 0.920 12.450 1.060 ;
        RECT 12.590 0.870 12.665 1.010 ;
        RECT 13.295 0.930 13.355 1.010 ;
        POLYGON 13.295 0.930 13.355 0.930 13.355 0.870 ;
        RECT 13.510 0.920 13.585 1.060 ;
        RECT 15.275 0.920 15.350 1.060 ;
        RECT 15.490 0.870 15.565 1.010 ;
        RECT 16.195 0.930 16.255 1.010 ;
        POLYGON 16.195 0.930 16.255 0.930 16.255 0.870 ;
        RECT 16.410 0.920 16.485 1.060 ;
        RECT 18.175 0.920 18.250 1.060 ;
        RECT 18.390 0.870 18.465 1.010 ;
        RECT 19.095 0.930 19.155 1.010 ;
        POLYGON 19.095 0.930 19.155 0.930 19.155 0.870 ;
        RECT 19.310 0.920 19.385 1.060 ;
        RECT 21.075 0.920 21.150 1.060 ;
        RECT 21.290 0.870 21.365 1.010 ;
        RECT 21.995 0.930 22.055 1.010 ;
        POLYGON 21.995 0.930 22.055 0.930 22.055 0.870 ;
        RECT 22.210 0.920 22.285 1.060 ;
        RECT 0.720 0.400 0.870 0.570 ;
        RECT 1.110 0.535 1.260 0.705 ;
        RECT 1.500 0.535 1.650 0.705 ;
        RECT 1.890 0.400 2.040 0.570 ;
        RECT 3.620 0.400 3.770 0.570 ;
        RECT 4.010 0.535 4.160 0.705 ;
        RECT 4.400 0.535 4.550 0.705 ;
        RECT 4.790 0.400 4.940 0.570 ;
        RECT 6.520 0.400 6.670 0.570 ;
        RECT 6.910 0.535 7.060 0.705 ;
        RECT 7.300 0.535 7.450 0.705 ;
        RECT 7.690 0.400 7.840 0.570 ;
        RECT 9.420 0.400 9.570 0.570 ;
        RECT 9.810 0.535 9.960 0.705 ;
        RECT 10.200 0.535 10.350 0.705 ;
        RECT 10.590 0.400 10.740 0.570 ;
        RECT 12.320 0.400 12.470 0.570 ;
        RECT 12.710 0.535 12.860 0.705 ;
        RECT 13.100 0.535 13.250 0.705 ;
        RECT 13.490 0.400 13.640 0.570 ;
        RECT 15.220 0.400 15.370 0.570 ;
        RECT 15.610 0.535 15.760 0.705 ;
        RECT 16.000 0.535 16.150 0.705 ;
        RECT 16.390 0.400 16.540 0.570 ;
        RECT 18.120 0.400 18.270 0.570 ;
        RECT 18.510 0.535 18.660 0.705 ;
        RECT 18.900 0.535 19.050 0.705 ;
        RECT 19.290 0.400 19.440 0.570 ;
        RECT 21.020 0.400 21.170 0.570 ;
        RECT 21.410 0.535 21.560 0.705 ;
        RECT 21.800 0.535 21.950 0.705 ;
        RECT 22.190 0.400 22.340 0.570 ;
        RECT 0.985 0.315 1.035 0.350 ;
        POLYGON 1.035 0.350 1.070 0.315 1.035 0.315 ;
        RECT 0.985 0.190 1.070 0.315 ;
        RECT 1.690 0.190 1.775 0.350 ;
        RECT 3.885 0.315 3.935 0.350 ;
        POLYGON 3.935 0.350 3.970 0.315 3.935 0.315 ;
        RECT 3.885 0.190 3.970 0.315 ;
        RECT 4.590 0.190 4.675 0.350 ;
        RECT 6.785 0.315 6.835 0.350 ;
        POLYGON 6.835 0.350 6.870 0.315 6.835 0.315 ;
        RECT 6.785 0.190 6.870 0.315 ;
        RECT 7.490 0.190 7.575 0.350 ;
        RECT 9.685 0.315 9.735 0.350 ;
        POLYGON 9.735 0.350 9.770 0.315 9.735 0.315 ;
        RECT 9.685 0.190 9.770 0.315 ;
        RECT 10.390 0.190 10.475 0.350 ;
        RECT 12.585 0.315 12.635 0.350 ;
        POLYGON 12.635 0.350 12.670 0.315 12.635 0.315 ;
        RECT 12.585 0.190 12.670 0.315 ;
        RECT 13.290 0.190 13.375 0.350 ;
        RECT 15.485 0.315 15.535 0.350 ;
        POLYGON 15.535 0.350 15.570 0.315 15.535 0.315 ;
        RECT 15.485 0.190 15.570 0.315 ;
        RECT 16.190 0.190 16.275 0.350 ;
        RECT 18.385 0.315 18.435 0.350 ;
        POLYGON 18.435 0.350 18.470 0.315 18.435 0.315 ;
        RECT 18.385 0.190 18.470 0.315 ;
        RECT 19.090 0.190 19.175 0.350 ;
        RECT 21.285 0.315 21.335 0.350 ;
        POLYGON 21.335 0.350 21.370 0.315 21.335 0.315 ;
        RECT 21.285 0.190 21.370 0.315 ;
        RECT 21.990 0.190 22.075 0.350 ;
      LAYER met1 ;
        RECT 0.000 20.030 23.060 20.100 ;
        RECT 0.000 18.680 23.060 18.750 ;
        RECT 0.000 17.330 23.060 17.400 ;
        RECT 0.000 15.980 23.060 16.050 ;
        RECT 0.000 14.630 23.060 14.700 ;
        RECT 0.000 13.280 23.060 13.350 ;
        RECT 0.000 11.930 23.060 12.000 ;
        RECT 0.000 10.580 23.060 10.650 ;
        RECT 0.000 9.230 23.060 9.300 ;
        RECT 0.000 7.880 23.060 7.950 ;
        RECT 0.000 6.530 23.060 6.600 ;
        RECT 0.000 5.180 23.060 5.250 ;
        RECT 0.000 3.830 23.060 3.900 ;
        RECT 0.000 2.480 23.060 2.550 ;
        RECT 0.000 1.130 23.060 1.200 ;
  END
END 10T_16x8_magic
END LIBRARY

