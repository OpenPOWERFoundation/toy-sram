magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< pwell >>
rect 10 76 526 458
<< nmos >>
rect 204 102 240 432
rect 296 102 332 432
<< ndiff >>
rect 148 420 204 432
rect 148 386 159 420
rect 193 386 204 420
rect 148 352 204 386
rect 148 318 159 352
rect 193 318 204 352
rect 148 284 204 318
rect 148 250 159 284
rect 193 250 204 284
rect 148 216 204 250
rect 148 182 159 216
rect 193 182 204 216
rect 148 148 204 182
rect 148 114 159 148
rect 193 114 204 148
rect 148 102 204 114
rect 240 420 296 432
rect 240 386 251 420
rect 285 386 296 420
rect 240 352 296 386
rect 240 318 251 352
rect 285 318 296 352
rect 240 284 296 318
rect 240 250 251 284
rect 285 250 296 284
rect 240 216 296 250
rect 240 182 251 216
rect 285 182 296 216
rect 240 148 296 182
rect 240 114 251 148
rect 285 114 296 148
rect 240 102 296 114
rect 332 420 388 432
rect 332 386 343 420
rect 377 386 388 420
rect 332 352 388 386
rect 332 318 343 352
rect 377 318 388 352
rect 332 284 388 318
rect 332 250 343 284
rect 377 250 388 284
rect 332 216 388 250
rect 332 182 343 216
rect 377 182 388 216
rect 332 148 388 182
rect 332 114 343 148
rect 377 114 388 148
rect 332 102 388 114
<< ndiffc >>
rect 159 386 193 420
rect 159 318 193 352
rect 159 250 193 284
rect 159 182 193 216
rect 159 114 193 148
rect 251 386 285 420
rect 251 318 285 352
rect 251 250 285 284
rect 251 182 285 216
rect 251 114 285 148
rect 343 386 377 420
rect 343 318 377 352
rect 343 250 377 284
rect 343 182 377 216
rect 343 114 377 148
<< psubdiff >>
rect 36 386 94 432
rect 36 352 48 386
rect 82 352 94 386
rect 36 318 94 352
rect 36 284 48 318
rect 82 284 94 318
rect 36 250 94 284
rect 36 216 48 250
rect 82 216 94 250
rect 36 182 94 216
rect 36 148 48 182
rect 82 148 94 182
rect 36 102 94 148
rect 442 386 500 432
rect 442 352 454 386
rect 488 352 500 386
rect 442 318 500 352
rect 442 284 454 318
rect 488 284 500 318
rect 442 250 500 284
rect 442 216 454 250
rect 488 216 500 250
rect 442 182 500 216
rect 442 148 454 182
rect 488 148 500 182
rect 442 102 500 148
<< psubdiffcont >>
rect 48 352 82 386
rect 48 284 82 318
rect 48 216 82 250
rect 48 148 82 182
rect 454 352 488 386
rect 454 284 488 318
rect 454 216 488 250
rect 454 148 488 182
<< poly >>
rect 167 504 369 524
rect 167 470 183 504
rect 217 470 251 504
rect 285 470 319 504
rect 353 470 369 504
rect 167 454 369 470
rect 204 432 240 454
rect 296 432 332 454
rect 204 80 240 102
rect 296 80 332 102
rect 167 64 369 80
rect 167 30 183 64
rect 217 30 251 64
rect 285 30 319 64
rect 353 30 369 64
rect 167 10 369 30
<< polycont >>
rect 183 470 217 504
rect 251 470 285 504
rect 319 470 353 504
rect 183 30 217 64
rect 251 30 285 64
rect 319 30 353 64
<< locali >>
rect 167 470 179 504
rect 217 470 251 504
rect 285 470 319 504
rect 357 470 369 504
rect 159 420 193 436
rect 48 392 82 402
rect 48 320 82 352
rect 48 250 82 284
rect 48 182 82 214
rect 48 132 82 142
rect 159 352 193 358
rect 159 284 193 286
rect 159 248 193 250
rect 159 176 193 182
rect 159 98 193 114
rect 251 420 285 436
rect 251 352 285 358
rect 251 284 285 286
rect 251 248 285 250
rect 251 176 285 182
rect 251 98 285 114
rect 343 420 377 436
rect 343 352 377 358
rect 343 284 377 286
rect 343 248 377 250
rect 343 176 377 182
rect 454 392 488 402
rect 454 320 488 352
rect 454 250 488 284
rect 454 182 488 214
rect 454 132 488 142
rect 343 98 377 114
rect 167 30 179 64
rect 217 30 251 64
rect 285 30 319 64
rect 357 30 369 64
<< viali >>
rect 179 470 183 504
rect 183 470 213 504
rect 251 470 285 504
rect 323 470 353 504
rect 353 470 357 504
rect 48 386 82 392
rect 48 358 82 386
rect 48 318 82 320
rect 48 286 82 318
rect 48 216 82 248
rect 48 214 82 216
rect 48 148 82 176
rect 48 142 82 148
rect 159 386 193 392
rect 159 358 193 386
rect 159 318 193 320
rect 159 286 193 318
rect 159 216 193 248
rect 159 214 193 216
rect 159 148 193 176
rect 159 142 193 148
rect 251 386 285 392
rect 251 358 285 386
rect 251 318 285 320
rect 251 286 285 318
rect 251 216 285 248
rect 251 214 285 216
rect 251 148 285 176
rect 251 142 285 148
rect 343 386 377 392
rect 343 358 377 386
rect 343 318 377 320
rect 343 286 377 318
rect 343 216 377 248
rect 343 214 377 216
rect 343 148 377 176
rect 343 142 377 148
rect 454 386 488 392
rect 454 358 488 386
rect 454 318 488 320
rect 454 286 488 318
rect 454 216 488 248
rect 454 214 488 216
rect 454 148 488 176
rect 454 142 488 148
rect 179 30 183 64
rect 183 30 213 64
rect 251 30 285 64
rect 323 30 353 64
rect 353 30 357 64
<< metal1 >>
rect 167 504 369 524
rect 167 470 179 504
rect 213 470 251 504
rect 285 470 323 504
rect 357 470 369 504
rect 167 458 369 470
rect 36 392 94 420
rect 36 358 48 392
rect 82 358 94 392
rect 36 320 94 358
rect 36 286 48 320
rect 82 286 94 320
rect 36 248 94 286
rect 36 214 48 248
rect 82 214 94 248
rect 36 176 94 214
rect 36 142 48 176
rect 82 142 94 176
rect 36 114 94 142
rect 150 392 202 420
rect 150 358 159 392
rect 193 358 202 392
rect 150 320 202 358
rect 150 286 159 320
rect 193 286 202 320
rect 150 248 202 286
rect 150 236 159 248
rect 193 236 202 248
rect 150 176 202 184
rect 150 172 159 176
rect 193 172 202 176
rect 150 114 202 120
rect 242 414 294 420
rect 242 358 251 362
rect 285 358 294 362
rect 242 350 294 358
rect 242 286 251 298
rect 285 286 294 298
rect 242 248 294 286
rect 242 214 251 248
rect 285 214 294 248
rect 242 176 294 214
rect 242 142 251 176
rect 285 142 294 176
rect 242 114 294 142
rect 334 392 386 420
rect 334 358 343 392
rect 377 358 386 392
rect 334 320 386 358
rect 334 286 343 320
rect 377 286 386 320
rect 334 248 386 286
rect 334 236 343 248
rect 377 236 386 248
rect 334 176 386 184
rect 334 172 343 176
rect 377 172 386 176
rect 334 114 386 120
rect 442 392 500 420
rect 442 358 454 392
rect 488 358 500 392
rect 442 320 500 358
rect 442 286 454 320
rect 488 286 500 320
rect 442 248 500 286
rect 442 214 454 248
rect 488 214 500 248
rect 442 176 500 214
rect 442 142 454 176
rect 488 142 500 176
rect 442 114 500 142
rect 167 64 369 76
rect 167 30 179 64
rect 213 30 251 64
rect 285 30 323 64
rect 357 30 369 64
rect 167 10 369 30
<< via1 >>
rect 150 214 159 236
rect 159 214 193 236
rect 193 214 202 236
rect 150 184 202 214
rect 150 142 159 172
rect 159 142 193 172
rect 193 142 202 172
rect 150 120 202 142
rect 242 392 294 414
rect 242 362 251 392
rect 251 362 285 392
rect 285 362 294 392
rect 242 320 294 350
rect 242 298 251 320
rect 251 298 285 320
rect 285 298 294 320
rect 334 214 343 236
rect 343 214 377 236
rect 377 214 386 236
rect 334 184 386 214
rect 334 142 343 172
rect 343 142 377 172
rect 377 142 386 172
rect 334 120 386 142
<< metal2 >>
rect 10 414 526 420
rect 10 362 242 414
rect 294 362 526 414
rect 10 350 526 362
rect 10 298 242 350
rect 294 298 526 350
rect 10 292 526 298
rect 10 236 526 242
rect 10 184 150 236
rect 202 184 334 236
rect 386 184 526 236
rect 10 172 526 184
rect 10 120 150 172
rect 202 120 334 172
rect 386 120 526 172
rect 10 114 526 120
<< labels >>
flabel metal2 s 10 114 30 242 7 FreeSans 300 180 0 0 SOURCE
port 3 nsew
flabel metal2 s 10 292 30 420 7 FreeSans 300 180 0 0 DRAIN
port 1 nsew
flabel metal1 s 36 114 94 130 3 FreeSans 300 90 0 0 SUBSTRATE
port 4 nsew
flabel metal1 s 442 114 500 130 3 FreeSans 300 90 0 0 SUBSTRATE
port 4 nsew
flabel metal1 s 167 10 369 76 0 FreeSans 300 0 0 0 GATE
port 2 nsew
flabel metal1 s 167 458 369 524 0 FreeSans 300 0 0 0 GATE
port 2 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 4001922
string GDS_START 3994322
<< end >>
