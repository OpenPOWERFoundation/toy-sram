magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< locali >>
rect 181 1150 193 1184
rect 227 1150 265 1184
rect 299 1150 337 1184
rect 371 1150 383 1184
rect 181 30 193 64
rect 227 30 265 64
rect 299 30 337 64
rect 371 30 383 64
<< viali >>
rect 193 1150 227 1184
rect 265 1150 299 1184
rect 337 1150 371 1184
rect 193 30 227 64
rect 265 30 299 64
rect 337 30 371 64
<< obsli1 >>
rect 48 1020 82 1058
rect 48 948 82 986
rect 48 876 82 914
rect 48 804 82 842
rect 48 732 82 770
rect 48 660 82 698
rect 48 588 82 626
rect 48 516 82 554
rect 48 444 82 482
rect 48 372 82 410
rect 48 300 82 338
rect 48 228 82 266
rect 48 122 82 194
rect 159 98 193 1116
rect 265 98 299 1116
rect 371 98 405 1116
rect 482 1020 516 1058
rect 482 948 516 986
rect 482 876 516 914
rect 482 804 516 842
rect 482 732 516 770
rect 482 660 516 698
rect 482 588 516 626
rect 482 516 516 554
rect 482 444 516 482
rect 482 372 516 410
rect 482 300 516 338
rect 482 228 516 266
rect 482 122 516 194
<< obsli1c >>
rect 48 1058 82 1092
rect 48 986 82 1020
rect 48 914 82 948
rect 48 842 82 876
rect 48 770 82 804
rect 48 698 82 732
rect 48 626 82 660
rect 48 554 82 588
rect 48 482 82 516
rect 48 410 82 444
rect 48 338 82 372
rect 48 266 82 300
rect 48 194 82 228
rect 482 1058 516 1092
rect 482 986 516 1020
rect 482 914 516 948
rect 482 842 516 876
rect 482 770 516 804
rect 482 698 516 732
rect 482 626 516 660
rect 482 554 516 588
rect 482 482 516 516
rect 482 410 516 444
rect 482 338 516 372
rect 482 266 516 300
rect 482 194 516 228
<< metal1 >>
rect 181 1184 383 1204
rect 181 1150 193 1184
rect 227 1150 265 1184
rect 299 1150 337 1184
rect 371 1150 383 1184
rect 181 1138 383 1150
rect 36 1092 94 1104
rect 36 1058 48 1092
rect 82 1058 94 1092
rect 36 1020 94 1058
rect 36 986 48 1020
rect 82 986 94 1020
rect 36 948 94 986
rect 36 914 48 948
rect 82 914 94 948
rect 36 876 94 914
rect 36 842 48 876
rect 82 842 94 876
rect 36 804 94 842
rect 36 770 48 804
rect 82 770 94 804
rect 36 732 94 770
rect 36 698 48 732
rect 82 698 94 732
rect 36 660 94 698
rect 36 626 48 660
rect 82 626 94 660
rect 36 588 94 626
rect 36 554 48 588
rect 82 554 94 588
rect 36 516 94 554
rect 36 482 48 516
rect 82 482 94 516
rect 36 444 94 482
rect 36 410 48 444
rect 82 410 94 444
rect 36 372 94 410
rect 36 338 48 372
rect 82 338 94 372
rect 36 300 94 338
rect 36 266 48 300
rect 82 266 94 300
rect 36 228 94 266
rect 36 194 48 228
rect 82 194 94 228
rect 36 110 94 194
rect 470 1092 528 1104
rect 470 1058 482 1092
rect 516 1058 528 1092
rect 470 1020 528 1058
rect 470 986 482 1020
rect 516 986 528 1020
rect 470 948 528 986
rect 470 914 482 948
rect 516 914 528 948
rect 470 876 528 914
rect 470 842 482 876
rect 516 842 528 876
rect 470 804 528 842
rect 470 770 482 804
rect 516 770 528 804
rect 470 732 528 770
rect 470 698 482 732
rect 516 698 528 732
rect 470 660 528 698
rect 470 626 482 660
rect 516 626 528 660
rect 470 588 528 626
rect 470 554 482 588
rect 516 554 528 588
rect 470 516 528 554
rect 470 482 482 516
rect 516 482 528 516
rect 470 444 528 482
rect 470 410 482 444
rect 516 410 528 444
rect 470 372 528 410
rect 470 338 482 372
rect 516 338 528 372
rect 470 300 528 338
rect 470 266 482 300
rect 516 266 528 300
rect 470 228 528 266
rect 470 194 482 228
rect 516 194 528 228
rect 470 110 528 194
rect 181 64 383 76
rect 181 30 193 64
rect 227 30 265 64
rect 299 30 337 64
rect 371 30 383 64
rect 181 10 383 30
<< obsm1 >>
rect 150 110 202 1104
rect 256 110 308 1104
rect 362 110 414 1104
<< metal2 >>
rect 10 632 554 1104
rect 10 110 554 582
<< labels >>
rlabel metal2 s 10 632 554 1104 6 DRAIN
port 1 nsew
rlabel viali s 337 1150 371 1184 6 GATE
port 2 nsew
rlabel viali s 337 30 371 64 6 GATE
port 2 nsew
rlabel viali s 265 1150 299 1184 6 GATE
port 2 nsew
rlabel viali s 265 30 299 64 6 GATE
port 2 nsew
rlabel viali s 193 1150 227 1184 6 GATE
port 2 nsew
rlabel viali s 193 30 227 64 6 GATE
port 2 nsew
rlabel locali s 181 1150 383 1184 6 GATE
port 2 nsew
rlabel locali s 181 30 383 64 6 GATE
port 2 nsew
rlabel metal1 s 181 1138 383 1204 6 GATE
port 2 nsew
rlabel metal1 s 181 10 383 76 6 GATE
port 2 nsew
rlabel metal2 s 10 110 554 582 6 SOURCE
port 3 nsew
rlabel metal1 s 36 110 94 1104 6 SUBSTRATE
port 4 nsew
rlabel metal1 s 470 110 528 1104 6 SUBSTRATE
port 4 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 10 10 554 1204
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 5276298
string GDS_START 5260890
<< end >>
