magic
tech sky130A
magscale 1 2
timestamp 1656023017
<< pwell >>
rect 74 -896 89 -868
rect 464 -896 479 -867
rect 0 -1042 15 -1000
rect 537 -1042 552 -1000
rect 580 -1042 595 -1000
<< ndiffc >>
rect 74 -896 89 -868
rect 464 -896 479 -867
rect 654 -896 669 -868
rect 1044 -896 1059 -867
rect 1234 -896 1249 -868
rect 1624 -896 1639 -867
rect 1814 -896 1829 -868
rect 2204 -896 2219 -867
rect 2394 -896 2409 -868
rect 2784 -896 2799 -867
rect 2974 -896 2989 -868
rect 3364 -896 3379 -867
rect 3554 -896 3569 -868
rect 3944 -896 3959 -867
rect 4134 -896 4149 -868
rect 4524 -896 4539 -867
rect 0 -1042 15 -1000
rect 537 -1042 552 -1000
rect 580 -1042 595 -1000
rect 1117 -1042 1132 -1000
rect 1160 -1042 1175 -1000
rect 1697 -1042 1712 -1000
rect 1740 -1042 1755 -1000
rect 2277 -1042 2292 -1000
rect 2320 -1042 2335 -1000
rect 2857 -1042 2872 -1000
rect 2900 -1042 2915 -1000
rect 3437 -1042 3452 -1000
rect 3480 -1042 3495 -1000
rect 4017 -1042 4032 -1000
rect 4060 -1042 4075 -1000
rect 4597 -1042 4612 -1000
<< poly >>
rect 0 1050 30 1080
rect 0 780 30 810
rect 0 510 30 540
rect 0 240 30 270
rect 0 -30 30 0
rect 0 -300 30 -270
rect 0 -570 30 -540
rect 0 -840 30 -810
<< metal1 >>
rect 0 1036 15 1050
rect 0 912 15 946
rect 0 810 15 824
rect 0 766 15 780
rect 0 642 15 676
rect 0 540 15 554
rect 0 496 15 510
rect 0 372 15 406
rect 0 270 15 284
rect 0 226 15 240
rect 0 102 15 136
rect 0 0 15 14
rect 0 -44 15 -30
rect 0 -168 15 -134
rect 0 -270 15 -256
rect 0 -314 15 -300
rect 0 -438 15 -404
rect 0 -540 15 -526
rect 0 -584 15 -570
rect 0 -708 15 -674
rect 0 -810 15 -796
rect 0 -854 15 -840
rect 0 -978 15 -944
rect 0 -1080 15 -1066
use 10T_1x8_magic  10T_1x8_magic_7
timestamp 1656019537
transform 1 0 0 0 1 -540
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_6
timestamp 1656019537
transform 1 0 0 0 1 -270
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_5
timestamp 1656019537
transform 1 0 0 0 1 -810
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_4
timestamp 1656019537
transform 1 0 0 0 1 -1080
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_1
timestamp 1656019537
transform 1 0 0 0 1 0
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_0
timestamp 1656019537
transform 1 0 0 0 1 270
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_2
timestamp 1656019537
transform 1 0 0 0 1 810
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_3
timestamp 1656019537
transform 1 0 0 0 1 540
box -7 -4 4631 312
<< labels >>
rlabel locali 0 -1042 15 -1000 1 RBL1_0
port 1 ns signal output
rlabel locali 537 -1042 552 -1000 1 RBL0_0
port 2 ns signal output
rlabel locali 580 -1042 595 -1000 1 RBL1_1
port 3 ns signal output
rlabel locali 1117 -1042 1132 -1000 1 RBL0_1
port 4 ns signal output
rlabel locali 1160 -1042 1175 -1000 1 RBL1_2
port 5 ns signal output
rlabel locali 1697 -1042 1712 -1000 1 RBL0_2
port 6 ns signal output
rlabel locali 1740 -1042 1755 -1000 1 RBL1_3
port 7 ns signal output
rlabel locali 2277 -1042 2292 -1000 1 RBL0_3
port 8 ns signal output
rlabel locali 2320 -1042 2335 -1000 1 RBL1_4
port 9 ns signal output
rlabel locali 2857 -1042 2872 -1000 1 RBL0_4
port 10 ns signal output
rlabel locali 2900 -1042 2915 -1000 1 RBL1_5
port 11 ns signal output
rlabel locali 3437 -1042 3452 -1000 1 RBL0_5
port 12 ns signal output
rlabel locali 3480 -1042 3495 -1000 1 RBL1_6
port 13 ns signal output
rlabel locali 4017 -1042 4032 -1000 1 RBL0_6
port 14 ns signal output
rlabel locali 4060 -1042 4075 -1000 1 RBL1_7
port 15 ns signal output
rlabel locali 4597 -1042 4612 -1000 1 RBL0_7
port 16 ns signal output
rlabel locali 464 -896 479 -867 1 WBL_0
port 17 ns signal input
rlabel locali 74 -896 89 -868 1 WBLb_0
port 18 ns signal input
rlabel locali 1044 -896 1059 -867 1 WBL_1
port 19 ns signal input
rlabel locali 654 -896 669 -868 1 WBLb_1
port 20 ns signal input
rlabel locali 1624 -896 1639 -867 1 WBL_2
port 21 ns signal input
rlabel locali 1234 -896 1249 -868 1 WBLb_2
port 22 ns signal input
rlabel locali 2204 -896 2219 -867 1 WBL_3
port 23 ns signal input
rlabel locali 1814 -896 1829 -868 1 WBLb_3
port 24 ns signal input
rlabel locali 2784 -896 2799 -867 1 WBL_4
port 25 ns signal input
rlabel locali 2394 -896 2409 -868 1 WBLb_4
port 26 ns signal input
rlabel locali 3364 -896 3379 -867 1 WBL_5
port 27 ns signal input
rlabel locali 2974 -896 2989 -868 1 WBLb_5
port 28 ns signal input
rlabel locali 3944 -896 3959 -867 1 WBL_6
port 29 ns signal input
rlabel locali 3554 -896 3569 -868 1 WBLb_6
port 30 ns signal input
rlabel locali 4524 -896 4539 -867 1 WBL_7
port 31 ns signal input
rlabel locali 4134 -896 4149 -868 1 WBLb_7
port 32 ns signal input
rlabel poly 0 1050 30 1080 1 WWL_0
port 33 ew signal input
rlabel metal1 0 912 15 946 1 RWL_0
port 34 ew signal input
rlabel poly 0 780 30 810 1 WWL_1
port 35 ew signal input
rlabel metal1 0 642 15 676 1 RWL_1
port 36 ew signal input
rlabel poly 0 510 30 540 1 WWL_2
port 37 ew signal input
rlabel metal1 0 372 15 406 1 RWL_2
port 38 ew signal input
rlabel poly 0 240 30 270 1 WWL_3
port 39 ew signal input
rlabel metal1 0 102 15 136 1 RWL_3
port 40 ew signal input
rlabel poly 0 -30 30 0 1 WWL_4
port 41 ew signal input
rlabel metal1 0 -168 15 -134 1 RWL_4
port 42 ew signal input
rlabel poly 0 -300 30 -270 1 WWL_5
port 43 ew signal input
rlabel metal1 0 -438 15 -404 1 RWL_5
port 44 ew signal input
rlabel poly 0 -570 30 -540 1 WWL_6
port 45 ew signal input
rlabel metal1 0 -708 15 -674 1 RWL_6
port 46 ew signal input
rlabel poly 0 -840 30 -810 1 WWL_7
port 47 ew signal input
rlabel metal1 0 -978 15 -944 1 RWL_7
port 48 ew signal input
rlabel metal1 0 1036 15 1050 1 VDD
port 49 ew power bidirectional abutment
rlabel metal1 0 810 15 824 1 GND
port 50 ew ground bidirectional abutment
rlabel metal1 0 496 15 510 1 VDD
rlabel metal1 0 226 15 240 1 VDD
rlabel metal1 0 766 15 780 1 VDD
rlabel metal1 0 -44 15 -30 1 VDD
rlabel metal1 0 -584 15 -570 1 VDD
rlabel metal1 0 -854 15 -840 1 VDD
rlabel metal1 0 -314 15 -300 1 VDD
rlabel metal1 0 0 15 14 1 GND
rlabel metal1 0 270 15 284 1 GND
rlabel metal1 0 540 15 554 1 GND
rlabel metal1 0 -270 15 -256 1 GND
rlabel metal1 0 -1080 15 -1066 1 GND
rlabel metal1 0 -810 15 -796 1 GND
rlabel metal1 0 -540 15 -526 1 GND
<< end >>
