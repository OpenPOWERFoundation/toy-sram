** sch_path: /home/rjridle/osu-toy-sram/xschem/10T_32x32_xschem.sch
.subckt 10T_32x32_xschem WWL_0 RWL_0 WWL_1 RWL_1 WWL_2 RWL_2 WWL_3 RWL_3 WWL_4 RWL_4 WWL_5 RWL_5
+ WWL_6 RWL_6 WWL_7 RWL_7 WWL_8 RWL_8 WWL_9 RWL_9 WWL_10 RWL_10 WWL_11 RWL_11 WWL_12 RWL_12 WWL_13 RWL_13
+ WWL_14 RWL_14 WWL_15 RWL_15 WWL_16 RWL_16 WWL_17 RWL_17 WWL_18 RWL_18 WWL_19 RWL_19 WWL_20 RWL_20 WWL_21
+ RWL_21 WWL_22 RWL_22 WWL_23 RWL_23 WWL_24 RWL_24 WWL_25 RWL_25 WWL_26 RWL_26 WWL_27 RWL_27 WWL_28 RWL_28
+ WWL_29 RWL_29 WWL_30 RWL_30 WWL_31 RWL_31 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL0_3 RBL1_3 RBL0_4
+ RBL1_4 RBL0_5 RBL1_5 RBL0_6 RBL1_6 RBL0_7 RBL1_7 RBL0_8 RBL1_8 RBL0_9 RBL1_9 RBL0_10 RBL1_10 RBL0_11
+ RBL1_11 RBL0_12 RBL1_12 RBL0_13 RBL1_13 RBL0_14 RBL1_14 RBL0_15 RBL1_15 RBL0_16 RBL1_16 RBL0_17 RBL1_17
+ RBL0_18 RBL1_18 RBL0_19 RBL1_19 RBL0_20 RBL1_20 RBL0_21 RBL0_22 RBL0_23 RBL1_21 RBL1_22 RBL1_23 RBL0_24
+ RBL1_24 RBL0_25 RBL1_25 RBL0_26 RBL1_26 RBL0_27 RBL1_27 RBL0_28 RBL1_28 RBL0_29 RBL1_29 RBL0_30 RBL1_30
+ RBL0_31 RBL1_31 WBL_0 WBLb_0 WBL_1 WBLb_1 WBL_2 WBLb_2 WBL_3 WBLb_3 WBL_4 WBLb_4 WBL_5 WBLb_5 WBL_6 WBLb_6
+ WBL_7 WBLb_7 WBL_8 WBLb_8 WBL_9 WBLb_9 WBL_10 WBLb_10 WBL_11 WBLb_11 WBL_12 WBLb_12 WBL_13 WBLb_13 WBL_14
+ WBLb_14 WBL_15 WBLb_15 WBL_16 WBLb_16 WBL_17 WBLb_17 WBL_18 WBLb_18 WBL_19 WBLb_19 WBL_20 WBLb_20 WBL_21
+ WBLb_21 WBL_22 WBLb_22 WBL_23 WBLb_23 WBL_24 WBLb_24 WBL_25 WBLb_25 WBLb_26 WBL_26 WBL_27 WBLb_27 WBL_28
+ WBLb_28 WBL_29 WBLb_29 WBL_30 WBLb_30 WBL_31 WBLb_31 VDD GND

x1 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_2 RWL_2 VDD GND 10T_1x32_xschem
x2 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_3 RWL_3 VDD GND 10T_1x32_xschem
x3 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_4 RWL_4 VDD GND 10T_1x32_xschem
x4 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_5 RWL_5 VDD GND 10T_1x32_xschem
x5 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_6 RWL_6 VDD GND 10T_1x32_xschem
x6 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_7 RWL_7 VDD GND 10T_1x32_xschem
x7 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_1 RWL_1 VDD GND 10T_1x32_xschem
x8 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_0 RWL_0 VDD GND 10T_1x32_xschem
x9 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_8 RWL_8 VDD GND 10T_1x32_xschem
x10 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_9 RWL_9 VDD GND 10T_1x32_xschem
x11 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_12 RWL_12 VDD GND 10T_1x32_xschem
x12 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_13 RWL_13 VDD GND 10T_1x32_xschem
x13 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_14 RWL_14 VDD GND 10T_1x32_xschem
x14 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_15 RWL_15 VDD GND 10T_1x32_xschem
x15 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_16 RWL_16 VDD GND 10T_1x32_xschem
x16 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_17 RWL_17 VDD GND 10T_1x32_xschem
x17 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_11 RWL_11 VDD GND 10T_1x32_xschem
x18 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_10 RWL_10 VDD GND 10T_1x32_xschem
x19 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_18 RWL_18 VDD GND 10T_1x32_xschem
x20 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_19 RWL_19 VDD GND 10T_1x32_xschem
x21 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_22 RWL_22 VDD GND 10T_1x32_xschem
x22 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_23 RWL_23 VDD GND 10T_1x32_xschem
x23 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_24 RWL_24 VDD GND 10T_1x32_xschem
x24 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_25 RWL_25 VDD GND 10T_1x32_xschem
x25 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_26 RWL_26 VDD GND 10T_1x32_xschem
x26 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_27 RWL_27 VDD GND 10T_1x32_xschem
x27 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_21 RWL_21 VDD GND 10T_1x32_xschem
x28 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_20 RWL_20 VDD GND 10T_1x32_xschem
x29 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_28 RWL_28 VDD GND 10T_1x32_xschem
x30 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_29 RWL_29 VDD GND 10T_1x32_xschem
x31 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_30 RWL_30 VDD GND 10T_1x32_xschem
x32 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_31 RWL_31 VDD GND 10T_1x32_xschem
.ends

.subckt 10T_1x32_xschem  RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18
+ RBL0_26 WBL_26 WBL_2 RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11
+ WBLb_30 WBLb_22 RBL0_31 RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13
+ RBL1_5 WBL_4 RBL1_20 WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27
+ RBL1_3 WBLb_5 WBLb_13 RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29
+ WBLb_18 RBL0_21 WBLb_10 RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9
+ WBLb_24 WBLb_16 RBL1_23 RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1
+ WBL_13 RBL0_9 RBL0_28 WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19
+ WBL_14 RBL0_11 WBL_6 RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31
+ WBLb_23 RBL0_16 RBL0_8 WBLb_15 RBL0_0 WBLb_7 WWL RWL VDD GND

x1 WWL RWL
+ WBL_0 WBL_1 WBL_2 WBL_3 WBL_4 WBL_5 WBL_6 WBL_7 
+ WBLb_0 WBLb_1 WBLb_2 WBLb_3 WBLb_4 WBLb_5 WBLb_6 WBLb_7
+ RBL0_0 RBL0_1 RBL0_2 RBL0_3 RBL0_4 RBL0_5 RBL0_6 RBL0_7 
+ RBL1_0 RBL1_1 RBL1_2 RBL1_3 RBL1_4 RBL1_5 RBL1_6 RBL1_7
+ VDD GND 10T_1x8_xschem

x2 WWL RWL
+ WBL_8 WBL_9 WBL_10 WBL_11 WBL_12 WBL_13 WBL_14 WBL_15 
+ WBLb_8 WBLb_9 WBLb_10 WBLb_11 WBLb_12 WBLb_13 WBLb_14 WBLb_15
+ RBL0_8 RBL0_9 RBL0_10 RBL0_11 RBL0_12 RBL0_13 RBL0_14 RBL0_15
+ RBL1_8 RBL1_9 RBL1_10 RBL1_11 RBL1_12 RBL1_13 RBL1_14 RBL1_15
+ VDD GND 10T_1x8_xschem

x3 WWL RWL
+ WBL_16 WBL_17 WBL_18 WBL_19 WBL_20 WBL_21 WBL_22 WBL_23 
+ WBLb_16 WBLb_17 WBLb_18 WBLb_19 WBLb_20 WBLb_21 WBLb_22 WBLb_23
+ RBL0_16 RBL0_17 RBL0_18 RBL0_19 RBL0_20 RBL0_21 RBL0_22 RBL0_23
+ RBL1_16 RBL1_17 RBL1_18 RBL1_19 RBL1_20 RBL1_21 RBL1_22 RBL1_23
+ VDD GND 10T_1x8_xschem

x4 WWL RWL
+ WBL_24 WBL_25 WBL_26 WBL_27 WBL_28 WBL_29 WBL_30 WBL_31 
+ WBLb_24 WBLb_25 WBLb_26 WBLb_27 WBLb_28 WBLb_29 WBLb_30 WBLb_31
+ RBL0_24 RBL0_25 RBL0_26 RBL0_27 RBL0_28 RBL0_29 RBL0_30 RBL0_31 
+ RBL1_24 RBL1_25 RBL1_26 RBL1_27 RBL1_28 RBL1_29 RBL1_30 RBL1_31
+ VDD GND 10T_1x8_xschem
.ends


* expanding   symbol:  10T_1x8_xschem.sym # of pins=34
** sym_path: /home/rjridle/osu-toy-sram/xschem/10T_1x8_xschem.sym
** sch_path: /home/rjridle/osu-toy-sram/xschem/10T_1x8_xschem.sch
.subckt 10T_1x8_xschem  WWL RWL
+ WBL_0 WBL_1 WBL_2 WBL_3 WBL_4 WBL_5 WBL_6 WBL_7 
+ WBLb_0 WBLb_1 WBLb_2 WBLb_3 WBLb_4 WBLb_5 WBLb_6 WBLb_7
+ RBL0_0 RBL0_1 RBL0_2 RBL0_3 RBL0_4 RBL0_5 RBL0_6 RBL0_7 
+ RBL1_0 RBL1_1 RBL1_2 RBL1_3 RBL1_4 RBL1_5 RBL1_6 RBL1_7
+ VDD GND

x1 WWL WBL_0 RBL0_0 RBL1_0 WBLb_0 RWL RWL VDD GND 10T_toy_xschem
x2 WWL WBL_1 RBL0_1 RBL1_1 WBLb_1 RWL RWL VDD GND 10T_toy_xschem
x3 WWL WBL_2 RBL0_2 RBL1_2 WBLb_2 RWL RWL VDD GND 10T_toy_xschem
x4 WWL WBL_3 RBL0_3 RBL1_3 WBLb_3 RWL RWL VDD GND 10T_toy_xschem
x5 WWL WBL_4 RBL0_4 RBL1_4 WBLb_4 RWL RWL VDD GND 10T_toy_xschem
x6 WWL WBL_5 RBL0_5 RBL1_5 WBLb_5 RWL RWL VDD GND 10T_toy_xschem
x7 WWL WBL_6 RBL0_6 RBL1_6 WBLb_6 RWL RWL VDD GND 10T_toy_xschem
x8 WWL WBL_7 RBL0_7 RBL1_7 WBLb_7 RWL RWL VDD GND 10T_toy_xschem
.ends


* expanding   symbol:  10T_toy_xschem.sym # of pins=7
** sym_path: /home/rjridle/osu-toy-sram/xschem/10T_toy_xschem.sym
** sch_path: /home/rjridle/osu-toy-sram/xschem/10T_toy_xschem.sch
.subckt 10T_toy_xschem  WWL WBL RBL0 RBL1 WBLb RWL0 RWL1  VDD  GND
*.PININFO WWL:I RWL0:I RWL1:I WBL:I WBLb:I RBL0:O RBL1:O
x1 net1 net2 VDD GND INVX1
x2 net2 net1 VDD GND INVX1
XM1 net2 WWL WBL GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 mult=1 m=1
XM2 WBLb WWL net1 GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 mult=1 m=1
XM3 net3 net2 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 mult=1 m=1 
XM4 RBL0 RWL0 net3 GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 mult=1 m=1 
XM5 net4 net1 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 mult=1 m=1 
XM6 RBL1 RWL1 net4 GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 mult=1 m=1
.ends


* expanding   symbol:  INVX1.sym # of pins=2
** sym_path: /home/rjridle/osu-toy-sram/xschem/INVX1.sym
** sch_path: /home/rjridle/osu-toy-sram/xschem/INVX1.sch
.subckt INVX1  Y A  VDD  GND
*.PININFO A:I Y:O
XM1 Y A GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 mult=1 m=1 
XM2 Y A VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 mult=1 m=1 
.ends

.end
