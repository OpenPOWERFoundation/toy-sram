../toysram.vh