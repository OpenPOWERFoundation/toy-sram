magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< locali >>
rect 238 1369 588 1388
rect 238 1263 252 1369
rect 574 1263 588 1369
rect 238 1249 588 1263
rect 238 125 588 139
rect 238 19 252 125
rect 574 19 588 125
rect 238 0 588 19
<< viali >>
rect 252 1263 574 1369
rect 252 19 574 125
<< obsli1 >>
rect 116 1225 182 1291
rect 644 1225 710 1291
rect 116 1203 160 1225
rect 666 1203 710 1225
rect 41 1179 160 1203
rect 41 1145 60 1179
rect 94 1145 160 1179
rect 41 1107 160 1145
rect 41 1073 60 1107
rect 94 1073 160 1107
rect 41 1035 160 1073
rect 41 1001 60 1035
rect 94 1001 160 1035
rect 41 963 160 1001
rect 41 929 60 963
rect 94 929 160 963
rect 41 891 160 929
rect 41 857 60 891
rect 94 857 160 891
rect 41 819 160 857
rect 41 785 60 819
rect 94 785 160 819
rect 41 747 160 785
rect 41 713 60 747
rect 94 713 160 747
rect 41 675 160 713
rect 41 641 60 675
rect 94 641 160 675
rect 41 603 160 641
rect 41 569 60 603
rect 94 569 160 603
rect 41 531 160 569
rect 41 497 60 531
rect 94 497 160 531
rect 41 459 160 497
rect 41 425 60 459
rect 94 425 160 459
rect 41 387 160 425
rect 41 353 60 387
rect 94 353 160 387
rect 41 315 160 353
rect 41 281 60 315
rect 94 281 160 315
rect 41 243 160 281
rect 41 209 60 243
rect 94 209 160 243
rect 41 185 160 209
rect 212 185 246 1203
rect 304 185 338 1203
rect 396 185 430 1203
rect 488 185 522 1203
rect 580 185 614 1203
rect 666 1179 785 1203
rect 666 1145 732 1179
rect 766 1145 785 1179
rect 666 1107 785 1145
rect 666 1073 732 1107
rect 766 1073 785 1107
rect 666 1035 785 1073
rect 666 1001 732 1035
rect 766 1001 785 1035
rect 666 963 785 1001
rect 666 929 732 963
rect 766 929 785 963
rect 666 891 785 929
rect 666 857 732 891
rect 766 857 785 891
rect 666 819 785 857
rect 666 785 732 819
rect 766 785 785 819
rect 666 747 785 785
rect 666 713 732 747
rect 766 713 785 747
rect 666 675 785 713
rect 666 641 732 675
rect 766 641 785 675
rect 666 603 785 641
rect 666 569 732 603
rect 766 569 785 603
rect 666 531 785 569
rect 666 497 732 531
rect 766 497 785 531
rect 666 459 785 497
rect 666 425 732 459
rect 766 425 785 459
rect 666 387 785 425
rect 666 353 732 387
rect 766 353 785 387
rect 666 315 785 353
rect 666 281 732 315
rect 766 281 785 315
rect 666 243 785 281
rect 666 209 732 243
rect 766 209 785 243
rect 666 185 785 209
rect 116 163 160 185
rect 666 163 710 185
rect 116 97 182 163
rect 644 97 710 163
<< obsli1c >>
rect 60 1145 94 1179
rect 60 1073 94 1107
rect 60 1001 94 1035
rect 60 929 94 963
rect 60 857 94 891
rect 60 785 94 819
rect 60 713 94 747
rect 60 641 94 675
rect 60 569 94 603
rect 60 497 94 531
rect 60 425 94 459
rect 60 353 94 387
rect 60 281 94 315
rect 60 209 94 243
rect 732 1145 766 1179
rect 732 1073 766 1107
rect 732 1001 766 1035
rect 732 929 766 963
rect 732 857 766 891
rect 732 785 766 819
rect 732 713 766 747
rect 732 641 766 675
rect 732 569 766 603
rect 732 497 766 531
rect 732 425 766 459
rect 732 353 766 387
rect 732 281 766 315
rect 732 209 766 243
<< metal1 >>
rect 236 1369 590 1388
rect 236 1263 252 1369
rect 574 1263 590 1369
rect 236 1251 590 1263
rect 41 1179 100 1191
rect 41 1145 60 1179
rect 94 1145 100 1179
rect 41 1107 100 1145
rect 41 1073 60 1107
rect 94 1073 100 1107
rect 41 1035 100 1073
rect 41 1001 60 1035
rect 94 1001 100 1035
rect 41 963 100 1001
rect 41 929 60 963
rect 94 929 100 963
rect 41 891 100 929
rect 41 857 60 891
rect 94 857 100 891
rect 41 819 100 857
rect 41 785 60 819
rect 94 785 100 819
rect 41 747 100 785
rect 41 713 60 747
rect 94 713 100 747
rect 41 675 100 713
rect 41 641 60 675
rect 94 641 100 675
rect 41 603 100 641
rect 41 569 60 603
rect 94 569 100 603
rect 41 531 100 569
rect 41 497 60 531
rect 94 497 100 531
rect 41 459 100 497
rect 41 425 60 459
rect 94 425 100 459
rect 41 387 100 425
rect 41 353 60 387
rect 94 353 100 387
rect 41 315 100 353
rect 41 281 60 315
rect 94 281 100 315
rect 41 243 100 281
rect 41 209 60 243
rect 94 209 100 243
rect 41 197 100 209
rect 726 1179 785 1191
rect 726 1145 732 1179
rect 766 1145 785 1179
rect 726 1107 785 1145
rect 726 1073 732 1107
rect 766 1073 785 1107
rect 726 1035 785 1073
rect 726 1001 732 1035
rect 766 1001 785 1035
rect 726 963 785 1001
rect 726 929 732 963
rect 766 929 785 963
rect 726 891 785 929
rect 726 857 732 891
rect 766 857 785 891
rect 726 819 785 857
rect 726 785 732 819
rect 766 785 785 819
rect 726 747 785 785
rect 726 713 732 747
rect 766 713 785 747
rect 726 675 785 713
rect 726 641 732 675
rect 766 641 785 675
rect 726 603 785 641
rect 726 569 732 603
rect 766 569 785 603
rect 726 531 785 569
rect 726 497 732 531
rect 766 497 785 531
rect 726 459 785 497
rect 726 425 732 459
rect 766 425 785 459
rect 726 387 785 425
rect 726 353 732 387
rect 766 353 785 387
rect 726 315 785 353
rect 726 281 732 315
rect 766 281 785 315
rect 726 243 785 281
rect 726 209 732 243
rect 766 209 785 243
rect 726 197 785 209
rect 236 125 590 137
rect 236 19 252 125
rect 574 19 590 125
rect 236 0 590 19
<< obsm1 >>
rect 203 197 255 1191
rect 295 197 347 1191
rect 387 197 439 1191
rect 479 197 531 1191
rect 571 197 623 1191
<< metal2 >>
rect 14 719 812 1191
rect 14 197 812 669
<< labels >>
rlabel metal2 s 14 719 812 1191 6 DRAIN
port 1 nsew
rlabel viali s 252 1263 574 1369 6 GATE
port 2 nsew
rlabel viali s 252 19 574 125 6 GATE
port 2 nsew
rlabel locali s 238 1249 588 1388 6 GATE
port 2 nsew
rlabel locali s 238 0 588 139 6 GATE
port 2 nsew
rlabel metal1 s 236 1251 590 1388 6 GATE
port 2 nsew
rlabel metal1 s 236 0 590 137 6 GATE
port 2 nsew
rlabel metal2 s 14 197 812 669 6 SOURCE
port 3 nsew
rlabel metal1 s 41 197 100 1191 6 SUBSTRATE
port 4 nsew
rlabel metal1 s 726 197 785 1191 6 SUBSTRATE
port 4 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 14 0 812 1388
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 5776730
string GDS_START 5748672
<< end >>
