magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< pwell >>
rect 112 708 768 730
rect 0 98 880 708
rect 112 76 768 98
<< nmos >>
rect 194 102 224 704
rect 348 102 378 704
rect 502 102 532 704
rect 656 102 686 704
<< ndiff >>
rect 138 692 194 704
rect 138 658 149 692
rect 183 658 194 692
rect 138 624 194 658
rect 138 590 149 624
rect 183 590 194 624
rect 138 556 194 590
rect 138 522 149 556
rect 183 522 194 556
rect 138 488 194 522
rect 138 454 149 488
rect 183 454 194 488
rect 138 420 194 454
rect 138 386 149 420
rect 183 386 194 420
rect 138 352 194 386
rect 138 318 149 352
rect 183 318 194 352
rect 138 284 194 318
rect 138 250 149 284
rect 183 250 194 284
rect 138 216 194 250
rect 138 182 149 216
rect 183 182 194 216
rect 138 148 194 182
rect 138 114 149 148
rect 183 114 194 148
rect 138 102 194 114
rect 224 692 348 704
rect 224 114 235 692
rect 337 114 348 692
rect 224 102 348 114
rect 378 692 502 704
rect 378 114 389 692
rect 491 114 502 692
rect 378 102 502 114
rect 532 692 656 704
rect 532 114 543 692
rect 645 114 656 692
rect 532 102 656 114
rect 686 692 742 704
rect 686 658 697 692
rect 731 658 742 692
rect 686 624 742 658
rect 686 590 697 624
rect 731 590 742 624
rect 686 556 742 590
rect 686 522 697 556
rect 731 522 742 556
rect 686 488 742 522
rect 686 454 697 488
rect 731 454 742 488
rect 686 420 742 454
rect 686 386 697 420
rect 731 386 742 420
rect 686 352 742 386
rect 686 318 697 352
rect 731 318 742 352
rect 686 284 742 318
rect 686 250 697 284
rect 731 250 742 284
rect 686 216 742 250
rect 686 182 697 216
rect 731 182 742 216
rect 686 148 742 182
rect 686 114 697 148
rect 731 114 742 148
rect 686 102 742 114
<< ndiffc >>
rect 149 658 183 692
rect 149 590 183 624
rect 149 522 183 556
rect 149 454 183 488
rect 149 386 183 420
rect 149 318 183 352
rect 149 250 183 284
rect 149 182 183 216
rect 149 114 183 148
rect 235 114 337 692
rect 389 114 491 692
rect 543 114 645 692
rect 697 658 731 692
rect 697 590 731 624
rect 697 522 731 556
rect 697 454 731 488
rect 697 386 731 420
rect 697 318 731 352
rect 697 250 731 284
rect 697 182 731 216
rect 697 114 731 148
<< psubdiff >>
rect 26 658 84 682
rect 26 624 38 658
rect 72 624 84 658
rect 26 590 84 624
rect 26 556 38 590
rect 72 556 84 590
rect 26 522 84 556
rect 26 488 38 522
rect 72 488 84 522
rect 26 454 84 488
rect 26 420 38 454
rect 72 420 84 454
rect 26 386 84 420
rect 26 352 38 386
rect 72 352 84 386
rect 26 318 84 352
rect 26 284 38 318
rect 72 284 84 318
rect 26 250 84 284
rect 26 216 38 250
rect 72 216 84 250
rect 26 182 84 216
rect 26 148 38 182
rect 72 148 84 182
rect 26 124 84 148
rect 796 658 854 682
rect 796 624 808 658
rect 842 624 854 658
rect 796 590 854 624
rect 796 556 808 590
rect 842 556 854 590
rect 796 522 854 556
rect 796 488 808 522
rect 842 488 854 522
rect 796 454 854 488
rect 796 420 808 454
rect 842 420 854 454
rect 796 386 854 420
rect 796 352 808 386
rect 842 352 854 386
rect 796 318 854 352
rect 796 284 808 318
rect 842 284 854 318
rect 796 250 854 284
rect 796 216 808 250
rect 842 216 854 250
rect 796 182 854 216
rect 796 148 808 182
rect 842 148 854 182
rect 796 124 854 148
<< psubdiffcont >>
rect 38 624 72 658
rect 38 556 72 590
rect 38 488 72 522
rect 38 420 72 454
rect 38 352 72 386
rect 38 284 72 318
rect 38 216 72 250
rect 38 148 72 182
rect 808 624 842 658
rect 808 556 842 590
rect 808 488 842 522
rect 808 420 842 454
rect 808 352 842 386
rect 808 284 842 318
rect 808 216 842 250
rect 808 148 842 182
<< poly >>
rect 168 786 710 802
rect 168 752 184 786
rect 218 752 252 786
rect 286 752 320 786
rect 354 752 388 786
rect 422 752 456 786
rect 490 752 524 786
rect 558 752 592 786
rect 626 752 660 786
rect 694 752 710 786
rect 168 736 710 752
rect 194 704 224 736
rect 348 704 378 736
rect 502 704 532 736
rect 656 704 686 736
rect 194 70 224 102
rect 348 70 378 102
rect 502 70 532 102
rect 656 70 686 102
rect 168 54 710 70
rect 168 20 184 54
rect 218 20 252 54
rect 286 20 320 54
rect 354 20 388 54
rect 422 20 456 54
rect 490 20 524 54
rect 558 20 592 54
rect 626 20 660 54
rect 694 20 710 54
rect 168 4 710 20
<< polycont >>
rect 184 752 218 786
rect 252 752 286 786
rect 320 752 354 786
rect 388 752 422 786
rect 456 752 490 786
rect 524 752 558 786
rect 592 752 626 786
rect 660 752 694 786
rect 184 20 218 54
rect 252 20 286 54
rect 320 20 354 54
rect 388 20 422 54
rect 456 20 490 54
rect 524 20 558 54
rect 592 20 626 54
rect 660 20 694 54
<< locali >>
rect 22 658 88 763
rect 168 752 170 786
rect 218 752 252 786
rect 300 752 320 786
rect 354 752 362 786
rect 422 752 456 786
rect 492 752 524 786
rect 588 752 592 786
rect 626 752 650 786
rect 694 752 710 786
rect 22 602 38 658
rect 72 602 88 658
rect 22 590 88 602
rect 22 530 38 590
rect 72 530 88 590
rect 22 522 88 530
rect 22 458 38 522
rect 72 458 88 522
rect 22 454 88 458
rect 22 352 38 454
rect 72 352 88 454
rect 22 348 88 352
rect 22 284 38 348
rect 72 284 88 348
rect 22 276 88 284
rect 22 216 38 276
rect 72 216 88 276
rect 22 204 88 216
rect 22 148 38 204
rect 72 148 88 204
rect 22 43 88 148
rect 138 692 183 708
rect 138 677 149 692
rect 138 643 147 677
rect 181 643 183 658
rect 138 624 183 643
rect 138 605 149 624
rect 138 571 147 605
rect 181 571 183 590
rect 138 556 183 571
rect 138 533 149 556
rect 138 499 147 533
rect 181 499 183 522
rect 138 488 183 499
rect 138 461 149 488
rect 138 427 147 461
rect 181 427 183 454
rect 138 420 183 427
rect 138 389 149 420
rect 138 355 147 389
rect 181 355 183 386
rect 138 352 183 355
rect 138 318 149 352
rect 138 317 183 318
rect 138 283 147 317
rect 181 284 183 317
rect 138 250 149 283
rect 138 245 183 250
rect 138 211 147 245
rect 181 216 183 245
rect 138 182 149 211
rect 138 173 183 182
rect 138 139 147 173
rect 181 148 183 173
rect 138 114 149 139
rect 138 98 183 114
rect 233 692 339 708
rect 233 677 235 692
rect 337 677 339 692
rect 233 114 235 139
rect 337 114 339 139
rect 233 98 339 114
rect 387 692 493 708
rect 387 667 389 692
rect 491 667 493 692
rect 387 114 389 129
rect 491 114 493 129
rect 387 98 493 114
rect 541 692 647 708
rect 541 677 543 692
rect 645 677 647 692
rect 541 114 543 139
rect 645 114 647 139
rect 541 98 647 114
rect 697 692 742 708
rect 731 677 742 692
rect 697 643 699 658
rect 733 643 742 677
rect 697 624 742 643
rect 731 605 742 624
rect 697 571 699 590
rect 733 571 742 605
rect 697 556 742 571
rect 731 533 742 556
rect 697 499 699 522
rect 733 499 742 533
rect 697 488 742 499
rect 731 461 742 488
rect 697 427 699 454
rect 733 427 742 461
rect 697 420 742 427
rect 731 389 742 420
rect 697 355 699 386
rect 733 355 742 389
rect 697 352 742 355
rect 731 318 742 352
rect 697 317 742 318
rect 697 284 699 317
rect 733 283 742 317
rect 731 250 742 283
rect 697 245 742 250
rect 697 216 699 245
rect 733 211 742 245
rect 731 182 742 211
rect 697 173 742 182
rect 697 148 699 173
rect 733 139 742 173
rect 731 114 742 139
rect 697 98 742 114
rect 792 658 858 763
rect 792 602 808 658
rect 842 602 858 658
rect 792 590 858 602
rect 792 530 808 590
rect 842 530 858 590
rect 792 522 858 530
rect 792 458 808 522
rect 842 458 858 522
rect 792 454 858 458
rect 792 352 808 454
rect 842 352 858 454
rect 792 348 858 352
rect 792 284 808 348
rect 842 284 858 348
rect 792 276 858 284
rect 792 216 808 276
rect 842 216 858 276
rect 792 204 858 216
rect 792 148 808 204
rect 842 148 858 204
rect 168 20 170 54
rect 218 20 252 54
rect 300 20 320 54
rect 354 20 362 54
rect 422 20 456 54
rect 492 20 524 54
rect 588 20 592 54
rect 626 20 650 54
rect 694 20 710 54
rect 792 43 858 148
<< viali >>
rect 170 752 184 786
rect 184 752 204 786
rect 266 752 286 786
rect 286 752 300 786
rect 362 752 388 786
rect 388 752 396 786
rect 458 752 490 786
rect 490 752 492 786
rect 554 752 558 786
rect 558 752 588 786
rect 650 752 660 786
rect 660 752 684 786
rect 38 624 72 636
rect 38 602 72 624
rect 38 556 72 564
rect 38 530 72 556
rect 38 488 72 492
rect 38 458 72 488
rect 38 386 72 420
rect 38 318 72 348
rect 38 314 72 318
rect 38 250 72 276
rect 38 242 72 250
rect 38 182 72 204
rect 38 170 72 182
rect 147 658 149 677
rect 149 658 181 677
rect 147 643 181 658
rect 147 590 149 605
rect 149 590 181 605
rect 147 571 181 590
rect 147 522 149 533
rect 149 522 181 533
rect 147 499 181 522
rect 147 454 149 461
rect 149 454 181 461
rect 147 427 181 454
rect 147 386 149 389
rect 149 386 181 389
rect 147 355 181 386
rect 147 284 181 317
rect 147 283 149 284
rect 149 283 181 284
rect 147 216 181 245
rect 147 211 149 216
rect 149 211 181 216
rect 147 148 181 173
rect 147 139 149 148
rect 149 139 181 148
rect 233 139 235 677
rect 235 139 337 677
rect 337 139 339 677
rect 387 129 389 667
rect 389 129 491 667
rect 491 129 493 667
rect 541 139 543 677
rect 543 139 645 677
rect 645 139 647 677
rect 699 658 731 677
rect 731 658 733 677
rect 699 643 733 658
rect 699 590 731 605
rect 731 590 733 605
rect 699 571 733 590
rect 699 522 731 533
rect 731 522 733 533
rect 699 499 733 522
rect 699 454 731 461
rect 731 454 733 461
rect 699 427 733 454
rect 699 386 731 389
rect 731 386 733 389
rect 699 355 733 386
rect 699 284 733 317
rect 699 283 731 284
rect 731 283 733 284
rect 699 216 733 245
rect 699 211 731 216
rect 731 211 733 216
rect 699 148 733 173
rect 699 139 731 148
rect 731 139 733 148
rect 808 624 842 636
rect 808 602 842 624
rect 808 556 842 564
rect 808 530 842 556
rect 808 488 842 492
rect 808 458 842 488
rect 808 386 842 420
rect 808 318 842 348
rect 808 314 842 318
rect 808 250 842 276
rect 808 242 842 250
rect 808 182 842 204
rect 808 170 842 182
rect 170 20 184 54
rect 184 20 204 54
rect 266 20 286 54
rect 286 20 300 54
rect 362 20 388 54
rect 388 20 396 54
rect 458 20 490 54
rect 490 20 492 54
rect 554 20 558 54
rect 558 20 588 54
rect 650 20 660 54
rect 660 20 684 54
<< metal1 >>
rect 164 786 690 798
rect 164 752 170 786
rect 204 752 266 786
rect 300 752 362 786
rect 396 752 458 786
rect 492 752 554 786
rect 588 752 650 786
rect 684 752 690 786
rect 164 740 690 752
rect 138 677 194 704
rect 138 643 147 677
rect 181 643 194 677
rect 26 636 84 642
rect 26 602 38 636
rect 72 602 84 636
rect 26 564 84 602
rect 26 530 38 564
rect 72 530 84 564
rect 26 492 84 530
rect 26 458 38 492
rect 72 458 84 492
rect 26 420 84 458
rect 26 386 38 420
rect 72 386 84 420
rect 26 348 84 386
rect 26 314 38 348
rect 72 314 84 348
rect 26 276 84 314
rect 26 242 38 276
rect 72 242 84 276
rect 26 204 84 242
rect 26 170 38 204
rect 72 170 84 204
rect 26 164 84 170
rect 138 605 194 643
rect 138 571 147 605
rect 181 571 194 605
rect 138 533 194 571
rect 138 499 147 533
rect 181 499 194 533
rect 138 461 194 499
rect 138 427 147 461
rect 181 427 194 461
rect 138 389 194 427
rect 138 360 147 389
rect 181 360 194 389
rect 138 308 140 360
rect 192 308 194 360
rect 138 296 147 308
rect 181 296 194 308
rect 138 244 140 296
rect 192 244 194 296
rect 138 232 147 244
rect 181 232 194 244
rect 138 180 140 232
rect 192 180 194 232
rect 138 173 194 180
rect 138 168 147 173
rect 181 168 194 173
rect 138 116 140 168
rect 192 116 194 168
rect 138 102 194 116
rect 223 690 349 704
rect 223 446 228 690
rect 344 446 349 690
rect 223 139 233 446
rect 339 139 349 446
rect 223 102 349 139
rect 377 667 503 704
rect 377 360 387 667
rect 493 360 503 667
rect 377 116 382 360
rect 498 116 503 360
rect 377 102 503 116
rect 531 690 657 704
rect 531 446 536 690
rect 652 446 657 690
rect 531 139 541 446
rect 647 139 657 446
rect 531 102 657 139
rect 686 677 742 704
rect 686 643 699 677
rect 733 643 742 677
rect 686 605 742 643
rect 686 571 699 605
rect 733 571 742 605
rect 686 533 742 571
rect 686 499 699 533
rect 733 499 742 533
rect 686 461 742 499
rect 686 427 699 461
rect 733 427 742 461
rect 686 389 742 427
rect 686 360 699 389
rect 733 360 742 389
rect 686 308 688 360
rect 740 308 742 360
rect 686 296 699 308
rect 733 296 742 308
rect 686 244 688 296
rect 740 244 742 296
rect 686 232 699 244
rect 733 232 742 244
rect 686 180 688 232
rect 740 180 742 232
rect 686 173 742 180
rect 686 168 699 173
rect 733 168 742 173
rect 686 116 688 168
rect 740 116 742 168
rect 796 636 854 642
rect 796 602 808 636
rect 842 602 854 636
rect 796 564 854 602
rect 796 530 808 564
rect 842 530 854 564
rect 796 492 854 530
rect 796 458 808 492
rect 842 458 854 492
rect 796 420 854 458
rect 796 386 808 420
rect 842 386 854 420
rect 796 348 854 386
rect 796 314 808 348
rect 842 314 854 348
rect 796 276 854 314
rect 796 242 808 276
rect 842 242 854 276
rect 796 204 854 242
rect 796 170 808 204
rect 842 170 854 204
rect 796 164 854 170
rect 686 102 742 116
rect 164 54 690 66
rect 164 20 170 54
rect 204 20 266 54
rect 300 20 362 54
rect 396 20 458 54
rect 492 20 554 54
rect 588 20 650 54
rect 684 20 690 54
rect 164 8 690 20
<< via1 >>
rect 140 355 147 360
rect 147 355 181 360
rect 181 355 192 360
rect 140 317 192 355
rect 140 308 147 317
rect 147 308 181 317
rect 181 308 192 317
rect 140 283 147 296
rect 147 283 181 296
rect 181 283 192 296
rect 140 245 192 283
rect 140 244 147 245
rect 147 244 181 245
rect 181 244 192 245
rect 140 211 147 232
rect 147 211 181 232
rect 181 211 192 232
rect 140 180 192 211
rect 140 139 147 168
rect 147 139 181 168
rect 181 139 192 168
rect 140 116 192 139
rect 228 677 344 690
rect 228 446 233 677
rect 233 446 339 677
rect 339 446 344 677
rect 382 129 387 360
rect 387 129 493 360
rect 493 129 498 360
rect 382 116 498 129
rect 536 677 652 690
rect 536 446 541 677
rect 541 446 647 677
rect 647 446 652 677
rect 688 355 699 360
rect 699 355 733 360
rect 733 355 740 360
rect 688 317 740 355
rect 688 308 699 317
rect 699 308 733 317
rect 733 308 740 317
rect 688 283 699 296
rect 699 283 733 296
rect 733 283 740 296
rect 688 245 740 283
rect 688 244 699 245
rect 699 244 733 245
rect 733 244 740 245
rect 688 211 699 232
rect 699 211 733 232
rect 733 211 740 232
rect 688 180 740 211
rect 688 139 699 168
rect 699 139 733 168
rect 733 139 740 168
rect 688 116 740 139
<< metal2 >>
rect 0 690 880 696
rect 0 446 228 690
rect 344 446 536 690
rect 652 446 880 690
rect 0 440 880 446
rect 0 360 880 366
rect 0 308 140 360
rect 192 308 382 360
rect 0 296 382 308
rect 0 244 140 296
rect 192 244 382 296
rect 0 232 382 244
rect 0 180 140 232
rect 192 180 382 232
rect 0 168 382 180
rect 0 116 140 168
rect 192 116 382 168
rect 498 308 688 360
rect 740 308 880 360
rect 498 296 880 308
rect 498 244 688 296
rect 740 244 880 296
rect 498 232 880 244
rect 498 180 688 232
rect 740 180 880 232
rect 498 168 880 180
rect 498 116 688 168
rect 740 116 880 168
rect 0 110 880 116
<< labels >>
flabel comment s 584 406 584 406 0 FreeSans 300 0 0 0 D
flabel comment s 166 389 166 389 0 FreeSans 300 0 0 0 S
flabel comment s 436 406 436 406 0 FreeSans 300 0 0 0 S
flabel comment s 276 406 276 406 0 FreeSans 300 0 0 0 D
flabel comment s 714 389 714 389 0 FreeSans 300 180 0 0 S
flabel metal1 s 36 370 62 437 0 FreeSans 400 90 0 0 SUBSTRATE
port 4 nsew
flabel metal1 s 416 22 502 47 0 FreeSans 400 0 0 0 GATE
port 2 nsew
flabel metal2 s 88 319 164 344 0 FreeSans 400 0 0 0 SOURCE
port 3 nsew
flabel metal2 s 84 627 173 659 0 FreeSans 400 0 0 0 DRAIN
port 1 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 7206420
string GDS_START 7186208
<< end >>
