VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO 10T_32x32_magic_flattened
  CLASS BLOCK ;
  FOREIGN 10T_32x32_magic_flattened ;
  ORIGIN 0.000 0.000 ;
  SIZE 92.660 BY 43.200 ;
  PIN RBL1_0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444800 ;
    PORT
      LAYER li1 ;
        RECT 0.000 42.040 0.075 42.250 ;
        RECT 0.000 40.690 0.075 40.900 ;
        RECT 0.000 39.340 0.075 39.550 ;
        RECT 0.000 37.990 0.075 38.200 ;
        RECT 0.000 36.640 0.075 36.850 ;
        RECT 0.000 35.290 0.075 35.500 ;
        RECT 0.000 33.940 0.075 34.150 ;
        RECT 0.000 32.590 0.075 32.800 ;
        RECT 0.000 31.240 0.075 31.450 ;
        RECT 0.000 29.890 0.075 30.100 ;
        RECT 0.000 28.540 0.075 28.750 ;
        RECT 0.000 27.190 0.075 27.400 ;
        RECT 0.000 25.840 0.075 26.050 ;
        RECT 0.000 24.490 0.075 24.700 ;
        RECT 0.000 23.140 0.075 23.350 ;
        RECT 0.000 21.790 0.075 22.000 ;
        RECT 0.000 20.440 0.075 20.650 ;
        RECT 0.000 19.090 0.075 19.300 ;
        RECT 0.000 17.740 0.075 17.950 ;
        RECT 0.000 16.390 0.075 16.600 ;
        RECT 0.000 15.040 0.075 15.250 ;
        RECT 0.000 13.690 0.075 13.900 ;
        RECT 0.000 12.340 0.075 12.550 ;
        RECT 0.000 10.990 0.075 11.200 ;
        RECT 0.000 9.640 0.075 9.850 ;
        RECT 0.000 8.290 0.075 8.500 ;
        RECT 0.000 6.940 0.075 7.150 ;
        RECT 0.000 5.590 0.075 5.800 ;
        RECT 0.000 4.240 0.075 4.450 ;
        RECT 0.000 2.890 0.075 3.100 ;
        RECT 0.000 1.540 0.075 1.750 ;
        RECT 0.000 0.190 0.075 0.400 ;
    END
  END RBL1_0
  PIN RBL0_0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444800 ;
    PORT
      LAYER li1 ;
        RECT 2.685 42.040 2.760 42.250 ;
        RECT 2.685 40.690 2.760 40.900 ;
        RECT 2.685 39.340 2.760 39.550 ;
        RECT 2.685 37.990 2.760 38.200 ;
        RECT 2.685 36.640 2.760 36.850 ;
        RECT 2.685 35.290 2.760 35.500 ;
        RECT 2.685 33.940 2.760 34.150 ;
        RECT 2.685 32.590 2.760 32.800 ;
        RECT 2.685 31.240 2.760 31.450 ;
        RECT 2.685 29.890 2.760 30.100 ;
        RECT 2.685 28.540 2.760 28.750 ;
        RECT 2.685 27.190 2.760 27.400 ;
        RECT 2.685 25.840 2.760 26.050 ;
        RECT 2.685 24.490 2.760 24.700 ;
        RECT 2.685 23.140 2.760 23.350 ;
        RECT 2.685 21.790 2.760 22.000 ;
        RECT 2.685 20.440 2.760 20.650 ;
        RECT 2.685 19.090 2.760 19.300 ;
        RECT 2.685 17.740 2.760 17.950 ;
        RECT 2.685 16.390 2.760 16.600 ;
        RECT 2.685 15.040 2.760 15.250 ;
        RECT 2.685 13.690 2.760 13.900 ;
        RECT 2.685 12.340 2.760 12.550 ;
        RECT 2.685 10.990 2.760 11.200 ;
        RECT 2.685 9.640 2.760 9.850 ;
        RECT 2.685 8.290 2.760 8.500 ;
        RECT 2.685 6.940 2.760 7.150 ;
        RECT 2.685 5.590 2.760 5.800 ;
        RECT 2.685 4.240 2.760 4.450 ;
        RECT 2.685 2.890 2.760 3.100 ;
        RECT 2.685 1.540 2.760 1.750 ;
        RECT 2.685 0.190 2.760 0.400 ;
    END
  END RBL0_0
  PIN RBL1_1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444800 ;
    PORT
      LAYER li1 ;
        RECT 2.900 42.040 2.975 42.250 ;
        RECT 2.900 40.690 2.975 40.900 ;
        RECT 2.900 39.340 2.975 39.550 ;
        RECT 2.900 37.990 2.975 38.200 ;
        RECT 2.900 36.640 2.975 36.850 ;
        RECT 2.900 35.290 2.975 35.500 ;
        RECT 2.900 33.940 2.975 34.150 ;
        RECT 2.900 32.590 2.975 32.800 ;
        RECT 2.900 31.240 2.975 31.450 ;
        RECT 2.900 29.890 2.975 30.100 ;
        RECT 2.900 28.540 2.975 28.750 ;
        RECT 2.900 27.190 2.975 27.400 ;
        RECT 2.900 25.840 2.975 26.050 ;
        RECT 2.900 24.490 2.975 24.700 ;
        RECT 2.900 23.140 2.975 23.350 ;
        RECT 2.900 21.790 2.975 22.000 ;
        RECT 2.900 20.440 2.975 20.650 ;
        RECT 2.900 19.090 2.975 19.300 ;
        RECT 2.900 17.740 2.975 17.950 ;
        RECT 2.900 16.390 2.975 16.600 ;
        RECT 2.900 15.040 2.975 15.250 ;
        RECT 2.900 13.690 2.975 13.900 ;
        RECT 2.900 12.340 2.975 12.550 ;
        RECT 2.900 10.990 2.975 11.200 ;
        RECT 2.900 9.640 2.975 9.850 ;
        RECT 2.900 8.290 2.975 8.500 ;
        RECT 2.900 6.940 2.975 7.150 ;
        RECT 2.900 5.590 2.975 5.800 ;
        RECT 2.900 4.240 2.975 4.450 ;
        RECT 2.900 2.890 2.975 3.100 ;
        RECT 2.900 1.540 2.975 1.750 ;
        RECT 2.900 0.190 2.975 0.400 ;
    END
  END RBL1_1
  PIN RBL0_1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444800 ;
    PORT
      LAYER li1 ;
        RECT 5.585 42.040 5.660 42.250 ;
        RECT 5.585 40.690 5.660 40.900 ;
        RECT 5.585 39.340 5.660 39.550 ;
        RECT 5.585 37.990 5.660 38.200 ;
        RECT 5.585 36.640 5.660 36.850 ;
        RECT 5.585 35.290 5.660 35.500 ;
        RECT 5.585 33.940 5.660 34.150 ;
        RECT 5.585 32.590 5.660 32.800 ;
        RECT 5.585 31.240 5.660 31.450 ;
        RECT 5.585 29.890 5.660 30.100 ;
        RECT 5.585 28.540 5.660 28.750 ;
        RECT 5.585 27.190 5.660 27.400 ;
        RECT 5.585 25.840 5.660 26.050 ;
        RECT 5.585 24.490 5.660 24.700 ;
        RECT 5.585 23.140 5.660 23.350 ;
        RECT 5.585 21.790 5.660 22.000 ;
        RECT 5.585 20.440 5.660 20.650 ;
        RECT 5.585 19.090 5.660 19.300 ;
        RECT 5.585 17.740 5.660 17.950 ;
        RECT 5.585 16.390 5.660 16.600 ;
        RECT 5.585 15.040 5.660 15.250 ;
        RECT 5.585 13.690 5.660 13.900 ;
        RECT 5.585 12.340 5.660 12.550 ;
        RECT 5.585 10.990 5.660 11.200 ;
        RECT 5.585 9.640 5.660 9.850 ;
        RECT 5.585 8.290 5.660 8.500 ;
        RECT 5.585 6.940 5.660 7.150 ;
        RECT 5.585 5.590 5.660 5.800 ;
        RECT 5.585 4.240 5.660 4.450 ;
        RECT 5.585 2.890 5.660 3.100 ;
        RECT 5.585 1.540 5.660 1.750 ;
        RECT 5.585 0.190 5.660 0.400 ;
    END
  END RBL0_1
  PIN RBL1_2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444800 ;
    PORT
      LAYER li1 ;
        RECT 5.800 42.040 5.875 42.250 ;
        RECT 5.800 40.690 5.875 40.900 ;
        RECT 5.800 39.340 5.875 39.550 ;
        RECT 5.800 37.990 5.875 38.200 ;
        RECT 5.800 36.640 5.875 36.850 ;
        RECT 5.800 35.290 5.875 35.500 ;
        RECT 5.800 33.940 5.875 34.150 ;
        RECT 5.800 32.590 5.875 32.800 ;
        RECT 5.800 31.240 5.875 31.450 ;
        RECT 5.800 29.890 5.875 30.100 ;
        RECT 5.800 28.540 5.875 28.750 ;
        RECT 5.800 27.190 5.875 27.400 ;
        RECT 5.800 25.840 5.875 26.050 ;
        RECT 5.800 24.490 5.875 24.700 ;
        RECT 5.800 23.140 5.875 23.350 ;
        RECT 5.800 21.790 5.875 22.000 ;
        RECT 5.800 20.440 5.875 20.650 ;
        RECT 5.800 19.090 5.875 19.300 ;
        RECT 5.800 17.740 5.875 17.950 ;
        RECT 5.800 16.390 5.875 16.600 ;
        RECT 5.800 15.040 5.875 15.250 ;
        RECT 5.800 13.690 5.875 13.900 ;
        RECT 5.800 12.340 5.875 12.550 ;
        RECT 5.800 10.990 5.875 11.200 ;
        RECT 5.800 9.640 5.875 9.850 ;
        RECT 5.800 8.290 5.875 8.500 ;
        RECT 5.800 6.940 5.875 7.150 ;
        RECT 5.800 5.590 5.875 5.800 ;
        RECT 5.800 4.240 5.875 4.450 ;
        RECT 5.800 2.890 5.875 3.100 ;
        RECT 5.800 1.540 5.875 1.750 ;
        RECT 5.800 0.190 5.875 0.400 ;
    END
  END RBL1_2
  PIN RBL0_2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444800 ;
    PORT
      LAYER li1 ;
        RECT 8.485 42.040 8.560 42.250 ;
        RECT 8.485 40.690 8.560 40.900 ;
        RECT 8.485 39.340 8.560 39.550 ;
        RECT 8.485 37.990 8.560 38.200 ;
        RECT 8.485 36.640 8.560 36.850 ;
        RECT 8.485 35.290 8.560 35.500 ;
        RECT 8.485 33.940 8.560 34.150 ;
        RECT 8.485 32.590 8.560 32.800 ;
        RECT 8.485 31.240 8.560 31.450 ;
        RECT 8.485 29.890 8.560 30.100 ;
        RECT 8.485 28.540 8.560 28.750 ;
        RECT 8.485 27.190 8.560 27.400 ;
        RECT 8.485 25.840 8.560 26.050 ;
        RECT 8.485 24.490 8.560 24.700 ;
        RECT 8.485 23.140 8.560 23.350 ;
        RECT 8.485 21.790 8.560 22.000 ;
        RECT 8.485 20.440 8.560 20.650 ;
        RECT 8.485 19.090 8.560 19.300 ;
        RECT 8.485 17.740 8.560 17.950 ;
        RECT 8.485 16.390 8.560 16.600 ;
        RECT 8.485 15.040 8.560 15.250 ;
        RECT 8.485 13.690 8.560 13.900 ;
        RECT 8.485 12.340 8.560 12.550 ;
        RECT 8.485 10.990 8.560 11.200 ;
        RECT 8.485 9.640 8.560 9.850 ;
        RECT 8.485 8.290 8.560 8.500 ;
        RECT 8.485 6.940 8.560 7.150 ;
        RECT 8.485 5.590 8.560 5.800 ;
        RECT 8.485 4.240 8.560 4.450 ;
        RECT 8.485 2.890 8.560 3.100 ;
        RECT 8.485 1.540 8.560 1.750 ;
        RECT 8.485 0.190 8.560 0.400 ;
    END
  END RBL0_2
  PIN RBL1_3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444800 ;
    PORT
      LAYER li1 ;
        RECT 8.700 42.040 8.775 42.250 ;
        RECT 8.700 40.690 8.775 40.900 ;
        RECT 8.700 39.340 8.775 39.550 ;
        RECT 8.700 37.990 8.775 38.200 ;
        RECT 8.700 36.640 8.775 36.850 ;
        RECT 8.700 35.290 8.775 35.500 ;
        RECT 8.700 33.940 8.775 34.150 ;
        RECT 8.700 32.590 8.775 32.800 ;
        RECT 8.700 31.240 8.775 31.450 ;
        RECT 8.700 29.890 8.775 30.100 ;
        RECT 8.700 28.540 8.775 28.750 ;
        RECT 8.700 27.190 8.775 27.400 ;
        RECT 8.700 25.840 8.775 26.050 ;
        RECT 8.700 24.490 8.775 24.700 ;
        RECT 8.700 23.140 8.775 23.350 ;
        RECT 8.700 21.790 8.775 22.000 ;
        RECT 8.700 20.440 8.775 20.650 ;
        RECT 8.700 19.090 8.775 19.300 ;
        RECT 8.700 17.740 8.775 17.950 ;
        RECT 8.700 16.390 8.775 16.600 ;
        RECT 8.700 15.040 8.775 15.250 ;
        RECT 8.700 13.690 8.775 13.900 ;
        RECT 8.700 12.340 8.775 12.550 ;
        RECT 8.700 10.990 8.775 11.200 ;
        RECT 8.700 9.640 8.775 9.850 ;
        RECT 8.700 8.290 8.775 8.500 ;
        RECT 8.700 6.940 8.775 7.150 ;
        RECT 8.700 5.590 8.775 5.800 ;
        RECT 8.700 4.240 8.775 4.450 ;
        RECT 8.700 2.890 8.775 3.100 ;
        RECT 8.700 1.540 8.775 1.750 ;
        RECT 8.700 0.190 8.775 0.400 ;
    END
  END RBL1_3
  PIN RBL0_3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444800 ;
    PORT
      LAYER li1 ;
        RECT 11.385 42.040 11.460 42.250 ;
        RECT 11.385 40.690 11.460 40.900 ;
        RECT 11.385 39.340 11.460 39.550 ;
        RECT 11.385 37.990 11.460 38.200 ;
        RECT 11.385 36.640 11.460 36.850 ;
        RECT 11.385 35.290 11.460 35.500 ;
        RECT 11.385 33.940 11.460 34.150 ;
        RECT 11.385 32.590 11.460 32.800 ;
        RECT 11.385 31.240 11.460 31.450 ;
        RECT 11.385 29.890 11.460 30.100 ;
        RECT 11.385 28.540 11.460 28.750 ;
        RECT 11.385 27.190 11.460 27.400 ;
        RECT 11.385 25.840 11.460 26.050 ;
        RECT 11.385 24.490 11.460 24.700 ;
        RECT 11.385 23.140 11.460 23.350 ;
        RECT 11.385 21.790 11.460 22.000 ;
        RECT 11.385 20.440 11.460 20.650 ;
        RECT 11.385 19.090 11.460 19.300 ;
        RECT 11.385 17.740 11.460 17.950 ;
        RECT 11.385 16.390 11.460 16.600 ;
        RECT 11.385 15.040 11.460 15.250 ;
        RECT 11.385 13.690 11.460 13.900 ;
        RECT 11.385 12.340 11.460 12.550 ;
        RECT 11.385 10.990 11.460 11.200 ;
        RECT 11.385 9.640 11.460 9.850 ;
        RECT 11.385 8.290 11.460 8.500 ;
        RECT 11.385 6.940 11.460 7.150 ;
        RECT 11.385 5.590 11.460 5.800 ;
        RECT 11.385 4.240 11.460 4.450 ;
        RECT 11.385 2.890 11.460 3.100 ;
        RECT 11.385 1.540 11.460 1.750 ;
        RECT 11.385 0.190 11.460 0.400 ;
    END
  END RBL0_3
  PIN RBL1_4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444800 ;
    PORT
      LAYER li1 ;
        RECT 11.600 42.040 11.675 42.250 ;
        RECT 11.600 40.690 11.675 40.900 ;
        RECT 11.600 39.340 11.675 39.550 ;
        RECT 11.600 37.990 11.675 38.200 ;
        RECT 11.600 36.640 11.675 36.850 ;
        RECT 11.600 35.290 11.675 35.500 ;
        RECT 11.600 33.940 11.675 34.150 ;
        RECT 11.600 32.590 11.675 32.800 ;
        RECT 11.600 31.240 11.675 31.450 ;
        RECT 11.600 29.890 11.675 30.100 ;
        RECT 11.600 28.540 11.675 28.750 ;
        RECT 11.600 27.190 11.675 27.400 ;
        RECT 11.600 25.840 11.675 26.050 ;
        RECT 11.600 24.490 11.675 24.700 ;
        RECT 11.600 23.140 11.675 23.350 ;
        RECT 11.600 21.790 11.675 22.000 ;
        RECT 11.600 20.440 11.675 20.650 ;
        RECT 11.600 19.090 11.675 19.300 ;
        RECT 11.600 17.740 11.675 17.950 ;
        RECT 11.600 16.390 11.675 16.600 ;
        RECT 11.600 15.040 11.675 15.250 ;
        RECT 11.600 13.690 11.675 13.900 ;
        RECT 11.600 12.340 11.675 12.550 ;
        RECT 11.600 10.990 11.675 11.200 ;
        RECT 11.600 9.640 11.675 9.850 ;
        RECT 11.600 8.290 11.675 8.500 ;
        RECT 11.600 6.940 11.675 7.150 ;
        RECT 11.600 5.590 11.675 5.800 ;
        RECT 11.600 4.240 11.675 4.450 ;
        RECT 11.600 2.890 11.675 3.100 ;
        RECT 11.600 1.540 11.675 1.750 ;
        RECT 11.600 0.190 11.675 0.400 ;
    END
  END RBL1_4
  PIN RBL0_4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444800 ;
    PORT
      LAYER li1 ;
        RECT 14.285 42.040 14.360 42.250 ;
        RECT 14.285 40.690 14.360 40.900 ;
        RECT 14.285 39.340 14.360 39.550 ;
        RECT 14.285 37.990 14.360 38.200 ;
        RECT 14.285 36.640 14.360 36.850 ;
        RECT 14.285 35.290 14.360 35.500 ;
        RECT 14.285 33.940 14.360 34.150 ;
        RECT 14.285 32.590 14.360 32.800 ;
        RECT 14.285 31.240 14.360 31.450 ;
        RECT 14.285 29.890 14.360 30.100 ;
        RECT 14.285 28.540 14.360 28.750 ;
        RECT 14.285 27.190 14.360 27.400 ;
        RECT 14.285 25.840 14.360 26.050 ;
        RECT 14.285 24.490 14.360 24.700 ;
        RECT 14.285 23.140 14.360 23.350 ;
        RECT 14.285 21.790 14.360 22.000 ;
        RECT 14.285 20.440 14.360 20.650 ;
        RECT 14.285 19.090 14.360 19.300 ;
        RECT 14.285 17.740 14.360 17.950 ;
        RECT 14.285 16.390 14.360 16.600 ;
        RECT 14.285 15.040 14.360 15.250 ;
        RECT 14.285 13.690 14.360 13.900 ;
        RECT 14.285 12.340 14.360 12.550 ;
        RECT 14.285 10.990 14.360 11.200 ;
        RECT 14.285 9.640 14.360 9.850 ;
        RECT 14.285 8.290 14.360 8.500 ;
        RECT 14.285 6.940 14.360 7.150 ;
        RECT 14.285 5.590 14.360 5.800 ;
        RECT 14.285 4.240 14.360 4.450 ;
        RECT 14.285 2.890 14.360 3.100 ;
        RECT 14.285 1.540 14.360 1.750 ;
        RECT 14.285 0.190 14.360 0.400 ;
    END
  END RBL0_4
  PIN RBL1_5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444800 ;
    PORT
      LAYER li1 ;
        RECT 14.500 42.040 14.575 42.250 ;
        RECT 14.500 40.690 14.575 40.900 ;
        RECT 14.500 39.340 14.575 39.550 ;
        RECT 14.500 37.990 14.575 38.200 ;
        RECT 14.500 36.640 14.575 36.850 ;
        RECT 14.500 35.290 14.575 35.500 ;
        RECT 14.500 33.940 14.575 34.150 ;
        RECT 14.500 32.590 14.575 32.800 ;
        RECT 14.500 31.240 14.575 31.450 ;
        RECT 14.500 29.890 14.575 30.100 ;
        RECT 14.500 28.540 14.575 28.750 ;
        RECT 14.500 27.190 14.575 27.400 ;
        RECT 14.500 25.840 14.575 26.050 ;
        RECT 14.500 24.490 14.575 24.700 ;
        RECT 14.500 23.140 14.575 23.350 ;
        RECT 14.500 21.790 14.575 22.000 ;
        RECT 14.500 20.440 14.575 20.650 ;
        RECT 14.500 19.090 14.575 19.300 ;
        RECT 14.500 17.740 14.575 17.950 ;
        RECT 14.500 16.390 14.575 16.600 ;
        RECT 14.500 15.040 14.575 15.250 ;
        RECT 14.500 13.690 14.575 13.900 ;
        RECT 14.500 12.340 14.575 12.550 ;
        RECT 14.500 10.990 14.575 11.200 ;
        RECT 14.500 9.640 14.575 9.850 ;
        RECT 14.500 8.290 14.575 8.500 ;
        RECT 14.500 6.940 14.575 7.150 ;
        RECT 14.500 5.590 14.575 5.800 ;
        RECT 14.500 4.240 14.575 4.450 ;
        RECT 14.500 2.890 14.575 3.100 ;
        RECT 14.500 1.540 14.575 1.750 ;
        RECT 14.500 0.190 14.575 0.400 ;
    END
  END RBL1_5
  PIN RBL0_5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444800 ;
    PORT
      LAYER li1 ;
        RECT 17.185 42.040 17.260 42.250 ;
        RECT 17.185 40.690 17.260 40.900 ;
        RECT 17.185 39.340 17.260 39.550 ;
        RECT 17.185 37.990 17.260 38.200 ;
        RECT 17.185 36.640 17.260 36.850 ;
        RECT 17.185 35.290 17.260 35.500 ;
        RECT 17.185 33.940 17.260 34.150 ;
        RECT 17.185 32.590 17.260 32.800 ;
        RECT 17.185 31.240 17.260 31.450 ;
        RECT 17.185 29.890 17.260 30.100 ;
        RECT 17.185 28.540 17.260 28.750 ;
        RECT 17.185 27.190 17.260 27.400 ;
        RECT 17.185 25.840 17.260 26.050 ;
        RECT 17.185 24.490 17.260 24.700 ;
        RECT 17.185 23.140 17.260 23.350 ;
        RECT 17.185 21.790 17.260 22.000 ;
        RECT 17.185 20.440 17.260 20.650 ;
        RECT 17.185 19.090 17.260 19.300 ;
        RECT 17.185 17.740 17.260 17.950 ;
        RECT 17.185 16.390 17.260 16.600 ;
        RECT 17.185 15.040 17.260 15.250 ;
        RECT 17.185 13.690 17.260 13.900 ;
        RECT 17.185 12.340 17.260 12.550 ;
        RECT 17.185 10.990 17.260 11.200 ;
        RECT 17.185 9.640 17.260 9.850 ;
        RECT 17.185 8.290 17.260 8.500 ;
        RECT 17.185 6.940 17.260 7.150 ;
        RECT 17.185 5.590 17.260 5.800 ;
        RECT 17.185 4.240 17.260 4.450 ;
        RECT 17.185 2.890 17.260 3.100 ;
        RECT 17.185 1.540 17.260 1.750 ;
        RECT 17.185 0.190 17.260 0.400 ;
    END
  END RBL0_5
  PIN RBL1_6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444800 ;
    PORT
      LAYER li1 ;
        RECT 17.400 42.040 17.475 42.250 ;
        RECT 17.400 40.690 17.475 40.900 ;
        RECT 17.400 39.340 17.475 39.550 ;
        RECT 17.400 37.990 17.475 38.200 ;
        RECT 17.400 36.640 17.475 36.850 ;
        RECT 17.400 35.290 17.475 35.500 ;
        RECT 17.400 33.940 17.475 34.150 ;
        RECT 17.400 32.590 17.475 32.800 ;
        RECT 17.400 31.240 17.475 31.450 ;
        RECT 17.400 29.890 17.475 30.100 ;
        RECT 17.400 28.540 17.475 28.750 ;
        RECT 17.400 27.190 17.475 27.400 ;
        RECT 17.400 25.840 17.475 26.050 ;
        RECT 17.400 24.490 17.475 24.700 ;
        RECT 17.400 23.140 17.475 23.350 ;
        RECT 17.400 21.790 17.475 22.000 ;
        RECT 17.400 20.440 17.475 20.650 ;
        RECT 17.400 19.090 17.475 19.300 ;
        RECT 17.400 17.740 17.475 17.950 ;
        RECT 17.400 16.390 17.475 16.600 ;
        RECT 17.400 15.040 17.475 15.250 ;
        RECT 17.400 13.690 17.475 13.900 ;
        RECT 17.400 12.340 17.475 12.550 ;
        RECT 17.400 10.990 17.475 11.200 ;
        RECT 17.400 9.640 17.475 9.850 ;
        RECT 17.400 8.290 17.475 8.500 ;
        RECT 17.400 6.940 17.475 7.150 ;
        RECT 17.400 5.590 17.475 5.800 ;
        RECT 17.400 4.240 17.475 4.450 ;
        RECT 17.400 2.890 17.475 3.100 ;
        RECT 17.400 1.540 17.475 1.750 ;
        RECT 17.400 0.190 17.475 0.400 ;
    END
  END RBL1_6
  PIN RBL0_6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444800 ;
    PORT
      LAYER li1 ;
        RECT 20.085 42.040 20.160 42.250 ;
        RECT 20.085 40.690 20.160 40.900 ;
        RECT 20.085 39.340 20.160 39.550 ;
        RECT 20.085 37.990 20.160 38.200 ;
        RECT 20.085 36.640 20.160 36.850 ;
        RECT 20.085 35.290 20.160 35.500 ;
        RECT 20.085 33.940 20.160 34.150 ;
        RECT 20.085 32.590 20.160 32.800 ;
        RECT 20.085 31.240 20.160 31.450 ;
        RECT 20.085 29.890 20.160 30.100 ;
        RECT 20.085 28.540 20.160 28.750 ;
        RECT 20.085 27.190 20.160 27.400 ;
        RECT 20.085 25.840 20.160 26.050 ;
        RECT 20.085 24.490 20.160 24.700 ;
        RECT 20.085 23.140 20.160 23.350 ;
        RECT 20.085 21.790 20.160 22.000 ;
        RECT 20.085 20.440 20.160 20.650 ;
        RECT 20.085 19.090 20.160 19.300 ;
        RECT 20.085 17.740 20.160 17.950 ;
        RECT 20.085 16.390 20.160 16.600 ;
        RECT 20.085 15.040 20.160 15.250 ;
        RECT 20.085 13.690 20.160 13.900 ;
        RECT 20.085 12.340 20.160 12.550 ;
        RECT 20.085 10.990 20.160 11.200 ;
        RECT 20.085 9.640 20.160 9.850 ;
        RECT 20.085 8.290 20.160 8.500 ;
        RECT 20.085 6.940 20.160 7.150 ;
        RECT 20.085 5.590 20.160 5.800 ;
        RECT 20.085 4.240 20.160 4.450 ;
        RECT 20.085 2.890 20.160 3.100 ;
        RECT 20.085 1.540 20.160 1.750 ;
        RECT 20.085 0.190 20.160 0.400 ;
    END
  END RBL0_6
  PIN RBL1_7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444800 ;
    PORT
      LAYER li1 ;
        RECT 20.300 42.040 20.375 42.250 ;
        RECT 20.300 40.690 20.375 40.900 ;
        RECT 20.300 39.340 20.375 39.550 ;
        RECT 20.300 37.990 20.375 38.200 ;
        RECT 20.300 36.640 20.375 36.850 ;
        RECT 20.300 35.290 20.375 35.500 ;
        RECT 20.300 33.940 20.375 34.150 ;
        RECT 20.300 32.590 20.375 32.800 ;
        RECT 20.300 31.240 20.375 31.450 ;
        RECT 20.300 29.890 20.375 30.100 ;
        RECT 20.300 28.540 20.375 28.750 ;
        RECT 20.300 27.190 20.375 27.400 ;
        RECT 20.300 25.840 20.375 26.050 ;
        RECT 20.300 24.490 20.375 24.700 ;
        RECT 20.300 23.140 20.375 23.350 ;
        RECT 20.300 21.790 20.375 22.000 ;
        RECT 20.300 20.440 20.375 20.650 ;
        RECT 20.300 19.090 20.375 19.300 ;
        RECT 20.300 17.740 20.375 17.950 ;
        RECT 20.300 16.390 20.375 16.600 ;
        RECT 20.300 15.040 20.375 15.250 ;
        RECT 20.300 13.690 20.375 13.900 ;
        RECT 20.300 12.340 20.375 12.550 ;
        RECT 20.300 10.990 20.375 11.200 ;
        RECT 20.300 9.640 20.375 9.850 ;
        RECT 20.300 8.290 20.375 8.500 ;
        RECT 20.300 6.940 20.375 7.150 ;
        RECT 20.300 5.590 20.375 5.800 ;
        RECT 20.300 4.240 20.375 4.450 ;
        RECT 20.300 2.890 20.375 3.100 ;
        RECT 20.300 1.540 20.375 1.750 ;
        RECT 20.300 0.190 20.375 0.400 ;
    END
  END RBL1_7
  PIN RBL0_7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444800 ;
    PORT
      LAYER li1 ;
        RECT 22.985 42.040 23.060 42.250 ;
        RECT 22.985 40.690 23.060 40.900 ;
        RECT 22.985 39.340 23.060 39.550 ;
        RECT 22.985 37.990 23.060 38.200 ;
        RECT 22.985 36.640 23.060 36.850 ;
        RECT 22.985 35.290 23.060 35.500 ;
        RECT 22.985 33.940 23.060 34.150 ;
        RECT 22.985 32.590 23.060 32.800 ;
        RECT 22.985 31.240 23.060 31.450 ;
        RECT 22.985 29.890 23.060 30.100 ;
        RECT 22.985 28.540 23.060 28.750 ;
        RECT 22.985 27.190 23.060 27.400 ;
        RECT 22.985 25.840 23.060 26.050 ;
        RECT 22.985 24.490 23.060 24.700 ;
        RECT 22.985 23.140 23.060 23.350 ;
        RECT 22.985 21.790 23.060 22.000 ;
        RECT 22.985 20.440 23.060 20.650 ;
        RECT 22.985 19.090 23.060 19.300 ;
        RECT 22.985 17.740 23.060 17.950 ;
        RECT 22.985 16.390 23.060 16.600 ;
        RECT 22.985 15.040 23.060 15.250 ;
        RECT 22.985 13.690 23.060 13.900 ;
        RECT 22.985 12.340 23.060 12.550 ;
        RECT 22.985 10.990 23.060 11.200 ;
        RECT 22.985 9.640 23.060 9.850 ;
        RECT 22.985 8.290 23.060 8.500 ;
        RECT 22.985 6.940 23.060 7.150 ;
        RECT 22.985 5.590 23.060 5.800 ;
        RECT 22.985 4.240 23.060 4.450 ;
        RECT 22.985 2.890 23.060 3.100 ;
        RECT 22.985 1.540 23.060 1.750 ;
        RECT 22.985 0.190 23.060 0.400 ;
    END
  END RBL0_7
  PIN RBL1_8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444800 ;
    PORT
      LAYER li1 ;
        RECT 23.200 42.040 23.275 42.250 ;
        RECT 23.200 40.690 23.275 40.900 ;
        RECT 23.200 39.340 23.275 39.550 ;
        RECT 23.200 37.990 23.275 38.200 ;
        RECT 23.200 36.640 23.275 36.850 ;
        RECT 23.200 35.290 23.275 35.500 ;
        RECT 23.200 33.940 23.275 34.150 ;
        RECT 23.200 32.590 23.275 32.800 ;
        RECT 23.200 31.240 23.275 31.450 ;
        RECT 23.200 29.890 23.275 30.100 ;
        RECT 23.200 28.540 23.275 28.750 ;
        RECT 23.200 27.190 23.275 27.400 ;
        RECT 23.200 25.840 23.275 26.050 ;
        RECT 23.200 24.490 23.275 24.700 ;
        RECT 23.200 23.140 23.275 23.350 ;
        RECT 23.200 21.790 23.275 22.000 ;
        RECT 23.200 20.440 23.275 20.650 ;
        RECT 23.200 19.090 23.275 19.300 ;
        RECT 23.200 17.740 23.275 17.950 ;
        RECT 23.200 16.390 23.275 16.600 ;
        RECT 23.200 15.040 23.275 15.250 ;
        RECT 23.200 13.690 23.275 13.900 ;
        RECT 23.200 12.340 23.275 12.550 ;
        RECT 23.200 10.990 23.275 11.200 ;
        RECT 23.200 9.640 23.275 9.850 ;
        RECT 23.200 8.290 23.275 8.500 ;
        RECT 23.200 6.940 23.275 7.150 ;
        RECT 23.200 5.590 23.275 5.800 ;
        RECT 23.200 4.240 23.275 4.450 ;
        RECT 23.200 2.890 23.275 3.100 ;
        RECT 23.200 1.545 23.275 1.755 ;
        RECT 23.200 0.195 23.275 0.405 ;
    END
  END RBL1_8
  PIN RBL0_8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.445175 ;
    PORT
      LAYER li1 ;
        RECT 25.885 42.040 25.960 42.250 ;
        RECT 25.885 40.690 25.960 40.900 ;
        RECT 25.885 39.340 25.960 39.550 ;
        RECT 25.885 37.990 25.960 38.200 ;
        RECT 25.885 36.640 25.960 36.850 ;
        RECT 25.885 35.290 25.960 35.500 ;
        RECT 25.885 33.940 25.960 34.150 ;
        RECT 25.885 32.590 25.960 32.800 ;
        RECT 25.885 31.240 25.960 31.450 ;
        RECT 25.885 29.890 25.960 30.100 ;
        RECT 25.885 28.540 25.960 28.750 ;
        RECT 25.885 27.190 25.960 27.400 ;
        RECT 25.885 25.840 25.960 26.050 ;
        RECT 25.885 24.490 25.960 24.700 ;
        RECT 25.885 23.140 25.960 23.350 ;
        RECT 25.885 21.790 25.960 22.000 ;
        RECT 25.885 20.440 25.960 20.650 ;
        RECT 25.885 19.090 25.960 19.300 ;
        RECT 25.885 17.740 25.960 17.950 ;
        RECT 25.885 16.390 25.960 16.600 ;
        RECT 25.885 15.040 25.960 15.250 ;
        RECT 25.885 13.690 25.960 13.900 ;
        RECT 25.885 12.340 25.960 12.550 ;
        RECT 25.885 10.990 25.960 11.200 ;
        RECT 25.885 9.640 25.960 9.850 ;
        RECT 25.885 8.290 25.960 8.500 ;
        RECT 25.885 6.940 25.960 7.150 ;
        RECT 25.885 5.590 25.960 5.800 ;
        RECT 25.885 4.240 25.960 4.450 ;
        RECT 25.885 2.890 25.960 3.100 ;
        RECT 25.885 1.545 25.960 1.755 ;
        RECT 25.885 0.190 25.960 0.405 ;
    END
  END RBL0_8
  PIN RBL1_9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.445175 ;
    PORT
      LAYER li1 ;
        RECT 26.100 42.040 26.175 42.250 ;
        RECT 26.100 40.690 26.175 40.900 ;
        RECT 26.100 39.340 26.175 39.550 ;
        RECT 26.100 37.990 26.175 38.200 ;
        RECT 26.100 36.640 26.175 36.850 ;
        RECT 26.100 35.290 26.175 35.500 ;
        RECT 26.100 33.940 26.175 34.150 ;
        RECT 26.100 32.590 26.175 32.800 ;
        RECT 26.100 31.240 26.175 31.450 ;
        RECT 26.100 29.890 26.175 30.100 ;
        RECT 26.100 28.540 26.175 28.750 ;
        RECT 26.100 27.190 26.175 27.400 ;
        RECT 26.100 25.840 26.175 26.050 ;
        RECT 26.100 24.490 26.175 24.700 ;
        RECT 26.100 23.140 26.175 23.350 ;
        RECT 26.100 21.790 26.175 22.000 ;
        RECT 26.100 20.440 26.175 20.650 ;
        RECT 26.100 19.090 26.175 19.300 ;
        RECT 26.100 17.740 26.175 17.950 ;
        RECT 26.100 16.390 26.175 16.600 ;
        RECT 26.100 15.040 26.175 15.250 ;
        RECT 26.100 13.690 26.175 13.900 ;
        RECT 26.100 12.340 26.175 12.550 ;
        RECT 26.100 10.990 26.175 11.200 ;
        RECT 26.100 9.640 26.175 9.850 ;
        RECT 26.100 8.290 26.175 8.500 ;
        RECT 26.100 6.940 26.175 7.150 ;
        RECT 26.100 5.590 26.175 5.800 ;
        RECT 26.100 4.240 26.175 4.450 ;
        RECT 26.100 2.890 26.175 3.100 ;
        RECT 26.100 1.545 26.175 1.755 ;
        RECT 26.100 0.190 26.175 0.405 ;
    END
  END RBL1_9
  PIN RBL0_9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.445175 ;
    PORT
      LAYER li1 ;
        RECT 28.785 42.040 28.860 42.250 ;
        RECT 28.785 40.690 28.860 40.900 ;
        RECT 28.785 39.340 28.860 39.550 ;
        RECT 28.785 37.990 28.860 38.200 ;
        RECT 28.785 36.640 28.860 36.850 ;
        RECT 28.785 35.290 28.860 35.500 ;
        RECT 28.785 33.940 28.860 34.150 ;
        RECT 28.785 32.590 28.860 32.800 ;
        RECT 28.785 31.240 28.860 31.450 ;
        RECT 28.785 29.890 28.860 30.100 ;
        RECT 28.785 28.540 28.860 28.750 ;
        RECT 28.785 27.190 28.860 27.400 ;
        RECT 28.785 25.840 28.860 26.050 ;
        RECT 28.785 24.490 28.860 24.700 ;
        RECT 28.785 23.140 28.860 23.350 ;
        RECT 28.785 21.790 28.860 22.000 ;
        RECT 28.785 20.440 28.860 20.650 ;
        RECT 28.785 19.090 28.860 19.300 ;
        RECT 28.785 17.740 28.860 17.950 ;
        RECT 28.785 16.390 28.860 16.600 ;
        RECT 28.785 15.040 28.860 15.250 ;
        RECT 28.785 13.690 28.860 13.900 ;
        RECT 28.785 12.340 28.860 12.550 ;
        RECT 28.785 10.990 28.860 11.200 ;
        RECT 28.785 9.640 28.860 9.850 ;
        RECT 28.785 8.290 28.860 8.500 ;
        RECT 28.785 6.940 28.860 7.150 ;
        RECT 28.785 5.590 28.860 5.800 ;
        RECT 28.785 4.240 28.860 4.450 ;
        RECT 28.785 2.890 28.860 3.100 ;
        RECT 28.785 1.545 28.860 1.755 ;
        RECT 28.785 0.190 28.860 0.405 ;
    END
  END RBL0_9
  PIN RBL1_10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.445175 ;
    PORT
      LAYER li1 ;
        RECT 29.000 42.040 29.075 42.250 ;
        RECT 29.000 40.690 29.075 40.900 ;
        RECT 29.000 39.340 29.075 39.550 ;
        RECT 29.000 37.990 29.075 38.200 ;
        RECT 29.000 36.640 29.075 36.850 ;
        RECT 29.000 35.290 29.075 35.500 ;
        RECT 29.000 33.940 29.075 34.150 ;
        RECT 29.000 32.590 29.075 32.800 ;
        RECT 29.000 31.240 29.075 31.450 ;
        RECT 29.000 29.890 29.075 30.100 ;
        RECT 29.000 28.540 29.075 28.750 ;
        RECT 29.000 27.190 29.075 27.400 ;
        RECT 29.000 25.840 29.075 26.050 ;
        RECT 29.000 24.490 29.075 24.700 ;
        RECT 29.000 23.140 29.075 23.350 ;
        RECT 29.000 21.790 29.075 22.000 ;
        RECT 29.000 20.440 29.075 20.650 ;
        RECT 29.000 19.090 29.075 19.300 ;
        RECT 29.000 17.740 29.075 17.950 ;
        RECT 29.000 16.390 29.075 16.600 ;
        RECT 29.000 15.040 29.075 15.250 ;
        RECT 29.000 13.690 29.075 13.900 ;
        RECT 29.000 12.340 29.075 12.550 ;
        RECT 29.000 10.990 29.075 11.200 ;
        RECT 29.000 9.640 29.075 9.850 ;
        RECT 29.000 8.290 29.075 8.500 ;
        RECT 29.000 6.940 29.075 7.150 ;
        RECT 29.000 5.590 29.075 5.800 ;
        RECT 29.000 4.240 29.075 4.450 ;
        RECT 29.000 2.890 29.075 3.100 ;
        RECT 29.000 1.545 29.075 1.755 ;
        RECT 29.000 0.190 29.075 0.405 ;
    END
  END RBL1_10
  PIN RBL0_10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.445175 ;
    PORT
      LAYER li1 ;
        RECT 31.685 42.040 31.760 42.250 ;
        RECT 31.685 40.690 31.760 40.900 ;
        RECT 31.685 39.340 31.760 39.550 ;
        RECT 31.685 37.990 31.760 38.200 ;
        RECT 31.685 36.640 31.760 36.850 ;
        RECT 31.685 35.290 31.760 35.500 ;
        RECT 31.685 33.940 31.760 34.150 ;
        RECT 31.685 32.590 31.760 32.800 ;
        RECT 31.685 31.240 31.760 31.450 ;
        RECT 31.685 29.890 31.760 30.100 ;
        RECT 31.685 28.540 31.760 28.750 ;
        RECT 31.685 27.190 31.760 27.400 ;
        RECT 31.685 25.840 31.760 26.050 ;
        RECT 31.685 24.490 31.760 24.700 ;
        RECT 31.685 23.140 31.760 23.350 ;
        RECT 31.685 21.790 31.760 22.000 ;
        RECT 31.685 20.440 31.760 20.650 ;
        RECT 31.685 19.090 31.760 19.300 ;
        RECT 31.685 17.740 31.760 17.950 ;
        RECT 31.685 16.390 31.760 16.600 ;
        RECT 31.685 15.040 31.760 15.250 ;
        RECT 31.685 13.690 31.760 13.900 ;
        RECT 31.685 12.340 31.760 12.550 ;
        RECT 31.685 10.990 31.760 11.200 ;
        RECT 31.685 9.640 31.760 9.850 ;
        RECT 31.685 8.290 31.760 8.500 ;
        RECT 31.685 6.940 31.760 7.150 ;
        RECT 31.685 5.590 31.760 5.800 ;
        RECT 31.685 4.240 31.760 4.450 ;
        RECT 31.685 2.890 31.760 3.100 ;
        RECT 31.685 1.545 31.760 1.755 ;
        RECT 31.685 0.190 31.760 0.405 ;
    END
  END RBL0_10
  PIN RBL1_11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.445175 ;
    PORT
      LAYER li1 ;
        RECT 31.900 42.040 31.975 42.250 ;
        RECT 31.900 40.690 31.975 40.900 ;
        RECT 31.900 39.340 31.975 39.550 ;
        RECT 31.900 37.990 31.975 38.200 ;
        RECT 31.900 36.640 31.975 36.850 ;
        RECT 31.900 35.290 31.975 35.500 ;
        RECT 31.900 33.940 31.975 34.150 ;
        RECT 31.900 32.590 31.975 32.800 ;
        RECT 31.900 31.240 31.975 31.450 ;
        RECT 31.900 29.890 31.975 30.100 ;
        RECT 31.900 28.540 31.975 28.750 ;
        RECT 31.900 27.190 31.975 27.400 ;
        RECT 31.900 25.840 31.975 26.050 ;
        RECT 31.900 24.490 31.975 24.700 ;
        RECT 31.900 23.140 31.975 23.350 ;
        RECT 31.900 21.790 31.975 22.000 ;
        RECT 31.900 20.440 31.975 20.650 ;
        RECT 31.900 19.090 31.975 19.300 ;
        RECT 31.900 17.740 31.975 17.950 ;
        RECT 31.900 16.390 31.975 16.600 ;
        RECT 31.900 15.040 31.975 15.250 ;
        RECT 31.900 13.690 31.975 13.900 ;
        RECT 31.900 12.340 31.975 12.550 ;
        RECT 31.900 10.990 31.975 11.200 ;
        RECT 31.900 9.640 31.975 9.850 ;
        RECT 31.900 8.290 31.975 8.500 ;
        RECT 31.900 6.940 31.975 7.150 ;
        RECT 31.900 5.590 31.975 5.800 ;
        RECT 31.900 4.240 31.975 4.450 ;
        RECT 31.900 2.890 31.975 3.100 ;
        RECT 31.900 1.545 31.975 1.755 ;
        RECT 31.900 0.190 31.975 0.405 ;
    END
  END RBL1_11
  PIN RBL0_11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.445175 ;
    PORT
      LAYER li1 ;
        RECT 34.585 42.040 34.660 42.250 ;
        RECT 34.585 40.690 34.660 40.900 ;
        RECT 34.585 39.340 34.660 39.550 ;
        RECT 34.585 37.990 34.660 38.200 ;
        RECT 34.585 36.640 34.660 36.850 ;
        RECT 34.585 35.290 34.660 35.500 ;
        RECT 34.585 33.940 34.660 34.150 ;
        RECT 34.585 32.590 34.660 32.800 ;
        RECT 34.585 31.240 34.660 31.450 ;
        RECT 34.585 29.890 34.660 30.100 ;
        RECT 34.585 28.540 34.660 28.750 ;
        RECT 34.585 27.190 34.660 27.400 ;
        RECT 34.585 25.840 34.660 26.050 ;
        RECT 34.585 24.490 34.660 24.700 ;
        RECT 34.585 23.140 34.660 23.350 ;
        RECT 34.585 21.790 34.660 22.000 ;
        RECT 34.585 20.440 34.660 20.650 ;
        RECT 34.585 19.090 34.660 19.300 ;
        RECT 34.585 17.740 34.660 17.950 ;
        RECT 34.585 16.390 34.660 16.600 ;
        RECT 34.585 15.040 34.660 15.250 ;
        RECT 34.585 13.690 34.660 13.900 ;
        RECT 34.585 12.340 34.660 12.550 ;
        RECT 34.585 10.990 34.660 11.200 ;
        RECT 34.585 9.640 34.660 9.850 ;
        RECT 34.585 8.290 34.660 8.500 ;
        RECT 34.585 6.940 34.660 7.150 ;
        RECT 34.585 5.590 34.660 5.800 ;
        RECT 34.585 4.240 34.660 4.450 ;
        RECT 34.585 2.890 34.660 3.100 ;
        RECT 34.585 1.545 34.660 1.755 ;
        RECT 34.585 0.190 34.660 0.405 ;
    END
  END RBL0_11
  PIN RBL1_12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.445175 ;
    PORT
      LAYER li1 ;
        RECT 34.800 42.040 34.875 42.250 ;
        RECT 34.800 40.690 34.875 40.900 ;
        RECT 34.800 39.340 34.875 39.550 ;
        RECT 34.800 37.990 34.875 38.200 ;
        RECT 34.800 36.640 34.875 36.850 ;
        RECT 34.800 35.290 34.875 35.500 ;
        RECT 34.800 33.940 34.875 34.150 ;
        RECT 34.800 32.590 34.875 32.800 ;
        RECT 34.800 31.240 34.875 31.450 ;
        RECT 34.800 29.890 34.875 30.100 ;
        RECT 34.800 28.540 34.875 28.750 ;
        RECT 34.800 27.190 34.875 27.400 ;
        RECT 34.800 25.840 34.875 26.050 ;
        RECT 34.800 24.490 34.875 24.700 ;
        RECT 34.800 23.140 34.875 23.350 ;
        RECT 34.800 21.790 34.875 22.000 ;
        RECT 34.800 20.440 34.875 20.650 ;
        RECT 34.800 19.090 34.875 19.300 ;
        RECT 34.800 17.740 34.875 17.950 ;
        RECT 34.800 16.390 34.875 16.600 ;
        RECT 34.800 15.040 34.875 15.250 ;
        RECT 34.800 13.690 34.875 13.900 ;
        RECT 34.800 12.340 34.875 12.550 ;
        RECT 34.800 10.990 34.875 11.200 ;
        RECT 34.800 9.640 34.875 9.850 ;
        RECT 34.800 8.290 34.875 8.500 ;
        RECT 34.800 6.940 34.875 7.150 ;
        RECT 34.800 5.590 34.875 5.800 ;
        RECT 34.800 4.240 34.875 4.450 ;
        RECT 34.800 2.890 34.875 3.100 ;
        RECT 34.800 1.545 34.875 1.755 ;
        RECT 34.800 0.190 34.875 0.405 ;
    END
  END RBL1_12
  PIN RBL0_12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.445175 ;
    PORT
      LAYER li1 ;
        RECT 37.485 42.040 37.560 42.250 ;
        RECT 37.485 40.690 37.560 40.900 ;
        RECT 37.485 39.340 37.560 39.550 ;
        RECT 37.485 37.990 37.560 38.200 ;
        RECT 37.485 36.640 37.560 36.850 ;
        RECT 37.485 35.290 37.560 35.500 ;
        RECT 37.485 33.940 37.560 34.150 ;
        RECT 37.485 32.590 37.560 32.800 ;
        RECT 37.485 31.240 37.560 31.450 ;
        RECT 37.485 29.890 37.560 30.100 ;
        RECT 37.485 28.540 37.560 28.750 ;
        RECT 37.485 27.190 37.560 27.400 ;
        RECT 37.485 25.840 37.560 26.050 ;
        RECT 37.485 24.490 37.560 24.700 ;
        RECT 37.485 23.140 37.560 23.350 ;
        RECT 37.485 21.790 37.560 22.000 ;
        RECT 37.485 20.440 37.560 20.650 ;
        RECT 37.485 19.090 37.560 19.300 ;
        RECT 37.485 17.740 37.560 17.950 ;
        RECT 37.485 16.390 37.560 16.600 ;
        RECT 37.485 15.040 37.560 15.250 ;
        RECT 37.485 13.690 37.560 13.900 ;
        RECT 37.485 12.340 37.560 12.550 ;
        RECT 37.485 10.990 37.560 11.200 ;
        RECT 37.485 9.640 37.560 9.850 ;
        RECT 37.485 8.290 37.560 8.500 ;
        RECT 37.485 6.940 37.560 7.150 ;
        RECT 37.485 5.590 37.560 5.800 ;
        RECT 37.485 4.240 37.560 4.450 ;
        RECT 37.485 2.890 37.560 3.100 ;
        RECT 37.485 1.545 37.560 1.755 ;
        RECT 37.485 0.190 37.560 0.405 ;
    END
  END RBL0_12
  PIN RBL1_13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.445175 ;
    PORT
      LAYER li1 ;
        RECT 37.700 42.040 37.775 42.250 ;
        RECT 37.700 40.690 37.775 40.900 ;
        RECT 37.700 39.340 37.775 39.550 ;
        RECT 37.700 37.990 37.775 38.200 ;
        RECT 37.700 36.640 37.775 36.850 ;
        RECT 37.700 35.290 37.775 35.500 ;
        RECT 37.700 33.940 37.775 34.150 ;
        RECT 37.700 32.590 37.775 32.800 ;
        RECT 37.700 31.240 37.775 31.450 ;
        RECT 37.700 29.890 37.775 30.100 ;
        RECT 37.700 28.540 37.775 28.750 ;
        RECT 37.700 27.190 37.775 27.400 ;
        RECT 37.700 25.840 37.775 26.050 ;
        RECT 37.700 24.490 37.775 24.700 ;
        RECT 37.700 23.140 37.775 23.350 ;
        RECT 37.700 21.790 37.775 22.000 ;
        RECT 37.700 20.440 37.775 20.650 ;
        RECT 37.700 19.090 37.775 19.300 ;
        RECT 37.700 17.740 37.775 17.950 ;
        RECT 37.700 16.390 37.775 16.600 ;
        RECT 37.700 15.040 37.775 15.250 ;
        RECT 37.700 13.690 37.775 13.900 ;
        RECT 37.700 12.340 37.775 12.550 ;
        RECT 37.700 10.990 37.775 11.200 ;
        RECT 37.700 9.640 37.775 9.850 ;
        RECT 37.700 8.290 37.775 8.500 ;
        RECT 37.700 6.940 37.775 7.150 ;
        RECT 37.700 5.590 37.775 5.800 ;
        RECT 37.700 4.240 37.775 4.450 ;
        RECT 37.700 2.890 37.775 3.100 ;
        RECT 37.700 1.545 37.775 1.755 ;
        RECT 37.700 0.190 37.775 0.405 ;
    END
  END RBL1_13
  PIN RBL0_13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.445175 ;
    PORT
      LAYER li1 ;
        RECT 40.385 42.040 40.460 42.250 ;
        RECT 40.385 40.690 40.460 40.900 ;
        RECT 40.385 39.340 40.460 39.550 ;
        RECT 40.385 37.990 40.460 38.200 ;
        RECT 40.385 36.640 40.460 36.850 ;
        RECT 40.385 35.290 40.460 35.500 ;
        RECT 40.385 33.940 40.460 34.150 ;
        RECT 40.385 32.590 40.460 32.800 ;
        RECT 40.385 31.240 40.460 31.450 ;
        RECT 40.385 29.890 40.460 30.100 ;
        RECT 40.385 28.540 40.460 28.750 ;
        RECT 40.385 27.190 40.460 27.400 ;
        RECT 40.385 25.840 40.460 26.050 ;
        RECT 40.385 24.490 40.460 24.700 ;
        RECT 40.385 23.140 40.460 23.350 ;
        RECT 40.385 21.790 40.460 22.000 ;
        RECT 40.385 20.440 40.460 20.650 ;
        RECT 40.385 19.090 40.460 19.300 ;
        RECT 40.385 17.740 40.460 17.950 ;
        RECT 40.385 16.390 40.460 16.600 ;
        RECT 40.385 15.040 40.460 15.250 ;
        RECT 40.385 13.690 40.460 13.900 ;
        RECT 40.385 12.340 40.460 12.550 ;
        RECT 40.385 10.990 40.460 11.200 ;
        RECT 40.385 9.640 40.460 9.850 ;
        RECT 40.385 8.290 40.460 8.500 ;
        RECT 40.385 6.940 40.460 7.150 ;
        RECT 40.385 5.590 40.460 5.800 ;
        RECT 40.385 4.240 40.460 4.450 ;
        RECT 40.385 2.890 40.460 3.100 ;
        RECT 40.385 1.545 40.460 1.755 ;
        RECT 40.385 0.190 40.460 0.405 ;
    END
  END RBL0_13
  PIN RBL1_14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.445175 ;
    PORT
      LAYER li1 ;
        RECT 40.600 42.040 40.675 42.250 ;
        RECT 40.600 40.690 40.675 40.900 ;
        RECT 40.600 39.340 40.675 39.550 ;
        RECT 40.600 37.990 40.675 38.200 ;
        RECT 40.600 36.640 40.675 36.850 ;
        RECT 40.600 35.290 40.675 35.500 ;
        RECT 40.600 33.940 40.675 34.150 ;
        RECT 40.600 32.590 40.675 32.800 ;
        RECT 40.600 31.240 40.675 31.450 ;
        RECT 40.600 29.890 40.675 30.100 ;
        RECT 40.600 28.540 40.675 28.750 ;
        RECT 40.600 27.190 40.675 27.400 ;
        RECT 40.600 25.840 40.675 26.050 ;
        RECT 40.600 24.490 40.675 24.700 ;
        RECT 40.600 23.140 40.675 23.350 ;
        RECT 40.600 21.790 40.675 22.000 ;
        RECT 40.600 20.440 40.675 20.650 ;
        RECT 40.600 19.090 40.675 19.300 ;
        RECT 40.600 17.740 40.675 17.950 ;
        RECT 40.600 16.390 40.675 16.600 ;
        RECT 40.600 15.040 40.675 15.250 ;
        RECT 40.600 13.690 40.675 13.900 ;
        RECT 40.600 12.340 40.675 12.550 ;
        RECT 40.600 10.990 40.675 11.200 ;
        RECT 40.600 9.640 40.675 9.850 ;
        RECT 40.600 8.290 40.675 8.500 ;
        RECT 40.600 6.940 40.675 7.150 ;
        RECT 40.600 5.590 40.675 5.800 ;
        RECT 40.600 4.240 40.675 4.450 ;
        RECT 40.600 2.890 40.675 3.100 ;
        RECT 40.600 1.545 40.675 1.755 ;
        RECT 40.600 0.190 40.675 0.405 ;
    END
  END RBL1_14
  PIN RBL0_14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.445175 ;
    PORT
      LAYER li1 ;
        RECT 43.285 42.040 43.360 42.250 ;
        RECT 43.285 40.690 43.360 40.900 ;
        RECT 43.285 39.340 43.360 39.550 ;
        RECT 43.285 37.990 43.360 38.200 ;
        RECT 43.285 36.640 43.360 36.850 ;
        RECT 43.285 35.290 43.360 35.500 ;
        RECT 43.285 33.940 43.360 34.150 ;
        RECT 43.285 32.590 43.360 32.800 ;
        RECT 43.285 31.240 43.360 31.450 ;
        RECT 43.285 29.890 43.360 30.100 ;
        RECT 43.285 28.540 43.360 28.750 ;
        RECT 43.285 27.190 43.360 27.400 ;
        RECT 43.285 25.840 43.360 26.050 ;
        RECT 43.285 24.490 43.360 24.700 ;
        RECT 43.285 23.140 43.360 23.350 ;
        RECT 43.285 21.790 43.360 22.000 ;
        RECT 43.285 20.440 43.360 20.650 ;
        RECT 43.285 19.090 43.360 19.300 ;
        RECT 43.285 17.740 43.360 17.950 ;
        RECT 43.285 16.390 43.360 16.600 ;
        RECT 43.285 15.040 43.360 15.250 ;
        RECT 43.285 13.690 43.360 13.900 ;
        RECT 43.285 12.340 43.360 12.550 ;
        RECT 43.285 10.990 43.360 11.200 ;
        RECT 43.285 9.640 43.360 9.850 ;
        RECT 43.285 8.290 43.360 8.500 ;
        RECT 43.285 6.940 43.360 7.150 ;
        RECT 43.285 5.590 43.360 5.800 ;
        RECT 43.285 4.240 43.360 4.450 ;
        RECT 43.285 2.890 43.360 3.100 ;
        RECT 43.285 1.545 43.360 1.755 ;
        RECT 43.285 0.190 43.360 0.405 ;
    END
  END RBL0_14
  PIN RBL1_15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.445175 ;
    PORT
      LAYER li1 ;
        RECT 43.500 42.040 43.575 42.250 ;
        RECT 43.500 40.690 43.575 40.900 ;
        RECT 43.500 39.340 43.575 39.550 ;
        RECT 43.500 37.990 43.575 38.200 ;
        RECT 43.500 36.640 43.575 36.850 ;
        RECT 43.500 35.290 43.575 35.500 ;
        RECT 43.500 33.940 43.575 34.150 ;
        RECT 43.500 32.590 43.575 32.800 ;
        RECT 43.500 31.240 43.575 31.450 ;
        RECT 43.500 29.890 43.575 30.100 ;
        RECT 43.500 28.540 43.575 28.750 ;
        RECT 43.500 27.190 43.575 27.400 ;
        RECT 43.500 25.840 43.575 26.050 ;
        RECT 43.500 24.490 43.575 24.700 ;
        RECT 43.500 23.140 43.575 23.350 ;
        RECT 43.500 21.790 43.575 22.000 ;
        RECT 43.500 20.440 43.575 20.650 ;
        RECT 43.500 19.090 43.575 19.300 ;
        RECT 43.500 17.740 43.575 17.950 ;
        RECT 43.500 16.390 43.575 16.600 ;
        RECT 43.500 15.040 43.575 15.250 ;
        RECT 43.500 13.690 43.575 13.900 ;
        RECT 43.500 12.340 43.575 12.550 ;
        RECT 43.500 10.990 43.575 11.200 ;
        RECT 43.500 9.640 43.575 9.850 ;
        RECT 43.500 8.290 43.575 8.500 ;
        RECT 43.500 6.940 43.575 7.150 ;
        RECT 43.500 5.590 43.575 5.800 ;
        RECT 43.500 4.240 43.575 4.450 ;
        RECT 43.500 2.890 43.575 3.100 ;
        RECT 43.500 1.545 43.575 1.755 ;
        RECT 43.500 0.190 43.575 0.405 ;
    END
  END RBL1_15
  PIN RBL0_15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.445175 ;
    PORT
      LAYER li1 ;
        RECT 46.185 42.040 46.260 42.250 ;
        RECT 46.185 40.690 46.260 40.900 ;
        RECT 46.185 39.340 46.260 39.550 ;
        RECT 46.185 37.990 46.260 38.200 ;
        RECT 46.185 36.640 46.260 36.850 ;
        RECT 46.185 35.290 46.260 35.500 ;
        RECT 46.185 33.940 46.260 34.150 ;
        RECT 46.185 32.590 46.260 32.800 ;
        RECT 46.185 31.240 46.260 31.450 ;
        RECT 46.185 29.890 46.260 30.100 ;
        RECT 46.185 28.540 46.260 28.750 ;
        RECT 46.185 27.190 46.260 27.400 ;
        RECT 46.185 25.840 46.260 26.050 ;
        RECT 46.185 24.490 46.260 24.700 ;
        RECT 46.185 23.140 46.260 23.350 ;
        RECT 46.185 21.790 46.260 22.000 ;
        RECT 46.185 20.440 46.260 20.650 ;
        RECT 46.185 19.090 46.260 19.300 ;
        RECT 46.185 17.740 46.260 17.950 ;
        RECT 46.185 16.390 46.260 16.600 ;
        RECT 46.185 15.040 46.260 15.250 ;
        RECT 46.185 13.690 46.260 13.900 ;
        RECT 46.185 12.340 46.260 12.550 ;
        RECT 46.185 10.990 46.260 11.200 ;
        RECT 46.185 9.640 46.260 9.850 ;
        RECT 46.185 8.290 46.260 8.500 ;
        RECT 46.185 6.940 46.260 7.150 ;
        RECT 46.185 5.590 46.260 5.800 ;
        RECT 46.185 4.240 46.260 4.450 ;
        RECT 46.185 2.890 46.260 3.100 ;
        RECT 46.185 1.545 46.260 1.755 ;
        RECT 46.185 0.190 46.260 0.405 ;
    END
  END RBL0_15
  PIN RWL_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 42.360 0.365 42.530 ;
        RECT 2.395 42.360 2.545 42.530 ;
        RECT 3.115 42.360 3.265 42.530 ;
        RECT 5.295 42.360 5.445 42.530 ;
        RECT 6.015 42.360 6.165 42.530 ;
        RECT 8.195 42.360 8.345 42.530 ;
        RECT 8.915 42.360 9.065 42.530 ;
        RECT 11.095 42.360 11.245 42.530 ;
        RECT 11.815 42.360 11.965 42.530 ;
        RECT 13.995 42.360 14.145 42.530 ;
        RECT 14.715 42.360 14.865 42.530 ;
        RECT 16.895 42.360 17.045 42.530 ;
        RECT 17.615 42.360 17.765 42.530 ;
        RECT 19.795 42.360 19.945 42.530 ;
        RECT 20.515 42.360 20.665 42.530 ;
        RECT 22.695 42.360 22.845 42.530 ;
        RECT 23.415 42.360 23.565 42.530 ;
        RECT 25.595 42.360 25.745 42.530 ;
        RECT 26.315 42.360 26.465 42.530 ;
        RECT 28.495 42.360 28.645 42.530 ;
        RECT 29.215 42.360 29.365 42.530 ;
        RECT 31.395 42.360 31.545 42.530 ;
        RECT 32.115 42.360 32.265 42.530 ;
        RECT 34.295 42.360 34.445 42.530 ;
        RECT 35.015 42.360 35.165 42.530 ;
        RECT 37.195 42.360 37.345 42.530 ;
        RECT 37.915 42.360 38.065 42.530 ;
        RECT 40.095 42.360 40.245 42.530 ;
        RECT 40.815 42.360 40.965 42.530 ;
        RECT 42.995 42.360 43.145 42.530 ;
        RECT 43.715 42.360 43.865 42.530 ;
        RECT 45.895 42.360 46.045 42.530 ;
        RECT 46.615 42.360 46.765 42.530 ;
        RECT 48.795 42.360 48.945 42.530 ;
        RECT 49.515 42.360 49.665 42.530 ;
        RECT 51.695 42.360 51.845 42.530 ;
        RECT 52.415 42.360 52.565 42.530 ;
        RECT 54.595 42.360 54.745 42.530 ;
        RECT 55.315 42.360 55.465 42.530 ;
        RECT 57.495 42.360 57.645 42.530 ;
        RECT 58.215 42.360 58.365 42.530 ;
        RECT 60.395 42.360 60.545 42.530 ;
        RECT 61.115 42.360 61.265 42.530 ;
        RECT 63.295 42.360 63.445 42.530 ;
        RECT 64.015 42.360 64.165 42.530 ;
        RECT 66.195 42.360 66.345 42.530 ;
        RECT 66.915 42.360 67.065 42.530 ;
        RECT 69.095 42.360 69.245 42.530 ;
        RECT 69.815 42.360 69.965 42.530 ;
        RECT 71.995 42.360 72.145 42.530 ;
        RECT 72.715 42.360 72.865 42.530 ;
        RECT 74.895 42.360 75.045 42.530 ;
        RECT 75.615 42.360 75.765 42.530 ;
        RECT 77.795 42.360 77.945 42.530 ;
        RECT 78.515 42.360 78.665 42.530 ;
        RECT 80.695 42.360 80.845 42.530 ;
        RECT 81.415 42.360 81.565 42.530 ;
        RECT 83.595 42.360 83.745 42.530 ;
        RECT 84.315 42.360 84.465 42.530 ;
        RECT 86.495 42.360 86.645 42.530 ;
        RECT 87.215 42.360 87.365 42.530 ;
        RECT 89.395 42.360 89.545 42.530 ;
        RECT 90.115 42.360 90.265 42.530 ;
        RECT 92.295 42.360 92.445 42.530 ;
      LAYER met1 ;
        RECT 0.000 42.360 92.445 42.530 ;
    END
  END RWL_0
  PIN RWL_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 41.010 0.365 41.180 ;
        RECT 2.395 41.010 2.545 41.180 ;
        RECT 3.115 41.010 3.265 41.180 ;
        RECT 5.295 41.010 5.445 41.180 ;
        RECT 6.015 41.010 6.165 41.180 ;
        RECT 8.195 41.010 8.345 41.180 ;
        RECT 8.915 41.010 9.065 41.180 ;
        RECT 11.095 41.010 11.245 41.180 ;
        RECT 11.815 41.010 11.965 41.180 ;
        RECT 13.995 41.010 14.145 41.180 ;
        RECT 14.715 41.010 14.865 41.180 ;
        RECT 16.895 41.010 17.045 41.180 ;
        RECT 17.615 41.010 17.765 41.180 ;
        RECT 19.795 41.010 19.945 41.180 ;
        RECT 20.515 41.010 20.665 41.180 ;
        RECT 22.695 41.010 22.845 41.180 ;
        RECT 23.415 41.010 23.565 41.180 ;
        RECT 25.595 41.010 25.745 41.180 ;
        RECT 26.315 41.010 26.465 41.180 ;
        RECT 28.495 41.010 28.645 41.180 ;
        RECT 29.215 41.010 29.365 41.180 ;
        RECT 31.395 41.010 31.545 41.180 ;
        RECT 32.115 41.010 32.265 41.180 ;
        RECT 34.295 41.010 34.445 41.180 ;
        RECT 35.015 41.010 35.165 41.180 ;
        RECT 37.195 41.010 37.345 41.180 ;
        RECT 37.915 41.010 38.065 41.180 ;
        RECT 40.095 41.010 40.245 41.180 ;
        RECT 40.815 41.010 40.965 41.180 ;
        RECT 42.995 41.010 43.145 41.180 ;
        RECT 43.715 41.010 43.865 41.180 ;
        RECT 45.895 41.010 46.045 41.180 ;
        RECT 46.615 41.010 46.765 41.180 ;
        RECT 48.795 41.010 48.945 41.180 ;
        RECT 49.515 41.010 49.665 41.180 ;
        RECT 51.695 41.010 51.845 41.180 ;
        RECT 52.415 41.010 52.565 41.180 ;
        RECT 54.595 41.010 54.745 41.180 ;
        RECT 55.315 41.010 55.465 41.180 ;
        RECT 57.495 41.010 57.645 41.180 ;
        RECT 58.215 41.010 58.365 41.180 ;
        RECT 60.395 41.010 60.545 41.180 ;
        RECT 61.115 41.010 61.265 41.180 ;
        RECT 63.295 41.010 63.445 41.180 ;
        RECT 64.015 41.010 64.165 41.180 ;
        RECT 66.195 41.010 66.345 41.180 ;
        RECT 66.915 41.010 67.065 41.180 ;
        RECT 69.095 41.010 69.245 41.180 ;
        RECT 69.815 41.010 69.965 41.180 ;
        RECT 71.995 41.010 72.145 41.180 ;
        RECT 72.715 41.010 72.865 41.180 ;
        RECT 74.895 41.010 75.045 41.180 ;
        RECT 75.615 41.010 75.765 41.180 ;
        RECT 77.795 41.010 77.945 41.180 ;
        RECT 78.515 41.010 78.665 41.180 ;
        RECT 80.695 41.010 80.845 41.180 ;
        RECT 81.415 41.010 81.565 41.180 ;
        RECT 83.595 41.010 83.745 41.180 ;
        RECT 84.315 41.010 84.465 41.180 ;
        RECT 86.495 41.010 86.645 41.180 ;
        RECT 87.215 41.010 87.365 41.180 ;
        RECT 89.395 41.010 89.545 41.180 ;
        RECT 90.115 41.010 90.265 41.180 ;
        RECT 92.295 41.010 92.445 41.180 ;
      LAYER met1 ;
        RECT 0.000 41.010 92.445 41.180 ;
    END
  END RWL_1
  PIN RWL_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 39.660 0.365 39.830 ;
        RECT 2.395 39.660 2.545 39.830 ;
        RECT 3.115 39.660 3.265 39.830 ;
        RECT 5.295 39.660 5.445 39.830 ;
        RECT 6.015 39.660 6.165 39.830 ;
        RECT 8.195 39.660 8.345 39.830 ;
        RECT 8.915 39.660 9.065 39.830 ;
        RECT 11.095 39.660 11.245 39.830 ;
        RECT 11.815 39.660 11.965 39.830 ;
        RECT 13.995 39.660 14.145 39.830 ;
        RECT 14.715 39.660 14.865 39.830 ;
        RECT 16.895 39.660 17.045 39.830 ;
        RECT 17.615 39.660 17.765 39.830 ;
        RECT 19.795 39.660 19.945 39.830 ;
        RECT 20.515 39.660 20.665 39.830 ;
        RECT 22.695 39.660 22.845 39.830 ;
        RECT 23.415 39.660 23.565 39.830 ;
        RECT 25.595 39.660 25.745 39.830 ;
        RECT 26.315 39.660 26.465 39.830 ;
        RECT 28.495 39.660 28.645 39.830 ;
        RECT 29.215 39.660 29.365 39.830 ;
        RECT 31.395 39.660 31.545 39.830 ;
        RECT 32.115 39.660 32.265 39.830 ;
        RECT 34.295 39.660 34.445 39.830 ;
        RECT 35.015 39.660 35.165 39.830 ;
        RECT 37.195 39.660 37.345 39.830 ;
        RECT 37.915 39.660 38.065 39.830 ;
        RECT 40.095 39.660 40.245 39.830 ;
        RECT 40.815 39.660 40.965 39.830 ;
        RECT 42.995 39.660 43.145 39.830 ;
        RECT 43.715 39.660 43.865 39.830 ;
        RECT 45.895 39.660 46.045 39.830 ;
        RECT 46.615 39.660 46.765 39.830 ;
        RECT 48.795 39.660 48.945 39.830 ;
        RECT 49.515 39.660 49.665 39.830 ;
        RECT 51.695 39.660 51.845 39.830 ;
        RECT 52.415 39.660 52.565 39.830 ;
        RECT 54.595 39.660 54.745 39.830 ;
        RECT 55.315 39.660 55.465 39.830 ;
        RECT 57.495 39.660 57.645 39.830 ;
        RECT 58.215 39.660 58.365 39.830 ;
        RECT 60.395 39.660 60.545 39.830 ;
        RECT 61.115 39.660 61.265 39.830 ;
        RECT 63.295 39.660 63.445 39.830 ;
        RECT 64.015 39.660 64.165 39.830 ;
        RECT 66.195 39.660 66.345 39.830 ;
        RECT 66.915 39.660 67.065 39.830 ;
        RECT 69.095 39.660 69.245 39.830 ;
        RECT 69.815 39.660 69.965 39.830 ;
        RECT 71.995 39.660 72.145 39.830 ;
        RECT 72.715 39.660 72.865 39.830 ;
        RECT 74.895 39.660 75.045 39.830 ;
        RECT 75.615 39.660 75.765 39.830 ;
        RECT 77.795 39.660 77.945 39.830 ;
        RECT 78.515 39.660 78.665 39.830 ;
        RECT 80.695 39.660 80.845 39.830 ;
        RECT 81.415 39.660 81.565 39.830 ;
        RECT 83.595 39.660 83.745 39.830 ;
        RECT 84.315 39.660 84.465 39.830 ;
        RECT 86.495 39.660 86.645 39.830 ;
        RECT 87.215 39.660 87.365 39.830 ;
        RECT 89.395 39.660 89.545 39.830 ;
        RECT 90.115 39.660 90.265 39.830 ;
        RECT 92.295 39.660 92.445 39.830 ;
      LAYER met1 ;
        RECT 0.000 39.660 92.445 39.830 ;
    END
  END RWL_2
  PIN RWL_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.504000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 38.310 0.365 38.480 ;
        RECT 2.395 38.310 2.545 38.480 ;
        RECT 3.115 38.310 3.265 38.480 ;
        RECT 5.295 38.310 5.445 38.480 ;
        RECT 6.015 38.310 6.165 38.480 ;
        RECT 8.195 38.310 8.345 38.480 ;
        RECT 8.915 38.310 9.065 38.480 ;
        RECT 11.095 38.310 11.245 38.480 ;
        RECT 11.815 38.310 11.965 38.480 ;
        RECT 13.995 38.310 14.145 38.480 ;
        RECT 14.715 38.310 14.865 38.480 ;
        RECT 16.895 38.310 17.045 38.480 ;
        RECT 17.615 38.310 17.765 38.480 ;
        RECT 19.795 38.310 19.945 38.480 ;
        RECT 20.515 38.310 20.665 38.480 ;
        RECT 22.695 38.310 22.845 38.480 ;
      LAYER met1 ;
        RECT 0.000 38.310 22.845 38.480 ;
    END
  END RWL_3
  PIN RWL_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 36.960 0.365 37.130 ;
        RECT 2.395 36.960 2.545 37.130 ;
        RECT 3.115 36.960 3.265 37.130 ;
        RECT 5.295 36.960 5.445 37.130 ;
        RECT 6.015 36.960 6.165 37.130 ;
        RECT 8.195 36.960 8.345 37.130 ;
        RECT 8.915 36.960 9.065 37.130 ;
        RECT 11.095 36.960 11.245 37.130 ;
        RECT 11.815 36.960 11.965 37.130 ;
        RECT 13.995 36.960 14.145 37.130 ;
        RECT 14.715 36.960 14.865 37.130 ;
        RECT 16.895 36.960 17.045 37.130 ;
        RECT 17.615 36.960 17.765 37.130 ;
        RECT 19.795 36.960 19.945 37.130 ;
        RECT 20.515 36.960 20.665 37.130 ;
        RECT 22.695 36.960 22.845 37.130 ;
        RECT 23.415 36.960 23.565 37.130 ;
        RECT 25.595 36.960 25.745 37.130 ;
        RECT 26.315 36.960 26.465 37.130 ;
        RECT 28.495 36.960 28.645 37.130 ;
        RECT 29.215 36.960 29.365 37.130 ;
        RECT 31.395 36.960 31.545 37.130 ;
        RECT 32.115 36.960 32.265 37.130 ;
        RECT 34.295 36.960 34.445 37.130 ;
        RECT 35.015 36.960 35.165 37.130 ;
        RECT 37.195 36.960 37.345 37.130 ;
        RECT 37.915 36.960 38.065 37.130 ;
        RECT 40.095 36.960 40.245 37.130 ;
        RECT 40.815 36.960 40.965 37.130 ;
        RECT 42.995 36.960 43.145 37.130 ;
        RECT 43.715 36.960 43.865 37.130 ;
        RECT 45.895 36.960 46.045 37.130 ;
        RECT 46.615 36.960 46.765 37.130 ;
        RECT 48.795 36.960 48.945 37.130 ;
        RECT 49.515 36.960 49.665 37.130 ;
        RECT 51.695 36.960 51.845 37.130 ;
        RECT 52.415 36.960 52.565 37.130 ;
        RECT 54.595 36.960 54.745 37.130 ;
        RECT 55.315 36.960 55.465 37.130 ;
        RECT 57.495 36.960 57.645 37.130 ;
        RECT 58.215 36.960 58.365 37.130 ;
        RECT 60.395 36.960 60.545 37.130 ;
        RECT 61.115 36.960 61.265 37.130 ;
        RECT 63.295 36.960 63.445 37.130 ;
        RECT 64.015 36.960 64.165 37.130 ;
        RECT 66.195 36.960 66.345 37.130 ;
        RECT 66.915 36.960 67.065 37.130 ;
        RECT 69.095 36.960 69.245 37.130 ;
        RECT 69.815 36.960 69.965 37.130 ;
        RECT 71.995 36.960 72.145 37.130 ;
        RECT 72.715 36.960 72.865 37.130 ;
        RECT 74.895 36.960 75.045 37.130 ;
        RECT 75.615 36.960 75.765 37.130 ;
        RECT 77.795 36.960 77.945 37.130 ;
        RECT 78.515 36.960 78.665 37.130 ;
        RECT 80.695 36.960 80.845 37.130 ;
        RECT 81.415 36.960 81.565 37.130 ;
        RECT 83.595 36.960 83.745 37.130 ;
        RECT 84.315 36.960 84.465 37.130 ;
        RECT 86.495 36.960 86.645 37.130 ;
        RECT 87.215 36.960 87.365 37.130 ;
        RECT 89.395 36.960 89.545 37.130 ;
        RECT 90.115 36.960 90.265 37.130 ;
        RECT 92.295 36.960 92.445 37.130 ;
      LAYER met1 ;
        RECT 0.000 36.960 92.445 37.130 ;
    END
  END RWL_4
  PIN RWL_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 35.610 0.365 35.780 ;
        RECT 2.395 35.610 2.545 35.780 ;
        RECT 3.115 35.610 3.265 35.780 ;
        RECT 5.295 35.610 5.445 35.780 ;
        RECT 6.015 35.610 6.165 35.780 ;
        RECT 8.195 35.610 8.345 35.780 ;
        RECT 8.915 35.610 9.065 35.780 ;
        RECT 11.095 35.610 11.245 35.780 ;
        RECT 11.815 35.610 11.965 35.780 ;
        RECT 13.995 35.610 14.145 35.780 ;
        RECT 14.715 35.610 14.865 35.780 ;
        RECT 16.895 35.610 17.045 35.780 ;
        RECT 17.615 35.610 17.765 35.780 ;
        RECT 19.795 35.610 19.945 35.780 ;
        RECT 20.515 35.610 20.665 35.780 ;
        RECT 22.695 35.610 22.845 35.780 ;
        RECT 23.415 35.610 23.565 35.780 ;
        RECT 25.595 35.610 25.745 35.780 ;
        RECT 26.315 35.610 26.465 35.780 ;
        RECT 28.495 35.610 28.645 35.780 ;
        RECT 29.215 35.610 29.365 35.780 ;
        RECT 31.395 35.610 31.545 35.780 ;
        RECT 32.115 35.610 32.265 35.780 ;
        RECT 34.295 35.610 34.445 35.780 ;
        RECT 35.015 35.610 35.165 35.780 ;
        RECT 37.195 35.610 37.345 35.780 ;
        RECT 37.915 35.610 38.065 35.780 ;
        RECT 40.095 35.610 40.245 35.780 ;
        RECT 40.815 35.610 40.965 35.780 ;
        RECT 42.995 35.610 43.145 35.780 ;
        RECT 43.715 35.610 43.865 35.780 ;
        RECT 45.895 35.610 46.045 35.780 ;
        RECT 46.615 35.610 46.765 35.780 ;
        RECT 48.795 35.610 48.945 35.780 ;
        RECT 49.515 35.610 49.665 35.780 ;
        RECT 51.695 35.610 51.845 35.780 ;
        RECT 52.415 35.610 52.565 35.780 ;
        RECT 54.595 35.610 54.745 35.780 ;
        RECT 55.315 35.610 55.465 35.780 ;
        RECT 57.495 35.610 57.645 35.780 ;
        RECT 58.215 35.610 58.365 35.780 ;
        RECT 60.395 35.610 60.545 35.780 ;
        RECT 61.115 35.610 61.265 35.780 ;
        RECT 63.295 35.610 63.445 35.780 ;
        RECT 64.015 35.610 64.165 35.780 ;
        RECT 66.195 35.610 66.345 35.780 ;
        RECT 66.915 35.610 67.065 35.780 ;
        RECT 69.095 35.610 69.245 35.780 ;
        RECT 69.815 35.610 69.965 35.780 ;
        RECT 71.995 35.610 72.145 35.780 ;
        RECT 72.715 35.610 72.865 35.780 ;
        RECT 74.895 35.610 75.045 35.780 ;
        RECT 75.615 35.610 75.765 35.780 ;
        RECT 77.795 35.610 77.945 35.780 ;
        RECT 78.515 35.610 78.665 35.780 ;
        RECT 80.695 35.610 80.845 35.780 ;
        RECT 81.415 35.610 81.565 35.780 ;
        RECT 83.595 35.610 83.745 35.780 ;
        RECT 84.315 35.610 84.465 35.780 ;
        RECT 86.495 35.610 86.645 35.780 ;
        RECT 87.215 35.610 87.365 35.780 ;
        RECT 89.395 35.610 89.545 35.780 ;
        RECT 90.115 35.610 90.265 35.780 ;
        RECT 92.295 35.610 92.445 35.780 ;
      LAYER met1 ;
        RECT 0.000 35.610 92.445 35.780 ;
    END
  END RWL_5
  PIN RWL_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 34.260 0.365 34.430 ;
        RECT 2.395 34.260 2.545 34.430 ;
        RECT 3.115 34.260 3.265 34.430 ;
        RECT 5.295 34.260 5.445 34.430 ;
        RECT 6.015 34.260 6.165 34.430 ;
        RECT 8.195 34.260 8.345 34.430 ;
        RECT 8.915 34.260 9.065 34.430 ;
        RECT 11.095 34.260 11.245 34.430 ;
        RECT 11.815 34.260 11.965 34.430 ;
        RECT 13.995 34.260 14.145 34.430 ;
        RECT 14.715 34.260 14.865 34.430 ;
        RECT 16.895 34.260 17.045 34.430 ;
        RECT 17.615 34.260 17.765 34.430 ;
        RECT 19.795 34.260 19.945 34.430 ;
        RECT 20.515 34.260 20.665 34.430 ;
        RECT 22.695 34.260 22.845 34.430 ;
        RECT 23.415 34.260 23.565 34.430 ;
        RECT 25.595 34.260 25.745 34.430 ;
        RECT 26.315 34.260 26.465 34.430 ;
        RECT 28.495 34.260 28.645 34.430 ;
        RECT 29.215 34.260 29.365 34.430 ;
        RECT 31.395 34.260 31.545 34.430 ;
        RECT 32.115 34.260 32.265 34.430 ;
        RECT 34.295 34.260 34.445 34.430 ;
        RECT 35.015 34.260 35.165 34.430 ;
        RECT 37.195 34.260 37.345 34.430 ;
        RECT 37.915 34.260 38.065 34.430 ;
        RECT 40.095 34.260 40.245 34.430 ;
        RECT 40.815 34.260 40.965 34.430 ;
        RECT 42.995 34.260 43.145 34.430 ;
        RECT 43.715 34.260 43.865 34.430 ;
        RECT 45.895 34.260 46.045 34.430 ;
        RECT 46.615 34.260 46.765 34.430 ;
        RECT 48.795 34.260 48.945 34.430 ;
        RECT 49.515 34.260 49.665 34.430 ;
        RECT 51.695 34.260 51.845 34.430 ;
        RECT 52.415 34.260 52.565 34.430 ;
        RECT 54.595 34.260 54.745 34.430 ;
        RECT 55.315 34.260 55.465 34.430 ;
        RECT 57.495 34.260 57.645 34.430 ;
        RECT 58.215 34.260 58.365 34.430 ;
        RECT 60.395 34.260 60.545 34.430 ;
        RECT 61.115 34.260 61.265 34.430 ;
        RECT 63.295 34.260 63.445 34.430 ;
        RECT 64.015 34.260 64.165 34.430 ;
        RECT 66.195 34.260 66.345 34.430 ;
        RECT 66.915 34.260 67.065 34.430 ;
        RECT 69.095 34.260 69.245 34.430 ;
        RECT 69.815 34.260 69.965 34.430 ;
        RECT 71.995 34.260 72.145 34.430 ;
        RECT 72.715 34.260 72.865 34.430 ;
        RECT 74.895 34.260 75.045 34.430 ;
        RECT 75.615 34.260 75.765 34.430 ;
        RECT 77.795 34.260 77.945 34.430 ;
        RECT 78.515 34.260 78.665 34.430 ;
        RECT 80.695 34.260 80.845 34.430 ;
        RECT 81.415 34.260 81.565 34.430 ;
        RECT 83.595 34.260 83.745 34.430 ;
        RECT 84.315 34.260 84.465 34.430 ;
        RECT 86.495 34.260 86.645 34.430 ;
        RECT 87.215 34.260 87.365 34.430 ;
        RECT 89.395 34.260 89.545 34.430 ;
        RECT 90.115 34.260 90.265 34.430 ;
        RECT 92.295 34.260 92.445 34.430 ;
      LAYER met1 ;
        RECT 0.000 34.260 92.445 34.430 ;
    END
  END RWL_6
  PIN RWL_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 32.910 0.365 33.080 ;
        RECT 2.395 32.910 2.545 33.080 ;
        RECT 3.115 32.910 3.265 33.080 ;
        RECT 5.295 32.910 5.445 33.080 ;
        RECT 6.015 32.910 6.165 33.080 ;
        RECT 8.195 32.910 8.345 33.080 ;
        RECT 8.915 32.910 9.065 33.080 ;
        RECT 11.095 32.910 11.245 33.080 ;
        RECT 11.815 32.910 11.965 33.080 ;
        RECT 13.995 32.910 14.145 33.080 ;
        RECT 14.715 32.910 14.865 33.080 ;
        RECT 16.895 32.910 17.045 33.080 ;
        RECT 17.615 32.910 17.765 33.080 ;
        RECT 19.795 32.910 19.945 33.080 ;
        RECT 20.515 32.910 20.665 33.080 ;
        RECT 22.695 32.910 22.845 33.080 ;
        RECT 23.415 32.910 23.565 33.080 ;
        RECT 25.595 32.910 25.745 33.080 ;
        RECT 26.315 32.910 26.465 33.080 ;
        RECT 28.495 32.910 28.645 33.080 ;
        RECT 29.215 32.910 29.365 33.080 ;
        RECT 31.395 32.910 31.545 33.080 ;
        RECT 32.115 32.910 32.265 33.080 ;
        RECT 34.295 32.910 34.445 33.080 ;
        RECT 35.015 32.910 35.165 33.080 ;
        RECT 37.195 32.910 37.345 33.080 ;
        RECT 37.915 32.910 38.065 33.080 ;
        RECT 40.095 32.910 40.245 33.080 ;
        RECT 40.815 32.910 40.965 33.080 ;
        RECT 42.995 32.910 43.145 33.080 ;
        RECT 43.715 32.910 43.865 33.080 ;
        RECT 45.895 32.910 46.045 33.080 ;
        RECT 46.615 32.910 46.765 33.080 ;
        RECT 48.795 32.910 48.945 33.080 ;
        RECT 49.515 32.910 49.665 33.080 ;
        RECT 51.695 32.910 51.845 33.080 ;
        RECT 52.415 32.910 52.565 33.080 ;
        RECT 54.595 32.910 54.745 33.080 ;
        RECT 55.315 32.910 55.465 33.080 ;
        RECT 57.495 32.910 57.645 33.080 ;
        RECT 58.215 32.910 58.365 33.080 ;
        RECT 60.395 32.910 60.545 33.080 ;
        RECT 61.115 32.910 61.265 33.080 ;
        RECT 63.295 32.910 63.445 33.080 ;
        RECT 64.015 32.910 64.165 33.080 ;
        RECT 66.195 32.910 66.345 33.080 ;
        RECT 66.915 32.910 67.065 33.080 ;
        RECT 69.095 32.910 69.245 33.080 ;
        RECT 69.815 32.910 69.965 33.080 ;
        RECT 71.995 32.910 72.145 33.080 ;
        RECT 72.715 32.910 72.865 33.080 ;
        RECT 74.895 32.910 75.045 33.080 ;
        RECT 75.615 32.910 75.765 33.080 ;
        RECT 77.795 32.910 77.945 33.080 ;
        RECT 78.515 32.910 78.665 33.080 ;
        RECT 80.695 32.910 80.845 33.080 ;
        RECT 81.415 32.910 81.565 33.080 ;
        RECT 83.595 32.910 83.745 33.080 ;
        RECT 84.315 32.910 84.465 33.080 ;
        RECT 86.495 32.910 86.645 33.080 ;
        RECT 87.215 32.910 87.365 33.080 ;
        RECT 89.395 32.910 89.545 33.080 ;
        RECT 90.115 32.910 90.265 33.080 ;
        RECT 92.295 32.910 92.445 33.080 ;
      LAYER met1 ;
        RECT 0.000 32.910 92.445 33.080 ;
    END
  END RWL_7
  PIN RWL_8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 31.560 0.365 31.730 ;
        RECT 2.395 31.560 2.545 31.730 ;
        RECT 3.115 31.560 3.265 31.730 ;
        RECT 5.295 31.560 5.445 31.730 ;
        RECT 6.015 31.560 6.165 31.730 ;
        RECT 8.195 31.560 8.345 31.730 ;
        RECT 8.915 31.560 9.065 31.730 ;
        RECT 11.095 31.560 11.245 31.730 ;
        RECT 11.815 31.560 11.965 31.730 ;
        RECT 13.995 31.560 14.145 31.730 ;
        RECT 14.715 31.560 14.865 31.730 ;
        RECT 16.895 31.560 17.045 31.730 ;
        RECT 17.615 31.560 17.765 31.730 ;
        RECT 19.795 31.560 19.945 31.730 ;
        RECT 20.515 31.560 20.665 31.730 ;
        RECT 22.695 31.560 22.845 31.730 ;
        RECT 23.415 31.560 23.565 31.730 ;
        RECT 25.595 31.560 25.745 31.730 ;
        RECT 26.315 31.560 26.465 31.730 ;
        RECT 28.495 31.560 28.645 31.730 ;
        RECT 29.215 31.560 29.365 31.730 ;
        RECT 31.395 31.560 31.545 31.730 ;
        RECT 32.115 31.560 32.265 31.730 ;
        RECT 34.295 31.560 34.445 31.730 ;
        RECT 35.015 31.560 35.165 31.730 ;
        RECT 37.195 31.560 37.345 31.730 ;
        RECT 37.915 31.560 38.065 31.730 ;
        RECT 40.095 31.560 40.245 31.730 ;
        RECT 40.815 31.560 40.965 31.730 ;
        RECT 42.995 31.560 43.145 31.730 ;
        RECT 43.715 31.560 43.865 31.730 ;
        RECT 45.895 31.560 46.045 31.730 ;
        RECT 46.615 31.560 46.765 31.730 ;
        RECT 48.795 31.560 48.945 31.730 ;
        RECT 49.515 31.560 49.665 31.730 ;
        RECT 51.695 31.560 51.845 31.730 ;
        RECT 52.415 31.560 52.565 31.730 ;
        RECT 54.595 31.560 54.745 31.730 ;
        RECT 55.315 31.560 55.465 31.730 ;
        RECT 57.495 31.560 57.645 31.730 ;
        RECT 58.215 31.560 58.365 31.730 ;
        RECT 60.395 31.560 60.545 31.730 ;
        RECT 61.115 31.560 61.265 31.730 ;
        RECT 63.295 31.560 63.445 31.730 ;
        RECT 64.015 31.560 64.165 31.730 ;
        RECT 66.195 31.560 66.345 31.730 ;
        RECT 66.915 31.560 67.065 31.730 ;
        RECT 69.095 31.560 69.245 31.730 ;
        RECT 69.815 31.560 69.965 31.730 ;
        RECT 71.995 31.560 72.145 31.730 ;
        RECT 72.715 31.560 72.865 31.730 ;
        RECT 74.895 31.560 75.045 31.730 ;
        RECT 75.615 31.560 75.765 31.730 ;
        RECT 77.795 31.560 77.945 31.730 ;
        RECT 78.515 31.560 78.665 31.730 ;
        RECT 80.695 31.560 80.845 31.730 ;
        RECT 81.415 31.560 81.565 31.730 ;
        RECT 83.595 31.560 83.745 31.730 ;
        RECT 84.315 31.560 84.465 31.730 ;
        RECT 86.495 31.560 86.645 31.730 ;
        RECT 87.215 31.560 87.365 31.730 ;
        RECT 89.395 31.560 89.545 31.730 ;
        RECT 90.115 31.560 90.265 31.730 ;
        RECT 92.295 31.560 92.445 31.730 ;
      LAYER met1 ;
        RECT 0.000 31.560 92.445 31.730 ;
    END
  END RWL_8
  PIN RWL_9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 30.210 0.365 30.380 ;
        RECT 2.395 30.210 2.545 30.380 ;
        RECT 3.115 30.210 3.265 30.380 ;
        RECT 5.295 30.210 5.445 30.380 ;
        RECT 6.015 30.210 6.165 30.380 ;
        RECT 8.195 30.210 8.345 30.380 ;
        RECT 8.915 30.210 9.065 30.380 ;
        RECT 11.095 30.210 11.245 30.380 ;
        RECT 11.815 30.210 11.965 30.380 ;
        RECT 13.995 30.210 14.145 30.380 ;
        RECT 14.715 30.210 14.865 30.380 ;
        RECT 16.895 30.210 17.045 30.380 ;
        RECT 17.615 30.210 17.765 30.380 ;
        RECT 19.795 30.210 19.945 30.380 ;
        RECT 20.515 30.210 20.665 30.380 ;
        RECT 22.695 30.210 22.845 30.380 ;
        RECT 23.415 30.210 23.565 30.380 ;
        RECT 25.595 30.210 25.745 30.380 ;
        RECT 26.315 30.210 26.465 30.380 ;
        RECT 28.495 30.210 28.645 30.380 ;
        RECT 29.215 30.210 29.365 30.380 ;
        RECT 31.395 30.210 31.545 30.380 ;
        RECT 32.115 30.210 32.265 30.380 ;
        RECT 34.295 30.210 34.445 30.380 ;
        RECT 35.015 30.210 35.165 30.380 ;
        RECT 37.195 30.210 37.345 30.380 ;
        RECT 37.915 30.210 38.065 30.380 ;
        RECT 40.095 30.210 40.245 30.380 ;
        RECT 40.815 30.210 40.965 30.380 ;
        RECT 42.995 30.210 43.145 30.380 ;
        RECT 43.715 30.210 43.865 30.380 ;
        RECT 45.895 30.210 46.045 30.380 ;
        RECT 46.615 30.210 46.765 30.380 ;
        RECT 48.795 30.210 48.945 30.380 ;
        RECT 49.515 30.210 49.665 30.380 ;
        RECT 51.695 30.210 51.845 30.380 ;
        RECT 52.415 30.210 52.565 30.380 ;
        RECT 54.595 30.210 54.745 30.380 ;
        RECT 55.315 30.210 55.465 30.380 ;
        RECT 57.495 30.210 57.645 30.380 ;
        RECT 58.215 30.210 58.365 30.380 ;
        RECT 60.395 30.210 60.545 30.380 ;
        RECT 61.115 30.210 61.265 30.380 ;
        RECT 63.295 30.210 63.445 30.380 ;
        RECT 64.015 30.210 64.165 30.380 ;
        RECT 66.195 30.210 66.345 30.380 ;
        RECT 66.915 30.210 67.065 30.380 ;
        RECT 69.095 30.210 69.245 30.380 ;
        RECT 69.815 30.210 69.965 30.380 ;
        RECT 71.995 30.210 72.145 30.380 ;
        RECT 72.715 30.210 72.865 30.380 ;
        RECT 74.895 30.210 75.045 30.380 ;
        RECT 75.615 30.210 75.765 30.380 ;
        RECT 77.795 30.210 77.945 30.380 ;
        RECT 78.515 30.210 78.665 30.380 ;
        RECT 80.695 30.210 80.845 30.380 ;
        RECT 81.415 30.210 81.565 30.380 ;
        RECT 83.595 30.210 83.745 30.380 ;
        RECT 84.315 30.210 84.465 30.380 ;
        RECT 86.495 30.210 86.645 30.380 ;
        RECT 87.215 30.210 87.365 30.380 ;
        RECT 89.395 30.210 89.545 30.380 ;
        RECT 90.115 30.210 90.265 30.380 ;
        RECT 92.295 30.210 92.445 30.380 ;
      LAYER met1 ;
        RECT 0.000 30.210 92.445 30.380 ;
    END
  END RWL_9
  PIN RWL_10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 28.860 0.365 29.030 ;
        RECT 2.395 28.860 2.545 29.030 ;
        RECT 3.115 28.860 3.265 29.030 ;
        RECT 5.295 28.860 5.445 29.030 ;
        RECT 6.015 28.860 6.165 29.030 ;
        RECT 8.195 28.860 8.345 29.030 ;
        RECT 8.915 28.860 9.065 29.030 ;
        RECT 11.095 28.860 11.245 29.030 ;
        RECT 11.815 28.860 11.965 29.030 ;
        RECT 13.995 28.860 14.145 29.030 ;
        RECT 14.715 28.860 14.865 29.030 ;
        RECT 16.895 28.860 17.045 29.030 ;
        RECT 17.615 28.860 17.765 29.030 ;
        RECT 19.795 28.860 19.945 29.030 ;
        RECT 20.515 28.860 20.665 29.030 ;
        RECT 22.695 28.860 22.845 29.030 ;
        RECT 23.415 28.860 23.565 29.030 ;
        RECT 25.595 28.860 25.745 29.030 ;
        RECT 26.315 28.860 26.465 29.030 ;
        RECT 28.495 28.860 28.645 29.030 ;
        RECT 29.215 28.860 29.365 29.030 ;
        RECT 31.395 28.860 31.545 29.030 ;
        RECT 32.115 28.860 32.265 29.030 ;
        RECT 34.295 28.860 34.445 29.030 ;
        RECT 35.015 28.860 35.165 29.030 ;
        RECT 37.195 28.860 37.345 29.030 ;
        RECT 37.915 28.860 38.065 29.030 ;
        RECT 40.095 28.860 40.245 29.030 ;
        RECT 40.815 28.860 40.965 29.030 ;
        RECT 42.995 28.860 43.145 29.030 ;
        RECT 43.715 28.860 43.865 29.030 ;
        RECT 45.895 28.860 46.045 29.030 ;
        RECT 46.615 28.860 46.765 29.030 ;
        RECT 48.795 28.860 48.945 29.030 ;
        RECT 49.515 28.860 49.665 29.030 ;
        RECT 51.695 28.860 51.845 29.030 ;
        RECT 52.415 28.860 52.565 29.030 ;
        RECT 54.595 28.860 54.745 29.030 ;
        RECT 55.315 28.860 55.465 29.030 ;
        RECT 57.495 28.860 57.645 29.030 ;
        RECT 58.215 28.860 58.365 29.030 ;
        RECT 60.395 28.860 60.545 29.030 ;
        RECT 61.115 28.860 61.265 29.030 ;
        RECT 63.295 28.860 63.445 29.030 ;
        RECT 64.015 28.860 64.165 29.030 ;
        RECT 66.195 28.860 66.345 29.030 ;
        RECT 66.915 28.860 67.065 29.030 ;
        RECT 69.095 28.860 69.245 29.030 ;
        RECT 69.815 28.860 69.965 29.030 ;
        RECT 71.995 28.860 72.145 29.030 ;
        RECT 72.715 28.860 72.865 29.030 ;
        RECT 74.895 28.860 75.045 29.030 ;
        RECT 75.615 28.860 75.765 29.030 ;
        RECT 77.795 28.860 77.945 29.030 ;
        RECT 78.515 28.860 78.665 29.030 ;
        RECT 80.695 28.860 80.845 29.030 ;
        RECT 81.415 28.860 81.565 29.030 ;
        RECT 83.595 28.860 83.745 29.030 ;
        RECT 84.315 28.860 84.465 29.030 ;
        RECT 86.495 28.860 86.645 29.030 ;
        RECT 87.215 28.860 87.365 29.030 ;
        RECT 89.395 28.860 89.545 29.030 ;
        RECT 90.115 28.860 90.265 29.030 ;
        RECT 92.295 28.860 92.445 29.030 ;
      LAYER met1 ;
        RECT 0.000 28.860 92.445 29.030 ;
    END
  END RWL_10
  PIN RWL_11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 27.510 0.365 27.680 ;
        RECT 2.395 27.510 2.545 27.680 ;
        RECT 3.115 27.510 3.265 27.680 ;
        RECT 5.295 27.510 5.445 27.680 ;
        RECT 6.015 27.510 6.165 27.680 ;
        RECT 8.195 27.510 8.345 27.680 ;
        RECT 8.915 27.510 9.065 27.680 ;
        RECT 11.095 27.510 11.245 27.680 ;
        RECT 11.815 27.510 11.965 27.680 ;
        RECT 13.995 27.510 14.145 27.680 ;
        RECT 14.715 27.510 14.865 27.680 ;
        RECT 16.895 27.510 17.045 27.680 ;
        RECT 17.615 27.510 17.765 27.680 ;
        RECT 19.795 27.510 19.945 27.680 ;
        RECT 20.515 27.510 20.665 27.680 ;
        RECT 22.695 27.510 22.845 27.680 ;
        RECT 23.415 27.510 23.565 27.680 ;
        RECT 25.595 27.510 25.745 27.680 ;
        RECT 26.315 27.510 26.465 27.680 ;
        RECT 28.495 27.510 28.645 27.680 ;
        RECT 29.215 27.510 29.365 27.680 ;
        RECT 31.395 27.510 31.545 27.680 ;
        RECT 32.115 27.510 32.265 27.680 ;
        RECT 34.295 27.510 34.445 27.680 ;
        RECT 35.015 27.510 35.165 27.680 ;
        RECT 37.195 27.510 37.345 27.680 ;
        RECT 37.915 27.510 38.065 27.680 ;
        RECT 40.095 27.510 40.245 27.680 ;
        RECT 40.815 27.510 40.965 27.680 ;
        RECT 42.995 27.510 43.145 27.680 ;
        RECT 43.715 27.510 43.865 27.680 ;
        RECT 45.895 27.510 46.045 27.680 ;
        RECT 46.615 27.510 46.765 27.680 ;
        RECT 48.795 27.510 48.945 27.680 ;
        RECT 49.515 27.510 49.665 27.680 ;
        RECT 51.695 27.510 51.845 27.680 ;
        RECT 52.415 27.510 52.565 27.680 ;
        RECT 54.595 27.510 54.745 27.680 ;
        RECT 55.315 27.510 55.465 27.680 ;
        RECT 57.495 27.510 57.645 27.680 ;
        RECT 58.215 27.510 58.365 27.680 ;
        RECT 60.395 27.510 60.545 27.680 ;
        RECT 61.115 27.510 61.265 27.680 ;
        RECT 63.295 27.510 63.445 27.680 ;
        RECT 64.015 27.510 64.165 27.680 ;
        RECT 66.195 27.510 66.345 27.680 ;
        RECT 66.915 27.510 67.065 27.680 ;
        RECT 69.095 27.510 69.245 27.680 ;
        RECT 69.815 27.510 69.965 27.680 ;
        RECT 71.995 27.510 72.145 27.680 ;
        RECT 72.715 27.510 72.865 27.680 ;
        RECT 74.895 27.510 75.045 27.680 ;
        RECT 75.615 27.510 75.765 27.680 ;
        RECT 77.795 27.510 77.945 27.680 ;
        RECT 78.515 27.510 78.665 27.680 ;
        RECT 80.695 27.510 80.845 27.680 ;
        RECT 81.415 27.510 81.565 27.680 ;
        RECT 83.595 27.510 83.745 27.680 ;
        RECT 84.315 27.510 84.465 27.680 ;
        RECT 86.495 27.510 86.645 27.680 ;
        RECT 87.215 27.510 87.365 27.680 ;
        RECT 89.395 27.510 89.545 27.680 ;
        RECT 90.115 27.510 90.265 27.680 ;
        RECT 92.295 27.510 92.445 27.680 ;
      LAYER met1 ;
        RECT 0.000 27.510 92.445 27.680 ;
    END
  END RWL_11
  PIN RWL_12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 26.160 0.365 26.330 ;
        RECT 2.395 26.160 2.545 26.330 ;
        RECT 3.115 26.160 3.265 26.330 ;
        RECT 5.295 26.160 5.445 26.330 ;
        RECT 6.015 26.160 6.165 26.330 ;
        RECT 8.195 26.160 8.345 26.330 ;
        RECT 8.915 26.160 9.065 26.330 ;
        RECT 11.095 26.160 11.245 26.330 ;
        RECT 11.815 26.160 11.965 26.330 ;
        RECT 13.995 26.160 14.145 26.330 ;
        RECT 14.715 26.160 14.865 26.330 ;
        RECT 16.895 26.160 17.045 26.330 ;
        RECT 17.615 26.160 17.765 26.330 ;
        RECT 19.795 26.160 19.945 26.330 ;
        RECT 20.515 26.160 20.665 26.330 ;
        RECT 22.695 26.160 22.845 26.330 ;
        RECT 23.415 26.160 23.565 26.330 ;
        RECT 25.595 26.160 25.745 26.330 ;
        RECT 26.315 26.160 26.465 26.330 ;
        RECT 28.495 26.160 28.645 26.330 ;
        RECT 29.215 26.160 29.365 26.330 ;
        RECT 31.395 26.160 31.545 26.330 ;
        RECT 32.115 26.160 32.265 26.330 ;
        RECT 34.295 26.160 34.445 26.330 ;
        RECT 35.015 26.160 35.165 26.330 ;
        RECT 37.195 26.160 37.345 26.330 ;
        RECT 37.915 26.160 38.065 26.330 ;
        RECT 40.095 26.160 40.245 26.330 ;
        RECT 40.815 26.160 40.965 26.330 ;
        RECT 42.995 26.160 43.145 26.330 ;
        RECT 43.715 26.160 43.865 26.330 ;
        RECT 45.895 26.160 46.045 26.330 ;
        RECT 46.615 26.160 46.765 26.330 ;
        RECT 48.795 26.160 48.945 26.330 ;
        RECT 49.515 26.160 49.665 26.330 ;
        RECT 51.695 26.160 51.845 26.330 ;
        RECT 52.415 26.160 52.565 26.330 ;
        RECT 54.595 26.160 54.745 26.330 ;
        RECT 55.315 26.160 55.465 26.330 ;
        RECT 57.495 26.160 57.645 26.330 ;
        RECT 58.215 26.160 58.365 26.330 ;
        RECT 60.395 26.160 60.545 26.330 ;
        RECT 61.115 26.160 61.265 26.330 ;
        RECT 63.295 26.160 63.445 26.330 ;
        RECT 64.015 26.160 64.165 26.330 ;
        RECT 66.195 26.160 66.345 26.330 ;
        RECT 66.915 26.160 67.065 26.330 ;
        RECT 69.095 26.160 69.245 26.330 ;
        RECT 69.815 26.160 69.965 26.330 ;
        RECT 71.995 26.160 72.145 26.330 ;
        RECT 72.715 26.160 72.865 26.330 ;
        RECT 74.895 26.160 75.045 26.330 ;
        RECT 75.615 26.160 75.765 26.330 ;
        RECT 77.795 26.160 77.945 26.330 ;
        RECT 78.515 26.160 78.665 26.330 ;
        RECT 80.695 26.160 80.845 26.330 ;
        RECT 81.415 26.160 81.565 26.330 ;
        RECT 83.595 26.160 83.745 26.330 ;
        RECT 84.315 26.160 84.465 26.330 ;
        RECT 86.495 26.160 86.645 26.330 ;
        RECT 87.215 26.160 87.365 26.330 ;
        RECT 89.395 26.160 89.545 26.330 ;
        RECT 90.115 26.160 90.265 26.330 ;
        RECT 92.295 26.160 92.445 26.330 ;
      LAYER met1 ;
        RECT 0.000 26.160 92.445 26.330 ;
    END
  END RWL_12
  PIN RWL_13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 24.810 0.365 24.980 ;
        RECT 2.395 24.810 2.545 24.980 ;
        RECT 3.115 24.810 3.265 24.980 ;
        RECT 5.295 24.810 5.445 24.980 ;
        RECT 6.015 24.810 6.165 24.980 ;
        RECT 8.195 24.810 8.345 24.980 ;
        RECT 8.915 24.810 9.065 24.980 ;
        RECT 11.095 24.810 11.245 24.980 ;
        RECT 11.815 24.810 11.965 24.980 ;
        RECT 13.995 24.810 14.145 24.980 ;
        RECT 14.715 24.810 14.865 24.980 ;
        RECT 16.895 24.810 17.045 24.980 ;
        RECT 17.615 24.810 17.765 24.980 ;
        RECT 19.795 24.810 19.945 24.980 ;
        RECT 20.515 24.810 20.665 24.980 ;
        RECT 22.695 24.810 22.845 24.980 ;
        RECT 23.415 24.810 23.565 24.980 ;
        RECT 25.595 24.810 25.745 24.980 ;
        RECT 26.315 24.810 26.465 24.980 ;
        RECT 28.495 24.810 28.645 24.980 ;
        RECT 29.215 24.810 29.365 24.980 ;
        RECT 31.395 24.810 31.545 24.980 ;
        RECT 32.115 24.810 32.265 24.980 ;
        RECT 34.295 24.810 34.445 24.980 ;
        RECT 35.015 24.810 35.165 24.980 ;
        RECT 37.195 24.810 37.345 24.980 ;
        RECT 37.915 24.810 38.065 24.980 ;
        RECT 40.095 24.810 40.245 24.980 ;
        RECT 40.815 24.810 40.965 24.980 ;
        RECT 42.995 24.810 43.145 24.980 ;
        RECT 43.715 24.810 43.865 24.980 ;
        RECT 45.895 24.810 46.045 24.980 ;
        RECT 46.615 24.810 46.765 24.980 ;
        RECT 48.795 24.810 48.945 24.980 ;
        RECT 49.515 24.810 49.665 24.980 ;
        RECT 51.695 24.810 51.845 24.980 ;
        RECT 52.415 24.810 52.565 24.980 ;
        RECT 54.595 24.810 54.745 24.980 ;
        RECT 55.315 24.810 55.465 24.980 ;
        RECT 57.495 24.810 57.645 24.980 ;
        RECT 58.215 24.810 58.365 24.980 ;
        RECT 60.395 24.810 60.545 24.980 ;
        RECT 61.115 24.810 61.265 24.980 ;
        RECT 63.295 24.810 63.445 24.980 ;
        RECT 64.015 24.810 64.165 24.980 ;
        RECT 66.195 24.810 66.345 24.980 ;
        RECT 66.915 24.810 67.065 24.980 ;
        RECT 69.095 24.810 69.245 24.980 ;
        RECT 69.815 24.810 69.965 24.980 ;
        RECT 71.995 24.810 72.145 24.980 ;
        RECT 72.715 24.810 72.865 24.980 ;
        RECT 74.895 24.810 75.045 24.980 ;
        RECT 75.615 24.810 75.765 24.980 ;
        RECT 77.795 24.810 77.945 24.980 ;
        RECT 78.515 24.810 78.665 24.980 ;
        RECT 80.695 24.810 80.845 24.980 ;
        RECT 81.415 24.810 81.565 24.980 ;
        RECT 83.595 24.810 83.745 24.980 ;
        RECT 84.315 24.810 84.465 24.980 ;
        RECT 86.495 24.810 86.645 24.980 ;
        RECT 87.215 24.810 87.365 24.980 ;
        RECT 89.395 24.810 89.545 24.980 ;
        RECT 90.115 24.810 90.265 24.980 ;
        RECT 92.295 24.810 92.445 24.980 ;
      LAYER met1 ;
        RECT 0.000 24.810 92.445 24.980 ;
    END
  END RWL_13
  PIN RWL_14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 23.460 0.365 23.630 ;
        RECT 2.395 23.460 2.545 23.630 ;
        RECT 3.115 23.460 3.265 23.630 ;
        RECT 5.295 23.460 5.445 23.630 ;
        RECT 6.015 23.460 6.165 23.630 ;
        RECT 8.195 23.460 8.345 23.630 ;
        RECT 8.915 23.460 9.065 23.630 ;
        RECT 11.095 23.460 11.245 23.630 ;
        RECT 11.815 23.460 11.965 23.630 ;
        RECT 13.995 23.460 14.145 23.630 ;
        RECT 14.715 23.460 14.865 23.630 ;
        RECT 16.895 23.460 17.045 23.630 ;
        RECT 17.615 23.460 17.765 23.630 ;
        RECT 19.795 23.460 19.945 23.630 ;
        RECT 20.515 23.460 20.665 23.630 ;
        RECT 22.695 23.460 22.845 23.630 ;
        RECT 23.415 23.460 23.565 23.630 ;
        RECT 25.595 23.460 25.745 23.630 ;
        RECT 26.315 23.460 26.465 23.630 ;
        RECT 28.495 23.460 28.645 23.630 ;
        RECT 29.215 23.460 29.365 23.630 ;
        RECT 31.395 23.460 31.545 23.630 ;
        RECT 32.115 23.460 32.265 23.630 ;
        RECT 34.295 23.460 34.445 23.630 ;
        RECT 35.015 23.460 35.165 23.630 ;
        RECT 37.195 23.460 37.345 23.630 ;
        RECT 37.915 23.460 38.065 23.630 ;
        RECT 40.095 23.460 40.245 23.630 ;
        RECT 40.815 23.460 40.965 23.630 ;
        RECT 42.995 23.460 43.145 23.630 ;
        RECT 43.715 23.460 43.865 23.630 ;
        RECT 45.895 23.460 46.045 23.630 ;
        RECT 46.615 23.460 46.765 23.630 ;
        RECT 48.795 23.460 48.945 23.630 ;
        RECT 49.515 23.460 49.665 23.630 ;
        RECT 51.695 23.460 51.845 23.630 ;
        RECT 52.415 23.460 52.565 23.630 ;
        RECT 54.595 23.460 54.745 23.630 ;
        RECT 55.315 23.460 55.465 23.630 ;
        RECT 57.495 23.460 57.645 23.630 ;
        RECT 58.215 23.460 58.365 23.630 ;
        RECT 60.395 23.460 60.545 23.630 ;
        RECT 61.115 23.460 61.265 23.630 ;
        RECT 63.295 23.460 63.445 23.630 ;
        RECT 64.015 23.460 64.165 23.630 ;
        RECT 66.195 23.460 66.345 23.630 ;
        RECT 66.915 23.460 67.065 23.630 ;
        RECT 69.095 23.460 69.245 23.630 ;
        RECT 69.815 23.460 69.965 23.630 ;
        RECT 71.995 23.460 72.145 23.630 ;
        RECT 72.715 23.460 72.865 23.630 ;
        RECT 74.895 23.460 75.045 23.630 ;
        RECT 75.615 23.460 75.765 23.630 ;
        RECT 77.795 23.460 77.945 23.630 ;
        RECT 78.515 23.460 78.665 23.630 ;
        RECT 80.695 23.460 80.845 23.630 ;
        RECT 81.415 23.460 81.565 23.630 ;
        RECT 83.595 23.460 83.745 23.630 ;
        RECT 84.315 23.460 84.465 23.630 ;
        RECT 86.495 23.460 86.645 23.630 ;
        RECT 87.215 23.460 87.365 23.630 ;
        RECT 89.395 23.460 89.545 23.630 ;
        RECT 90.115 23.460 90.265 23.630 ;
        RECT 92.295 23.460 92.445 23.630 ;
      LAYER met1 ;
        RECT 0.000 23.460 92.445 23.630 ;
    END
  END RWL_14
  PIN RWL_15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 22.110 0.365 22.280 ;
        RECT 2.395 22.110 2.545 22.280 ;
        RECT 3.115 22.110 3.265 22.280 ;
        RECT 5.295 22.110 5.445 22.280 ;
        RECT 6.015 22.110 6.165 22.280 ;
        RECT 8.195 22.110 8.345 22.280 ;
        RECT 8.915 22.110 9.065 22.280 ;
        RECT 11.095 22.110 11.245 22.280 ;
        RECT 11.815 22.110 11.965 22.280 ;
        RECT 13.995 22.110 14.145 22.280 ;
        RECT 14.715 22.110 14.865 22.280 ;
        RECT 16.895 22.110 17.045 22.280 ;
        RECT 17.615 22.110 17.765 22.280 ;
        RECT 19.795 22.110 19.945 22.280 ;
        RECT 20.515 22.110 20.665 22.280 ;
        RECT 22.695 22.110 22.845 22.280 ;
        RECT 23.415 22.110 23.565 22.280 ;
        RECT 25.595 22.110 25.745 22.280 ;
        RECT 26.315 22.110 26.465 22.280 ;
        RECT 28.495 22.110 28.645 22.280 ;
        RECT 29.215 22.110 29.365 22.280 ;
        RECT 31.395 22.110 31.545 22.280 ;
        RECT 32.115 22.110 32.265 22.280 ;
        RECT 34.295 22.110 34.445 22.280 ;
        RECT 35.015 22.110 35.165 22.280 ;
        RECT 37.195 22.110 37.345 22.280 ;
        RECT 37.915 22.110 38.065 22.280 ;
        RECT 40.095 22.110 40.245 22.280 ;
        RECT 40.815 22.110 40.965 22.280 ;
        RECT 42.995 22.110 43.145 22.280 ;
        RECT 43.715 22.110 43.865 22.280 ;
        RECT 45.895 22.110 46.045 22.280 ;
        RECT 46.615 22.110 46.765 22.280 ;
        RECT 48.795 22.110 48.945 22.280 ;
        RECT 49.515 22.110 49.665 22.280 ;
        RECT 51.695 22.110 51.845 22.280 ;
        RECT 52.415 22.110 52.565 22.280 ;
        RECT 54.595 22.110 54.745 22.280 ;
        RECT 55.315 22.110 55.465 22.280 ;
        RECT 57.495 22.110 57.645 22.280 ;
        RECT 58.215 22.110 58.365 22.280 ;
        RECT 60.395 22.110 60.545 22.280 ;
        RECT 61.115 22.110 61.265 22.280 ;
        RECT 63.295 22.110 63.445 22.280 ;
        RECT 64.015 22.110 64.165 22.280 ;
        RECT 66.195 22.110 66.345 22.280 ;
        RECT 66.915 22.110 67.065 22.280 ;
        RECT 69.095 22.110 69.245 22.280 ;
        RECT 69.815 22.110 69.965 22.280 ;
        RECT 71.995 22.110 72.145 22.280 ;
        RECT 72.715 22.110 72.865 22.280 ;
        RECT 74.895 22.110 75.045 22.280 ;
        RECT 75.615 22.110 75.765 22.280 ;
        RECT 77.795 22.110 77.945 22.280 ;
        RECT 78.515 22.110 78.665 22.280 ;
        RECT 80.695 22.110 80.845 22.280 ;
        RECT 81.415 22.110 81.565 22.280 ;
        RECT 83.595 22.110 83.745 22.280 ;
        RECT 84.315 22.110 84.465 22.280 ;
        RECT 86.495 22.110 86.645 22.280 ;
        RECT 87.215 22.110 87.365 22.280 ;
        RECT 89.395 22.110 89.545 22.280 ;
        RECT 90.115 22.110 90.265 22.280 ;
        RECT 92.295 22.110 92.445 22.280 ;
      LAYER met1 ;
        RECT 0.000 22.110 92.445 22.280 ;
    END
  END RWL_15
  PIN RWL_16
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 20.760 0.365 20.930 ;
        RECT 2.395 20.760 2.545 20.930 ;
        RECT 3.115 20.760 3.265 20.930 ;
        RECT 5.295 20.760 5.445 20.930 ;
        RECT 6.015 20.760 6.165 20.930 ;
        RECT 8.195 20.760 8.345 20.930 ;
        RECT 8.915 20.760 9.065 20.930 ;
        RECT 11.095 20.760 11.245 20.930 ;
        RECT 11.815 20.760 11.965 20.930 ;
        RECT 13.995 20.760 14.145 20.930 ;
        RECT 14.715 20.760 14.865 20.930 ;
        RECT 16.895 20.760 17.045 20.930 ;
        RECT 17.615 20.760 17.765 20.930 ;
        RECT 19.795 20.760 19.945 20.930 ;
        RECT 20.515 20.760 20.665 20.930 ;
        RECT 22.695 20.760 22.845 20.930 ;
        RECT 23.415 20.760 23.565 20.930 ;
        RECT 25.595 20.760 25.745 20.930 ;
        RECT 26.315 20.760 26.465 20.930 ;
        RECT 28.495 20.760 28.645 20.930 ;
        RECT 29.215 20.760 29.365 20.930 ;
        RECT 31.395 20.760 31.545 20.930 ;
        RECT 32.115 20.760 32.265 20.930 ;
        RECT 34.295 20.760 34.445 20.930 ;
        RECT 35.015 20.760 35.165 20.930 ;
        RECT 37.195 20.760 37.345 20.930 ;
        RECT 37.915 20.760 38.065 20.930 ;
        RECT 40.095 20.760 40.245 20.930 ;
        RECT 40.815 20.760 40.965 20.930 ;
        RECT 42.995 20.760 43.145 20.930 ;
        RECT 43.715 20.760 43.865 20.930 ;
        RECT 45.895 20.760 46.045 20.930 ;
        RECT 46.615 20.760 46.765 20.930 ;
        RECT 48.795 20.760 48.945 20.930 ;
        RECT 49.515 20.760 49.665 20.930 ;
        RECT 51.695 20.760 51.845 20.930 ;
        RECT 52.415 20.760 52.565 20.930 ;
        RECT 54.595 20.760 54.745 20.930 ;
        RECT 55.315 20.760 55.465 20.930 ;
        RECT 57.495 20.760 57.645 20.930 ;
        RECT 58.215 20.760 58.365 20.930 ;
        RECT 60.395 20.760 60.545 20.930 ;
        RECT 61.115 20.760 61.265 20.930 ;
        RECT 63.295 20.760 63.445 20.930 ;
        RECT 64.015 20.760 64.165 20.930 ;
        RECT 66.195 20.760 66.345 20.930 ;
        RECT 66.915 20.760 67.065 20.930 ;
        RECT 69.095 20.760 69.245 20.930 ;
        RECT 69.815 20.760 69.965 20.930 ;
        RECT 71.995 20.760 72.145 20.930 ;
        RECT 72.715 20.760 72.865 20.930 ;
        RECT 74.895 20.760 75.045 20.930 ;
        RECT 75.615 20.760 75.765 20.930 ;
        RECT 77.795 20.760 77.945 20.930 ;
        RECT 78.515 20.760 78.665 20.930 ;
        RECT 80.695 20.760 80.845 20.930 ;
        RECT 81.415 20.760 81.565 20.930 ;
        RECT 83.595 20.760 83.745 20.930 ;
        RECT 84.315 20.760 84.465 20.930 ;
        RECT 86.495 20.760 86.645 20.930 ;
        RECT 87.215 20.760 87.365 20.930 ;
        RECT 89.395 20.760 89.545 20.930 ;
        RECT 90.115 20.760 90.265 20.930 ;
        RECT 92.295 20.760 92.445 20.930 ;
      LAYER met1 ;
        RECT 0.000 20.760 92.445 20.930 ;
    END
  END RWL_16
  PIN RWL_17
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 19.410 0.365 19.580 ;
        RECT 2.395 19.410 2.545 19.580 ;
        RECT 3.115 19.410 3.265 19.580 ;
        RECT 5.295 19.410 5.445 19.580 ;
        RECT 6.015 19.410 6.165 19.580 ;
        RECT 8.195 19.410 8.345 19.580 ;
        RECT 8.915 19.410 9.065 19.580 ;
        RECT 11.095 19.410 11.245 19.580 ;
        RECT 11.815 19.410 11.965 19.580 ;
        RECT 13.995 19.410 14.145 19.580 ;
        RECT 14.715 19.410 14.865 19.580 ;
        RECT 16.895 19.410 17.045 19.580 ;
        RECT 17.615 19.410 17.765 19.580 ;
        RECT 19.795 19.410 19.945 19.580 ;
        RECT 20.515 19.410 20.665 19.580 ;
        RECT 22.695 19.410 22.845 19.580 ;
        RECT 23.415 19.410 23.565 19.580 ;
        RECT 25.595 19.410 25.745 19.580 ;
        RECT 26.315 19.410 26.465 19.580 ;
        RECT 28.495 19.410 28.645 19.580 ;
        RECT 29.215 19.410 29.365 19.580 ;
        RECT 31.395 19.410 31.545 19.580 ;
        RECT 32.115 19.410 32.265 19.580 ;
        RECT 34.295 19.410 34.445 19.580 ;
        RECT 35.015 19.410 35.165 19.580 ;
        RECT 37.195 19.410 37.345 19.580 ;
        RECT 37.915 19.410 38.065 19.580 ;
        RECT 40.095 19.410 40.245 19.580 ;
        RECT 40.815 19.410 40.965 19.580 ;
        RECT 42.995 19.410 43.145 19.580 ;
        RECT 43.715 19.410 43.865 19.580 ;
        RECT 45.895 19.410 46.045 19.580 ;
        RECT 46.615 19.410 46.765 19.580 ;
        RECT 48.795 19.410 48.945 19.580 ;
        RECT 49.515 19.410 49.665 19.580 ;
        RECT 51.695 19.410 51.845 19.580 ;
        RECT 52.415 19.410 52.565 19.580 ;
        RECT 54.595 19.410 54.745 19.580 ;
        RECT 55.315 19.410 55.465 19.580 ;
        RECT 57.495 19.410 57.645 19.580 ;
        RECT 58.215 19.410 58.365 19.580 ;
        RECT 60.395 19.410 60.545 19.580 ;
        RECT 61.115 19.410 61.265 19.580 ;
        RECT 63.295 19.410 63.445 19.580 ;
        RECT 64.015 19.410 64.165 19.580 ;
        RECT 66.195 19.410 66.345 19.580 ;
        RECT 66.915 19.410 67.065 19.580 ;
        RECT 69.095 19.410 69.245 19.580 ;
        RECT 69.815 19.410 69.965 19.580 ;
        RECT 71.995 19.410 72.145 19.580 ;
        RECT 72.715 19.410 72.865 19.580 ;
        RECT 74.895 19.410 75.045 19.580 ;
        RECT 75.615 19.410 75.765 19.580 ;
        RECT 77.795 19.410 77.945 19.580 ;
        RECT 78.515 19.410 78.665 19.580 ;
        RECT 80.695 19.410 80.845 19.580 ;
        RECT 81.415 19.410 81.565 19.580 ;
        RECT 83.595 19.410 83.745 19.580 ;
        RECT 84.315 19.410 84.465 19.580 ;
        RECT 86.495 19.410 86.645 19.580 ;
        RECT 87.215 19.410 87.365 19.580 ;
        RECT 89.395 19.410 89.545 19.580 ;
        RECT 90.115 19.410 90.265 19.580 ;
        RECT 92.295 19.410 92.445 19.580 ;
      LAYER met1 ;
        RECT 0.000 19.410 92.445 19.580 ;
    END
  END RWL_17
  PIN RWL_18
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 18.060 0.365 18.230 ;
        RECT 2.395 18.060 2.545 18.230 ;
        RECT 3.115 18.060 3.265 18.230 ;
        RECT 5.295 18.060 5.445 18.230 ;
        RECT 6.015 18.060 6.165 18.230 ;
        RECT 8.195 18.060 8.345 18.230 ;
        RECT 8.915 18.060 9.065 18.230 ;
        RECT 11.095 18.060 11.245 18.230 ;
        RECT 11.815 18.060 11.965 18.230 ;
        RECT 13.995 18.060 14.145 18.230 ;
        RECT 14.715 18.060 14.865 18.230 ;
        RECT 16.895 18.060 17.045 18.230 ;
        RECT 17.615 18.060 17.765 18.230 ;
        RECT 19.795 18.060 19.945 18.230 ;
        RECT 20.515 18.060 20.665 18.230 ;
        RECT 22.695 18.060 22.845 18.230 ;
        RECT 23.415 18.060 23.565 18.230 ;
        RECT 25.595 18.060 25.745 18.230 ;
        RECT 26.315 18.060 26.465 18.230 ;
        RECT 28.495 18.060 28.645 18.230 ;
        RECT 29.215 18.060 29.365 18.230 ;
        RECT 31.395 18.060 31.545 18.230 ;
        RECT 32.115 18.060 32.265 18.230 ;
        RECT 34.295 18.060 34.445 18.230 ;
        RECT 35.015 18.060 35.165 18.230 ;
        RECT 37.195 18.060 37.345 18.230 ;
        RECT 37.915 18.060 38.065 18.230 ;
        RECT 40.095 18.060 40.245 18.230 ;
        RECT 40.815 18.060 40.965 18.230 ;
        RECT 42.995 18.060 43.145 18.230 ;
        RECT 43.715 18.060 43.865 18.230 ;
        RECT 45.895 18.060 46.045 18.230 ;
        RECT 46.615 18.060 46.765 18.230 ;
        RECT 48.795 18.060 48.945 18.230 ;
        RECT 49.515 18.060 49.665 18.230 ;
        RECT 51.695 18.060 51.845 18.230 ;
        RECT 52.415 18.060 52.565 18.230 ;
        RECT 54.595 18.060 54.745 18.230 ;
        RECT 55.315 18.060 55.465 18.230 ;
        RECT 57.495 18.060 57.645 18.230 ;
        RECT 58.215 18.060 58.365 18.230 ;
        RECT 60.395 18.060 60.545 18.230 ;
        RECT 61.115 18.060 61.265 18.230 ;
        RECT 63.295 18.060 63.445 18.230 ;
        RECT 64.015 18.060 64.165 18.230 ;
        RECT 66.195 18.060 66.345 18.230 ;
        RECT 66.915 18.060 67.065 18.230 ;
        RECT 69.095 18.060 69.245 18.230 ;
        RECT 69.815 18.060 69.965 18.230 ;
        RECT 71.995 18.060 72.145 18.230 ;
        RECT 72.715 18.060 72.865 18.230 ;
        RECT 74.895 18.060 75.045 18.230 ;
        RECT 75.615 18.060 75.765 18.230 ;
        RECT 77.795 18.060 77.945 18.230 ;
        RECT 78.515 18.060 78.665 18.230 ;
        RECT 80.695 18.060 80.845 18.230 ;
        RECT 81.415 18.060 81.565 18.230 ;
        RECT 83.595 18.060 83.745 18.230 ;
        RECT 84.315 18.060 84.465 18.230 ;
        RECT 86.495 18.060 86.645 18.230 ;
        RECT 87.215 18.060 87.365 18.230 ;
        RECT 89.395 18.060 89.545 18.230 ;
        RECT 90.115 18.060 90.265 18.230 ;
        RECT 92.295 18.060 92.445 18.230 ;
      LAYER met1 ;
        RECT 0.000 18.060 92.445 18.230 ;
    END
  END RWL_18
  PIN RWL_19
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 16.710 0.365 16.880 ;
        RECT 2.395 16.710 2.545 16.880 ;
        RECT 3.115 16.710 3.265 16.880 ;
        RECT 5.295 16.710 5.445 16.880 ;
        RECT 6.015 16.710 6.165 16.880 ;
        RECT 8.195 16.710 8.345 16.880 ;
        RECT 8.915 16.710 9.065 16.880 ;
        RECT 11.095 16.710 11.245 16.880 ;
        RECT 11.815 16.710 11.965 16.880 ;
        RECT 13.995 16.710 14.145 16.880 ;
        RECT 14.715 16.710 14.865 16.880 ;
        RECT 16.895 16.710 17.045 16.880 ;
        RECT 17.615 16.710 17.765 16.880 ;
        RECT 19.795 16.710 19.945 16.880 ;
        RECT 20.515 16.710 20.665 16.880 ;
        RECT 22.695 16.710 22.845 16.880 ;
        RECT 23.415 16.710 23.565 16.880 ;
        RECT 25.595 16.710 25.745 16.880 ;
        RECT 26.315 16.710 26.465 16.880 ;
        RECT 28.495 16.710 28.645 16.880 ;
        RECT 29.215 16.710 29.365 16.880 ;
        RECT 31.395 16.710 31.545 16.880 ;
        RECT 32.115 16.710 32.265 16.880 ;
        RECT 34.295 16.710 34.445 16.880 ;
        RECT 35.015 16.710 35.165 16.880 ;
        RECT 37.195 16.710 37.345 16.880 ;
        RECT 37.915 16.710 38.065 16.880 ;
        RECT 40.095 16.710 40.245 16.880 ;
        RECT 40.815 16.710 40.965 16.880 ;
        RECT 42.995 16.710 43.145 16.880 ;
        RECT 43.715 16.710 43.865 16.880 ;
        RECT 45.895 16.710 46.045 16.880 ;
        RECT 46.615 16.710 46.765 16.880 ;
        RECT 48.795 16.710 48.945 16.880 ;
        RECT 49.515 16.710 49.665 16.880 ;
        RECT 51.695 16.710 51.845 16.880 ;
        RECT 52.415 16.710 52.565 16.880 ;
        RECT 54.595 16.710 54.745 16.880 ;
        RECT 55.315 16.710 55.465 16.880 ;
        RECT 57.495 16.710 57.645 16.880 ;
        RECT 58.215 16.710 58.365 16.880 ;
        RECT 60.395 16.710 60.545 16.880 ;
        RECT 61.115 16.710 61.265 16.880 ;
        RECT 63.295 16.710 63.445 16.880 ;
        RECT 64.015 16.710 64.165 16.880 ;
        RECT 66.195 16.710 66.345 16.880 ;
        RECT 66.915 16.710 67.065 16.880 ;
        RECT 69.095 16.710 69.245 16.880 ;
        RECT 69.815 16.710 69.965 16.880 ;
        RECT 71.995 16.710 72.145 16.880 ;
        RECT 72.715 16.710 72.865 16.880 ;
        RECT 74.895 16.710 75.045 16.880 ;
        RECT 75.615 16.710 75.765 16.880 ;
        RECT 77.795 16.710 77.945 16.880 ;
        RECT 78.515 16.710 78.665 16.880 ;
        RECT 80.695 16.710 80.845 16.880 ;
        RECT 81.415 16.710 81.565 16.880 ;
        RECT 83.595 16.710 83.745 16.880 ;
        RECT 84.315 16.710 84.465 16.880 ;
        RECT 86.495 16.710 86.645 16.880 ;
        RECT 87.215 16.710 87.365 16.880 ;
        RECT 89.395 16.710 89.545 16.880 ;
        RECT 90.115 16.710 90.265 16.880 ;
        RECT 92.295 16.710 92.445 16.880 ;
      LAYER met1 ;
        RECT 0.000 16.710 92.445 16.880 ;
    END
  END RWL_19
  PIN RWL_20
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 15.360 0.365 15.530 ;
        RECT 2.395 15.360 2.545 15.530 ;
        RECT 3.115 15.360 3.265 15.530 ;
        RECT 5.295 15.360 5.445 15.530 ;
        RECT 6.015 15.360 6.165 15.530 ;
        RECT 8.195 15.360 8.345 15.530 ;
        RECT 8.915 15.360 9.065 15.530 ;
        RECT 11.095 15.360 11.245 15.530 ;
        RECT 11.815 15.360 11.965 15.530 ;
        RECT 13.995 15.360 14.145 15.530 ;
        RECT 14.715 15.360 14.865 15.530 ;
        RECT 16.895 15.360 17.045 15.530 ;
        RECT 17.615 15.360 17.765 15.530 ;
        RECT 19.795 15.360 19.945 15.530 ;
        RECT 20.515 15.360 20.665 15.530 ;
        RECT 22.695 15.360 22.845 15.530 ;
        RECT 23.415 15.360 23.565 15.530 ;
        RECT 25.595 15.360 25.745 15.530 ;
        RECT 26.315 15.360 26.465 15.530 ;
        RECT 28.495 15.360 28.645 15.530 ;
        RECT 29.215 15.360 29.365 15.530 ;
        RECT 31.395 15.360 31.545 15.530 ;
        RECT 32.115 15.360 32.265 15.530 ;
        RECT 34.295 15.360 34.445 15.530 ;
        RECT 35.015 15.360 35.165 15.530 ;
        RECT 37.195 15.360 37.345 15.530 ;
        RECT 37.915 15.360 38.065 15.530 ;
        RECT 40.095 15.360 40.245 15.530 ;
        RECT 40.815 15.360 40.965 15.530 ;
        RECT 42.995 15.360 43.145 15.530 ;
        RECT 43.715 15.360 43.865 15.530 ;
        RECT 45.895 15.360 46.045 15.530 ;
        RECT 46.615 15.360 46.765 15.530 ;
        RECT 48.795 15.360 48.945 15.530 ;
        RECT 49.515 15.360 49.665 15.530 ;
        RECT 51.695 15.360 51.845 15.530 ;
        RECT 52.415 15.360 52.565 15.530 ;
        RECT 54.595 15.360 54.745 15.530 ;
        RECT 55.315 15.360 55.465 15.530 ;
        RECT 57.495 15.360 57.645 15.530 ;
        RECT 58.215 15.360 58.365 15.530 ;
        RECT 60.395 15.360 60.545 15.530 ;
        RECT 61.115 15.360 61.265 15.530 ;
        RECT 63.295 15.360 63.445 15.530 ;
        RECT 64.015 15.360 64.165 15.530 ;
        RECT 66.195 15.360 66.345 15.530 ;
        RECT 66.915 15.360 67.065 15.530 ;
        RECT 69.095 15.360 69.245 15.530 ;
        RECT 69.815 15.360 69.965 15.530 ;
        RECT 71.995 15.360 72.145 15.530 ;
        RECT 72.715 15.360 72.865 15.530 ;
        RECT 74.895 15.360 75.045 15.530 ;
        RECT 75.615 15.360 75.765 15.530 ;
        RECT 77.795 15.360 77.945 15.530 ;
        RECT 78.515 15.360 78.665 15.530 ;
        RECT 80.695 15.360 80.845 15.530 ;
        RECT 81.415 15.360 81.565 15.530 ;
        RECT 83.595 15.360 83.745 15.530 ;
        RECT 84.315 15.360 84.465 15.530 ;
        RECT 86.495 15.360 86.645 15.530 ;
        RECT 87.215 15.360 87.365 15.530 ;
        RECT 89.395 15.360 89.545 15.530 ;
        RECT 90.115 15.360 90.265 15.530 ;
        RECT 92.295 15.360 92.445 15.530 ;
      LAYER met1 ;
        RECT 0.000 15.360 92.445 15.530 ;
    END
  END RWL_20
  PIN RWL_21
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 14.010 0.365 14.180 ;
        RECT 2.395 14.010 2.545 14.180 ;
        RECT 3.115 14.010 3.265 14.180 ;
        RECT 5.295 14.010 5.445 14.180 ;
        RECT 6.015 14.010 6.165 14.180 ;
        RECT 8.195 14.010 8.345 14.180 ;
        RECT 8.915 14.010 9.065 14.180 ;
        RECT 11.095 14.010 11.245 14.180 ;
        RECT 11.815 14.010 11.965 14.180 ;
        RECT 13.995 14.010 14.145 14.180 ;
        RECT 14.715 14.010 14.865 14.180 ;
        RECT 16.895 14.010 17.045 14.180 ;
        RECT 17.615 14.010 17.765 14.180 ;
        RECT 19.795 14.010 19.945 14.180 ;
        RECT 20.515 14.010 20.665 14.180 ;
        RECT 22.695 14.010 22.845 14.180 ;
        RECT 23.415 14.010 23.565 14.180 ;
        RECT 25.595 14.010 25.745 14.180 ;
        RECT 26.315 14.010 26.465 14.180 ;
        RECT 28.495 14.010 28.645 14.180 ;
        RECT 29.215 14.010 29.365 14.180 ;
        RECT 31.395 14.010 31.545 14.180 ;
        RECT 32.115 14.010 32.265 14.180 ;
        RECT 34.295 14.010 34.445 14.180 ;
        RECT 35.015 14.010 35.165 14.180 ;
        RECT 37.195 14.010 37.345 14.180 ;
        RECT 37.915 14.010 38.065 14.180 ;
        RECT 40.095 14.010 40.245 14.180 ;
        RECT 40.815 14.010 40.965 14.180 ;
        RECT 42.995 14.010 43.145 14.180 ;
        RECT 43.715 14.010 43.865 14.180 ;
        RECT 45.895 14.010 46.045 14.180 ;
        RECT 46.615 14.010 46.765 14.180 ;
        RECT 48.795 14.010 48.945 14.180 ;
        RECT 49.515 14.010 49.665 14.180 ;
        RECT 51.695 14.010 51.845 14.180 ;
        RECT 52.415 14.010 52.565 14.180 ;
        RECT 54.595 14.010 54.745 14.180 ;
        RECT 55.315 14.010 55.465 14.180 ;
        RECT 57.495 14.010 57.645 14.180 ;
        RECT 58.215 14.010 58.365 14.180 ;
        RECT 60.395 14.010 60.545 14.180 ;
        RECT 61.115 14.010 61.265 14.180 ;
        RECT 63.295 14.010 63.445 14.180 ;
        RECT 64.015 14.010 64.165 14.180 ;
        RECT 66.195 14.010 66.345 14.180 ;
        RECT 66.915 14.010 67.065 14.180 ;
        RECT 69.095 14.010 69.245 14.180 ;
        RECT 69.815 14.010 69.965 14.180 ;
        RECT 71.995 14.010 72.145 14.180 ;
        RECT 72.715 14.010 72.865 14.180 ;
        RECT 74.895 14.010 75.045 14.180 ;
        RECT 75.615 14.010 75.765 14.180 ;
        RECT 77.795 14.010 77.945 14.180 ;
        RECT 78.515 14.010 78.665 14.180 ;
        RECT 80.695 14.010 80.845 14.180 ;
        RECT 81.415 14.010 81.565 14.180 ;
        RECT 83.595 14.010 83.745 14.180 ;
        RECT 84.315 14.010 84.465 14.180 ;
        RECT 86.495 14.010 86.645 14.180 ;
        RECT 87.215 14.010 87.365 14.180 ;
        RECT 89.395 14.010 89.545 14.180 ;
        RECT 90.115 14.010 90.265 14.180 ;
        RECT 92.295 14.010 92.445 14.180 ;
      LAYER met1 ;
        RECT 0.000 14.010 92.445 14.180 ;
    END
  END RWL_21
  PIN RWL_22
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 12.660 0.365 12.830 ;
        RECT 2.395 12.660 2.545 12.830 ;
        RECT 3.115 12.660 3.265 12.830 ;
        RECT 5.295 12.660 5.445 12.830 ;
        RECT 6.015 12.660 6.165 12.830 ;
        RECT 8.195 12.660 8.345 12.830 ;
        RECT 8.915 12.660 9.065 12.830 ;
        RECT 11.095 12.660 11.245 12.830 ;
        RECT 11.815 12.660 11.965 12.830 ;
        RECT 13.995 12.660 14.145 12.830 ;
        RECT 14.715 12.660 14.865 12.830 ;
        RECT 16.895 12.660 17.045 12.830 ;
        RECT 17.615 12.660 17.765 12.830 ;
        RECT 19.795 12.660 19.945 12.830 ;
        RECT 20.515 12.660 20.665 12.830 ;
        RECT 22.695 12.660 22.845 12.830 ;
        RECT 23.415 12.660 23.565 12.830 ;
        RECT 25.595 12.660 25.745 12.830 ;
        RECT 26.315 12.660 26.465 12.830 ;
        RECT 28.495 12.660 28.645 12.830 ;
        RECT 29.215 12.660 29.365 12.830 ;
        RECT 31.395 12.660 31.545 12.830 ;
        RECT 32.115 12.660 32.265 12.830 ;
        RECT 34.295 12.660 34.445 12.830 ;
        RECT 35.015 12.660 35.165 12.830 ;
        RECT 37.195 12.660 37.345 12.830 ;
        RECT 37.915 12.660 38.065 12.830 ;
        RECT 40.095 12.660 40.245 12.830 ;
        RECT 40.815 12.660 40.965 12.830 ;
        RECT 42.995 12.660 43.145 12.830 ;
        RECT 43.715 12.660 43.865 12.830 ;
        RECT 45.895 12.660 46.045 12.830 ;
        RECT 46.615 12.660 46.765 12.830 ;
        RECT 48.795 12.660 48.945 12.830 ;
        RECT 49.515 12.660 49.665 12.830 ;
        RECT 51.695 12.660 51.845 12.830 ;
        RECT 52.415 12.660 52.565 12.830 ;
        RECT 54.595 12.660 54.745 12.830 ;
        RECT 55.315 12.660 55.465 12.830 ;
        RECT 57.495 12.660 57.645 12.830 ;
        RECT 58.215 12.660 58.365 12.830 ;
        RECT 60.395 12.660 60.545 12.830 ;
        RECT 61.115 12.660 61.265 12.830 ;
        RECT 63.295 12.660 63.445 12.830 ;
        RECT 64.015 12.660 64.165 12.830 ;
        RECT 66.195 12.660 66.345 12.830 ;
        RECT 66.915 12.660 67.065 12.830 ;
        RECT 69.095 12.660 69.245 12.830 ;
        RECT 69.815 12.660 69.965 12.830 ;
        RECT 71.995 12.660 72.145 12.830 ;
        RECT 72.715 12.660 72.865 12.830 ;
        RECT 74.895 12.660 75.045 12.830 ;
        RECT 75.615 12.660 75.765 12.830 ;
        RECT 77.795 12.660 77.945 12.830 ;
        RECT 78.515 12.660 78.665 12.830 ;
        RECT 80.695 12.660 80.845 12.830 ;
        RECT 81.415 12.660 81.565 12.830 ;
        RECT 83.595 12.660 83.745 12.830 ;
        RECT 84.315 12.660 84.465 12.830 ;
        RECT 86.495 12.660 86.645 12.830 ;
        RECT 87.215 12.660 87.365 12.830 ;
        RECT 89.395 12.660 89.545 12.830 ;
        RECT 90.115 12.660 90.265 12.830 ;
        RECT 92.295 12.660 92.445 12.830 ;
      LAYER met1 ;
        RECT 0.000 12.660 92.445 12.830 ;
    END
  END RWL_22
  PIN RWL_23
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 11.310 0.365 11.480 ;
        RECT 2.395 11.310 2.545 11.480 ;
        RECT 3.115 11.310 3.265 11.480 ;
        RECT 5.295 11.310 5.445 11.480 ;
        RECT 6.015 11.310 6.165 11.480 ;
        RECT 8.195 11.310 8.345 11.480 ;
        RECT 8.915 11.310 9.065 11.480 ;
        RECT 11.095 11.310 11.245 11.480 ;
        RECT 11.815 11.310 11.965 11.480 ;
        RECT 13.995 11.310 14.145 11.480 ;
        RECT 14.715 11.310 14.865 11.480 ;
        RECT 16.895 11.310 17.045 11.480 ;
        RECT 17.615 11.310 17.765 11.480 ;
        RECT 19.795 11.310 19.945 11.480 ;
        RECT 20.515 11.310 20.665 11.480 ;
        RECT 22.695 11.310 22.845 11.480 ;
        RECT 23.415 11.310 23.565 11.480 ;
        RECT 25.595 11.310 25.745 11.480 ;
        RECT 26.315 11.310 26.465 11.480 ;
        RECT 28.495 11.310 28.645 11.480 ;
        RECT 29.215 11.310 29.365 11.480 ;
        RECT 31.395 11.310 31.545 11.480 ;
        RECT 32.115 11.310 32.265 11.480 ;
        RECT 34.295 11.310 34.445 11.480 ;
        RECT 35.015 11.310 35.165 11.480 ;
        RECT 37.195 11.310 37.345 11.480 ;
        RECT 37.915 11.310 38.065 11.480 ;
        RECT 40.095 11.310 40.245 11.480 ;
        RECT 40.815 11.310 40.965 11.480 ;
        RECT 42.995 11.310 43.145 11.480 ;
        RECT 43.715 11.310 43.865 11.480 ;
        RECT 45.895 11.310 46.045 11.480 ;
        RECT 46.615 11.310 46.765 11.480 ;
        RECT 48.795 11.310 48.945 11.480 ;
        RECT 49.515 11.310 49.665 11.480 ;
        RECT 51.695 11.310 51.845 11.480 ;
        RECT 52.415 11.310 52.565 11.480 ;
        RECT 54.595 11.310 54.745 11.480 ;
        RECT 55.315 11.310 55.465 11.480 ;
        RECT 57.495 11.310 57.645 11.480 ;
        RECT 58.215 11.310 58.365 11.480 ;
        RECT 60.395 11.310 60.545 11.480 ;
        RECT 61.115 11.310 61.265 11.480 ;
        RECT 63.295 11.310 63.445 11.480 ;
        RECT 64.015 11.310 64.165 11.480 ;
        RECT 66.195 11.310 66.345 11.480 ;
        RECT 66.915 11.310 67.065 11.480 ;
        RECT 69.095 11.310 69.245 11.480 ;
        RECT 69.815 11.310 69.965 11.480 ;
        RECT 71.995 11.310 72.145 11.480 ;
        RECT 72.715 11.310 72.865 11.480 ;
        RECT 74.895 11.310 75.045 11.480 ;
        RECT 75.615 11.310 75.765 11.480 ;
        RECT 77.795 11.310 77.945 11.480 ;
        RECT 78.515 11.310 78.665 11.480 ;
        RECT 80.695 11.310 80.845 11.480 ;
        RECT 81.415 11.310 81.565 11.480 ;
        RECT 83.595 11.310 83.745 11.480 ;
        RECT 84.315 11.310 84.465 11.480 ;
        RECT 86.495 11.310 86.645 11.480 ;
        RECT 87.215 11.310 87.365 11.480 ;
        RECT 89.395 11.310 89.545 11.480 ;
        RECT 90.115 11.310 90.265 11.480 ;
        RECT 92.295 11.310 92.445 11.480 ;
      LAYER met1 ;
        RECT 0.000 11.310 92.445 11.480 ;
    END
  END RWL_23
  PIN RWL_24
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 9.960 0.365 10.130 ;
        RECT 2.395 9.960 2.545 10.130 ;
        RECT 3.115 9.960 3.265 10.130 ;
        RECT 5.295 9.960 5.445 10.130 ;
        RECT 6.015 9.960 6.165 10.130 ;
        RECT 8.195 9.960 8.345 10.130 ;
        RECT 8.915 9.960 9.065 10.130 ;
        RECT 11.095 9.960 11.245 10.130 ;
        RECT 11.815 9.960 11.965 10.130 ;
        RECT 13.995 9.960 14.145 10.130 ;
        RECT 14.715 9.960 14.865 10.130 ;
        RECT 16.895 9.960 17.045 10.130 ;
        RECT 17.615 9.960 17.765 10.130 ;
        RECT 19.795 9.960 19.945 10.130 ;
        RECT 20.515 9.960 20.665 10.130 ;
        RECT 22.695 9.960 22.845 10.130 ;
        RECT 23.415 9.960 23.565 10.130 ;
        RECT 25.595 9.960 25.745 10.130 ;
        RECT 26.315 9.960 26.465 10.130 ;
        RECT 28.495 9.960 28.645 10.130 ;
        RECT 29.215 9.960 29.365 10.130 ;
        RECT 31.395 9.960 31.545 10.130 ;
        RECT 32.115 9.960 32.265 10.130 ;
        RECT 34.295 9.960 34.445 10.130 ;
        RECT 35.015 9.960 35.165 10.130 ;
        RECT 37.195 9.960 37.345 10.130 ;
        RECT 37.915 9.960 38.065 10.130 ;
        RECT 40.095 9.960 40.245 10.130 ;
        RECT 40.815 9.960 40.965 10.130 ;
        RECT 42.995 9.960 43.145 10.130 ;
        RECT 43.715 9.960 43.865 10.130 ;
        RECT 45.895 9.960 46.045 10.130 ;
        RECT 46.615 9.960 46.765 10.130 ;
        RECT 48.795 9.960 48.945 10.130 ;
        RECT 49.515 9.960 49.665 10.130 ;
        RECT 51.695 9.960 51.845 10.130 ;
        RECT 52.415 9.960 52.565 10.130 ;
        RECT 54.595 9.960 54.745 10.130 ;
        RECT 55.315 9.960 55.465 10.130 ;
        RECT 57.495 9.960 57.645 10.130 ;
        RECT 58.215 9.960 58.365 10.130 ;
        RECT 60.395 9.960 60.545 10.130 ;
        RECT 61.115 9.960 61.265 10.130 ;
        RECT 63.295 9.960 63.445 10.130 ;
        RECT 64.015 9.960 64.165 10.130 ;
        RECT 66.195 9.960 66.345 10.130 ;
        RECT 66.915 9.960 67.065 10.130 ;
        RECT 69.095 9.960 69.245 10.130 ;
        RECT 69.815 9.960 69.965 10.130 ;
        RECT 71.995 9.960 72.145 10.130 ;
        RECT 72.715 9.960 72.865 10.130 ;
        RECT 74.895 9.960 75.045 10.130 ;
        RECT 75.615 9.960 75.765 10.130 ;
        RECT 77.795 9.960 77.945 10.130 ;
        RECT 78.515 9.960 78.665 10.130 ;
        RECT 80.695 9.960 80.845 10.130 ;
        RECT 81.415 9.960 81.565 10.130 ;
        RECT 83.595 9.960 83.745 10.130 ;
        RECT 84.315 9.960 84.465 10.130 ;
        RECT 86.495 9.960 86.645 10.130 ;
        RECT 87.215 9.960 87.365 10.130 ;
        RECT 89.395 9.960 89.545 10.130 ;
        RECT 90.115 9.960 90.265 10.130 ;
        RECT 92.295 9.960 92.445 10.130 ;
      LAYER met1 ;
        RECT 0.000 9.960 92.445 10.130 ;
    END
  END RWL_24
  PIN RWL_25
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 8.610 0.365 8.780 ;
        RECT 2.395 8.610 2.545 8.780 ;
        RECT 3.115 8.610 3.265 8.780 ;
        RECT 5.295 8.610 5.445 8.780 ;
        RECT 6.015 8.610 6.165 8.780 ;
        RECT 8.195 8.610 8.345 8.780 ;
        RECT 8.915 8.610 9.065 8.780 ;
        RECT 11.095 8.610 11.245 8.780 ;
        RECT 11.815 8.610 11.965 8.780 ;
        RECT 13.995 8.610 14.145 8.780 ;
        RECT 14.715 8.610 14.865 8.780 ;
        RECT 16.895 8.610 17.045 8.780 ;
        RECT 17.615 8.610 17.765 8.780 ;
        RECT 19.795 8.610 19.945 8.780 ;
        RECT 20.515 8.610 20.665 8.780 ;
        RECT 22.695 8.610 22.845 8.780 ;
        RECT 23.415 8.610 23.565 8.780 ;
        RECT 25.595 8.610 25.745 8.780 ;
        RECT 26.315 8.610 26.465 8.780 ;
        RECT 28.495 8.610 28.645 8.780 ;
        RECT 29.215 8.610 29.365 8.780 ;
        RECT 31.395 8.610 31.545 8.780 ;
        RECT 32.115 8.610 32.265 8.780 ;
        RECT 34.295 8.610 34.445 8.780 ;
        RECT 35.015 8.610 35.165 8.780 ;
        RECT 37.195 8.610 37.345 8.780 ;
        RECT 37.915 8.610 38.065 8.780 ;
        RECT 40.095 8.610 40.245 8.780 ;
        RECT 40.815 8.610 40.965 8.780 ;
        RECT 42.995 8.610 43.145 8.780 ;
        RECT 43.715 8.610 43.865 8.780 ;
        RECT 45.895 8.610 46.045 8.780 ;
        RECT 46.615 8.610 46.765 8.780 ;
        RECT 48.795 8.610 48.945 8.780 ;
        RECT 49.515 8.610 49.665 8.780 ;
        RECT 51.695 8.610 51.845 8.780 ;
        RECT 52.415 8.610 52.565 8.780 ;
        RECT 54.595 8.610 54.745 8.780 ;
        RECT 55.315 8.610 55.465 8.780 ;
        RECT 57.495 8.610 57.645 8.780 ;
        RECT 58.215 8.610 58.365 8.780 ;
        RECT 60.395 8.610 60.545 8.780 ;
        RECT 61.115 8.610 61.265 8.780 ;
        RECT 63.295 8.610 63.445 8.780 ;
        RECT 64.015 8.610 64.165 8.780 ;
        RECT 66.195 8.610 66.345 8.780 ;
        RECT 66.915 8.610 67.065 8.780 ;
        RECT 69.095 8.610 69.245 8.780 ;
        RECT 69.815 8.610 69.965 8.780 ;
        RECT 71.995 8.610 72.145 8.780 ;
        RECT 72.715 8.610 72.865 8.780 ;
        RECT 74.895 8.610 75.045 8.780 ;
        RECT 75.615 8.610 75.765 8.780 ;
        RECT 77.795 8.610 77.945 8.780 ;
        RECT 78.515 8.610 78.665 8.780 ;
        RECT 80.695 8.610 80.845 8.780 ;
        RECT 81.415 8.610 81.565 8.780 ;
        RECT 83.595 8.610 83.745 8.780 ;
        RECT 84.315 8.610 84.465 8.780 ;
        RECT 86.495 8.610 86.645 8.780 ;
        RECT 87.215 8.610 87.365 8.780 ;
        RECT 89.395 8.610 89.545 8.780 ;
        RECT 90.115 8.610 90.265 8.780 ;
        RECT 92.295 8.610 92.445 8.780 ;
      LAYER met1 ;
        RECT 0.000 8.610 92.445 8.780 ;
    END
  END RWL_25
  PIN RWL_26
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 7.260 0.365 7.430 ;
        RECT 2.395 7.260 2.545 7.430 ;
        RECT 3.115 7.260 3.265 7.430 ;
        RECT 5.295 7.260 5.445 7.430 ;
        RECT 6.015 7.260 6.165 7.430 ;
        RECT 8.195 7.260 8.345 7.430 ;
        RECT 8.915 7.260 9.065 7.430 ;
        RECT 11.095 7.260 11.245 7.430 ;
        RECT 11.815 7.260 11.965 7.430 ;
        RECT 13.995 7.260 14.145 7.430 ;
        RECT 14.715 7.260 14.865 7.430 ;
        RECT 16.895 7.260 17.045 7.430 ;
        RECT 17.615 7.260 17.765 7.430 ;
        RECT 19.795 7.260 19.945 7.430 ;
        RECT 20.515 7.260 20.665 7.430 ;
        RECT 22.695 7.260 22.845 7.430 ;
        RECT 23.415 7.260 23.565 7.430 ;
        RECT 25.595 7.260 25.745 7.430 ;
        RECT 26.315 7.260 26.465 7.430 ;
        RECT 28.495 7.260 28.645 7.430 ;
        RECT 29.215 7.260 29.365 7.430 ;
        RECT 31.395 7.260 31.545 7.430 ;
        RECT 32.115 7.260 32.265 7.430 ;
        RECT 34.295 7.260 34.445 7.430 ;
        RECT 35.015 7.260 35.165 7.430 ;
        RECT 37.195 7.260 37.345 7.430 ;
        RECT 37.915 7.260 38.065 7.430 ;
        RECT 40.095 7.260 40.245 7.430 ;
        RECT 40.815 7.260 40.965 7.430 ;
        RECT 42.995 7.260 43.145 7.430 ;
        RECT 43.715 7.260 43.865 7.430 ;
        RECT 45.895 7.260 46.045 7.430 ;
        RECT 46.615 7.260 46.765 7.430 ;
        RECT 48.795 7.260 48.945 7.430 ;
        RECT 49.515 7.260 49.665 7.430 ;
        RECT 51.695 7.260 51.845 7.430 ;
        RECT 52.415 7.260 52.565 7.430 ;
        RECT 54.595 7.260 54.745 7.430 ;
        RECT 55.315 7.260 55.465 7.430 ;
        RECT 57.495 7.260 57.645 7.430 ;
        RECT 58.215 7.260 58.365 7.430 ;
        RECT 60.395 7.260 60.545 7.430 ;
        RECT 61.115 7.260 61.265 7.430 ;
        RECT 63.295 7.260 63.445 7.430 ;
        RECT 64.015 7.260 64.165 7.430 ;
        RECT 66.195 7.260 66.345 7.430 ;
        RECT 66.915 7.260 67.065 7.430 ;
        RECT 69.095 7.260 69.245 7.430 ;
        RECT 69.815 7.260 69.965 7.430 ;
        RECT 71.995 7.260 72.145 7.430 ;
        RECT 72.715 7.260 72.865 7.430 ;
        RECT 74.895 7.260 75.045 7.430 ;
        RECT 75.615 7.260 75.765 7.430 ;
        RECT 77.795 7.260 77.945 7.430 ;
        RECT 78.515 7.260 78.665 7.430 ;
        RECT 80.695 7.260 80.845 7.430 ;
        RECT 81.415 7.260 81.565 7.430 ;
        RECT 83.595 7.260 83.745 7.430 ;
        RECT 84.315 7.260 84.465 7.430 ;
        RECT 86.495 7.260 86.645 7.430 ;
        RECT 87.215 7.260 87.365 7.430 ;
        RECT 89.395 7.260 89.545 7.430 ;
        RECT 90.115 7.260 90.265 7.430 ;
        RECT 92.295 7.260 92.445 7.430 ;
      LAYER met1 ;
        RECT 0.000 7.260 92.445 7.430 ;
    END
  END RWL_26
  PIN RWL_27
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 5.910 0.365 6.080 ;
        RECT 2.395 5.910 2.545 6.080 ;
        RECT 3.115 5.910 3.265 6.080 ;
        RECT 5.295 5.910 5.445 6.080 ;
        RECT 6.015 5.910 6.165 6.080 ;
        RECT 8.195 5.910 8.345 6.080 ;
        RECT 8.915 5.910 9.065 6.080 ;
        RECT 11.095 5.910 11.245 6.080 ;
        RECT 11.815 5.910 11.965 6.080 ;
        RECT 13.995 5.910 14.145 6.080 ;
        RECT 14.715 5.910 14.865 6.080 ;
        RECT 16.895 5.910 17.045 6.080 ;
        RECT 17.615 5.910 17.765 6.080 ;
        RECT 19.795 5.910 19.945 6.080 ;
        RECT 20.515 5.910 20.665 6.080 ;
        RECT 22.695 5.910 22.845 6.080 ;
        RECT 23.415 5.910 23.565 6.080 ;
        RECT 25.595 5.910 25.745 6.080 ;
        RECT 26.315 5.910 26.465 6.080 ;
        RECT 28.495 5.910 28.645 6.080 ;
        RECT 29.215 5.910 29.365 6.080 ;
        RECT 31.395 5.910 31.545 6.080 ;
        RECT 32.115 5.910 32.265 6.080 ;
        RECT 34.295 5.910 34.445 6.080 ;
        RECT 35.015 5.910 35.165 6.080 ;
        RECT 37.195 5.910 37.345 6.080 ;
        RECT 37.915 5.910 38.065 6.080 ;
        RECT 40.095 5.910 40.245 6.080 ;
        RECT 40.815 5.910 40.965 6.080 ;
        RECT 42.995 5.910 43.145 6.080 ;
        RECT 43.715 5.910 43.865 6.080 ;
        RECT 45.895 5.910 46.045 6.080 ;
        RECT 46.615 5.910 46.765 6.080 ;
        RECT 48.795 5.910 48.945 6.080 ;
        RECT 49.515 5.910 49.665 6.080 ;
        RECT 51.695 5.910 51.845 6.080 ;
        RECT 52.415 5.910 52.565 6.080 ;
        RECT 54.595 5.910 54.745 6.080 ;
        RECT 55.315 5.910 55.465 6.080 ;
        RECT 57.495 5.910 57.645 6.080 ;
        RECT 58.215 5.910 58.365 6.080 ;
        RECT 60.395 5.910 60.545 6.080 ;
        RECT 61.115 5.910 61.265 6.080 ;
        RECT 63.295 5.910 63.445 6.080 ;
        RECT 64.015 5.910 64.165 6.080 ;
        RECT 66.195 5.910 66.345 6.080 ;
        RECT 66.915 5.910 67.065 6.080 ;
        RECT 69.095 5.910 69.245 6.080 ;
        RECT 69.815 5.910 69.965 6.080 ;
        RECT 71.995 5.910 72.145 6.080 ;
        RECT 72.715 5.910 72.865 6.080 ;
        RECT 74.895 5.910 75.045 6.080 ;
        RECT 75.615 5.910 75.765 6.080 ;
        RECT 77.795 5.910 77.945 6.080 ;
        RECT 78.515 5.910 78.665 6.080 ;
        RECT 80.695 5.910 80.845 6.080 ;
        RECT 81.415 5.910 81.565 6.080 ;
        RECT 83.595 5.910 83.745 6.080 ;
        RECT 84.315 5.910 84.465 6.080 ;
        RECT 86.495 5.910 86.645 6.080 ;
        RECT 87.215 5.910 87.365 6.080 ;
        RECT 89.395 5.910 89.545 6.080 ;
        RECT 90.115 5.910 90.265 6.080 ;
        RECT 92.295 5.910 92.445 6.080 ;
      LAYER met1 ;
        RECT 0.000 5.910 92.445 6.080 ;
    END
  END RWL_27
  PIN RWL_28
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 4.560 0.365 4.730 ;
        RECT 2.395 4.560 2.545 4.730 ;
        RECT 3.115 4.560 3.265 4.730 ;
        RECT 5.295 4.560 5.445 4.730 ;
        RECT 6.015 4.560 6.165 4.730 ;
        RECT 8.195 4.560 8.345 4.730 ;
        RECT 8.915 4.560 9.065 4.730 ;
        RECT 11.095 4.560 11.245 4.730 ;
        RECT 11.815 4.560 11.965 4.730 ;
        RECT 13.995 4.560 14.145 4.730 ;
        RECT 14.715 4.560 14.865 4.730 ;
        RECT 16.895 4.560 17.045 4.730 ;
        RECT 17.615 4.560 17.765 4.730 ;
        RECT 19.795 4.560 19.945 4.730 ;
        RECT 20.515 4.560 20.665 4.730 ;
        RECT 22.695 4.560 22.845 4.730 ;
        RECT 23.415 4.560 23.565 4.730 ;
        RECT 25.595 4.560 25.745 4.730 ;
        RECT 26.315 4.560 26.465 4.730 ;
        RECT 28.495 4.560 28.645 4.730 ;
        RECT 29.215 4.560 29.365 4.730 ;
        RECT 31.395 4.560 31.545 4.730 ;
        RECT 32.115 4.560 32.265 4.730 ;
        RECT 34.295 4.560 34.445 4.730 ;
        RECT 35.015 4.560 35.165 4.730 ;
        RECT 37.195 4.560 37.345 4.730 ;
        RECT 37.915 4.560 38.065 4.730 ;
        RECT 40.095 4.560 40.245 4.730 ;
        RECT 40.815 4.560 40.965 4.730 ;
        RECT 42.995 4.560 43.145 4.730 ;
        RECT 43.715 4.560 43.865 4.730 ;
        RECT 45.895 4.560 46.045 4.730 ;
        RECT 46.615 4.560 46.765 4.730 ;
        RECT 48.795 4.560 48.945 4.730 ;
        RECT 49.515 4.560 49.665 4.730 ;
        RECT 51.695 4.560 51.845 4.730 ;
        RECT 52.415 4.560 52.565 4.730 ;
        RECT 54.595 4.560 54.745 4.730 ;
        RECT 55.315 4.560 55.465 4.730 ;
        RECT 57.495 4.560 57.645 4.730 ;
        RECT 58.215 4.560 58.365 4.730 ;
        RECT 60.395 4.560 60.545 4.730 ;
        RECT 61.115 4.560 61.265 4.730 ;
        RECT 63.295 4.560 63.445 4.730 ;
        RECT 64.015 4.560 64.165 4.730 ;
        RECT 66.195 4.560 66.345 4.730 ;
        RECT 66.915 4.560 67.065 4.730 ;
        RECT 69.095 4.560 69.245 4.730 ;
        RECT 69.815 4.560 69.965 4.730 ;
        RECT 71.995 4.560 72.145 4.730 ;
        RECT 72.715 4.560 72.865 4.730 ;
        RECT 74.895 4.560 75.045 4.730 ;
        RECT 75.615 4.560 75.765 4.730 ;
        RECT 77.795 4.560 77.945 4.730 ;
        RECT 78.515 4.560 78.665 4.730 ;
        RECT 80.695 4.560 80.845 4.730 ;
        RECT 81.415 4.560 81.565 4.730 ;
        RECT 83.595 4.560 83.745 4.730 ;
        RECT 84.315 4.560 84.465 4.730 ;
        RECT 86.495 4.560 86.645 4.730 ;
        RECT 87.215 4.560 87.365 4.730 ;
        RECT 89.395 4.560 89.545 4.730 ;
        RECT 90.115 4.560 90.265 4.730 ;
        RECT 92.295 4.560 92.445 4.730 ;
      LAYER met1 ;
        RECT 0.000 4.560 92.445 4.730 ;
    END
  END RWL_28
  PIN RWL_29
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 3.210 0.365 3.380 ;
        RECT 2.395 3.210 2.545 3.380 ;
        RECT 3.115 3.210 3.265 3.380 ;
        RECT 5.295 3.210 5.445 3.380 ;
        RECT 6.015 3.210 6.165 3.380 ;
        RECT 8.195 3.210 8.345 3.380 ;
        RECT 8.915 3.210 9.065 3.380 ;
        RECT 11.095 3.210 11.245 3.380 ;
        RECT 11.815 3.210 11.965 3.380 ;
        RECT 13.995 3.210 14.145 3.380 ;
        RECT 14.715 3.210 14.865 3.380 ;
        RECT 16.895 3.210 17.045 3.380 ;
        RECT 17.615 3.210 17.765 3.380 ;
        RECT 19.795 3.210 19.945 3.380 ;
        RECT 20.515 3.210 20.665 3.380 ;
        RECT 22.695 3.210 22.845 3.380 ;
        RECT 23.415 3.210 23.565 3.380 ;
        RECT 25.595 3.210 25.745 3.380 ;
        RECT 26.315 3.210 26.465 3.380 ;
        RECT 28.495 3.210 28.645 3.380 ;
        RECT 29.215 3.210 29.365 3.380 ;
        RECT 31.395 3.210 31.545 3.380 ;
        RECT 32.115 3.210 32.265 3.380 ;
        RECT 34.295 3.210 34.445 3.380 ;
        RECT 35.015 3.210 35.165 3.380 ;
        RECT 37.195 3.210 37.345 3.380 ;
        RECT 37.915 3.210 38.065 3.380 ;
        RECT 40.095 3.210 40.245 3.380 ;
        RECT 40.815 3.210 40.965 3.380 ;
        RECT 42.995 3.210 43.145 3.380 ;
        RECT 43.715 3.210 43.865 3.380 ;
        RECT 45.895 3.210 46.045 3.380 ;
        RECT 46.615 3.210 46.765 3.380 ;
        RECT 48.795 3.210 48.945 3.380 ;
        RECT 49.515 3.210 49.665 3.380 ;
        RECT 51.695 3.210 51.845 3.380 ;
        RECT 52.415 3.210 52.565 3.380 ;
        RECT 54.595 3.210 54.745 3.380 ;
        RECT 55.315 3.210 55.465 3.380 ;
        RECT 57.495 3.210 57.645 3.380 ;
        RECT 58.215 3.210 58.365 3.380 ;
        RECT 60.395 3.210 60.545 3.380 ;
        RECT 61.115 3.210 61.265 3.380 ;
        RECT 63.295 3.210 63.445 3.380 ;
        RECT 64.015 3.210 64.165 3.380 ;
        RECT 66.195 3.210 66.345 3.380 ;
        RECT 66.915 3.210 67.065 3.380 ;
        RECT 69.095 3.210 69.245 3.380 ;
        RECT 69.815 3.210 69.965 3.380 ;
        RECT 71.995 3.210 72.145 3.380 ;
        RECT 72.715 3.210 72.865 3.380 ;
        RECT 74.895 3.210 75.045 3.380 ;
        RECT 75.615 3.210 75.765 3.380 ;
        RECT 77.795 3.210 77.945 3.380 ;
        RECT 78.515 3.210 78.665 3.380 ;
        RECT 80.695 3.210 80.845 3.380 ;
        RECT 81.415 3.210 81.565 3.380 ;
        RECT 83.595 3.210 83.745 3.380 ;
        RECT 84.315 3.210 84.465 3.380 ;
        RECT 86.495 3.210 86.645 3.380 ;
        RECT 87.215 3.210 87.365 3.380 ;
        RECT 89.395 3.210 89.545 3.380 ;
        RECT 90.115 3.210 90.265 3.380 ;
        RECT 92.295 3.210 92.445 3.380 ;
      LAYER met1 ;
        RECT 0.000 3.210 92.445 3.380 ;
    END
  END RWL_29
  PIN RWL_30
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 1.860 0.365 2.030 ;
        RECT 2.395 1.860 2.545 2.030 ;
        RECT 3.115 1.860 3.265 2.030 ;
        RECT 5.295 1.860 5.445 2.030 ;
        RECT 6.015 1.860 6.165 2.030 ;
        RECT 8.195 1.860 8.345 2.030 ;
        RECT 8.915 1.860 9.065 2.030 ;
        RECT 11.095 1.860 11.245 2.030 ;
        RECT 11.815 1.860 11.965 2.030 ;
        RECT 13.995 1.860 14.145 2.030 ;
        RECT 14.715 1.860 14.865 2.030 ;
        RECT 16.895 1.860 17.045 2.030 ;
        RECT 17.615 1.860 17.765 2.030 ;
        RECT 19.795 1.860 19.945 2.030 ;
        RECT 20.515 1.860 20.665 2.030 ;
        RECT 22.695 1.860 22.845 2.030 ;
        RECT 23.415 1.865 23.565 2.035 ;
        RECT 25.595 1.865 25.745 2.035 ;
        RECT 26.315 1.865 26.465 2.035 ;
        RECT 28.495 1.865 28.645 2.035 ;
        RECT 29.215 1.865 29.365 2.035 ;
        RECT 31.395 1.865 31.545 2.035 ;
        RECT 32.115 1.865 32.265 2.035 ;
        RECT 34.295 1.865 34.445 2.035 ;
        RECT 35.015 1.865 35.165 2.035 ;
        RECT 37.195 1.865 37.345 2.035 ;
        RECT 37.915 1.865 38.065 2.035 ;
        RECT 40.095 1.865 40.245 2.035 ;
        RECT 40.815 1.865 40.965 2.035 ;
        RECT 42.995 1.865 43.145 2.035 ;
        RECT 43.715 1.865 43.865 2.035 ;
        RECT 45.895 1.865 46.045 2.035 ;
        RECT 46.615 1.865 46.765 2.035 ;
        RECT 48.795 1.865 48.945 2.035 ;
        RECT 49.515 1.865 49.665 2.035 ;
        RECT 51.695 1.865 51.845 2.035 ;
        RECT 52.415 1.865 52.565 2.035 ;
        RECT 54.595 1.865 54.745 2.035 ;
        RECT 55.315 1.865 55.465 2.035 ;
        RECT 57.495 1.865 57.645 2.035 ;
        RECT 58.215 1.865 58.365 2.035 ;
        RECT 60.395 1.865 60.545 2.035 ;
        RECT 61.115 1.865 61.265 2.035 ;
        RECT 63.295 1.865 63.445 2.035 ;
        RECT 64.015 1.865 64.165 2.035 ;
        RECT 66.195 1.865 66.345 2.035 ;
        RECT 66.915 1.865 67.065 2.035 ;
        RECT 69.095 1.865 69.245 2.035 ;
        RECT 69.815 1.865 69.965 2.035 ;
        RECT 71.995 1.865 72.145 2.035 ;
        RECT 72.715 1.865 72.865 2.035 ;
        RECT 74.895 1.865 75.045 2.035 ;
        RECT 75.615 1.865 75.765 2.035 ;
        RECT 77.795 1.865 77.945 2.035 ;
        RECT 78.515 1.865 78.665 2.035 ;
        RECT 80.695 1.865 80.845 2.035 ;
        RECT 81.415 1.865 81.565 2.035 ;
        RECT 83.595 1.865 83.745 2.035 ;
        RECT 84.315 1.865 84.465 2.035 ;
        RECT 86.495 1.865 86.645 2.035 ;
        RECT 87.215 1.865 87.365 2.035 ;
        RECT 89.395 1.865 89.545 2.035 ;
        RECT 90.115 1.865 90.265 2.035 ;
        RECT 92.295 1.865 92.445 2.035 ;
      LAYER met1 ;
        RECT 23.200 2.030 69.245 2.035 ;
        RECT 69.600 2.030 92.445 2.035 ;
        RECT 0.000 1.865 92.445 2.030 ;
        RECT 0.000 1.860 23.415 1.865 ;
        RECT 68.925 1.860 69.815 1.865 ;
        RECT 0.000 1.855 0.075 1.860 ;
    END
  END RWL_30
  PIN RWL_31
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 0.510 0.365 0.680 ;
        RECT 2.395 0.510 2.545 0.680 ;
        RECT 3.115 0.510 3.265 0.680 ;
        RECT 5.295 0.510 5.445 0.680 ;
        RECT 6.015 0.510 6.165 0.680 ;
        RECT 8.195 0.510 8.345 0.680 ;
        RECT 8.915 0.510 9.065 0.680 ;
        RECT 11.095 0.510 11.245 0.680 ;
        RECT 11.815 0.510 11.965 0.680 ;
        RECT 13.995 0.510 14.145 0.680 ;
        RECT 14.715 0.510 14.865 0.680 ;
        RECT 16.895 0.510 17.045 0.680 ;
        RECT 17.615 0.510 17.765 0.680 ;
        RECT 19.795 0.510 19.945 0.680 ;
        RECT 20.515 0.510 20.665 0.680 ;
        RECT 22.695 0.510 22.845 0.680 ;
        RECT 23.415 0.515 23.565 0.685 ;
        RECT 25.595 0.515 25.745 0.685 ;
        RECT 26.315 0.515 26.465 0.685 ;
        RECT 28.495 0.515 28.645 0.685 ;
        RECT 29.215 0.515 29.365 0.685 ;
        RECT 31.395 0.515 31.545 0.685 ;
        RECT 32.115 0.515 32.265 0.685 ;
        RECT 34.295 0.515 34.445 0.685 ;
        RECT 35.015 0.515 35.165 0.685 ;
        RECT 37.195 0.515 37.345 0.685 ;
        RECT 37.915 0.515 38.065 0.685 ;
        RECT 40.095 0.515 40.245 0.685 ;
        RECT 40.815 0.515 40.965 0.685 ;
        RECT 42.995 0.515 43.145 0.685 ;
        RECT 43.715 0.515 43.865 0.685 ;
        RECT 45.895 0.515 46.045 0.685 ;
        RECT 46.615 0.515 46.765 0.685 ;
        RECT 48.795 0.515 48.945 0.685 ;
        RECT 49.515 0.515 49.665 0.685 ;
        RECT 51.695 0.515 51.845 0.685 ;
        RECT 52.415 0.515 52.565 0.685 ;
        RECT 54.595 0.515 54.745 0.685 ;
        RECT 55.315 0.515 55.465 0.685 ;
        RECT 57.495 0.515 57.645 0.685 ;
        RECT 58.215 0.515 58.365 0.685 ;
        RECT 60.395 0.515 60.545 0.685 ;
        RECT 61.115 0.515 61.265 0.685 ;
        RECT 63.295 0.515 63.445 0.685 ;
        RECT 64.015 0.515 64.165 0.685 ;
        RECT 66.195 0.515 66.345 0.685 ;
        RECT 66.915 0.515 67.065 0.685 ;
        RECT 69.095 0.515 69.245 0.685 ;
        RECT 69.815 0.515 69.965 0.685 ;
        RECT 71.995 0.515 72.145 0.685 ;
        RECT 72.715 0.515 72.865 0.685 ;
        RECT 74.895 0.515 75.045 0.685 ;
        RECT 75.615 0.515 75.765 0.685 ;
        RECT 77.795 0.515 77.945 0.685 ;
        RECT 78.515 0.515 78.665 0.685 ;
        RECT 80.695 0.515 80.845 0.685 ;
        RECT 81.415 0.515 81.565 0.685 ;
        RECT 83.595 0.515 83.745 0.685 ;
        RECT 84.315 0.515 84.465 0.685 ;
        RECT 86.495 0.515 86.645 0.685 ;
        RECT 87.215 0.515 87.365 0.685 ;
        RECT 89.395 0.515 89.545 0.685 ;
        RECT 90.115 0.515 90.265 0.685 ;
        RECT 92.295 0.515 92.445 0.685 ;
      LAYER met1 ;
        RECT 23.155 0.680 92.445 0.685 ;
        RECT 0.000 0.515 92.445 0.680 ;
        RECT 0.000 0.510 23.155 0.515 ;
    END
  END RWL_31
  PIN RBL1_16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444800 ;
    PORT
      LAYER li1 ;
        RECT 46.400 42.040 46.475 42.250 ;
        RECT 46.400 40.690 46.475 40.900 ;
        RECT 46.400 39.340 46.475 39.550 ;
        RECT 46.400 37.990 46.475 38.200 ;
        RECT 46.400 36.640 46.475 36.850 ;
        RECT 46.400 35.290 46.475 35.500 ;
        RECT 46.400 33.940 46.475 34.150 ;
        RECT 46.400 32.590 46.475 32.800 ;
        RECT 46.400 31.240 46.475 31.450 ;
        RECT 46.400 29.890 46.475 30.100 ;
        RECT 46.400 28.540 46.475 28.750 ;
        RECT 46.400 27.190 46.475 27.400 ;
        RECT 46.400 25.840 46.475 26.050 ;
        RECT 46.400 24.490 46.475 24.700 ;
        RECT 46.400 23.140 46.475 23.350 ;
        RECT 46.400 21.790 46.475 22.000 ;
        RECT 46.400 20.440 46.475 20.650 ;
        RECT 46.400 19.090 46.475 19.300 ;
        RECT 46.400 17.740 46.475 17.950 ;
        RECT 46.400 16.390 46.475 16.600 ;
        RECT 46.400 15.040 46.475 15.250 ;
        RECT 46.400 13.690 46.475 13.900 ;
        RECT 46.400 12.340 46.475 12.550 ;
        RECT 46.400 10.990 46.475 11.200 ;
        RECT 46.400 9.640 46.475 9.850 ;
        RECT 46.400 8.290 46.475 8.500 ;
        RECT 46.400 6.940 46.475 7.150 ;
        RECT 46.400 5.590 46.475 5.800 ;
        RECT 46.400 4.240 46.475 4.450 ;
        RECT 46.400 2.890 46.475 3.100 ;
        RECT 46.400 1.545 46.475 1.755 ;
        RECT 46.400 0.195 46.475 0.405 ;
    END
  END RBL1_16
  PIN RBL0_16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444800 ;
    PORT
      LAYER li1 ;
        RECT 49.085 42.040 49.160 42.250 ;
        RECT 49.085 40.690 49.160 40.900 ;
        RECT 49.085 39.340 49.160 39.550 ;
        RECT 49.085 37.990 49.160 38.200 ;
        RECT 49.085 36.640 49.160 36.850 ;
        RECT 49.085 35.290 49.160 35.500 ;
        RECT 49.085 33.940 49.160 34.150 ;
        RECT 49.085 32.590 49.160 32.800 ;
        RECT 49.085 31.240 49.160 31.450 ;
        RECT 49.085 29.890 49.160 30.100 ;
        RECT 49.085 28.540 49.160 28.750 ;
        RECT 49.085 27.190 49.160 27.400 ;
        RECT 49.085 25.840 49.160 26.050 ;
        RECT 49.085 24.490 49.160 24.700 ;
        RECT 49.085 23.140 49.160 23.350 ;
        RECT 49.085 21.790 49.160 22.000 ;
        RECT 49.085 20.440 49.160 20.650 ;
        RECT 49.085 19.090 49.160 19.300 ;
        RECT 49.085 17.740 49.160 17.950 ;
        RECT 49.085 16.390 49.160 16.600 ;
        RECT 49.085 15.040 49.160 15.250 ;
        RECT 49.085 13.690 49.160 13.900 ;
        RECT 49.085 12.340 49.160 12.550 ;
        RECT 49.085 10.990 49.160 11.200 ;
        RECT 49.085 9.640 49.160 9.850 ;
        RECT 49.085 8.290 49.160 8.500 ;
        RECT 49.085 6.940 49.160 7.150 ;
        RECT 49.085 5.590 49.160 5.800 ;
        RECT 49.085 4.240 49.160 4.450 ;
        RECT 49.085 2.890 49.160 3.100 ;
        RECT 49.085 1.545 49.160 1.755 ;
        RECT 49.085 0.195 49.160 0.405 ;
    END
  END RBL0_16
  PIN RBL1_17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444800 ;
    PORT
      LAYER li1 ;
        RECT 49.300 42.040 49.375 42.250 ;
        RECT 49.300 40.690 49.375 40.900 ;
        RECT 49.300 39.340 49.375 39.550 ;
        RECT 49.300 37.990 49.375 38.200 ;
        RECT 49.300 36.640 49.375 36.850 ;
        RECT 49.300 35.290 49.375 35.500 ;
        RECT 49.300 33.940 49.375 34.150 ;
        RECT 49.300 32.590 49.375 32.800 ;
        RECT 49.300 31.240 49.375 31.450 ;
        RECT 49.300 29.890 49.375 30.100 ;
        RECT 49.300 28.540 49.375 28.750 ;
        RECT 49.300 27.190 49.375 27.400 ;
        RECT 49.300 25.840 49.375 26.050 ;
        RECT 49.300 24.490 49.375 24.700 ;
        RECT 49.300 23.140 49.375 23.350 ;
        RECT 49.300 21.790 49.375 22.000 ;
        RECT 49.300 20.440 49.375 20.650 ;
        RECT 49.300 19.090 49.375 19.300 ;
        RECT 49.300 17.740 49.375 17.950 ;
        RECT 49.300 16.390 49.375 16.600 ;
        RECT 49.300 15.040 49.375 15.250 ;
        RECT 49.300 13.690 49.375 13.900 ;
        RECT 49.300 12.340 49.375 12.550 ;
        RECT 49.300 10.990 49.375 11.200 ;
        RECT 49.300 9.640 49.375 9.850 ;
        RECT 49.300 8.290 49.375 8.500 ;
        RECT 49.300 6.940 49.375 7.150 ;
        RECT 49.300 5.590 49.375 5.800 ;
        RECT 49.300 4.240 49.375 4.450 ;
        RECT 49.300 2.890 49.375 3.100 ;
        RECT 49.300 1.545 49.375 1.755 ;
        RECT 49.300 0.195 49.375 0.405 ;
    END
  END RBL1_17
  PIN RBL0_17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444800 ;
    PORT
      LAYER li1 ;
        RECT 51.985 42.040 52.060 42.250 ;
        RECT 51.985 40.690 52.060 40.900 ;
        RECT 51.985 39.340 52.060 39.550 ;
        RECT 51.985 37.990 52.060 38.200 ;
        RECT 51.985 36.640 52.060 36.850 ;
        RECT 51.985 35.290 52.060 35.500 ;
        RECT 51.985 33.940 52.060 34.150 ;
        RECT 51.985 32.590 52.060 32.800 ;
        RECT 51.985 31.240 52.060 31.450 ;
        RECT 51.985 29.890 52.060 30.100 ;
        RECT 51.985 28.540 52.060 28.750 ;
        RECT 51.985 27.190 52.060 27.400 ;
        RECT 51.985 25.840 52.060 26.050 ;
        RECT 51.985 24.490 52.060 24.700 ;
        RECT 51.985 23.140 52.060 23.350 ;
        RECT 51.985 21.790 52.060 22.000 ;
        RECT 51.985 20.440 52.060 20.650 ;
        RECT 51.985 19.090 52.060 19.300 ;
        RECT 51.985 17.740 52.060 17.950 ;
        RECT 51.985 16.390 52.060 16.600 ;
        RECT 51.985 15.040 52.060 15.250 ;
        RECT 51.985 13.690 52.060 13.900 ;
        RECT 51.985 12.340 52.060 12.550 ;
        RECT 51.985 10.990 52.060 11.200 ;
        RECT 51.985 9.640 52.060 9.850 ;
        RECT 51.985 8.290 52.060 8.500 ;
        RECT 51.985 6.940 52.060 7.150 ;
        RECT 51.985 5.590 52.060 5.800 ;
        RECT 51.985 4.240 52.060 4.450 ;
        RECT 51.985 2.890 52.060 3.100 ;
        RECT 51.985 1.545 52.060 1.755 ;
        RECT 51.985 0.195 52.060 0.405 ;
    END
  END RBL0_17
  PIN RBL1_18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444800 ;
    PORT
      LAYER li1 ;
        RECT 52.200 42.040 52.275 42.250 ;
        RECT 52.200 40.690 52.275 40.900 ;
        RECT 52.200 39.340 52.275 39.550 ;
        RECT 52.200 37.990 52.275 38.200 ;
        RECT 52.200 36.640 52.275 36.850 ;
        RECT 52.200 35.290 52.275 35.500 ;
        RECT 52.200 33.940 52.275 34.150 ;
        RECT 52.200 32.590 52.275 32.800 ;
        RECT 52.200 31.240 52.275 31.450 ;
        RECT 52.200 29.890 52.275 30.100 ;
        RECT 52.200 28.540 52.275 28.750 ;
        RECT 52.200 27.190 52.275 27.400 ;
        RECT 52.200 25.840 52.275 26.050 ;
        RECT 52.200 24.490 52.275 24.700 ;
        RECT 52.200 23.140 52.275 23.350 ;
        RECT 52.200 21.790 52.275 22.000 ;
        RECT 52.200 20.440 52.275 20.650 ;
        RECT 52.200 19.090 52.275 19.300 ;
        RECT 52.200 17.740 52.275 17.950 ;
        RECT 52.200 16.390 52.275 16.600 ;
        RECT 52.200 15.040 52.275 15.250 ;
        RECT 52.200 13.690 52.275 13.900 ;
        RECT 52.200 12.340 52.275 12.550 ;
        RECT 52.200 10.990 52.275 11.200 ;
        RECT 52.200 9.640 52.275 9.850 ;
        RECT 52.200 8.290 52.275 8.500 ;
        RECT 52.200 6.940 52.275 7.150 ;
        RECT 52.200 5.590 52.275 5.800 ;
        RECT 52.200 4.240 52.275 4.450 ;
        RECT 52.200 2.890 52.275 3.100 ;
        RECT 52.200 1.545 52.275 1.755 ;
        RECT 52.200 0.195 52.275 0.405 ;
    END
  END RBL1_18
  PIN RBL0_18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444800 ;
    PORT
      LAYER li1 ;
        RECT 54.885 42.040 54.960 42.250 ;
        RECT 54.885 40.690 54.960 40.900 ;
        RECT 54.885 39.340 54.960 39.550 ;
        RECT 54.885 37.990 54.960 38.200 ;
        RECT 54.885 36.640 54.960 36.850 ;
        RECT 54.885 35.290 54.960 35.500 ;
        RECT 54.885 33.940 54.960 34.150 ;
        RECT 54.885 32.590 54.960 32.800 ;
        RECT 54.885 31.240 54.960 31.450 ;
        RECT 54.885 29.890 54.960 30.100 ;
        RECT 54.885 28.540 54.960 28.750 ;
        RECT 54.885 27.190 54.960 27.400 ;
        RECT 54.885 25.840 54.960 26.050 ;
        RECT 54.885 24.490 54.960 24.700 ;
        RECT 54.885 23.140 54.960 23.350 ;
        RECT 54.885 21.790 54.960 22.000 ;
        RECT 54.885 20.440 54.960 20.650 ;
        RECT 54.885 19.090 54.960 19.300 ;
        RECT 54.885 17.740 54.960 17.950 ;
        RECT 54.885 16.390 54.960 16.600 ;
        RECT 54.885 15.040 54.960 15.250 ;
        RECT 54.885 13.690 54.960 13.900 ;
        RECT 54.885 12.340 54.960 12.550 ;
        RECT 54.885 10.990 54.960 11.200 ;
        RECT 54.885 9.640 54.960 9.850 ;
        RECT 54.885 8.290 54.960 8.500 ;
        RECT 54.885 6.940 54.960 7.150 ;
        RECT 54.885 5.590 54.960 5.800 ;
        RECT 54.885 4.240 54.960 4.450 ;
        RECT 54.885 2.890 54.960 3.100 ;
        RECT 54.885 1.545 54.960 1.755 ;
        RECT 54.885 0.195 54.960 0.405 ;
    END
  END RBL0_18
  PIN RBL1_19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444800 ;
    PORT
      LAYER li1 ;
        RECT 55.100 42.040 55.175 42.250 ;
        RECT 55.100 40.690 55.175 40.900 ;
        RECT 55.100 39.340 55.175 39.550 ;
        RECT 55.100 37.990 55.175 38.200 ;
        RECT 55.100 36.640 55.175 36.850 ;
        RECT 55.100 35.290 55.175 35.500 ;
        RECT 55.100 33.940 55.175 34.150 ;
        RECT 55.100 32.590 55.175 32.800 ;
        RECT 55.100 31.240 55.175 31.450 ;
        RECT 55.100 29.890 55.175 30.100 ;
        RECT 55.100 28.540 55.175 28.750 ;
        RECT 55.100 27.190 55.175 27.400 ;
        RECT 55.100 25.840 55.175 26.050 ;
        RECT 55.100 24.490 55.175 24.700 ;
        RECT 55.100 23.140 55.175 23.350 ;
        RECT 55.100 21.790 55.175 22.000 ;
        RECT 55.100 20.440 55.175 20.650 ;
        RECT 55.100 19.090 55.175 19.300 ;
        RECT 55.100 17.740 55.175 17.950 ;
        RECT 55.100 16.390 55.175 16.600 ;
        RECT 55.100 15.040 55.175 15.250 ;
        RECT 55.100 13.690 55.175 13.900 ;
        RECT 55.100 12.340 55.175 12.550 ;
        RECT 55.100 10.990 55.175 11.200 ;
        RECT 55.100 9.640 55.175 9.850 ;
        RECT 55.100 8.290 55.175 8.500 ;
        RECT 55.100 6.940 55.175 7.150 ;
        RECT 55.100 5.590 55.175 5.800 ;
        RECT 55.100 4.240 55.175 4.450 ;
        RECT 55.100 2.890 55.175 3.100 ;
        RECT 55.100 1.545 55.175 1.755 ;
        RECT 55.100 0.195 55.175 0.405 ;
    END
  END RBL1_19
  PIN RBL0_19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444800 ;
    PORT
      LAYER li1 ;
        RECT 57.785 42.040 57.860 42.250 ;
        RECT 57.785 40.690 57.860 40.900 ;
        RECT 57.785 39.340 57.860 39.550 ;
        RECT 57.785 37.990 57.860 38.200 ;
        RECT 57.785 36.640 57.860 36.850 ;
        RECT 57.785 35.290 57.860 35.500 ;
        RECT 57.785 33.940 57.860 34.150 ;
        RECT 57.785 32.590 57.860 32.800 ;
        RECT 57.785 31.240 57.860 31.450 ;
        RECT 57.785 29.890 57.860 30.100 ;
        RECT 57.785 28.540 57.860 28.750 ;
        RECT 57.785 27.190 57.860 27.400 ;
        RECT 57.785 25.840 57.860 26.050 ;
        RECT 57.785 24.490 57.860 24.700 ;
        RECT 57.785 23.140 57.860 23.350 ;
        RECT 57.785 21.790 57.860 22.000 ;
        RECT 57.785 20.440 57.860 20.650 ;
        RECT 57.785 19.090 57.860 19.300 ;
        RECT 57.785 17.740 57.860 17.950 ;
        RECT 57.785 16.390 57.860 16.600 ;
        RECT 57.785 15.040 57.860 15.250 ;
        RECT 57.785 13.690 57.860 13.900 ;
        RECT 57.785 12.340 57.860 12.550 ;
        RECT 57.785 10.990 57.860 11.200 ;
        RECT 57.785 9.640 57.860 9.850 ;
        RECT 57.785 8.290 57.860 8.500 ;
        RECT 57.785 6.940 57.860 7.150 ;
        RECT 57.785 5.590 57.860 5.800 ;
        RECT 57.785 4.240 57.860 4.450 ;
        RECT 57.785 2.890 57.860 3.100 ;
        RECT 57.785 1.545 57.860 1.755 ;
        RECT 57.785 0.195 57.860 0.405 ;
    END
  END RBL0_19
  PIN RBL1_20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444800 ;
    PORT
      LAYER li1 ;
        RECT 58.000 42.040 58.075 42.250 ;
        RECT 58.000 40.690 58.075 40.900 ;
        RECT 58.000 39.340 58.075 39.550 ;
        RECT 58.000 37.990 58.075 38.200 ;
        RECT 58.000 36.640 58.075 36.850 ;
        RECT 58.000 35.290 58.075 35.500 ;
        RECT 58.000 33.940 58.075 34.150 ;
        RECT 58.000 32.590 58.075 32.800 ;
        RECT 58.000 31.240 58.075 31.450 ;
        RECT 58.000 29.890 58.075 30.100 ;
        RECT 58.000 28.540 58.075 28.750 ;
        RECT 58.000 27.190 58.075 27.400 ;
        RECT 58.000 25.840 58.075 26.050 ;
        RECT 58.000 24.490 58.075 24.700 ;
        RECT 58.000 23.140 58.075 23.350 ;
        RECT 58.000 21.790 58.075 22.000 ;
        RECT 58.000 20.440 58.075 20.650 ;
        RECT 58.000 19.090 58.075 19.300 ;
        RECT 58.000 17.740 58.075 17.950 ;
        RECT 58.000 16.390 58.075 16.600 ;
        RECT 58.000 15.040 58.075 15.250 ;
        RECT 58.000 13.690 58.075 13.900 ;
        RECT 58.000 12.340 58.075 12.550 ;
        RECT 58.000 10.990 58.075 11.200 ;
        RECT 58.000 9.640 58.075 9.850 ;
        RECT 58.000 8.290 58.075 8.500 ;
        RECT 58.000 6.940 58.075 7.150 ;
        RECT 58.000 5.590 58.075 5.800 ;
        RECT 58.000 4.240 58.075 4.450 ;
        RECT 58.000 2.890 58.075 3.100 ;
        RECT 58.000 1.545 58.075 1.755 ;
        RECT 58.000 0.195 58.075 0.405 ;
    END
  END RBL1_20
  PIN RBL0_20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444800 ;
    PORT
      LAYER li1 ;
        RECT 60.685 42.040 60.760 42.250 ;
        RECT 60.685 40.690 60.760 40.900 ;
        RECT 60.685 39.340 60.760 39.550 ;
        RECT 60.685 37.990 60.760 38.200 ;
        RECT 60.685 36.640 60.760 36.850 ;
        RECT 60.685 35.290 60.760 35.500 ;
        RECT 60.685 33.940 60.760 34.150 ;
        RECT 60.685 32.590 60.760 32.800 ;
        RECT 60.685 31.240 60.760 31.450 ;
        RECT 60.685 29.890 60.760 30.100 ;
        RECT 60.685 28.540 60.760 28.750 ;
        RECT 60.685 27.190 60.760 27.400 ;
        RECT 60.685 25.840 60.760 26.050 ;
        RECT 60.685 24.490 60.760 24.700 ;
        RECT 60.685 23.140 60.760 23.350 ;
        RECT 60.685 21.790 60.760 22.000 ;
        RECT 60.685 20.440 60.760 20.650 ;
        RECT 60.685 19.090 60.760 19.300 ;
        RECT 60.685 17.740 60.760 17.950 ;
        RECT 60.685 16.390 60.760 16.600 ;
        RECT 60.685 15.040 60.760 15.250 ;
        RECT 60.685 13.690 60.760 13.900 ;
        RECT 60.685 12.340 60.760 12.550 ;
        RECT 60.685 10.990 60.760 11.200 ;
        RECT 60.685 9.640 60.760 9.850 ;
        RECT 60.685 8.290 60.760 8.500 ;
        RECT 60.685 6.940 60.760 7.150 ;
        RECT 60.685 5.590 60.760 5.800 ;
        RECT 60.685 4.240 60.760 4.450 ;
        RECT 60.685 2.890 60.760 3.100 ;
        RECT 60.685 1.545 60.760 1.755 ;
        RECT 60.685 0.195 60.760 0.405 ;
    END
  END RBL0_20
  PIN RBL1_21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444800 ;
    PORT
      LAYER li1 ;
        RECT 60.900 42.040 60.975 42.250 ;
        RECT 60.900 40.690 60.975 40.900 ;
        RECT 60.900 39.340 60.975 39.550 ;
        RECT 60.900 37.990 60.975 38.200 ;
        RECT 60.900 36.640 60.975 36.850 ;
        RECT 60.900 35.290 60.975 35.500 ;
        RECT 60.900 33.940 60.975 34.150 ;
        RECT 60.900 32.590 60.975 32.800 ;
        RECT 60.900 31.240 60.975 31.450 ;
        RECT 60.900 29.890 60.975 30.100 ;
        RECT 60.900 28.540 60.975 28.750 ;
        RECT 60.900 27.190 60.975 27.400 ;
        RECT 60.900 25.840 60.975 26.050 ;
        RECT 60.900 24.490 60.975 24.700 ;
        RECT 60.900 23.140 60.975 23.350 ;
        RECT 60.900 21.790 60.975 22.000 ;
        RECT 60.900 20.440 60.975 20.650 ;
        RECT 60.900 19.090 60.975 19.300 ;
        RECT 60.900 17.740 60.975 17.950 ;
        RECT 60.900 16.390 60.975 16.600 ;
        RECT 60.900 15.040 60.975 15.250 ;
        RECT 60.900 13.690 60.975 13.900 ;
        RECT 60.900 12.340 60.975 12.550 ;
        RECT 60.900 10.990 60.975 11.200 ;
        RECT 60.900 9.640 60.975 9.850 ;
        RECT 60.900 8.290 60.975 8.500 ;
        RECT 60.900 6.940 60.975 7.150 ;
        RECT 60.900 5.590 60.975 5.800 ;
        RECT 60.900 4.240 60.975 4.450 ;
        RECT 60.900 2.890 60.975 3.100 ;
        RECT 60.900 1.545 60.975 1.755 ;
        RECT 60.900 0.195 60.975 0.405 ;
    END
  END RBL1_21
  PIN RBL0_21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444800 ;
    PORT
      LAYER li1 ;
        RECT 63.585 42.040 63.660 42.250 ;
        RECT 63.585 40.690 63.660 40.900 ;
        RECT 63.585 39.340 63.660 39.550 ;
        RECT 63.585 37.990 63.660 38.200 ;
        RECT 63.585 36.640 63.660 36.850 ;
        RECT 63.585 35.290 63.660 35.500 ;
        RECT 63.585 33.940 63.660 34.150 ;
        RECT 63.585 32.590 63.660 32.800 ;
        RECT 63.585 31.240 63.660 31.450 ;
        RECT 63.585 29.890 63.660 30.100 ;
        RECT 63.585 28.540 63.660 28.750 ;
        RECT 63.585 27.190 63.660 27.400 ;
        RECT 63.585 25.840 63.660 26.050 ;
        RECT 63.585 24.490 63.660 24.700 ;
        RECT 63.585 23.140 63.660 23.350 ;
        RECT 63.585 21.790 63.660 22.000 ;
        RECT 63.585 20.440 63.660 20.650 ;
        RECT 63.585 19.090 63.660 19.300 ;
        RECT 63.585 17.740 63.660 17.950 ;
        RECT 63.585 16.390 63.660 16.600 ;
        RECT 63.585 15.040 63.660 15.250 ;
        RECT 63.585 13.690 63.660 13.900 ;
        RECT 63.585 12.340 63.660 12.550 ;
        RECT 63.585 10.990 63.660 11.200 ;
        RECT 63.585 9.640 63.660 9.850 ;
        RECT 63.585 8.290 63.660 8.500 ;
        RECT 63.585 6.940 63.660 7.150 ;
        RECT 63.585 5.590 63.660 5.800 ;
        RECT 63.585 4.240 63.660 4.450 ;
        RECT 63.585 2.890 63.660 3.100 ;
        RECT 63.585 1.545 63.660 1.755 ;
        RECT 63.585 0.195 63.660 0.405 ;
    END
  END RBL0_21
  PIN RBL1_22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444800 ;
    PORT
      LAYER li1 ;
        RECT 63.800 42.040 63.875 42.250 ;
        RECT 63.800 40.690 63.875 40.900 ;
        RECT 63.800 39.340 63.875 39.550 ;
        RECT 63.800 37.990 63.875 38.200 ;
        RECT 63.800 36.640 63.875 36.850 ;
        RECT 63.800 35.290 63.875 35.500 ;
        RECT 63.800 33.940 63.875 34.150 ;
        RECT 63.800 32.590 63.875 32.800 ;
        RECT 63.800 31.240 63.875 31.450 ;
        RECT 63.800 29.890 63.875 30.100 ;
        RECT 63.800 28.540 63.875 28.750 ;
        RECT 63.800 27.190 63.875 27.400 ;
        RECT 63.800 25.840 63.875 26.050 ;
        RECT 63.800 24.490 63.875 24.700 ;
        RECT 63.800 23.140 63.875 23.350 ;
        RECT 63.800 21.790 63.875 22.000 ;
        RECT 63.800 20.440 63.875 20.650 ;
        RECT 63.800 19.090 63.875 19.300 ;
        RECT 63.800 17.740 63.875 17.950 ;
        RECT 63.800 16.390 63.875 16.600 ;
        RECT 63.800 15.040 63.875 15.250 ;
        RECT 63.800 13.690 63.875 13.900 ;
        RECT 63.800 12.340 63.875 12.550 ;
        RECT 63.800 10.990 63.875 11.200 ;
        RECT 63.800 9.640 63.875 9.850 ;
        RECT 63.800 8.290 63.875 8.500 ;
        RECT 63.800 6.940 63.875 7.150 ;
        RECT 63.800 5.590 63.875 5.800 ;
        RECT 63.800 4.240 63.875 4.450 ;
        RECT 63.800 2.890 63.875 3.100 ;
        RECT 63.800 1.545 63.875 1.755 ;
        RECT 63.800 0.195 63.875 0.405 ;
    END
  END RBL1_22
  PIN RBL0_22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444800 ;
    PORT
      LAYER li1 ;
        RECT 66.485 42.040 66.560 42.250 ;
        RECT 66.485 40.690 66.560 40.900 ;
        RECT 66.485 39.340 66.560 39.550 ;
        RECT 66.485 37.990 66.560 38.200 ;
        RECT 66.485 36.640 66.560 36.850 ;
        RECT 66.485 35.290 66.560 35.500 ;
        RECT 66.485 33.940 66.560 34.150 ;
        RECT 66.485 32.590 66.560 32.800 ;
        RECT 66.485 31.240 66.560 31.450 ;
        RECT 66.485 29.890 66.560 30.100 ;
        RECT 66.485 28.540 66.560 28.750 ;
        RECT 66.485 27.190 66.560 27.400 ;
        RECT 66.485 25.840 66.560 26.050 ;
        RECT 66.485 24.490 66.560 24.700 ;
        RECT 66.485 23.140 66.560 23.350 ;
        RECT 66.485 21.790 66.560 22.000 ;
        RECT 66.485 20.440 66.560 20.650 ;
        RECT 66.485 19.090 66.560 19.300 ;
        RECT 66.485 17.740 66.560 17.950 ;
        RECT 66.485 16.390 66.560 16.600 ;
        RECT 66.485 15.040 66.560 15.250 ;
        RECT 66.485 13.690 66.560 13.900 ;
        RECT 66.485 12.340 66.560 12.550 ;
        RECT 66.485 10.990 66.560 11.200 ;
        RECT 66.485 9.640 66.560 9.850 ;
        RECT 66.485 8.290 66.560 8.500 ;
        RECT 66.485 6.940 66.560 7.150 ;
        RECT 66.485 5.590 66.560 5.800 ;
        RECT 66.485 4.240 66.560 4.450 ;
        RECT 66.485 2.890 66.560 3.100 ;
        RECT 66.485 1.545 66.560 1.755 ;
        RECT 66.485 0.195 66.560 0.405 ;
    END
  END RBL0_22
  PIN RBL1_23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444800 ;
    PORT
      LAYER li1 ;
        RECT 66.700 42.040 66.775 42.250 ;
        RECT 66.700 40.690 66.775 40.900 ;
        RECT 66.700 39.340 66.775 39.550 ;
        RECT 66.700 37.990 66.775 38.200 ;
        RECT 66.700 36.640 66.775 36.850 ;
        RECT 66.700 35.290 66.775 35.500 ;
        RECT 66.700 33.940 66.775 34.150 ;
        RECT 66.700 32.590 66.775 32.800 ;
        RECT 66.700 31.240 66.775 31.450 ;
        RECT 66.700 29.890 66.775 30.100 ;
        RECT 66.700 28.540 66.775 28.750 ;
        RECT 66.700 27.190 66.775 27.400 ;
        RECT 66.700 25.840 66.775 26.050 ;
        RECT 66.700 24.490 66.775 24.700 ;
        RECT 66.700 23.140 66.775 23.350 ;
        RECT 66.700 21.790 66.775 22.000 ;
        RECT 66.700 20.440 66.775 20.650 ;
        RECT 66.700 19.090 66.775 19.300 ;
        RECT 66.700 17.740 66.775 17.950 ;
        RECT 66.700 16.390 66.775 16.600 ;
        RECT 66.700 15.040 66.775 15.250 ;
        RECT 66.700 13.690 66.775 13.900 ;
        RECT 66.700 12.340 66.775 12.550 ;
        RECT 66.700 10.990 66.775 11.200 ;
        RECT 66.700 9.640 66.775 9.850 ;
        RECT 66.700 8.290 66.775 8.500 ;
        RECT 66.700 6.940 66.775 7.150 ;
        RECT 66.700 5.590 66.775 5.800 ;
        RECT 66.700 4.240 66.775 4.450 ;
        RECT 66.700 2.890 66.775 3.100 ;
        RECT 66.700 1.545 66.775 1.755 ;
        RECT 66.700 0.195 66.775 0.405 ;
    END
  END RBL1_23
  PIN RBL0_23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444800 ;
    PORT
      LAYER li1 ;
        RECT 69.385 42.040 69.460 42.250 ;
        RECT 69.385 40.690 69.460 40.900 ;
        RECT 69.385 39.340 69.460 39.550 ;
        RECT 69.385 37.990 69.460 38.200 ;
        RECT 69.385 36.640 69.460 36.850 ;
        RECT 69.385 35.290 69.460 35.500 ;
        RECT 69.385 33.940 69.460 34.150 ;
        RECT 69.385 32.590 69.460 32.800 ;
        RECT 69.385 31.240 69.460 31.450 ;
        RECT 69.385 29.890 69.460 30.100 ;
        RECT 69.385 28.540 69.460 28.750 ;
        RECT 69.385 27.190 69.460 27.400 ;
        RECT 69.385 25.840 69.460 26.050 ;
        RECT 69.385 24.490 69.460 24.700 ;
        RECT 69.385 23.140 69.460 23.350 ;
        RECT 69.385 21.790 69.460 22.000 ;
        RECT 69.385 20.440 69.460 20.650 ;
        RECT 69.385 19.090 69.460 19.300 ;
        RECT 69.385 17.740 69.460 17.950 ;
        RECT 69.385 16.390 69.460 16.600 ;
        RECT 69.385 15.040 69.460 15.250 ;
        RECT 69.385 13.690 69.460 13.900 ;
        RECT 69.385 12.340 69.460 12.550 ;
        RECT 69.385 10.990 69.460 11.200 ;
        RECT 69.385 9.640 69.460 9.850 ;
        RECT 69.385 8.290 69.460 8.500 ;
        RECT 69.385 6.940 69.460 7.150 ;
        RECT 69.385 5.590 69.460 5.800 ;
        RECT 69.385 4.240 69.460 4.450 ;
        RECT 69.385 2.890 69.460 3.100 ;
        RECT 69.385 1.545 69.460 1.755 ;
        RECT 69.385 0.195 69.460 0.405 ;
    END
  END RBL0_23
  PIN RBL1_24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.444800 ;
    PORT
      LAYER li1 ;
        RECT 69.600 42.040 69.675 42.250 ;
        RECT 69.600 40.690 69.675 40.900 ;
        RECT 69.600 39.340 69.675 39.550 ;
        RECT 69.600 37.990 69.675 38.200 ;
        RECT 69.600 36.640 69.675 36.850 ;
        RECT 69.600 35.290 69.675 35.500 ;
        RECT 69.600 33.940 69.675 34.150 ;
        RECT 69.600 32.590 69.675 32.800 ;
        RECT 69.600 31.240 69.675 31.450 ;
        RECT 69.600 29.890 69.675 30.100 ;
        RECT 69.600 28.540 69.675 28.750 ;
        RECT 69.600 27.190 69.675 27.400 ;
        RECT 69.600 25.840 69.675 26.050 ;
        RECT 69.600 24.490 69.675 24.700 ;
        RECT 69.600 23.140 69.675 23.350 ;
        RECT 69.600 21.790 69.675 22.000 ;
        RECT 69.600 20.440 69.675 20.650 ;
        RECT 69.600 19.090 69.675 19.300 ;
        RECT 69.600 17.740 69.675 17.950 ;
        RECT 69.600 16.390 69.675 16.600 ;
        RECT 69.600 15.040 69.675 15.250 ;
        RECT 69.600 13.690 69.675 13.900 ;
        RECT 69.600 12.340 69.675 12.550 ;
        RECT 69.600 10.990 69.675 11.200 ;
        RECT 69.600 9.640 69.675 9.850 ;
        RECT 69.600 8.290 69.675 8.500 ;
        RECT 69.600 6.940 69.675 7.150 ;
        RECT 69.600 5.590 69.675 5.800 ;
        RECT 69.600 4.240 69.675 4.450 ;
        RECT 69.600 2.890 69.675 3.100 ;
        RECT 69.600 1.545 69.675 1.755 ;
        RECT 69.600 0.195 69.675 0.405 ;
    END
  END RBL1_24
  PIN RBL0_24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.445175 ;
    PORT
      LAYER li1 ;
        RECT 72.285 42.040 72.360 42.250 ;
        RECT 72.285 40.690 72.360 40.900 ;
        RECT 72.285 39.340 72.360 39.550 ;
        RECT 72.285 37.990 72.360 38.200 ;
        RECT 72.285 36.640 72.360 36.850 ;
        RECT 72.285 35.290 72.360 35.500 ;
        RECT 72.285 33.940 72.360 34.150 ;
        RECT 72.285 32.590 72.360 32.800 ;
        RECT 72.285 31.240 72.360 31.450 ;
        RECT 72.285 29.890 72.360 30.100 ;
        RECT 72.285 28.540 72.360 28.750 ;
        RECT 72.285 27.190 72.360 27.400 ;
        RECT 72.285 25.840 72.360 26.050 ;
        RECT 72.285 24.490 72.360 24.700 ;
        RECT 72.285 23.140 72.360 23.350 ;
        RECT 72.285 21.790 72.360 22.000 ;
        RECT 72.285 20.440 72.360 20.650 ;
        RECT 72.285 19.090 72.360 19.300 ;
        RECT 72.285 17.740 72.360 17.950 ;
        RECT 72.285 16.390 72.360 16.600 ;
        RECT 72.285 15.040 72.360 15.250 ;
        RECT 72.285 13.690 72.360 13.900 ;
        RECT 72.285 12.340 72.360 12.550 ;
        RECT 72.285 10.990 72.360 11.200 ;
        RECT 72.285 9.640 72.360 9.850 ;
        RECT 72.285 8.290 72.360 8.500 ;
        RECT 72.285 6.940 72.360 7.150 ;
        RECT 72.285 5.590 72.360 5.800 ;
        RECT 72.285 4.240 72.360 4.450 ;
        RECT 72.285 2.890 72.360 3.100 ;
        RECT 72.285 1.545 72.360 1.755 ;
        RECT 72.285 0.190 72.360 0.405 ;
    END
  END RBL0_24
  PIN RBL1_25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.445175 ;
    PORT
      LAYER li1 ;
        RECT 72.500 42.040 72.575 42.250 ;
        RECT 72.500 40.690 72.575 40.900 ;
        RECT 72.500 39.340 72.575 39.550 ;
        RECT 72.500 37.990 72.575 38.200 ;
        RECT 72.500 36.640 72.575 36.850 ;
        RECT 72.500 35.290 72.575 35.500 ;
        RECT 72.500 33.940 72.575 34.150 ;
        RECT 72.500 32.590 72.575 32.800 ;
        RECT 72.500 31.240 72.575 31.450 ;
        RECT 72.500 29.890 72.575 30.100 ;
        RECT 72.500 28.540 72.575 28.750 ;
        RECT 72.500 27.190 72.575 27.400 ;
        RECT 72.500 25.840 72.575 26.050 ;
        RECT 72.500 24.490 72.575 24.700 ;
        RECT 72.500 23.140 72.575 23.350 ;
        RECT 72.500 21.790 72.575 22.000 ;
        RECT 72.500 20.440 72.575 20.650 ;
        RECT 72.500 19.090 72.575 19.300 ;
        RECT 72.500 17.740 72.575 17.950 ;
        RECT 72.500 16.390 72.575 16.600 ;
        RECT 72.500 15.040 72.575 15.250 ;
        RECT 72.500 13.690 72.575 13.900 ;
        RECT 72.500 12.340 72.575 12.550 ;
        RECT 72.500 10.990 72.575 11.200 ;
        RECT 72.500 9.640 72.575 9.850 ;
        RECT 72.500 8.290 72.575 8.500 ;
        RECT 72.500 6.940 72.575 7.150 ;
        RECT 72.500 5.590 72.575 5.800 ;
        RECT 72.500 4.240 72.575 4.450 ;
        RECT 72.500 2.890 72.575 3.100 ;
        RECT 72.500 1.545 72.575 1.755 ;
        RECT 72.500 0.190 72.575 0.405 ;
    END
  END RBL1_25
  PIN RBL0_25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.445175 ;
    PORT
      LAYER li1 ;
        RECT 75.185 42.040 75.260 42.250 ;
        RECT 75.185 40.690 75.260 40.900 ;
        RECT 75.185 39.340 75.260 39.550 ;
        RECT 75.185 37.990 75.260 38.200 ;
        RECT 75.185 36.640 75.260 36.850 ;
        RECT 75.185 35.290 75.260 35.500 ;
        RECT 75.185 33.940 75.260 34.150 ;
        RECT 75.185 32.590 75.260 32.800 ;
        RECT 75.185 31.240 75.260 31.450 ;
        RECT 75.185 29.890 75.260 30.100 ;
        RECT 75.185 28.540 75.260 28.750 ;
        RECT 75.185 27.190 75.260 27.400 ;
        RECT 75.185 25.840 75.260 26.050 ;
        RECT 75.185 24.490 75.260 24.700 ;
        RECT 75.185 23.140 75.260 23.350 ;
        RECT 75.185 21.790 75.260 22.000 ;
        RECT 75.185 20.440 75.260 20.650 ;
        RECT 75.185 19.090 75.260 19.300 ;
        RECT 75.185 17.740 75.260 17.950 ;
        RECT 75.185 16.390 75.260 16.600 ;
        RECT 75.185 15.040 75.260 15.250 ;
        RECT 75.185 13.690 75.260 13.900 ;
        RECT 75.185 12.340 75.260 12.550 ;
        RECT 75.185 10.990 75.260 11.200 ;
        RECT 75.185 9.640 75.260 9.850 ;
        RECT 75.185 8.290 75.260 8.500 ;
        RECT 75.185 6.940 75.260 7.150 ;
        RECT 75.185 5.590 75.260 5.800 ;
        RECT 75.185 4.240 75.260 4.450 ;
        RECT 75.185 2.890 75.260 3.100 ;
        RECT 75.185 1.545 75.260 1.755 ;
        RECT 75.185 0.190 75.260 0.405 ;
    END
  END RBL0_25
  PIN RBL1_26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.445175 ;
    PORT
      LAYER li1 ;
        RECT 75.400 42.040 75.475 42.250 ;
        RECT 75.400 40.690 75.475 40.900 ;
        RECT 75.400 39.340 75.475 39.550 ;
        RECT 75.400 37.990 75.475 38.200 ;
        RECT 75.400 36.640 75.475 36.850 ;
        RECT 75.400 35.290 75.475 35.500 ;
        RECT 75.400 33.940 75.475 34.150 ;
        RECT 75.400 32.590 75.475 32.800 ;
        RECT 75.400 31.240 75.475 31.450 ;
        RECT 75.400 29.890 75.475 30.100 ;
        RECT 75.400 28.540 75.475 28.750 ;
        RECT 75.400 27.190 75.475 27.400 ;
        RECT 75.400 25.840 75.475 26.050 ;
        RECT 75.400 24.490 75.475 24.700 ;
        RECT 75.400 23.140 75.475 23.350 ;
        RECT 75.400 21.790 75.475 22.000 ;
        RECT 75.400 20.440 75.475 20.650 ;
        RECT 75.400 19.090 75.475 19.300 ;
        RECT 75.400 17.740 75.475 17.950 ;
        RECT 75.400 16.390 75.475 16.600 ;
        RECT 75.400 15.040 75.475 15.250 ;
        RECT 75.400 13.690 75.475 13.900 ;
        RECT 75.400 12.340 75.475 12.550 ;
        RECT 75.400 10.990 75.475 11.200 ;
        RECT 75.400 9.640 75.475 9.850 ;
        RECT 75.400 8.290 75.475 8.500 ;
        RECT 75.400 6.940 75.475 7.150 ;
        RECT 75.400 5.590 75.475 5.800 ;
        RECT 75.400 4.240 75.475 4.450 ;
        RECT 75.400 2.890 75.475 3.100 ;
        RECT 75.400 1.545 75.475 1.755 ;
        RECT 75.400 0.190 75.475 0.405 ;
    END
  END RBL1_26
  PIN RBL0_26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.445175 ;
    PORT
      LAYER li1 ;
        RECT 78.085 42.040 78.160 42.250 ;
        RECT 78.085 40.690 78.160 40.900 ;
        RECT 78.085 39.340 78.160 39.550 ;
        RECT 78.085 37.990 78.160 38.200 ;
        RECT 78.085 36.640 78.160 36.850 ;
        RECT 78.085 35.290 78.160 35.500 ;
        RECT 78.085 33.940 78.160 34.150 ;
        RECT 78.085 32.590 78.160 32.800 ;
        RECT 78.085 31.240 78.160 31.450 ;
        RECT 78.085 29.890 78.160 30.100 ;
        RECT 78.085 28.540 78.160 28.750 ;
        RECT 78.085 27.190 78.160 27.400 ;
        RECT 78.085 25.840 78.160 26.050 ;
        RECT 78.085 24.490 78.160 24.700 ;
        RECT 78.085 23.140 78.160 23.350 ;
        RECT 78.085 21.790 78.160 22.000 ;
        RECT 78.085 20.440 78.160 20.650 ;
        RECT 78.085 19.090 78.160 19.300 ;
        RECT 78.085 17.740 78.160 17.950 ;
        RECT 78.085 16.390 78.160 16.600 ;
        RECT 78.085 15.040 78.160 15.250 ;
        RECT 78.085 13.690 78.160 13.900 ;
        RECT 78.085 12.340 78.160 12.550 ;
        RECT 78.085 10.990 78.160 11.200 ;
        RECT 78.085 9.640 78.160 9.850 ;
        RECT 78.085 8.290 78.160 8.500 ;
        RECT 78.085 6.940 78.160 7.150 ;
        RECT 78.085 5.590 78.160 5.800 ;
        RECT 78.085 4.240 78.160 4.450 ;
        RECT 78.085 2.890 78.160 3.100 ;
        RECT 78.085 1.545 78.160 1.755 ;
        RECT 78.085 0.190 78.160 0.405 ;
    END
  END RBL0_26
  PIN RBL1_27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.445175 ;
    PORT
      LAYER li1 ;
        RECT 78.300 42.040 78.375 42.250 ;
        RECT 78.300 40.690 78.375 40.900 ;
        RECT 78.300 39.340 78.375 39.550 ;
        RECT 78.300 37.990 78.375 38.200 ;
        RECT 78.300 36.640 78.375 36.850 ;
        RECT 78.300 35.290 78.375 35.500 ;
        RECT 78.300 33.940 78.375 34.150 ;
        RECT 78.300 32.590 78.375 32.800 ;
        RECT 78.300 31.240 78.375 31.450 ;
        RECT 78.300 29.890 78.375 30.100 ;
        RECT 78.300 28.540 78.375 28.750 ;
        RECT 78.300 27.190 78.375 27.400 ;
        RECT 78.300 25.840 78.375 26.050 ;
        RECT 78.300 24.490 78.375 24.700 ;
        RECT 78.300 23.140 78.375 23.350 ;
        RECT 78.300 21.790 78.375 22.000 ;
        RECT 78.300 20.440 78.375 20.650 ;
        RECT 78.300 19.090 78.375 19.300 ;
        RECT 78.300 17.740 78.375 17.950 ;
        RECT 78.300 16.390 78.375 16.600 ;
        RECT 78.300 15.040 78.375 15.250 ;
        RECT 78.300 13.690 78.375 13.900 ;
        RECT 78.300 12.340 78.375 12.550 ;
        RECT 78.300 10.990 78.375 11.200 ;
        RECT 78.300 9.640 78.375 9.850 ;
        RECT 78.300 8.290 78.375 8.500 ;
        RECT 78.300 6.940 78.375 7.150 ;
        RECT 78.300 5.590 78.375 5.800 ;
        RECT 78.300 4.240 78.375 4.450 ;
        RECT 78.300 2.890 78.375 3.100 ;
        RECT 78.300 1.545 78.375 1.755 ;
        RECT 78.300 0.190 78.375 0.405 ;
    END
  END RBL1_27
  PIN RBL0_27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.445175 ;
    PORT
      LAYER li1 ;
        RECT 80.985 42.040 81.060 42.250 ;
        RECT 80.985 40.690 81.060 40.900 ;
        RECT 80.985 39.340 81.060 39.550 ;
        RECT 80.985 37.990 81.060 38.200 ;
        RECT 80.985 36.640 81.060 36.850 ;
        RECT 80.985 35.290 81.060 35.500 ;
        RECT 80.985 33.940 81.060 34.150 ;
        RECT 80.985 32.590 81.060 32.800 ;
        RECT 80.985 31.240 81.060 31.450 ;
        RECT 80.985 29.890 81.060 30.100 ;
        RECT 80.985 28.540 81.060 28.750 ;
        RECT 80.985 27.190 81.060 27.400 ;
        RECT 80.985 25.840 81.060 26.050 ;
        RECT 80.985 24.490 81.060 24.700 ;
        RECT 80.985 23.140 81.060 23.350 ;
        RECT 80.985 21.790 81.060 22.000 ;
        RECT 80.985 20.440 81.060 20.650 ;
        RECT 80.985 19.090 81.060 19.300 ;
        RECT 80.985 17.740 81.060 17.950 ;
        RECT 80.985 16.390 81.060 16.600 ;
        RECT 80.985 15.040 81.060 15.250 ;
        RECT 80.985 13.690 81.060 13.900 ;
        RECT 80.985 12.340 81.060 12.550 ;
        RECT 80.985 10.990 81.060 11.200 ;
        RECT 80.985 9.640 81.060 9.850 ;
        RECT 80.985 8.290 81.060 8.500 ;
        RECT 80.985 6.940 81.060 7.150 ;
        RECT 80.985 5.590 81.060 5.800 ;
        RECT 80.985 4.240 81.060 4.450 ;
        RECT 80.985 2.890 81.060 3.100 ;
        RECT 80.985 1.545 81.060 1.755 ;
        RECT 80.985 0.190 81.060 0.405 ;
    END
  END RBL0_27
  PIN RBL1_28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.445175 ;
    PORT
      LAYER li1 ;
        RECT 81.200 42.040 81.275 42.250 ;
        RECT 81.200 40.690 81.275 40.900 ;
        RECT 81.200 39.340 81.275 39.550 ;
        RECT 81.200 37.990 81.275 38.200 ;
        RECT 81.200 36.640 81.275 36.850 ;
        RECT 81.200 35.290 81.275 35.500 ;
        RECT 81.200 33.940 81.275 34.150 ;
        RECT 81.200 32.590 81.275 32.800 ;
        RECT 81.200 31.240 81.275 31.450 ;
        RECT 81.200 29.890 81.275 30.100 ;
        RECT 81.200 28.540 81.275 28.750 ;
        RECT 81.200 27.190 81.275 27.400 ;
        RECT 81.200 25.840 81.275 26.050 ;
        RECT 81.200 24.490 81.275 24.700 ;
        RECT 81.200 23.140 81.275 23.350 ;
        RECT 81.200 21.790 81.275 22.000 ;
        RECT 81.200 20.440 81.275 20.650 ;
        RECT 81.200 19.090 81.275 19.300 ;
        RECT 81.200 17.740 81.275 17.950 ;
        RECT 81.200 16.390 81.275 16.600 ;
        RECT 81.200 15.040 81.275 15.250 ;
        RECT 81.200 13.690 81.275 13.900 ;
        RECT 81.200 12.340 81.275 12.550 ;
        RECT 81.200 10.990 81.275 11.200 ;
        RECT 81.200 9.640 81.275 9.850 ;
        RECT 81.200 8.290 81.275 8.500 ;
        RECT 81.200 6.940 81.275 7.150 ;
        RECT 81.200 5.590 81.275 5.800 ;
        RECT 81.200 4.240 81.275 4.450 ;
        RECT 81.200 2.890 81.275 3.100 ;
        RECT 81.200 1.545 81.275 1.755 ;
        RECT 81.200 0.190 81.275 0.405 ;
    END
  END RBL1_28
  PIN RBL0_28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.445175 ;
    PORT
      LAYER li1 ;
        RECT 83.885 42.040 83.960 42.250 ;
        RECT 83.885 40.690 83.960 40.900 ;
        RECT 83.885 39.340 83.960 39.550 ;
        RECT 83.885 37.990 83.960 38.200 ;
        RECT 83.885 36.640 83.960 36.850 ;
        RECT 83.885 35.290 83.960 35.500 ;
        RECT 83.885 33.940 83.960 34.150 ;
        RECT 83.885 32.590 83.960 32.800 ;
        RECT 83.885 31.240 83.960 31.450 ;
        RECT 83.885 29.890 83.960 30.100 ;
        RECT 83.885 28.540 83.960 28.750 ;
        RECT 83.885 27.190 83.960 27.400 ;
        RECT 83.885 25.840 83.960 26.050 ;
        RECT 83.885 24.490 83.960 24.700 ;
        RECT 83.885 23.140 83.960 23.350 ;
        RECT 83.885 21.790 83.960 22.000 ;
        RECT 83.885 20.440 83.960 20.650 ;
        RECT 83.885 19.090 83.960 19.300 ;
        RECT 83.885 17.740 83.960 17.950 ;
        RECT 83.885 16.390 83.960 16.600 ;
        RECT 83.885 15.040 83.960 15.250 ;
        RECT 83.885 13.690 83.960 13.900 ;
        RECT 83.885 12.340 83.960 12.550 ;
        RECT 83.885 10.990 83.960 11.200 ;
        RECT 83.885 9.640 83.960 9.850 ;
        RECT 83.885 8.290 83.960 8.500 ;
        RECT 83.885 6.940 83.960 7.150 ;
        RECT 83.885 5.590 83.960 5.800 ;
        RECT 83.885 4.240 83.960 4.450 ;
        RECT 83.885 2.890 83.960 3.100 ;
        RECT 83.885 1.545 83.960 1.755 ;
        RECT 83.885 0.190 83.960 0.405 ;
    END
  END RBL0_28
  PIN RBL1_29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.445175 ;
    PORT
      LAYER li1 ;
        RECT 84.100 42.040 84.175 42.250 ;
        RECT 84.100 40.690 84.175 40.900 ;
        RECT 84.100 39.340 84.175 39.550 ;
        RECT 84.100 37.990 84.175 38.200 ;
        RECT 84.100 36.640 84.175 36.850 ;
        RECT 84.100 35.290 84.175 35.500 ;
        RECT 84.100 33.940 84.175 34.150 ;
        RECT 84.100 32.590 84.175 32.800 ;
        RECT 84.100 31.240 84.175 31.450 ;
        RECT 84.100 29.890 84.175 30.100 ;
        RECT 84.100 28.540 84.175 28.750 ;
        RECT 84.100 27.190 84.175 27.400 ;
        RECT 84.100 25.840 84.175 26.050 ;
        RECT 84.100 24.490 84.175 24.700 ;
        RECT 84.100 23.140 84.175 23.350 ;
        RECT 84.100 21.790 84.175 22.000 ;
        RECT 84.100 20.440 84.175 20.650 ;
        RECT 84.100 19.090 84.175 19.300 ;
        RECT 84.100 17.740 84.175 17.950 ;
        RECT 84.100 16.390 84.175 16.600 ;
        RECT 84.100 15.040 84.175 15.250 ;
        RECT 84.100 13.690 84.175 13.900 ;
        RECT 84.100 12.340 84.175 12.550 ;
        RECT 84.100 10.990 84.175 11.200 ;
        RECT 84.100 9.640 84.175 9.850 ;
        RECT 84.100 8.290 84.175 8.500 ;
        RECT 84.100 6.940 84.175 7.150 ;
        RECT 84.100 5.590 84.175 5.800 ;
        RECT 84.100 4.240 84.175 4.450 ;
        RECT 84.100 2.890 84.175 3.100 ;
        RECT 84.100 1.545 84.175 1.755 ;
        RECT 84.100 0.190 84.175 0.405 ;
    END
  END RBL1_29
  PIN RBL0_29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.445175 ;
    PORT
      LAYER li1 ;
        RECT 86.785 42.040 86.860 42.250 ;
        RECT 86.785 40.690 86.860 40.900 ;
        RECT 86.785 39.340 86.860 39.550 ;
        RECT 86.785 37.990 86.860 38.200 ;
        RECT 86.785 36.640 86.860 36.850 ;
        RECT 86.785 35.290 86.860 35.500 ;
        RECT 86.785 33.940 86.860 34.150 ;
        RECT 86.785 32.590 86.860 32.800 ;
        RECT 86.785 31.240 86.860 31.450 ;
        RECT 86.785 29.890 86.860 30.100 ;
        RECT 86.785 28.540 86.860 28.750 ;
        RECT 86.785 27.190 86.860 27.400 ;
        RECT 86.785 25.840 86.860 26.050 ;
        RECT 86.785 24.490 86.860 24.700 ;
        RECT 86.785 23.140 86.860 23.350 ;
        RECT 86.785 21.790 86.860 22.000 ;
        RECT 86.785 20.440 86.860 20.650 ;
        RECT 86.785 19.090 86.860 19.300 ;
        RECT 86.785 17.740 86.860 17.950 ;
        RECT 86.785 16.390 86.860 16.600 ;
        RECT 86.785 15.040 86.860 15.250 ;
        RECT 86.785 13.690 86.860 13.900 ;
        RECT 86.785 12.340 86.860 12.550 ;
        RECT 86.785 10.990 86.860 11.200 ;
        RECT 86.785 9.640 86.860 9.850 ;
        RECT 86.785 8.290 86.860 8.500 ;
        RECT 86.785 6.940 86.860 7.150 ;
        RECT 86.785 5.590 86.860 5.800 ;
        RECT 86.785 4.240 86.860 4.450 ;
        RECT 86.785 2.890 86.860 3.100 ;
        RECT 86.785 1.545 86.860 1.755 ;
        RECT 86.785 0.190 86.860 0.405 ;
    END
  END RBL0_29
  PIN RBL1_30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.445175 ;
    PORT
      LAYER li1 ;
        RECT 87.000 42.040 87.075 42.250 ;
        RECT 87.000 40.690 87.075 40.900 ;
        RECT 87.000 39.340 87.075 39.550 ;
        RECT 87.000 37.990 87.075 38.200 ;
        RECT 87.000 36.640 87.075 36.850 ;
        RECT 87.000 35.290 87.075 35.500 ;
        RECT 87.000 33.940 87.075 34.150 ;
        RECT 87.000 32.590 87.075 32.800 ;
        RECT 87.000 31.240 87.075 31.450 ;
        RECT 87.000 29.890 87.075 30.100 ;
        RECT 87.000 28.540 87.075 28.750 ;
        RECT 87.000 27.190 87.075 27.400 ;
        RECT 87.000 25.840 87.075 26.050 ;
        RECT 87.000 24.490 87.075 24.700 ;
        RECT 87.000 23.140 87.075 23.350 ;
        RECT 87.000 21.790 87.075 22.000 ;
        RECT 87.000 20.440 87.075 20.650 ;
        RECT 87.000 19.090 87.075 19.300 ;
        RECT 87.000 17.740 87.075 17.950 ;
        RECT 87.000 16.390 87.075 16.600 ;
        RECT 87.000 15.040 87.075 15.250 ;
        RECT 87.000 13.690 87.075 13.900 ;
        RECT 87.000 12.340 87.075 12.550 ;
        RECT 87.000 10.990 87.075 11.200 ;
        RECT 87.000 9.640 87.075 9.850 ;
        RECT 87.000 8.290 87.075 8.500 ;
        RECT 87.000 6.940 87.075 7.150 ;
        RECT 87.000 5.590 87.075 5.800 ;
        RECT 87.000 4.240 87.075 4.450 ;
        RECT 87.000 2.890 87.075 3.100 ;
        RECT 87.000 1.545 87.075 1.755 ;
        RECT 87.000 0.190 87.075 0.405 ;
    END
  END RBL1_30
  PIN RBL0_30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.445175 ;
    PORT
      LAYER li1 ;
        RECT 89.685 42.040 89.760 42.250 ;
        RECT 89.685 40.690 89.760 40.900 ;
        RECT 89.685 39.340 89.760 39.550 ;
        RECT 89.685 37.990 89.760 38.200 ;
        RECT 89.685 36.640 89.760 36.850 ;
        RECT 89.685 35.290 89.760 35.500 ;
        RECT 89.685 33.940 89.760 34.150 ;
        RECT 89.685 32.590 89.760 32.800 ;
        RECT 89.685 31.240 89.760 31.450 ;
        RECT 89.685 29.890 89.760 30.100 ;
        RECT 89.685 28.540 89.760 28.750 ;
        RECT 89.685 27.190 89.760 27.400 ;
        RECT 89.685 25.840 89.760 26.050 ;
        RECT 89.685 24.490 89.760 24.700 ;
        RECT 89.685 23.140 89.760 23.350 ;
        RECT 89.685 21.790 89.760 22.000 ;
        RECT 89.685 20.440 89.760 20.650 ;
        RECT 89.685 19.090 89.760 19.300 ;
        RECT 89.685 17.740 89.760 17.950 ;
        RECT 89.685 16.390 89.760 16.600 ;
        RECT 89.685 15.040 89.760 15.250 ;
        RECT 89.685 13.690 89.760 13.900 ;
        RECT 89.685 12.340 89.760 12.550 ;
        RECT 89.685 10.990 89.760 11.200 ;
        RECT 89.685 9.640 89.760 9.850 ;
        RECT 89.685 8.290 89.760 8.500 ;
        RECT 89.685 6.940 89.760 7.150 ;
        RECT 89.685 5.590 89.760 5.800 ;
        RECT 89.685 4.240 89.760 4.450 ;
        RECT 89.685 2.890 89.760 3.100 ;
        RECT 89.685 1.545 89.760 1.755 ;
        RECT 89.685 0.190 89.760 0.405 ;
    END
  END RBL0_30
  PIN RBL1_31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.445175 ;
    PORT
      LAYER li1 ;
        RECT 89.900 42.040 89.975 42.250 ;
        RECT 89.900 40.690 89.975 40.900 ;
        RECT 89.900 39.340 89.975 39.550 ;
        RECT 89.900 37.990 89.975 38.200 ;
        RECT 89.900 36.640 89.975 36.850 ;
        RECT 89.900 35.290 89.975 35.500 ;
        RECT 89.900 33.940 89.975 34.150 ;
        RECT 89.900 32.590 89.975 32.800 ;
        RECT 89.900 31.240 89.975 31.450 ;
        RECT 89.900 29.890 89.975 30.100 ;
        RECT 89.900 28.540 89.975 28.750 ;
        RECT 89.900 27.190 89.975 27.400 ;
        RECT 89.900 25.840 89.975 26.050 ;
        RECT 89.900 24.490 89.975 24.700 ;
        RECT 89.900 23.140 89.975 23.350 ;
        RECT 89.900 21.790 89.975 22.000 ;
        RECT 89.900 20.440 89.975 20.650 ;
        RECT 89.900 19.090 89.975 19.300 ;
        RECT 89.900 17.740 89.975 17.950 ;
        RECT 89.900 16.390 89.975 16.600 ;
        RECT 89.900 15.040 89.975 15.250 ;
        RECT 89.900 13.690 89.975 13.900 ;
        RECT 89.900 12.340 89.975 12.550 ;
        RECT 89.900 10.990 89.975 11.200 ;
        RECT 89.900 9.640 89.975 9.850 ;
        RECT 89.900 8.290 89.975 8.500 ;
        RECT 89.900 6.940 89.975 7.150 ;
        RECT 89.900 5.590 89.975 5.800 ;
        RECT 89.900 4.240 89.975 4.450 ;
        RECT 89.900 2.890 89.975 3.100 ;
        RECT 89.900 1.545 89.975 1.755 ;
        RECT 89.900 0.190 89.975 0.405 ;
    END
  END RBL1_31
  PIN RBL0_31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.445175 ;
    PORT
      LAYER li1 ;
        RECT 92.585 42.040 92.660 42.250 ;
        RECT 92.585 40.690 92.660 40.900 ;
        RECT 92.585 39.340 92.660 39.550 ;
        RECT 92.585 37.990 92.660 38.200 ;
        RECT 92.585 36.640 92.660 36.850 ;
        RECT 92.585 35.290 92.660 35.500 ;
        RECT 92.585 33.940 92.660 34.150 ;
        RECT 92.585 32.590 92.660 32.800 ;
        RECT 92.585 31.240 92.660 31.450 ;
        RECT 92.585 29.890 92.660 30.100 ;
        RECT 92.585 28.540 92.660 28.750 ;
        RECT 92.585 27.190 92.660 27.400 ;
        RECT 92.585 25.840 92.660 26.050 ;
        RECT 92.585 24.490 92.660 24.700 ;
        RECT 92.585 23.140 92.660 23.350 ;
        RECT 92.585 21.790 92.660 22.000 ;
        RECT 92.585 20.440 92.660 20.650 ;
        RECT 92.585 19.090 92.660 19.300 ;
        RECT 92.585 17.740 92.660 17.950 ;
        RECT 92.585 16.390 92.660 16.600 ;
        RECT 92.585 15.040 92.660 15.250 ;
        RECT 92.585 13.690 92.660 13.900 ;
        RECT 92.585 12.340 92.660 12.550 ;
        RECT 92.585 10.990 92.660 11.200 ;
        RECT 92.585 9.640 92.660 9.850 ;
        RECT 92.585 8.290 92.660 8.500 ;
        RECT 92.585 6.940 92.660 7.150 ;
        RECT 92.585 5.590 92.660 5.800 ;
        RECT 92.585 4.240 92.660 4.450 ;
        RECT 92.585 2.890 92.660 3.100 ;
        RECT 92.585 1.545 92.660 1.755 ;
        RECT 92.585 0.190 92.660 0.405 ;
    END
  END RBL0_31
  PIN WBL_16
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.773600 ;
    PORT
      LAYER li1 ;
        RECT 48.720 42.770 48.795 42.915 ;
        RECT 48.720 41.420 48.795 41.565 ;
        RECT 48.720 40.070 48.795 40.215 ;
        RECT 48.720 38.720 48.795 38.865 ;
        RECT 48.720 37.370 48.795 37.515 ;
        RECT 48.720 36.020 48.795 36.165 ;
        RECT 48.720 34.670 48.795 34.815 ;
        RECT 48.720 33.320 48.795 33.465 ;
        RECT 48.720 31.970 48.795 32.115 ;
        RECT 48.720 30.620 48.795 30.765 ;
        RECT 48.720 29.270 48.795 29.415 ;
        RECT 48.720 27.920 48.795 28.065 ;
        RECT 48.720 26.570 48.795 26.715 ;
        RECT 48.720 25.220 48.795 25.365 ;
        RECT 48.720 23.870 48.795 24.015 ;
        RECT 48.720 22.520 48.795 22.665 ;
        RECT 48.720 21.170 48.795 21.315 ;
        RECT 48.720 19.820 48.795 19.965 ;
        RECT 48.720 18.470 48.795 18.615 ;
        RECT 48.720 17.120 48.795 17.265 ;
        RECT 48.720 15.770 48.795 15.915 ;
        RECT 48.720 14.420 48.795 14.565 ;
        RECT 48.720 13.070 48.795 13.215 ;
        RECT 48.720 11.720 48.795 11.865 ;
        RECT 48.720 10.370 48.795 10.515 ;
        RECT 48.720 9.020 48.795 9.165 ;
        RECT 48.720 7.670 48.795 7.815 ;
        RECT 48.720 6.320 48.795 6.465 ;
        RECT 48.720 4.970 48.795 5.115 ;
        RECT 48.720 3.620 48.795 3.765 ;
        RECT 48.720 2.275 48.795 2.420 ;
        RECT 48.720 0.925 48.795 1.070 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.320 42.770 2.395 42.915 ;
        RECT 2.320 41.420 2.395 41.565 ;
        RECT 2.320 40.070 2.395 40.215 ;
        RECT 2.320 38.720 2.395 38.865 ;
        RECT 2.320 37.370 2.395 37.515 ;
        RECT 2.320 36.020 2.395 36.165 ;
        RECT 2.320 34.670 2.395 34.815 ;
        RECT 2.320 33.320 2.395 33.465 ;
        RECT 2.320 31.970 2.395 32.115 ;
        RECT 2.320 30.620 2.395 30.765 ;
        RECT 2.320 29.270 2.395 29.415 ;
        RECT 2.320 27.920 2.395 28.065 ;
        RECT 2.320 26.570 2.395 26.715 ;
        RECT 2.320 25.220 2.395 25.365 ;
        RECT 2.320 23.870 2.395 24.015 ;
        RECT 2.320 22.520 2.395 22.665 ;
        RECT 2.320 21.170 2.395 21.315 ;
        RECT 2.320 19.820 2.395 19.965 ;
        RECT 2.320 18.470 2.395 18.615 ;
        RECT 2.320 17.120 2.395 17.265 ;
        RECT 2.320 15.770 2.395 15.915 ;
        RECT 2.320 14.420 2.395 14.565 ;
        RECT 2.320 13.070 2.395 13.215 ;
        RECT 2.320 11.720 2.395 11.865 ;
        RECT 2.320 10.370 2.395 10.515 ;
        RECT 2.320 9.020 2.395 9.165 ;
        RECT 2.320 7.670 2.395 7.815 ;
        RECT 2.320 6.320 2.395 6.465 ;
        RECT 2.320 4.970 2.395 5.115 ;
        RECT 2.320 3.620 2.395 3.765 ;
        RECT 2.320 2.270 2.395 2.415 ;
        RECT 2.320 0.920 2.395 1.065 ;
    END
  END WBL_16
  PIN WBLb_16
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.739200 ;
    PORT
      LAYER li1 ;
        RECT 46.770 42.770 46.845 42.910 ;
        RECT 46.770 41.420 46.845 41.560 ;
        RECT 46.770 40.070 46.845 40.210 ;
        RECT 46.770 38.720 46.845 38.860 ;
        RECT 46.770 37.370 46.845 37.510 ;
        RECT 46.770 36.020 46.845 36.160 ;
        RECT 46.770 34.670 46.845 34.810 ;
        RECT 46.770 33.320 46.845 33.460 ;
        RECT 46.770 31.970 46.845 32.110 ;
        RECT 46.770 30.620 46.845 30.760 ;
        RECT 46.770 29.270 46.845 29.410 ;
        RECT 46.770 27.920 46.845 28.060 ;
        RECT 46.770 26.570 46.845 26.710 ;
        RECT 46.770 25.220 46.845 25.360 ;
        RECT 46.770 23.870 46.845 24.010 ;
        RECT 46.770 22.520 46.845 22.660 ;
        RECT 46.770 21.170 46.845 21.310 ;
        RECT 46.770 19.820 46.845 19.960 ;
        RECT 46.770 18.470 46.845 18.610 ;
        RECT 46.770 17.120 46.845 17.260 ;
        RECT 46.770 15.770 46.845 15.910 ;
        RECT 46.770 14.420 46.845 14.560 ;
        RECT 46.770 13.070 46.845 13.210 ;
        RECT 46.770 11.720 46.845 11.860 ;
        RECT 46.770 10.370 46.845 10.510 ;
        RECT 46.770 9.020 46.845 9.160 ;
        RECT 46.770 7.670 46.845 7.810 ;
        RECT 46.770 6.320 46.845 6.460 ;
        RECT 46.770 4.970 46.845 5.110 ;
        RECT 46.770 3.620 46.845 3.760 ;
        RECT 46.770 2.275 46.845 2.415 ;
        RECT 46.770 0.925 46.845 1.065 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.370 42.770 0.445 42.910 ;
        RECT 0.370 41.420 0.445 41.560 ;
        RECT 0.370 40.070 0.445 40.210 ;
        RECT 0.370 38.720 0.445 38.860 ;
        RECT 0.370 37.370 0.445 37.510 ;
        RECT 0.370 36.020 0.445 36.160 ;
        RECT 0.370 34.670 0.445 34.810 ;
        RECT 0.370 33.320 0.445 33.460 ;
        RECT 0.370 31.970 0.445 32.110 ;
        RECT 0.370 30.620 0.445 30.760 ;
        RECT 0.370 29.270 0.445 29.410 ;
        RECT 0.370 27.920 0.445 28.060 ;
        RECT 0.370 26.570 0.445 26.710 ;
        RECT 0.370 25.220 0.445 25.360 ;
        RECT 0.370 23.870 0.445 24.010 ;
        RECT 0.370 22.520 0.445 22.660 ;
        RECT 0.370 21.170 0.445 21.310 ;
        RECT 0.370 19.820 0.445 19.960 ;
        RECT 0.370 18.470 0.445 18.610 ;
        RECT 0.370 17.120 0.445 17.260 ;
        RECT 0.370 15.770 0.445 15.910 ;
        RECT 0.370 14.420 0.445 14.560 ;
        RECT 0.370 13.070 0.445 13.210 ;
        RECT 0.370 11.720 0.445 11.860 ;
        RECT 0.370 10.370 0.445 10.510 ;
        RECT 0.370 9.020 0.445 9.160 ;
        RECT 0.370 7.670 0.445 7.810 ;
        RECT 0.370 6.320 0.445 6.460 ;
        RECT 0.370 4.970 0.445 5.110 ;
        RECT 0.370 3.620 0.445 3.760 ;
        RECT 0.370 2.270 0.445 2.410 ;
        RECT 0.370 0.920 0.445 1.060 ;
    END
  END WBLb_16
  PIN WBL_17
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.773600 ;
    PORT
      LAYER li1 ;
        RECT 51.620 42.770 51.695 42.915 ;
        RECT 51.620 41.420 51.695 41.565 ;
        RECT 51.620 40.070 51.695 40.215 ;
        RECT 51.620 38.720 51.695 38.865 ;
        RECT 51.620 37.370 51.695 37.515 ;
        RECT 51.620 36.020 51.695 36.165 ;
        RECT 51.620 34.670 51.695 34.815 ;
        RECT 51.620 33.320 51.695 33.465 ;
        RECT 51.620 31.970 51.695 32.115 ;
        RECT 51.620 30.620 51.695 30.765 ;
        RECT 51.620 29.270 51.695 29.415 ;
        RECT 51.620 27.920 51.695 28.065 ;
        RECT 51.620 26.570 51.695 26.715 ;
        RECT 51.620 25.220 51.695 25.365 ;
        RECT 51.620 23.870 51.695 24.015 ;
        RECT 51.620 22.520 51.695 22.665 ;
        RECT 51.620 21.170 51.695 21.315 ;
        RECT 51.620 19.820 51.695 19.965 ;
        RECT 51.620 18.470 51.695 18.615 ;
        RECT 51.620 17.120 51.695 17.265 ;
        RECT 51.620 15.770 51.695 15.915 ;
        RECT 51.620 14.420 51.695 14.565 ;
        RECT 51.620 13.070 51.695 13.215 ;
        RECT 51.620 11.720 51.695 11.865 ;
        RECT 51.620 10.370 51.695 10.515 ;
        RECT 51.620 9.020 51.695 9.165 ;
        RECT 51.620 7.670 51.695 7.815 ;
        RECT 51.620 6.320 51.695 6.465 ;
        RECT 51.620 4.970 51.695 5.115 ;
        RECT 51.620 3.620 51.695 3.765 ;
        RECT 51.620 2.275 51.695 2.420 ;
        RECT 51.620 0.925 51.695 1.070 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.220 42.770 5.295 42.915 ;
        RECT 5.220 41.420 5.295 41.565 ;
        RECT 5.220 40.070 5.295 40.215 ;
        RECT 5.220 38.720 5.295 38.865 ;
        RECT 5.220 37.370 5.295 37.515 ;
        RECT 5.220 36.020 5.295 36.165 ;
        RECT 5.220 34.670 5.295 34.815 ;
        RECT 5.220 33.320 5.295 33.465 ;
        RECT 5.220 31.970 5.295 32.115 ;
        RECT 5.220 30.620 5.295 30.765 ;
        RECT 5.220 29.270 5.295 29.415 ;
        RECT 5.220 27.920 5.295 28.065 ;
        RECT 5.220 26.570 5.295 26.715 ;
        RECT 5.220 25.220 5.295 25.365 ;
        RECT 5.220 23.870 5.295 24.015 ;
        RECT 5.220 22.520 5.295 22.665 ;
        RECT 5.220 21.170 5.295 21.315 ;
        RECT 5.220 19.820 5.295 19.965 ;
        RECT 5.220 18.470 5.295 18.615 ;
        RECT 5.220 17.120 5.295 17.265 ;
        RECT 5.220 15.770 5.295 15.915 ;
        RECT 5.220 14.420 5.295 14.565 ;
        RECT 5.220 13.070 5.295 13.215 ;
        RECT 5.220 11.720 5.295 11.865 ;
        RECT 5.220 10.370 5.295 10.515 ;
        RECT 5.220 9.020 5.295 9.165 ;
        RECT 5.220 7.670 5.295 7.815 ;
        RECT 5.220 6.320 5.295 6.465 ;
        RECT 5.220 4.970 5.295 5.115 ;
        RECT 5.220 3.620 5.295 3.765 ;
        RECT 5.220 2.270 5.295 2.415 ;
        RECT 5.220 0.920 5.295 1.065 ;
    END
  END WBL_17
  PIN WBLb_17
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.739200 ;
    PORT
      LAYER li1 ;
        RECT 49.670 42.770 49.745 42.910 ;
        RECT 49.670 41.420 49.745 41.560 ;
        RECT 49.670 40.070 49.745 40.210 ;
        RECT 49.670 38.720 49.745 38.860 ;
        RECT 49.670 37.370 49.745 37.510 ;
        RECT 49.670 36.020 49.745 36.160 ;
        RECT 49.670 34.670 49.745 34.810 ;
        RECT 49.670 33.320 49.745 33.460 ;
        RECT 49.670 31.970 49.745 32.110 ;
        RECT 49.670 30.620 49.745 30.760 ;
        RECT 49.670 29.270 49.745 29.410 ;
        RECT 49.670 27.920 49.745 28.060 ;
        RECT 49.670 26.570 49.745 26.710 ;
        RECT 49.670 25.220 49.745 25.360 ;
        RECT 49.670 23.870 49.745 24.010 ;
        RECT 49.670 22.520 49.745 22.660 ;
        RECT 49.670 21.170 49.745 21.310 ;
        RECT 49.670 19.820 49.745 19.960 ;
        RECT 49.670 18.470 49.745 18.610 ;
        RECT 49.670 17.120 49.745 17.260 ;
        RECT 49.670 15.770 49.745 15.910 ;
        RECT 49.670 14.420 49.745 14.560 ;
        RECT 49.670 13.070 49.745 13.210 ;
        RECT 49.670 11.720 49.745 11.860 ;
        RECT 49.670 10.370 49.745 10.510 ;
        RECT 49.670 9.020 49.745 9.160 ;
        RECT 49.670 7.670 49.745 7.810 ;
        RECT 49.670 6.320 49.745 6.460 ;
        RECT 49.670 4.970 49.745 5.110 ;
        RECT 49.670 3.620 49.745 3.760 ;
        RECT 49.670 2.275 49.745 2.415 ;
        RECT 49.670 0.925 49.745 1.065 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.270 42.770 3.345 42.910 ;
        RECT 3.270 41.420 3.345 41.560 ;
        RECT 3.270 40.070 3.345 40.210 ;
        RECT 3.270 38.720 3.345 38.860 ;
        RECT 3.270 37.370 3.345 37.510 ;
        RECT 3.270 36.020 3.345 36.160 ;
        RECT 3.270 34.670 3.345 34.810 ;
        RECT 3.270 33.320 3.345 33.460 ;
        RECT 3.270 31.970 3.345 32.110 ;
        RECT 3.270 30.620 3.345 30.760 ;
        RECT 3.270 29.270 3.345 29.410 ;
        RECT 3.270 27.920 3.345 28.060 ;
        RECT 3.270 26.570 3.345 26.710 ;
        RECT 3.270 25.220 3.345 25.360 ;
        RECT 3.270 23.870 3.345 24.010 ;
        RECT 3.270 22.520 3.345 22.660 ;
        RECT 3.270 21.170 3.345 21.310 ;
        RECT 3.270 19.820 3.345 19.960 ;
        RECT 3.270 18.470 3.345 18.610 ;
        RECT 3.270 17.120 3.345 17.260 ;
        RECT 3.270 15.770 3.345 15.910 ;
        RECT 3.270 14.420 3.345 14.560 ;
        RECT 3.270 13.070 3.345 13.210 ;
        RECT 3.270 11.720 3.345 11.860 ;
        RECT 3.270 10.370 3.345 10.510 ;
        RECT 3.270 9.020 3.345 9.160 ;
        RECT 3.270 7.670 3.345 7.810 ;
        RECT 3.270 6.320 3.345 6.460 ;
        RECT 3.270 4.970 3.345 5.110 ;
        RECT 3.270 3.620 3.345 3.760 ;
        RECT 3.270 2.270 3.345 2.410 ;
        RECT 3.270 0.920 3.345 1.060 ;
    END
  END WBLb_17
  PIN WBL_18
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.773600 ;
    PORT
      LAYER li1 ;
        RECT 54.520 42.770 54.595 42.915 ;
        RECT 54.520 41.420 54.595 41.565 ;
        RECT 54.520 40.070 54.595 40.215 ;
        RECT 54.520 38.720 54.595 38.865 ;
        RECT 54.520 37.370 54.595 37.515 ;
        RECT 54.520 36.020 54.595 36.165 ;
        RECT 54.520 34.670 54.595 34.815 ;
        RECT 54.520 33.320 54.595 33.465 ;
        RECT 54.520 31.970 54.595 32.115 ;
        RECT 54.520 30.620 54.595 30.765 ;
        RECT 54.520 29.270 54.595 29.415 ;
        RECT 54.520 27.920 54.595 28.065 ;
        RECT 54.520 26.570 54.595 26.715 ;
        RECT 54.520 25.220 54.595 25.365 ;
        RECT 54.520 23.870 54.595 24.015 ;
        RECT 54.520 22.520 54.595 22.665 ;
        RECT 54.520 21.170 54.595 21.315 ;
        RECT 54.520 19.820 54.595 19.965 ;
        RECT 54.520 18.470 54.595 18.615 ;
        RECT 54.520 17.120 54.595 17.265 ;
        RECT 54.520 15.770 54.595 15.915 ;
        RECT 54.520 14.420 54.595 14.565 ;
        RECT 54.520 13.070 54.595 13.215 ;
        RECT 54.520 11.720 54.595 11.865 ;
        RECT 54.520 10.370 54.595 10.515 ;
        RECT 54.520 9.020 54.595 9.165 ;
        RECT 54.520 7.670 54.595 7.815 ;
        RECT 54.520 6.320 54.595 6.465 ;
        RECT 54.520 4.970 54.595 5.115 ;
        RECT 54.520 3.620 54.595 3.765 ;
        RECT 54.520 2.275 54.595 2.420 ;
        RECT 54.520 0.925 54.595 1.070 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.120 42.770 8.195 42.915 ;
        RECT 8.120 41.420 8.195 41.565 ;
        RECT 8.120 40.070 8.195 40.215 ;
        RECT 8.120 38.720 8.195 38.865 ;
        RECT 8.120 37.370 8.195 37.515 ;
        RECT 8.120 36.020 8.195 36.165 ;
        RECT 8.120 34.670 8.195 34.815 ;
        RECT 8.120 33.320 8.195 33.465 ;
        RECT 8.120 31.970 8.195 32.115 ;
        RECT 8.120 30.620 8.195 30.765 ;
        RECT 8.120 29.270 8.195 29.415 ;
        RECT 8.120 27.920 8.195 28.065 ;
        RECT 8.120 26.570 8.195 26.715 ;
        RECT 8.120 25.220 8.195 25.365 ;
        RECT 8.120 23.870 8.195 24.015 ;
        RECT 8.120 22.520 8.195 22.665 ;
        RECT 8.120 21.170 8.195 21.315 ;
        RECT 8.120 19.820 8.195 19.965 ;
        RECT 8.120 18.470 8.195 18.615 ;
        RECT 8.120 17.120 8.195 17.265 ;
        RECT 8.120 15.770 8.195 15.915 ;
        RECT 8.120 14.420 8.195 14.565 ;
        RECT 8.120 13.070 8.195 13.215 ;
        RECT 8.120 11.720 8.195 11.865 ;
        RECT 8.120 10.370 8.195 10.515 ;
        RECT 8.120 9.020 8.195 9.165 ;
        RECT 8.120 7.670 8.195 7.815 ;
        RECT 8.120 6.320 8.195 6.465 ;
        RECT 8.120 4.970 8.195 5.115 ;
        RECT 8.120 3.620 8.195 3.765 ;
        RECT 8.120 2.270 8.195 2.415 ;
        RECT 8.120 0.920 8.195 1.065 ;
    END
  END WBL_18
  PIN WBLb_18
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.739200 ;
    PORT
      LAYER li1 ;
        RECT 52.570 42.770 52.645 42.910 ;
        RECT 52.570 41.420 52.645 41.560 ;
        RECT 52.570 40.070 52.645 40.210 ;
        RECT 52.570 38.720 52.645 38.860 ;
        RECT 52.570 37.370 52.645 37.510 ;
        RECT 52.570 36.020 52.645 36.160 ;
        RECT 52.570 34.670 52.645 34.810 ;
        RECT 52.570 33.320 52.645 33.460 ;
        RECT 52.570 31.970 52.645 32.110 ;
        RECT 52.570 30.620 52.645 30.760 ;
        RECT 52.570 29.270 52.645 29.410 ;
        RECT 52.570 27.920 52.645 28.060 ;
        RECT 52.570 26.570 52.645 26.710 ;
        RECT 52.570 25.220 52.645 25.360 ;
        RECT 52.570 23.870 52.645 24.010 ;
        RECT 52.570 22.520 52.645 22.660 ;
        RECT 52.570 21.170 52.645 21.310 ;
        RECT 52.570 19.820 52.645 19.960 ;
        RECT 52.570 18.470 52.645 18.610 ;
        RECT 52.570 17.120 52.645 17.260 ;
        RECT 52.570 15.770 52.645 15.910 ;
        RECT 52.570 14.420 52.645 14.560 ;
        RECT 52.570 13.070 52.645 13.210 ;
        RECT 52.570 11.720 52.645 11.860 ;
        RECT 52.570 10.370 52.645 10.510 ;
        RECT 52.570 9.020 52.645 9.160 ;
        RECT 52.570 7.670 52.645 7.810 ;
        RECT 52.570 6.320 52.645 6.460 ;
        RECT 52.570 4.970 52.645 5.110 ;
        RECT 52.570 3.620 52.645 3.760 ;
        RECT 52.570 2.275 52.645 2.415 ;
        RECT 52.570 0.925 52.645 1.065 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.170 42.770 6.245 42.910 ;
        RECT 6.170 41.420 6.245 41.560 ;
        RECT 6.170 40.070 6.245 40.210 ;
        RECT 6.170 38.720 6.245 38.860 ;
        RECT 6.170 37.370 6.245 37.510 ;
        RECT 6.170 36.020 6.245 36.160 ;
        RECT 6.170 34.670 6.245 34.810 ;
        RECT 6.170 33.320 6.245 33.460 ;
        RECT 6.170 31.970 6.245 32.110 ;
        RECT 6.170 30.620 6.245 30.760 ;
        RECT 6.170 29.270 6.245 29.410 ;
        RECT 6.170 27.920 6.245 28.060 ;
        RECT 6.170 26.570 6.245 26.710 ;
        RECT 6.170 25.220 6.245 25.360 ;
        RECT 6.170 23.870 6.245 24.010 ;
        RECT 6.170 22.520 6.245 22.660 ;
        RECT 6.170 21.170 6.245 21.310 ;
        RECT 6.170 19.820 6.245 19.960 ;
        RECT 6.170 18.470 6.245 18.610 ;
        RECT 6.170 17.120 6.245 17.260 ;
        RECT 6.170 15.770 6.245 15.910 ;
        RECT 6.170 14.420 6.245 14.560 ;
        RECT 6.170 13.070 6.245 13.210 ;
        RECT 6.170 11.720 6.245 11.860 ;
        RECT 6.170 10.370 6.245 10.510 ;
        RECT 6.170 9.020 6.245 9.160 ;
        RECT 6.170 7.670 6.245 7.810 ;
        RECT 6.170 6.320 6.245 6.460 ;
        RECT 6.170 4.970 6.245 5.110 ;
        RECT 6.170 3.620 6.245 3.760 ;
        RECT 6.170 2.270 6.245 2.410 ;
        RECT 6.170 0.920 6.245 1.060 ;
    END
  END WBLb_18
  PIN WBL_19
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.773600 ;
    PORT
      LAYER li1 ;
        RECT 57.420 42.770 57.495 42.915 ;
        RECT 57.420 41.420 57.495 41.565 ;
        RECT 57.420 40.070 57.495 40.215 ;
        RECT 57.420 38.720 57.495 38.865 ;
        RECT 57.420 37.370 57.495 37.515 ;
        RECT 57.420 36.020 57.495 36.165 ;
        RECT 57.420 34.670 57.495 34.815 ;
        RECT 57.420 33.320 57.495 33.465 ;
        RECT 57.420 31.970 57.495 32.115 ;
        RECT 57.420 30.620 57.495 30.765 ;
        RECT 57.420 29.270 57.495 29.415 ;
        RECT 57.420 27.920 57.495 28.065 ;
        RECT 57.420 26.570 57.495 26.715 ;
        RECT 57.420 25.220 57.495 25.365 ;
        RECT 57.420 23.870 57.495 24.015 ;
        RECT 57.420 22.520 57.495 22.665 ;
        RECT 57.420 21.170 57.495 21.315 ;
        RECT 57.420 19.820 57.495 19.965 ;
        RECT 57.420 18.470 57.495 18.615 ;
        RECT 57.420 17.120 57.495 17.265 ;
        RECT 57.420 15.770 57.495 15.915 ;
        RECT 57.420 14.420 57.495 14.565 ;
        RECT 57.420 13.070 57.495 13.215 ;
        RECT 57.420 11.720 57.495 11.865 ;
        RECT 57.420 10.370 57.495 10.515 ;
        RECT 57.420 9.020 57.495 9.165 ;
        RECT 57.420 7.670 57.495 7.815 ;
        RECT 57.420 6.320 57.495 6.465 ;
        RECT 57.420 4.970 57.495 5.115 ;
        RECT 57.420 3.620 57.495 3.765 ;
        RECT 57.420 2.275 57.495 2.420 ;
        RECT 57.420 0.925 57.495 1.070 ;
    END
    PORT
      LAYER li1 ;
        RECT 11.020 42.770 11.095 42.915 ;
        RECT 11.020 41.420 11.095 41.565 ;
        RECT 11.020 40.070 11.095 40.215 ;
        RECT 11.020 38.720 11.095 38.865 ;
        RECT 11.020 37.370 11.095 37.515 ;
        RECT 11.020 36.020 11.095 36.165 ;
        RECT 11.020 34.670 11.095 34.815 ;
        RECT 11.020 33.320 11.095 33.465 ;
        RECT 11.020 31.970 11.095 32.115 ;
        RECT 11.020 30.620 11.095 30.765 ;
        RECT 11.020 29.270 11.095 29.415 ;
        RECT 11.020 27.920 11.095 28.065 ;
        RECT 11.020 26.570 11.095 26.715 ;
        RECT 11.020 25.220 11.095 25.365 ;
        RECT 11.020 23.870 11.095 24.015 ;
        RECT 11.020 22.520 11.095 22.665 ;
        RECT 11.020 21.170 11.095 21.315 ;
        RECT 11.020 19.820 11.095 19.965 ;
        RECT 11.020 18.470 11.095 18.615 ;
        RECT 11.020 17.120 11.095 17.265 ;
        RECT 11.020 15.770 11.095 15.915 ;
        RECT 11.020 14.420 11.095 14.565 ;
        RECT 11.020 13.070 11.095 13.215 ;
        RECT 11.020 11.720 11.095 11.865 ;
        RECT 11.020 10.370 11.095 10.515 ;
        RECT 11.020 9.020 11.095 9.165 ;
        RECT 11.020 7.670 11.095 7.815 ;
        RECT 11.020 6.320 11.095 6.465 ;
        RECT 11.020 4.970 11.095 5.115 ;
        RECT 11.020 3.620 11.095 3.765 ;
        RECT 11.020 2.270 11.095 2.415 ;
        RECT 11.020 0.920 11.095 1.065 ;
    END
  END WBL_19
  PIN WBLb_19
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.739200 ;
    PORT
      LAYER li1 ;
        RECT 55.470 42.770 55.545 42.910 ;
        RECT 55.470 41.420 55.545 41.560 ;
        RECT 55.470 40.070 55.545 40.210 ;
        RECT 55.470 38.720 55.545 38.860 ;
        RECT 55.470 37.370 55.545 37.510 ;
        RECT 55.470 36.020 55.545 36.160 ;
        RECT 55.470 34.670 55.545 34.810 ;
        RECT 55.470 33.320 55.545 33.460 ;
        RECT 55.470 31.970 55.545 32.110 ;
        RECT 55.470 30.620 55.545 30.760 ;
        RECT 55.470 29.270 55.545 29.410 ;
        RECT 55.470 27.920 55.545 28.060 ;
        RECT 55.470 26.570 55.545 26.710 ;
        RECT 55.470 25.220 55.545 25.360 ;
        RECT 55.470 23.870 55.545 24.010 ;
        RECT 55.470 22.520 55.545 22.660 ;
        RECT 55.470 21.170 55.545 21.310 ;
        RECT 55.470 19.820 55.545 19.960 ;
        RECT 55.470 18.470 55.545 18.610 ;
        RECT 55.470 17.120 55.545 17.260 ;
        RECT 55.470 15.770 55.545 15.910 ;
        RECT 55.470 14.420 55.545 14.560 ;
        RECT 55.470 13.070 55.545 13.210 ;
        RECT 55.470 11.720 55.545 11.860 ;
        RECT 55.470 10.370 55.545 10.510 ;
        RECT 55.470 9.020 55.545 9.160 ;
        RECT 55.470 7.670 55.545 7.810 ;
        RECT 55.470 6.320 55.545 6.460 ;
        RECT 55.470 4.970 55.545 5.110 ;
        RECT 55.470 3.620 55.545 3.760 ;
        RECT 55.470 2.275 55.545 2.415 ;
        RECT 55.470 0.925 55.545 1.065 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.070 42.770 9.145 42.910 ;
        RECT 9.070 41.420 9.145 41.560 ;
        RECT 9.070 40.070 9.145 40.210 ;
        RECT 9.070 38.720 9.145 38.860 ;
        RECT 9.070 37.370 9.145 37.510 ;
        RECT 9.070 36.020 9.145 36.160 ;
        RECT 9.070 34.670 9.145 34.810 ;
        RECT 9.070 33.320 9.145 33.460 ;
        RECT 9.070 31.970 9.145 32.110 ;
        RECT 9.070 30.620 9.145 30.760 ;
        RECT 9.070 29.270 9.145 29.410 ;
        RECT 9.070 27.920 9.145 28.060 ;
        RECT 9.070 26.570 9.145 26.710 ;
        RECT 9.070 25.220 9.145 25.360 ;
        RECT 9.070 23.870 9.145 24.010 ;
        RECT 9.070 22.520 9.145 22.660 ;
        RECT 9.070 21.170 9.145 21.310 ;
        RECT 9.070 19.820 9.145 19.960 ;
        RECT 9.070 18.470 9.145 18.610 ;
        RECT 9.070 17.120 9.145 17.260 ;
        RECT 9.070 15.770 9.145 15.910 ;
        RECT 9.070 14.420 9.145 14.560 ;
        RECT 9.070 13.070 9.145 13.210 ;
        RECT 9.070 11.720 9.145 11.860 ;
        RECT 9.070 10.370 9.145 10.510 ;
        RECT 9.070 9.020 9.145 9.160 ;
        RECT 9.070 7.670 9.145 7.810 ;
        RECT 9.070 6.320 9.145 6.460 ;
        RECT 9.070 4.970 9.145 5.110 ;
        RECT 9.070 3.620 9.145 3.760 ;
        RECT 9.070 2.270 9.145 2.410 ;
        RECT 9.070 0.920 9.145 1.060 ;
    END
  END WBLb_19
  PIN WBL_20
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.773600 ;
    PORT
      LAYER li1 ;
        RECT 60.320 42.770 60.395 42.915 ;
        RECT 60.320 41.420 60.395 41.565 ;
        RECT 60.320 40.070 60.395 40.215 ;
        RECT 60.320 38.720 60.395 38.865 ;
        RECT 60.320 37.370 60.395 37.515 ;
        RECT 60.320 36.020 60.395 36.165 ;
        RECT 60.320 34.670 60.395 34.815 ;
        RECT 60.320 33.320 60.395 33.465 ;
        RECT 60.320 31.970 60.395 32.115 ;
        RECT 60.320 30.620 60.395 30.765 ;
        RECT 60.320 29.270 60.395 29.415 ;
        RECT 60.320 27.920 60.395 28.065 ;
        RECT 60.320 26.570 60.395 26.715 ;
        RECT 60.320 25.220 60.395 25.365 ;
        RECT 60.320 23.870 60.395 24.015 ;
        RECT 60.320 22.520 60.395 22.665 ;
        RECT 60.320 21.170 60.395 21.315 ;
        RECT 60.320 19.820 60.395 19.965 ;
        RECT 60.320 18.470 60.395 18.615 ;
        RECT 60.320 17.120 60.395 17.265 ;
        RECT 60.320 15.770 60.395 15.915 ;
        RECT 60.320 14.420 60.395 14.565 ;
        RECT 60.320 13.070 60.395 13.215 ;
        RECT 60.320 11.720 60.395 11.865 ;
        RECT 60.320 10.370 60.395 10.515 ;
        RECT 60.320 9.020 60.395 9.165 ;
        RECT 60.320 7.670 60.395 7.815 ;
        RECT 60.320 6.320 60.395 6.465 ;
        RECT 60.320 4.970 60.395 5.115 ;
        RECT 60.320 3.620 60.395 3.765 ;
        RECT 60.320 2.275 60.395 2.420 ;
        RECT 60.320 0.925 60.395 1.070 ;
    END
    PORT
      LAYER li1 ;
        RECT 13.920 42.770 13.995 42.915 ;
        RECT 13.920 41.420 13.995 41.565 ;
        RECT 13.920 40.070 13.995 40.215 ;
        RECT 13.920 38.720 13.995 38.865 ;
        RECT 13.920 37.370 13.995 37.515 ;
        RECT 13.920 36.020 13.995 36.165 ;
        RECT 13.920 34.670 13.995 34.815 ;
        RECT 13.920 33.320 13.995 33.465 ;
        RECT 13.920 31.970 13.995 32.115 ;
        RECT 13.920 30.620 13.995 30.765 ;
        RECT 13.920 29.270 13.995 29.415 ;
        RECT 13.920 27.920 13.995 28.065 ;
        RECT 13.920 26.570 13.995 26.715 ;
        RECT 13.920 25.220 13.995 25.365 ;
        RECT 13.920 23.870 13.995 24.015 ;
        RECT 13.920 22.520 13.995 22.665 ;
        RECT 13.920 21.170 13.995 21.315 ;
        RECT 13.920 19.820 13.995 19.965 ;
        RECT 13.920 18.470 13.995 18.615 ;
        RECT 13.920 17.120 13.995 17.265 ;
        RECT 13.920 15.770 13.995 15.915 ;
        RECT 13.920 14.420 13.995 14.565 ;
        RECT 13.920 13.070 13.995 13.215 ;
        RECT 13.920 11.720 13.995 11.865 ;
        RECT 13.920 10.370 13.995 10.515 ;
        RECT 13.920 9.020 13.995 9.165 ;
        RECT 13.920 7.670 13.995 7.815 ;
        RECT 13.920 6.320 13.995 6.465 ;
        RECT 13.920 4.970 13.995 5.115 ;
        RECT 13.920 3.620 13.995 3.765 ;
        RECT 13.920 2.270 13.995 2.415 ;
        RECT 13.920 0.920 13.995 1.065 ;
    END
  END WBL_20
  PIN WBLb_20
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.739200 ;
    PORT
      LAYER li1 ;
        RECT 58.370 42.770 58.445 42.910 ;
        RECT 58.370 41.420 58.445 41.560 ;
        RECT 58.370 40.070 58.445 40.210 ;
        RECT 58.370 38.720 58.445 38.860 ;
        RECT 58.370 37.370 58.445 37.510 ;
        RECT 58.370 36.020 58.445 36.160 ;
        RECT 58.370 34.670 58.445 34.810 ;
        RECT 58.370 33.320 58.445 33.460 ;
        RECT 58.370 31.970 58.445 32.110 ;
        RECT 58.370 30.620 58.445 30.760 ;
        RECT 58.370 29.270 58.445 29.410 ;
        RECT 58.370 27.920 58.445 28.060 ;
        RECT 58.370 26.570 58.445 26.710 ;
        RECT 58.370 25.220 58.445 25.360 ;
        RECT 58.370 23.870 58.445 24.010 ;
        RECT 58.370 22.520 58.445 22.660 ;
        RECT 58.370 21.170 58.445 21.310 ;
        RECT 58.370 19.820 58.445 19.960 ;
        RECT 58.370 18.470 58.445 18.610 ;
        RECT 58.370 17.120 58.445 17.260 ;
        RECT 58.370 15.770 58.445 15.910 ;
        RECT 58.370 14.420 58.445 14.560 ;
        RECT 58.370 13.070 58.445 13.210 ;
        RECT 58.370 11.720 58.445 11.860 ;
        RECT 58.370 10.370 58.445 10.510 ;
        RECT 58.370 9.020 58.445 9.160 ;
        RECT 58.370 7.670 58.445 7.810 ;
        RECT 58.370 6.320 58.445 6.460 ;
        RECT 58.370 4.970 58.445 5.110 ;
        RECT 58.370 3.620 58.445 3.760 ;
        RECT 58.370 2.275 58.445 2.415 ;
        RECT 58.370 0.925 58.445 1.065 ;
    END
    PORT
      LAYER li1 ;
        RECT 11.970 42.770 12.045 42.910 ;
        RECT 11.970 41.420 12.045 41.560 ;
        RECT 11.970 40.070 12.045 40.210 ;
        RECT 11.970 38.720 12.045 38.860 ;
        RECT 11.970 37.370 12.045 37.510 ;
        RECT 11.970 36.020 12.045 36.160 ;
        RECT 11.970 34.670 12.045 34.810 ;
        RECT 11.970 33.320 12.045 33.460 ;
        RECT 11.970 31.970 12.045 32.110 ;
        RECT 11.970 30.620 12.045 30.760 ;
        RECT 11.970 29.270 12.045 29.410 ;
        RECT 11.970 27.920 12.045 28.060 ;
        RECT 11.970 26.570 12.045 26.710 ;
        RECT 11.970 25.220 12.045 25.360 ;
        RECT 11.970 23.870 12.045 24.010 ;
        RECT 11.970 22.520 12.045 22.660 ;
        RECT 11.970 21.170 12.045 21.310 ;
        RECT 11.970 19.820 12.045 19.960 ;
        RECT 11.970 18.470 12.045 18.610 ;
        RECT 11.970 17.120 12.045 17.260 ;
        RECT 11.970 15.770 12.045 15.910 ;
        RECT 11.970 14.420 12.045 14.560 ;
        RECT 11.970 13.070 12.045 13.210 ;
        RECT 11.970 11.720 12.045 11.860 ;
        RECT 11.970 10.370 12.045 10.510 ;
        RECT 11.970 9.020 12.045 9.160 ;
        RECT 11.970 7.670 12.045 7.810 ;
        RECT 11.970 6.320 12.045 6.460 ;
        RECT 11.970 4.970 12.045 5.110 ;
        RECT 11.970 3.620 12.045 3.760 ;
        RECT 11.970 2.270 12.045 2.410 ;
        RECT 11.970 0.920 12.045 1.060 ;
    END
  END WBLb_20
  PIN WBL_21
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.773600 ;
    PORT
      LAYER li1 ;
        RECT 63.220 42.770 63.295 42.915 ;
        RECT 63.220 41.420 63.295 41.565 ;
        RECT 63.220 40.070 63.295 40.215 ;
        RECT 63.220 38.720 63.295 38.865 ;
        RECT 63.220 37.370 63.295 37.515 ;
        RECT 63.220 36.020 63.295 36.165 ;
        RECT 63.220 34.670 63.295 34.815 ;
        RECT 63.220 33.320 63.295 33.465 ;
        RECT 63.220 31.970 63.295 32.115 ;
        RECT 63.220 30.620 63.295 30.765 ;
        RECT 63.220 29.270 63.295 29.415 ;
        RECT 63.220 27.920 63.295 28.065 ;
        RECT 63.220 26.570 63.295 26.715 ;
        RECT 63.220 25.220 63.295 25.365 ;
        RECT 63.220 23.870 63.295 24.015 ;
        RECT 63.220 22.520 63.295 22.665 ;
        RECT 63.220 21.170 63.295 21.315 ;
        RECT 63.220 19.820 63.295 19.965 ;
        RECT 63.220 18.470 63.295 18.615 ;
        RECT 63.220 17.120 63.295 17.265 ;
        RECT 63.220 15.770 63.295 15.915 ;
        RECT 63.220 14.420 63.295 14.565 ;
        RECT 63.220 13.070 63.295 13.215 ;
        RECT 63.220 11.720 63.295 11.865 ;
        RECT 63.220 10.370 63.295 10.515 ;
        RECT 63.220 9.020 63.295 9.165 ;
        RECT 63.220 7.670 63.295 7.815 ;
        RECT 63.220 6.320 63.295 6.465 ;
        RECT 63.220 4.970 63.295 5.115 ;
        RECT 63.220 3.620 63.295 3.765 ;
        RECT 63.220 2.275 63.295 2.420 ;
        RECT 63.220 0.925 63.295 1.070 ;
    END
    PORT
      LAYER li1 ;
        RECT 16.820 42.770 16.895 42.915 ;
        RECT 16.820 41.420 16.895 41.565 ;
        RECT 16.820 40.070 16.895 40.215 ;
        RECT 16.820 38.720 16.895 38.865 ;
        RECT 16.820 37.370 16.895 37.515 ;
        RECT 16.820 36.020 16.895 36.165 ;
        RECT 16.820 34.670 16.895 34.815 ;
        RECT 16.820 33.320 16.895 33.465 ;
        RECT 16.820 31.970 16.895 32.115 ;
        RECT 16.820 30.620 16.895 30.765 ;
        RECT 16.820 29.270 16.895 29.415 ;
        RECT 16.820 27.920 16.895 28.065 ;
        RECT 16.820 26.570 16.895 26.715 ;
        RECT 16.820 25.220 16.895 25.365 ;
        RECT 16.820 23.870 16.895 24.015 ;
        RECT 16.820 22.520 16.895 22.665 ;
        RECT 16.820 21.170 16.895 21.315 ;
        RECT 16.820 19.820 16.895 19.965 ;
        RECT 16.820 18.470 16.895 18.615 ;
        RECT 16.820 17.120 16.895 17.265 ;
        RECT 16.820 15.770 16.895 15.915 ;
        RECT 16.820 14.420 16.895 14.565 ;
        RECT 16.820 13.070 16.895 13.215 ;
        RECT 16.820 11.720 16.895 11.865 ;
        RECT 16.820 10.370 16.895 10.515 ;
        RECT 16.820 9.020 16.895 9.165 ;
        RECT 16.820 7.670 16.895 7.815 ;
        RECT 16.820 6.320 16.895 6.465 ;
        RECT 16.820 4.970 16.895 5.115 ;
        RECT 16.820 3.620 16.895 3.765 ;
        RECT 16.820 2.270 16.895 2.415 ;
        RECT 16.820 0.920 16.895 1.065 ;
    END
  END WBL_21
  PIN WBLb_21
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.739200 ;
    PORT
      LAYER li1 ;
        RECT 61.270 42.770 61.345 42.910 ;
        RECT 61.270 41.420 61.345 41.560 ;
        RECT 61.270 40.070 61.345 40.210 ;
        RECT 61.270 38.720 61.345 38.860 ;
        RECT 61.270 37.370 61.345 37.510 ;
        RECT 61.270 36.020 61.345 36.160 ;
        RECT 61.270 34.670 61.345 34.810 ;
        RECT 61.270 33.320 61.345 33.460 ;
        RECT 61.270 31.970 61.345 32.110 ;
        RECT 61.270 30.620 61.345 30.760 ;
        RECT 61.270 29.270 61.345 29.410 ;
        RECT 61.270 27.920 61.345 28.060 ;
        RECT 61.270 26.570 61.345 26.710 ;
        RECT 61.270 25.220 61.345 25.360 ;
        RECT 61.270 23.870 61.345 24.010 ;
        RECT 61.270 22.520 61.345 22.660 ;
        RECT 61.270 21.170 61.345 21.310 ;
        RECT 61.270 19.820 61.345 19.960 ;
        RECT 61.270 18.470 61.345 18.610 ;
        RECT 61.270 17.120 61.345 17.260 ;
        RECT 61.270 15.770 61.345 15.910 ;
        RECT 61.270 14.420 61.345 14.560 ;
        RECT 61.270 13.070 61.345 13.210 ;
        RECT 61.270 11.720 61.345 11.860 ;
        RECT 61.270 10.370 61.345 10.510 ;
        RECT 61.270 9.020 61.345 9.160 ;
        RECT 61.270 7.670 61.345 7.810 ;
        RECT 61.270 6.320 61.345 6.460 ;
        RECT 61.270 4.970 61.345 5.110 ;
        RECT 61.270 3.620 61.345 3.760 ;
        RECT 61.270 2.275 61.345 2.415 ;
        RECT 61.270 0.925 61.345 1.065 ;
    END
    PORT
      LAYER li1 ;
        RECT 14.870 42.770 14.945 42.910 ;
        RECT 14.870 41.420 14.945 41.560 ;
        RECT 14.870 40.070 14.945 40.210 ;
        RECT 14.870 38.720 14.945 38.860 ;
        RECT 14.870 37.370 14.945 37.510 ;
        RECT 14.870 36.020 14.945 36.160 ;
        RECT 14.870 34.670 14.945 34.810 ;
        RECT 14.870 33.320 14.945 33.460 ;
        RECT 14.870 31.970 14.945 32.110 ;
        RECT 14.870 30.620 14.945 30.760 ;
        RECT 14.870 29.270 14.945 29.410 ;
        RECT 14.870 27.920 14.945 28.060 ;
        RECT 14.870 26.570 14.945 26.710 ;
        RECT 14.870 25.220 14.945 25.360 ;
        RECT 14.870 23.870 14.945 24.010 ;
        RECT 14.870 22.520 14.945 22.660 ;
        RECT 14.870 21.170 14.945 21.310 ;
        RECT 14.870 19.820 14.945 19.960 ;
        RECT 14.870 18.470 14.945 18.610 ;
        RECT 14.870 17.120 14.945 17.260 ;
        RECT 14.870 15.770 14.945 15.910 ;
        RECT 14.870 14.420 14.945 14.560 ;
        RECT 14.870 13.070 14.945 13.210 ;
        RECT 14.870 11.720 14.945 11.860 ;
        RECT 14.870 10.370 14.945 10.510 ;
        RECT 14.870 9.020 14.945 9.160 ;
        RECT 14.870 7.670 14.945 7.810 ;
        RECT 14.870 6.320 14.945 6.460 ;
        RECT 14.870 4.970 14.945 5.110 ;
        RECT 14.870 3.620 14.945 3.760 ;
        RECT 14.870 2.270 14.945 2.410 ;
        RECT 14.870 0.920 14.945 1.060 ;
    END
  END WBLb_21
  PIN WBL_22
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.773600 ;
    PORT
      LAYER li1 ;
        RECT 66.120 42.770 66.195 42.915 ;
        RECT 66.120 41.420 66.195 41.565 ;
        RECT 66.120 40.070 66.195 40.215 ;
        RECT 66.120 38.720 66.195 38.865 ;
        RECT 66.120 37.370 66.195 37.515 ;
        RECT 66.120 36.020 66.195 36.165 ;
        RECT 66.120 34.670 66.195 34.815 ;
        RECT 66.120 33.320 66.195 33.465 ;
        RECT 66.120 31.970 66.195 32.115 ;
        RECT 66.120 30.620 66.195 30.765 ;
        RECT 66.120 29.270 66.195 29.415 ;
        RECT 66.120 27.920 66.195 28.065 ;
        RECT 66.120 26.570 66.195 26.715 ;
        RECT 66.120 25.220 66.195 25.365 ;
        RECT 66.120 23.870 66.195 24.015 ;
        RECT 66.120 22.520 66.195 22.665 ;
        RECT 66.120 21.170 66.195 21.315 ;
        RECT 66.120 19.820 66.195 19.965 ;
        RECT 66.120 18.470 66.195 18.615 ;
        RECT 66.120 17.120 66.195 17.265 ;
        RECT 66.120 15.770 66.195 15.915 ;
        RECT 66.120 14.420 66.195 14.565 ;
        RECT 66.120 13.070 66.195 13.215 ;
        RECT 66.120 11.720 66.195 11.865 ;
        RECT 66.120 10.370 66.195 10.515 ;
        RECT 66.120 9.020 66.195 9.165 ;
        RECT 66.120 7.670 66.195 7.815 ;
        RECT 66.120 6.320 66.195 6.465 ;
        RECT 66.120 4.970 66.195 5.115 ;
        RECT 66.120 3.620 66.195 3.765 ;
        RECT 66.120 2.275 66.195 2.420 ;
        RECT 66.120 0.925 66.195 1.070 ;
    END
    PORT
      LAYER li1 ;
        RECT 19.720 42.770 19.795 42.915 ;
        RECT 19.720 41.420 19.795 41.565 ;
        RECT 19.720 40.070 19.795 40.215 ;
        RECT 19.720 38.720 19.795 38.865 ;
        RECT 19.720 37.370 19.795 37.515 ;
        RECT 19.720 36.020 19.795 36.165 ;
        RECT 19.720 34.670 19.795 34.815 ;
        RECT 19.720 33.320 19.795 33.465 ;
        RECT 19.720 31.970 19.795 32.115 ;
        RECT 19.720 30.620 19.795 30.765 ;
        RECT 19.720 29.270 19.795 29.415 ;
        RECT 19.720 27.920 19.795 28.065 ;
        RECT 19.720 26.570 19.795 26.715 ;
        RECT 19.720 25.220 19.795 25.365 ;
        RECT 19.720 23.870 19.795 24.015 ;
        RECT 19.720 22.520 19.795 22.665 ;
        RECT 19.720 21.170 19.795 21.315 ;
        RECT 19.720 19.820 19.795 19.965 ;
        RECT 19.720 18.470 19.795 18.615 ;
        RECT 19.720 17.120 19.795 17.265 ;
        RECT 19.720 15.770 19.795 15.915 ;
        RECT 19.720 14.420 19.795 14.565 ;
        RECT 19.720 13.070 19.795 13.215 ;
        RECT 19.720 11.720 19.795 11.865 ;
        RECT 19.720 10.370 19.795 10.515 ;
        RECT 19.720 9.020 19.795 9.165 ;
        RECT 19.720 7.670 19.795 7.815 ;
        RECT 19.720 6.320 19.795 6.465 ;
        RECT 19.720 4.970 19.795 5.115 ;
        RECT 19.720 3.620 19.795 3.765 ;
        RECT 19.720 2.270 19.795 2.415 ;
        RECT 19.720 0.920 19.795 1.065 ;
    END
  END WBL_22
  PIN WBLb_22
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.739200 ;
    PORT
      LAYER li1 ;
        RECT 64.170 42.770 64.245 42.910 ;
        RECT 64.170 41.420 64.245 41.560 ;
        RECT 64.170 40.070 64.245 40.210 ;
        RECT 64.170 38.720 64.245 38.860 ;
        RECT 64.170 37.370 64.245 37.510 ;
        RECT 64.170 36.020 64.245 36.160 ;
        RECT 64.170 34.670 64.245 34.810 ;
        RECT 64.170 33.320 64.245 33.460 ;
        RECT 64.170 31.970 64.245 32.110 ;
        RECT 64.170 30.620 64.245 30.760 ;
        RECT 64.170 29.270 64.245 29.410 ;
        RECT 64.170 27.920 64.245 28.060 ;
        RECT 64.170 26.570 64.245 26.710 ;
        RECT 64.170 25.220 64.245 25.360 ;
        RECT 64.170 23.870 64.245 24.010 ;
        RECT 64.170 22.520 64.245 22.660 ;
        RECT 64.170 21.170 64.245 21.310 ;
        RECT 64.170 19.820 64.245 19.960 ;
        RECT 64.170 18.470 64.245 18.610 ;
        RECT 64.170 17.120 64.245 17.260 ;
        RECT 64.170 15.770 64.245 15.910 ;
        RECT 64.170 14.420 64.245 14.560 ;
        RECT 64.170 13.070 64.245 13.210 ;
        RECT 64.170 11.720 64.245 11.860 ;
        RECT 64.170 10.370 64.245 10.510 ;
        RECT 64.170 9.020 64.245 9.160 ;
        RECT 64.170 7.670 64.245 7.810 ;
        RECT 64.170 6.320 64.245 6.460 ;
        RECT 64.170 4.970 64.245 5.110 ;
        RECT 64.170 3.620 64.245 3.760 ;
        RECT 64.170 2.275 64.245 2.415 ;
        RECT 64.170 0.925 64.245 1.065 ;
    END
    PORT
      LAYER li1 ;
        RECT 17.770 42.770 17.845 42.910 ;
        RECT 17.770 41.420 17.845 41.560 ;
        RECT 17.770 40.070 17.845 40.210 ;
        RECT 17.770 38.720 17.845 38.860 ;
        RECT 17.770 37.370 17.845 37.510 ;
        RECT 17.770 36.020 17.845 36.160 ;
        RECT 17.770 34.670 17.845 34.810 ;
        RECT 17.770 33.320 17.845 33.460 ;
        RECT 17.770 31.970 17.845 32.110 ;
        RECT 17.770 30.620 17.845 30.760 ;
        RECT 17.770 29.270 17.845 29.410 ;
        RECT 17.770 27.920 17.845 28.060 ;
        RECT 17.770 26.570 17.845 26.710 ;
        RECT 17.770 25.220 17.845 25.360 ;
        RECT 17.770 23.870 17.845 24.010 ;
        RECT 17.770 22.520 17.845 22.660 ;
        RECT 17.770 21.170 17.845 21.310 ;
        RECT 17.770 19.820 17.845 19.960 ;
        RECT 17.770 18.470 17.845 18.610 ;
        RECT 17.770 17.120 17.845 17.260 ;
        RECT 17.770 15.770 17.845 15.910 ;
        RECT 17.770 14.420 17.845 14.560 ;
        RECT 17.770 13.070 17.845 13.210 ;
        RECT 17.770 11.720 17.845 11.860 ;
        RECT 17.770 10.370 17.845 10.510 ;
        RECT 17.770 9.020 17.845 9.160 ;
        RECT 17.770 7.670 17.845 7.810 ;
        RECT 17.770 6.320 17.845 6.460 ;
        RECT 17.770 4.970 17.845 5.110 ;
        RECT 17.770 3.620 17.845 3.760 ;
        RECT 17.770 2.270 17.845 2.410 ;
        RECT 17.770 0.920 17.845 1.060 ;
    END
  END WBLb_22
  PIN WBL_23
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.773600 ;
    PORT
      LAYER li1 ;
        RECT 69.020 42.770 69.095 42.915 ;
        RECT 69.020 41.420 69.095 41.565 ;
        RECT 69.020 40.070 69.095 40.215 ;
        RECT 69.020 38.720 69.095 38.865 ;
        RECT 69.020 37.370 69.095 37.515 ;
        RECT 69.020 36.020 69.095 36.165 ;
        RECT 69.020 34.670 69.095 34.815 ;
        RECT 69.020 33.320 69.095 33.465 ;
        RECT 69.020 31.970 69.095 32.115 ;
        RECT 69.020 30.620 69.095 30.765 ;
        RECT 69.020 29.270 69.095 29.415 ;
        RECT 69.020 27.920 69.095 28.065 ;
        RECT 69.020 26.570 69.095 26.715 ;
        RECT 69.020 25.220 69.095 25.365 ;
        RECT 69.020 23.870 69.095 24.015 ;
        RECT 69.020 22.520 69.095 22.665 ;
        RECT 69.020 21.170 69.095 21.315 ;
        RECT 69.020 19.820 69.095 19.965 ;
        RECT 69.020 18.470 69.095 18.615 ;
        RECT 69.020 17.120 69.095 17.265 ;
        RECT 69.020 15.770 69.095 15.915 ;
        RECT 69.020 14.420 69.095 14.565 ;
        RECT 69.020 13.070 69.095 13.215 ;
        RECT 69.020 11.720 69.095 11.865 ;
        RECT 69.020 10.370 69.095 10.515 ;
        RECT 69.020 9.020 69.095 9.165 ;
        RECT 69.020 7.670 69.095 7.815 ;
        RECT 69.020 6.320 69.095 6.465 ;
        RECT 69.020 4.970 69.095 5.115 ;
        RECT 69.020 3.620 69.095 3.765 ;
        RECT 69.020 2.275 69.095 2.420 ;
        RECT 69.020 0.925 69.095 1.070 ;
    END
    PORT
      LAYER li1 ;
        RECT 22.620 42.770 22.695 42.915 ;
        RECT 22.620 41.420 22.695 41.565 ;
        RECT 22.620 40.070 22.695 40.215 ;
        RECT 22.620 38.720 22.695 38.865 ;
        RECT 22.620 37.370 22.695 37.515 ;
        RECT 22.620 36.020 22.695 36.165 ;
        RECT 22.620 34.670 22.695 34.815 ;
        RECT 22.620 33.320 22.695 33.465 ;
        RECT 22.620 31.970 22.695 32.115 ;
        RECT 22.620 30.620 22.695 30.765 ;
        RECT 22.620 29.270 22.695 29.415 ;
        RECT 22.620 27.920 22.695 28.065 ;
        RECT 22.620 26.570 22.695 26.715 ;
        RECT 22.620 25.220 22.695 25.365 ;
        RECT 22.620 23.870 22.695 24.015 ;
        RECT 22.620 22.520 22.695 22.665 ;
        RECT 22.620 21.170 22.695 21.315 ;
        RECT 22.620 19.820 22.695 19.965 ;
        RECT 22.620 18.470 22.695 18.615 ;
        RECT 22.620 17.120 22.695 17.265 ;
        RECT 22.620 15.770 22.695 15.915 ;
        RECT 22.620 14.420 22.695 14.565 ;
        RECT 22.620 13.070 22.695 13.215 ;
        RECT 22.620 11.720 22.695 11.865 ;
        RECT 22.620 10.370 22.695 10.515 ;
        RECT 22.620 9.020 22.695 9.165 ;
        RECT 22.620 7.670 22.695 7.815 ;
        RECT 22.620 6.320 22.695 6.465 ;
        RECT 22.620 4.970 22.695 5.115 ;
        RECT 22.620 3.620 22.695 3.765 ;
        RECT 22.620 2.270 22.695 2.415 ;
        RECT 22.620 0.920 22.695 1.065 ;
    END
  END WBL_23
  PIN WBLb_23
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.739200 ;
    PORT
      LAYER li1 ;
        RECT 67.070 42.770 67.145 42.910 ;
        RECT 67.070 41.420 67.145 41.560 ;
        RECT 67.070 40.070 67.145 40.210 ;
        RECT 67.070 38.720 67.145 38.860 ;
        RECT 67.070 37.370 67.145 37.510 ;
        RECT 67.070 36.020 67.145 36.160 ;
        RECT 67.070 34.670 67.145 34.810 ;
        RECT 67.070 33.320 67.145 33.460 ;
        RECT 67.070 31.970 67.145 32.110 ;
        RECT 67.070 30.620 67.145 30.760 ;
        RECT 67.070 29.270 67.145 29.410 ;
        RECT 67.070 27.920 67.145 28.060 ;
        RECT 67.070 26.570 67.145 26.710 ;
        RECT 67.070 25.220 67.145 25.360 ;
        RECT 67.070 23.870 67.145 24.010 ;
        RECT 67.070 22.520 67.145 22.660 ;
        RECT 67.070 21.170 67.145 21.310 ;
        RECT 67.070 19.820 67.145 19.960 ;
        RECT 67.070 18.470 67.145 18.610 ;
        RECT 67.070 17.120 67.145 17.260 ;
        RECT 67.070 15.770 67.145 15.910 ;
        RECT 67.070 14.420 67.145 14.560 ;
        RECT 67.070 13.070 67.145 13.210 ;
        RECT 67.070 11.720 67.145 11.860 ;
        RECT 67.070 10.370 67.145 10.510 ;
        RECT 67.070 9.020 67.145 9.160 ;
        RECT 67.070 7.670 67.145 7.810 ;
        RECT 67.070 6.320 67.145 6.460 ;
        RECT 67.070 4.970 67.145 5.110 ;
        RECT 67.070 3.620 67.145 3.760 ;
        RECT 67.070 2.275 67.145 2.415 ;
        RECT 67.070 0.925 67.145 1.065 ;
    END
    PORT
      LAYER li1 ;
        RECT 20.670 42.770 20.745 42.910 ;
        RECT 20.670 41.420 20.745 41.560 ;
        RECT 20.670 40.070 20.745 40.210 ;
        RECT 20.670 38.720 20.745 38.860 ;
        RECT 20.670 37.370 20.745 37.510 ;
        RECT 20.670 36.020 20.745 36.160 ;
        RECT 20.670 34.670 20.745 34.810 ;
        RECT 20.670 33.320 20.745 33.460 ;
        RECT 20.670 31.970 20.745 32.110 ;
        RECT 20.670 30.620 20.745 30.760 ;
        RECT 20.670 29.270 20.745 29.410 ;
        RECT 20.670 27.920 20.745 28.060 ;
        RECT 20.670 26.570 20.745 26.710 ;
        RECT 20.670 25.220 20.745 25.360 ;
        RECT 20.670 23.870 20.745 24.010 ;
        RECT 20.670 22.520 20.745 22.660 ;
        RECT 20.670 21.170 20.745 21.310 ;
        RECT 20.670 19.820 20.745 19.960 ;
        RECT 20.670 18.470 20.745 18.610 ;
        RECT 20.670 17.120 20.745 17.260 ;
        RECT 20.670 15.770 20.745 15.910 ;
        RECT 20.670 14.420 20.745 14.560 ;
        RECT 20.670 13.070 20.745 13.210 ;
        RECT 20.670 11.720 20.745 11.860 ;
        RECT 20.670 10.370 20.745 10.510 ;
        RECT 20.670 9.020 20.745 9.160 ;
        RECT 20.670 7.670 20.745 7.810 ;
        RECT 20.670 6.320 20.745 6.460 ;
        RECT 20.670 4.970 20.745 5.110 ;
        RECT 20.670 3.620 20.745 3.760 ;
        RECT 20.670 2.270 20.745 2.410 ;
        RECT 20.670 0.920 20.745 1.060 ;
    END
  END WBLb_23
  PIN WBL_8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.773975 ;
    PORT
      LAYER li1 ;
        RECT 25.520 42.770 25.595 42.915 ;
        RECT 25.520 41.420 25.595 41.565 ;
        RECT 25.520 40.070 25.595 40.215 ;
        RECT 25.520 38.720 25.595 38.865 ;
        RECT 25.520 37.370 25.595 37.515 ;
        RECT 25.520 36.020 25.595 36.165 ;
        RECT 25.520 34.670 25.595 34.815 ;
        RECT 25.520 33.320 25.595 33.465 ;
        RECT 25.520 31.970 25.595 32.115 ;
        RECT 25.520 30.620 25.595 30.765 ;
        RECT 25.520 29.270 25.595 29.415 ;
        RECT 25.520 27.920 25.595 28.065 ;
        RECT 25.520 26.570 25.595 26.715 ;
        RECT 25.520 25.220 25.595 25.365 ;
        RECT 25.520 23.870 25.595 24.015 ;
        RECT 25.520 22.520 25.595 22.665 ;
        RECT 25.520 21.170 25.595 21.315 ;
        RECT 25.520 19.820 25.595 19.965 ;
        RECT 25.520 18.470 25.595 18.615 ;
        RECT 25.520 17.120 25.595 17.265 ;
        RECT 25.520 15.770 25.595 15.915 ;
        RECT 25.520 14.420 25.595 14.565 ;
        RECT 25.520 13.070 25.595 13.215 ;
        RECT 25.520 11.720 25.595 11.865 ;
        RECT 25.520 10.370 25.595 10.515 ;
        RECT 25.520 9.020 25.595 9.165 ;
        RECT 25.520 7.670 25.595 7.815 ;
        RECT 25.520 6.320 25.595 6.465 ;
        RECT 25.520 4.970 25.595 5.115 ;
        RECT 25.520 3.620 25.595 3.765 ;
        RECT 25.520 2.275 25.595 2.420 ;
        RECT 25.520 0.920 25.595 1.070 ;
    END
    PORT
      LAYER li1 ;
        RECT 71.920 42.770 71.995 42.915 ;
        RECT 71.920 41.420 71.995 41.565 ;
        RECT 71.920 40.070 71.995 40.215 ;
        RECT 71.920 38.720 71.995 38.865 ;
        RECT 71.920 37.370 71.995 37.515 ;
        RECT 71.920 36.020 71.995 36.165 ;
        RECT 71.920 34.670 71.995 34.815 ;
        RECT 71.920 33.320 71.995 33.465 ;
        RECT 71.920 31.970 71.995 32.115 ;
        RECT 71.920 30.620 71.995 30.765 ;
        RECT 71.920 29.270 71.995 29.415 ;
        RECT 71.920 27.920 71.995 28.065 ;
        RECT 71.920 26.570 71.995 26.715 ;
        RECT 71.920 25.220 71.995 25.365 ;
        RECT 71.920 23.870 71.995 24.015 ;
        RECT 71.920 22.520 71.995 22.665 ;
        RECT 71.920 21.170 71.995 21.315 ;
        RECT 71.920 19.820 71.995 19.965 ;
        RECT 71.920 18.470 71.995 18.615 ;
        RECT 71.920 17.120 71.995 17.265 ;
        RECT 71.920 15.770 71.995 15.915 ;
        RECT 71.920 14.420 71.995 14.565 ;
        RECT 71.920 13.070 71.995 13.215 ;
        RECT 71.920 11.720 71.995 11.865 ;
        RECT 71.920 10.370 71.995 10.515 ;
        RECT 71.920 9.020 71.995 9.165 ;
        RECT 71.920 7.670 71.995 7.815 ;
        RECT 71.920 6.320 71.995 6.465 ;
        RECT 71.920 4.970 71.995 5.115 ;
        RECT 71.920 3.620 71.995 3.765 ;
        RECT 71.920 2.275 71.995 2.420 ;
        RECT 71.920 0.925 71.995 1.070 ;
    END
  END WBL_8
  PIN WBLb_8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.739200 ;
    PORT
      LAYER li1 ;
        RECT 23.570 42.770 23.645 42.910 ;
        RECT 23.570 41.420 23.645 41.560 ;
        RECT 23.570 40.070 23.645 40.210 ;
        RECT 23.570 38.720 23.645 38.860 ;
        RECT 23.570 37.370 23.645 37.510 ;
        RECT 23.570 36.020 23.645 36.160 ;
        RECT 23.570 34.670 23.645 34.810 ;
        RECT 23.570 33.320 23.645 33.460 ;
        RECT 23.570 31.970 23.645 32.110 ;
        RECT 23.570 30.620 23.645 30.760 ;
        RECT 23.570 29.270 23.645 29.410 ;
        RECT 23.570 27.920 23.645 28.060 ;
        RECT 23.570 26.570 23.645 26.710 ;
        RECT 23.570 25.220 23.645 25.360 ;
        RECT 23.570 23.870 23.645 24.010 ;
        RECT 23.570 22.520 23.645 22.660 ;
        RECT 23.570 21.170 23.645 21.310 ;
        RECT 23.570 19.820 23.645 19.960 ;
        RECT 23.570 18.470 23.645 18.610 ;
        RECT 23.570 17.120 23.645 17.260 ;
        RECT 23.570 15.770 23.645 15.910 ;
        RECT 23.570 14.420 23.645 14.560 ;
        RECT 23.570 13.070 23.645 13.210 ;
        RECT 23.570 11.720 23.645 11.860 ;
        RECT 23.570 10.370 23.645 10.510 ;
        RECT 23.570 9.020 23.645 9.160 ;
        RECT 23.570 7.670 23.645 7.810 ;
        RECT 23.570 6.320 23.645 6.460 ;
        RECT 23.570 4.970 23.645 5.110 ;
        RECT 23.570 3.620 23.645 3.760 ;
        RECT 23.570 2.275 23.645 2.415 ;
        RECT 23.570 0.925 23.645 1.065 ;
    END
    PORT
      LAYER li1 ;
        RECT 69.970 42.770 70.045 42.910 ;
        RECT 69.970 41.420 70.045 41.560 ;
        RECT 69.970 40.070 70.045 40.210 ;
        RECT 69.970 38.720 70.045 38.860 ;
        RECT 69.970 37.370 70.045 37.510 ;
        RECT 69.970 36.020 70.045 36.160 ;
        RECT 69.970 34.670 70.045 34.810 ;
        RECT 69.970 33.320 70.045 33.460 ;
        RECT 69.970 31.970 70.045 32.110 ;
        RECT 69.970 30.620 70.045 30.760 ;
        RECT 69.970 29.270 70.045 29.410 ;
        RECT 69.970 27.920 70.045 28.060 ;
        RECT 69.970 26.570 70.045 26.710 ;
        RECT 69.970 25.220 70.045 25.360 ;
        RECT 69.970 23.870 70.045 24.010 ;
        RECT 69.970 22.520 70.045 22.660 ;
        RECT 69.970 21.170 70.045 21.310 ;
        RECT 69.970 19.820 70.045 19.960 ;
        RECT 69.970 18.470 70.045 18.610 ;
        RECT 69.970 17.120 70.045 17.260 ;
        RECT 69.970 15.770 70.045 15.910 ;
        RECT 69.970 14.420 70.045 14.560 ;
        RECT 69.970 13.070 70.045 13.210 ;
        RECT 69.970 11.720 70.045 11.860 ;
        RECT 69.970 10.370 70.045 10.510 ;
        RECT 69.970 9.020 70.045 9.160 ;
        RECT 69.970 7.670 70.045 7.810 ;
        RECT 69.970 6.320 70.045 6.460 ;
        RECT 69.970 4.970 70.045 5.110 ;
        RECT 69.970 3.620 70.045 3.760 ;
        RECT 69.970 2.275 70.045 2.415 ;
        RECT 69.970 0.925 70.045 1.065 ;
    END
  END WBLb_8
  PIN WBL_9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.773975 ;
    PORT
      LAYER li1 ;
        RECT 28.420 42.770 28.495 42.915 ;
        RECT 28.420 41.420 28.495 41.565 ;
        RECT 28.420 40.070 28.495 40.215 ;
        RECT 28.420 38.720 28.495 38.865 ;
        RECT 28.420 37.370 28.495 37.515 ;
        RECT 28.420 36.020 28.495 36.165 ;
        RECT 28.420 34.670 28.495 34.815 ;
        RECT 28.420 33.320 28.495 33.465 ;
        RECT 28.420 31.970 28.495 32.115 ;
        RECT 28.420 30.620 28.495 30.765 ;
        RECT 28.420 29.270 28.495 29.415 ;
        RECT 28.420 27.920 28.495 28.065 ;
        RECT 28.420 26.570 28.495 26.715 ;
        RECT 28.420 25.220 28.495 25.365 ;
        RECT 28.420 23.870 28.495 24.015 ;
        RECT 28.420 22.520 28.495 22.665 ;
        RECT 28.420 21.170 28.495 21.315 ;
        RECT 28.420 19.820 28.495 19.965 ;
        RECT 28.420 18.470 28.495 18.615 ;
        RECT 28.420 17.120 28.495 17.265 ;
        RECT 28.420 15.770 28.495 15.915 ;
        RECT 28.420 14.420 28.495 14.565 ;
        RECT 28.420 13.070 28.495 13.215 ;
        RECT 28.420 11.720 28.495 11.865 ;
        RECT 28.420 10.370 28.495 10.515 ;
        RECT 28.420 9.020 28.495 9.165 ;
        RECT 28.420 7.670 28.495 7.815 ;
        RECT 28.420 6.320 28.495 6.465 ;
        RECT 28.420 4.970 28.495 5.115 ;
        RECT 28.420 3.620 28.495 3.765 ;
        RECT 28.420 2.275 28.495 2.420 ;
        RECT 28.420 0.920 28.495 1.070 ;
    END
    PORT
      LAYER li1 ;
        RECT 74.820 42.770 74.895 42.915 ;
        RECT 74.820 41.420 74.895 41.565 ;
        RECT 74.820 40.070 74.895 40.215 ;
        RECT 74.820 38.720 74.895 38.865 ;
        RECT 74.820 37.370 74.895 37.515 ;
        RECT 74.820 36.020 74.895 36.165 ;
        RECT 74.820 34.670 74.895 34.815 ;
        RECT 74.820 33.320 74.895 33.465 ;
        RECT 74.820 31.970 74.895 32.115 ;
        RECT 74.820 30.620 74.895 30.765 ;
        RECT 74.820 29.270 74.895 29.415 ;
        RECT 74.820 27.920 74.895 28.065 ;
        RECT 74.820 26.570 74.895 26.715 ;
        RECT 74.820 25.220 74.895 25.365 ;
        RECT 74.820 23.870 74.895 24.015 ;
        RECT 74.820 22.520 74.895 22.665 ;
        RECT 74.820 21.170 74.895 21.315 ;
        RECT 74.820 19.820 74.895 19.965 ;
        RECT 74.820 18.470 74.895 18.615 ;
        RECT 74.820 17.120 74.895 17.265 ;
        RECT 74.820 15.770 74.895 15.915 ;
        RECT 74.820 14.420 74.895 14.565 ;
        RECT 74.820 13.070 74.895 13.215 ;
        RECT 74.820 11.720 74.895 11.865 ;
        RECT 74.820 10.370 74.895 10.515 ;
        RECT 74.820 9.020 74.895 9.165 ;
        RECT 74.820 7.670 74.895 7.815 ;
        RECT 74.820 6.320 74.895 6.465 ;
        RECT 74.820 4.970 74.895 5.115 ;
        RECT 74.820 3.620 74.895 3.765 ;
        RECT 74.820 2.275 74.895 2.420 ;
        RECT 74.820 0.925 74.895 1.070 ;
    END
  END WBL_9
  PIN WBLb_9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.739575 ;
    PORT
      LAYER li1 ;
        RECT 26.470 42.770 26.545 42.910 ;
        RECT 26.470 41.420 26.545 41.560 ;
        RECT 26.470 40.070 26.545 40.210 ;
        RECT 26.470 38.720 26.545 38.860 ;
        RECT 26.470 37.370 26.545 37.510 ;
        RECT 26.470 36.020 26.545 36.160 ;
        RECT 26.470 34.670 26.545 34.810 ;
        RECT 26.470 33.320 26.545 33.460 ;
        RECT 26.470 31.970 26.545 32.110 ;
        RECT 26.470 30.620 26.545 30.760 ;
        RECT 26.470 29.270 26.545 29.410 ;
        RECT 26.470 27.920 26.545 28.060 ;
        RECT 26.470 26.570 26.545 26.710 ;
        RECT 26.470 25.220 26.545 25.360 ;
        RECT 26.470 23.870 26.545 24.010 ;
        RECT 26.470 22.520 26.545 22.660 ;
        RECT 26.470 21.170 26.545 21.310 ;
        RECT 26.470 19.820 26.545 19.960 ;
        RECT 26.470 18.470 26.545 18.610 ;
        RECT 26.470 17.120 26.545 17.260 ;
        RECT 26.470 15.770 26.545 15.910 ;
        RECT 26.470 14.420 26.545 14.560 ;
        RECT 26.470 13.070 26.545 13.210 ;
        RECT 26.470 11.720 26.545 11.860 ;
        RECT 26.470 10.370 26.545 10.510 ;
        RECT 26.470 9.020 26.545 9.160 ;
        RECT 26.470 7.670 26.545 7.810 ;
        RECT 26.470 6.320 26.545 6.460 ;
        RECT 26.470 4.970 26.545 5.110 ;
        RECT 26.470 3.620 26.545 3.760 ;
        RECT 26.470 2.275 26.545 2.415 ;
        RECT 26.470 0.920 26.545 1.065 ;
    END
    PORT
      LAYER li1 ;
        RECT 72.870 42.770 72.945 42.910 ;
        RECT 72.870 41.420 72.945 41.560 ;
        RECT 72.870 40.070 72.945 40.210 ;
        RECT 72.870 38.720 72.945 38.860 ;
        RECT 72.870 37.370 72.945 37.510 ;
        RECT 72.870 36.020 72.945 36.160 ;
        RECT 72.870 34.670 72.945 34.810 ;
        RECT 72.870 33.320 72.945 33.460 ;
        RECT 72.870 31.970 72.945 32.110 ;
        RECT 72.870 30.620 72.945 30.760 ;
        RECT 72.870 29.270 72.945 29.410 ;
        RECT 72.870 27.920 72.945 28.060 ;
        RECT 72.870 26.570 72.945 26.710 ;
        RECT 72.870 25.220 72.945 25.360 ;
        RECT 72.870 23.870 72.945 24.010 ;
        RECT 72.870 22.520 72.945 22.660 ;
        RECT 72.870 21.170 72.945 21.310 ;
        RECT 72.870 19.820 72.945 19.960 ;
        RECT 72.870 18.470 72.945 18.610 ;
        RECT 72.870 17.120 72.945 17.260 ;
        RECT 72.870 15.770 72.945 15.910 ;
        RECT 72.870 14.420 72.945 14.560 ;
        RECT 72.870 13.070 72.945 13.210 ;
        RECT 72.870 11.720 72.945 11.860 ;
        RECT 72.870 10.370 72.945 10.510 ;
        RECT 72.870 9.020 72.945 9.160 ;
        RECT 72.870 7.670 72.945 7.810 ;
        RECT 72.870 6.320 72.945 6.460 ;
        RECT 72.870 4.970 72.945 5.110 ;
        RECT 72.870 3.620 72.945 3.760 ;
        RECT 72.870 2.275 72.945 2.415 ;
        RECT 72.870 0.925 72.945 1.065 ;
    END
  END WBLb_9
  PIN WBL_10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.773975 ;
    PORT
      LAYER li1 ;
        RECT 31.320 42.770 31.395 42.915 ;
        RECT 31.320 41.420 31.395 41.565 ;
        RECT 31.320 40.070 31.395 40.215 ;
        RECT 31.320 38.720 31.395 38.865 ;
        RECT 31.320 37.370 31.395 37.515 ;
        RECT 31.320 36.020 31.395 36.165 ;
        RECT 31.320 34.670 31.395 34.815 ;
        RECT 31.320 33.320 31.395 33.465 ;
        RECT 31.320 31.970 31.395 32.115 ;
        RECT 31.320 30.620 31.395 30.765 ;
        RECT 31.320 29.270 31.395 29.415 ;
        RECT 31.320 27.920 31.395 28.065 ;
        RECT 31.320 26.570 31.395 26.715 ;
        RECT 31.320 25.220 31.395 25.365 ;
        RECT 31.320 23.870 31.395 24.015 ;
        RECT 31.320 22.520 31.395 22.665 ;
        RECT 31.320 21.170 31.395 21.315 ;
        RECT 31.320 19.820 31.395 19.965 ;
        RECT 31.320 18.470 31.395 18.615 ;
        RECT 31.320 17.120 31.395 17.265 ;
        RECT 31.320 15.770 31.395 15.915 ;
        RECT 31.320 14.420 31.395 14.565 ;
        RECT 31.320 13.070 31.395 13.215 ;
        RECT 31.320 11.720 31.395 11.865 ;
        RECT 31.320 10.370 31.395 10.515 ;
        RECT 31.320 9.020 31.395 9.165 ;
        RECT 31.320 7.670 31.395 7.815 ;
        RECT 31.320 6.320 31.395 6.465 ;
        RECT 31.320 4.970 31.395 5.115 ;
        RECT 31.320 3.620 31.395 3.765 ;
        RECT 31.320 2.275 31.395 2.420 ;
        RECT 31.320 0.920 31.395 1.070 ;
    END
    PORT
      LAYER li1 ;
        RECT 77.720 42.770 77.795 42.915 ;
        RECT 77.720 41.420 77.795 41.565 ;
        RECT 77.720 40.070 77.795 40.215 ;
        RECT 77.720 38.720 77.795 38.865 ;
        RECT 77.720 37.370 77.795 37.515 ;
        RECT 77.720 36.020 77.795 36.165 ;
        RECT 77.720 34.670 77.795 34.815 ;
        RECT 77.720 33.320 77.795 33.465 ;
        RECT 77.720 31.970 77.795 32.115 ;
        RECT 77.720 30.620 77.795 30.765 ;
        RECT 77.720 29.270 77.795 29.415 ;
        RECT 77.720 27.920 77.795 28.065 ;
        RECT 77.720 26.570 77.795 26.715 ;
        RECT 77.720 25.220 77.795 25.365 ;
        RECT 77.720 23.870 77.795 24.015 ;
        RECT 77.720 22.520 77.795 22.665 ;
        RECT 77.720 21.170 77.795 21.315 ;
        RECT 77.720 19.820 77.795 19.965 ;
        RECT 77.720 18.470 77.795 18.615 ;
        RECT 77.720 17.120 77.795 17.265 ;
        RECT 77.720 15.770 77.795 15.915 ;
        RECT 77.720 14.420 77.795 14.565 ;
        RECT 77.720 13.070 77.795 13.215 ;
        RECT 77.720 11.720 77.795 11.865 ;
        RECT 77.720 10.370 77.795 10.515 ;
        RECT 77.720 9.020 77.795 9.165 ;
        RECT 77.720 7.670 77.795 7.815 ;
        RECT 77.720 6.320 77.795 6.465 ;
        RECT 77.720 4.970 77.795 5.115 ;
        RECT 77.720 3.620 77.795 3.765 ;
        RECT 77.720 2.275 77.795 2.420 ;
        RECT 77.720 0.925 77.795 1.070 ;
    END
  END WBL_10
  PIN WBLb_10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.739575 ;
    PORT
      LAYER li1 ;
        RECT 29.370 42.770 29.445 42.910 ;
        RECT 29.370 41.420 29.445 41.560 ;
        RECT 29.370 40.070 29.445 40.210 ;
        RECT 29.370 38.720 29.445 38.860 ;
        RECT 29.370 37.370 29.445 37.510 ;
        RECT 29.370 36.020 29.445 36.160 ;
        RECT 29.370 34.670 29.445 34.810 ;
        RECT 29.370 33.320 29.445 33.460 ;
        RECT 29.370 31.970 29.445 32.110 ;
        RECT 29.370 30.620 29.445 30.760 ;
        RECT 29.370 29.270 29.445 29.410 ;
        RECT 29.370 27.920 29.445 28.060 ;
        RECT 29.370 26.570 29.445 26.710 ;
        RECT 29.370 25.220 29.445 25.360 ;
        RECT 29.370 23.870 29.445 24.010 ;
        RECT 29.370 22.520 29.445 22.660 ;
        RECT 29.370 21.170 29.445 21.310 ;
        RECT 29.370 19.820 29.445 19.960 ;
        RECT 29.370 18.470 29.445 18.610 ;
        RECT 29.370 17.120 29.445 17.260 ;
        RECT 29.370 15.770 29.445 15.910 ;
        RECT 29.370 14.420 29.445 14.560 ;
        RECT 29.370 13.070 29.445 13.210 ;
        RECT 29.370 11.720 29.445 11.860 ;
        RECT 29.370 10.370 29.445 10.510 ;
        RECT 29.370 9.020 29.445 9.160 ;
        RECT 29.370 7.670 29.445 7.810 ;
        RECT 29.370 6.320 29.445 6.460 ;
        RECT 29.370 4.970 29.445 5.110 ;
        RECT 29.370 3.620 29.445 3.760 ;
        RECT 29.370 2.275 29.445 2.415 ;
        RECT 29.370 0.920 29.445 1.065 ;
    END
    PORT
      LAYER li1 ;
        RECT 75.770 42.770 75.845 42.910 ;
        RECT 75.770 41.420 75.845 41.560 ;
        RECT 75.770 40.070 75.845 40.210 ;
        RECT 75.770 38.720 75.845 38.860 ;
        RECT 75.770 37.370 75.845 37.510 ;
        RECT 75.770 36.020 75.845 36.160 ;
        RECT 75.770 34.670 75.845 34.810 ;
        RECT 75.770 33.320 75.845 33.460 ;
        RECT 75.770 31.970 75.845 32.110 ;
        RECT 75.770 30.620 75.845 30.760 ;
        RECT 75.770 29.270 75.845 29.410 ;
        RECT 75.770 27.920 75.845 28.060 ;
        RECT 75.770 26.570 75.845 26.710 ;
        RECT 75.770 25.220 75.845 25.360 ;
        RECT 75.770 23.870 75.845 24.010 ;
        RECT 75.770 22.520 75.845 22.660 ;
        RECT 75.770 21.170 75.845 21.310 ;
        RECT 75.770 19.820 75.845 19.960 ;
        RECT 75.770 18.470 75.845 18.610 ;
        RECT 75.770 17.120 75.845 17.260 ;
        RECT 75.770 15.770 75.845 15.910 ;
        RECT 75.770 14.420 75.845 14.560 ;
        RECT 75.770 13.070 75.845 13.210 ;
        RECT 75.770 11.720 75.845 11.860 ;
        RECT 75.770 10.370 75.845 10.510 ;
        RECT 75.770 9.020 75.845 9.160 ;
        RECT 75.770 7.670 75.845 7.810 ;
        RECT 75.770 6.320 75.845 6.460 ;
        RECT 75.770 4.970 75.845 5.110 ;
        RECT 75.770 3.620 75.845 3.760 ;
        RECT 75.770 2.275 75.845 2.415 ;
        RECT 75.770 0.925 75.845 1.065 ;
    END
  END WBLb_10
  PIN WBL_11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.773975 ;
    PORT
      LAYER li1 ;
        RECT 34.220 42.770 34.295 42.915 ;
        RECT 34.220 41.420 34.295 41.565 ;
        RECT 34.220 40.070 34.295 40.215 ;
        RECT 34.220 38.720 34.295 38.865 ;
        RECT 34.220 37.370 34.295 37.515 ;
        RECT 34.220 36.020 34.295 36.165 ;
        RECT 34.220 34.670 34.295 34.815 ;
        RECT 34.220 33.320 34.295 33.465 ;
        RECT 34.220 31.970 34.295 32.115 ;
        RECT 34.220 30.620 34.295 30.765 ;
        RECT 34.220 29.270 34.295 29.415 ;
        RECT 34.220 27.920 34.295 28.065 ;
        RECT 34.220 26.570 34.295 26.715 ;
        RECT 34.220 25.220 34.295 25.365 ;
        RECT 34.220 23.870 34.295 24.015 ;
        RECT 34.220 22.520 34.295 22.665 ;
        RECT 34.220 21.170 34.295 21.315 ;
        RECT 34.220 19.820 34.295 19.965 ;
        RECT 34.220 18.470 34.295 18.615 ;
        RECT 34.220 17.120 34.295 17.265 ;
        RECT 34.220 15.770 34.295 15.915 ;
        RECT 34.220 14.420 34.295 14.565 ;
        RECT 34.220 13.070 34.295 13.215 ;
        RECT 34.220 11.720 34.295 11.865 ;
        RECT 34.220 10.370 34.295 10.515 ;
        RECT 34.220 9.020 34.295 9.165 ;
        RECT 34.220 7.670 34.295 7.815 ;
        RECT 34.220 6.320 34.295 6.465 ;
        RECT 34.220 4.970 34.295 5.115 ;
        RECT 34.220 3.620 34.295 3.765 ;
        RECT 34.220 2.275 34.295 2.420 ;
        RECT 34.220 0.920 34.295 1.070 ;
    END
    PORT
      LAYER li1 ;
        RECT 80.620 42.770 80.695 42.915 ;
        RECT 80.620 41.420 80.695 41.565 ;
        RECT 80.620 40.070 80.695 40.215 ;
        RECT 80.620 38.720 80.695 38.865 ;
        RECT 80.620 37.370 80.695 37.515 ;
        RECT 80.620 36.020 80.695 36.165 ;
        RECT 80.620 34.670 80.695 34.815 ;
        RECT 80.620 33.320 80.695 33.465 ;
        RECT 80.620 31.970 80.695 32.115 ;
        RECT 80.620 30.620 80.695 30.765 ;
        RECT 80.620 29.270 80.695 29.415 ;
        RECT 80.620 27.920 80.695 28.065 ;
        RECT 80.620 26.570 80.695 26.715 ;
        RECT 80.620 25.220 80.695 25.365 ;
        RECT 80.620 23.870 80.695 24.015 ;
        RECT 80.620 22.520 80.695 22.665 ;
        RECT 80.620 21.170 80.695 21.315 ;
        RECT 80.620 19.820 80.695 19.965 ;
        RECT 80.620 18.470 80.695 18.615 ;
        RECT 80.620 17.120 80.695 17.265 ;
        RECT 80.620 15.770 80.695 15.915 ;
        RECT 80.620 14.420 80.695 14.565 ;
        RECT 80.620 13.070 80.695 13.215 ;
        RECT 80.620 11.720 80.695 11.865 ;
        RECT 80.620 10.370 80.695 10.515 ;
        RECT 80.620 9.020 80.695 9.165 ;
        RECT 80.620 7.670 80.695 7.815 ;
        RECT 80.620 6.320 80.695 6.465 ;
        RECT 80.620 4.970 80.695 5.115 ;
        RECT 80.620 3.620 80.695 3.765 ;
        RECT 80.620 2.275 80.695 2.420 ;
        RECT 80.620 0.925 80.695 1.070 ;
    END
  END WBL_11
  PIN WBLb_11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.739575 ;
    PORT
      LAYER li1 ;
        RECT 32.270 42.770 32.345 42.910 ;
        RECT 32.270 41.420 32.345 41.560 ;
        RECT 32.270 40.070 32.345 40.210 ;
        RECT 32.270 38.720 32.345 38.860 ;
        RECT 32.270 37.370 32.345 37.510 ;
        RECT 32.270 36.020 32.345 36.160 ;
        RECT 32.270 34.670 32.345 34.810 ;
        RECT 32.270 33.320 32.345 33.460 ;
        RECT 32.270 31.970 32.345 32.110 ;
        RECT 32.270 30.620 32.345 30.760 ;
        RECT 32.270 29.270 32.345 29.410 ;
        RECT 32.270 27.920 32.345 28.060 ;
        RECT 32.270 26.570 32.345 26.710 ;
        RECT 32.270 25.220 32.345 25.360 ;
        RECT 32.270 23.870 32.345 24.010 ;
        RECT 32.270 22.520 32.345 22.660 ;
        RECT 32.270 21.170 32.345 21.310 ;
        RECT 32.270 19.820 32.345 19.960 ;
        RECT 32.270 18.470 32.345 18.610 ;
        RECT 32.270 17.120 32.345 17.260 ;
        RECT 32.270 15.770 32.345 15.910 ;
        RECT 32.270 14.420 32.345 14.560 ;
        RECT 32.270 13.070 32.345 13.210 ;
        RECT 32.270 11.720 32.345 11.860 ;
        RECT 32.270 10.370 32.345 10.510 ;
        RECT 32.270 9.020 32.345 9.160 ;
        RECT 32.270 7.670 32.345 7.810 ;
        RECT 32.270 6.320 32.345 6.460 ;
        RECT 32.270 4.970 32.345 5.110 ;
        RECT 32.270 3.620 32.345 3.760 ;
        RECT 32.270 2.275 32.345 2.415 ;
        RECT 32.270 0.920 32.345 1.065 ;
    END
    PORT
      LAYER li1 ;
        RECT 78.670 42.770 78.745 42.910 ;
        RECT 78.670 41.420 78.745 41.560 ;
        RECT 78.670 40.070 78.745 40.210 ;
        RECT 78.670 38.720 78.745 38.860 ;
        RECT 78.670 37.370 78.745 37.510 ;
        RECT 78.670 36.020 78.745 36.160 ;
        RECT 78.670 34.670 78.745 34.810 ;
        RECT 78.670 33.320 78.745 33.460 ;
        RECT 78.670 31.970 78.745 32.110 ;
        RECT 78.670 30.620 78.745 30.760 ;
        RECT 78.670 29.270 78.745 29.410 ;
        RECT 78.670 27.920 78.745 28.060 ;
        RECT 78.670 26.570 78.745 26.710 ;
        RECT 78.670 25.220 78.745 25.360 ;
        RECT 78.670 23.870 78.745 24.010 ;
        RECT 78.670 22.520 78.745 22.660 ;
        RECT 78.670 21.170 78.745 21.310 ;
        RECT 78.670 19.820 78.745 19.960 ;
        RECT 78.670 18.470 78.745 18.610 ;
        RECT 78.670 17.120 78.745 17.260 ;
        RECT 78.670 15.770 78.745 15.910 ;
        RECT 78.670 14.420 78.745 14.560 ;
        RECT 78.670 13.070 78.745 13.210 ;
        RECT 78.670 11.720 78.745 11.860 ;
        RECT 78.670 10.370 78.745 10.510 ;
        RECT 78.670 9.020 78.745 9.160 ;
        RECT 78.670 7.670 78.745 7.810 ;
        RECT 78.670 6.320 78.745 6.460 ;
        RECT 78.670 4.970 78.745 5.110 ;
        RECT 78.670 3.620 78.745 3.760 ;
        RECT 78.670 2.275 78.745 2.415 ;
        RECT 78.670 0.925 78.745 1.065 ;
    END
  END WBLb_11
  PIN WBL_12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.773975 ;
    PORT
      LAYER li1 ;
        RECT 37.120 42.770 37.195 42.915 ;
        RECT 37.120 41.420 37.195 41.565 ;
        RECT 37.120 40.070 37.195 40.215 ;
        RECT 37.120 38.720 37.195 38.865 ;
        RECT 37.120 37.370 37.195 37.515 ;
        RECT 37.120 36.020 37.195 36.165 ;
        RECT 37.120 34.670 37.195 34.815 ;
        RECT 37.120 33.320 37.195 33.465 ;
        RECT 37.120 31.970 37.195 32.115 ;
        RECT 37.120 30.620 37.195 30.765 ;
        RECT 37.120 29.270 37.195 29.415 ;
        RECT 37.120 27.920 37.195 28.065 ;
        RECT 37.120 26.570 37.195 26.715 ;
        RECT 37.120 25.220 37.195 25.365 ;
        RECT 37.120 23.870 37.195 24.015 ;
        RECT 37.120 22.520 37.195 22.665 ;
        RECT 37.120 21.170 37.195 21.315 ;
        RECT 37.120 19.820 37.195 19.965 ;
        RECT 37.120 18.470 37.195 18.615 ;
        RECT 37.120 17.120 37.195 17.265 ;
        RECT 37.120 15.770 37.195 15.915 ;
        RECT 37.120 14.420 37.195 14.565 ;
        RECT 37.120 13.070 37.195 13.215 ;
        RECT 37.120 11.720 37.195 11.865 ;
        RECT 37.120 10.370 37.195 10.515 ;
        RECT 37.120 9.020 37.195 9.165 ;
        RECT 37.120 7.670 37.195 7.815 ;
        RECT 37.120 6.320 37.195 6.465 ;
        RECT 37.120 4.970 37.195 5.115 ;
        RECT 37.120 3.620 37.195 3.765 ;
        RECT 37.120 2.275 37.195 2.420 ;
        RECT 37.120 0.920 37.195 1.070 ;
    END
    PORT
      LAYER li1 ;
        RECT 83.520 42.770 83.595 42.915 ;
        RECT 83.520 41.420 83.595 41.565 ;
        RECT 83.520 40.070 83.595 40.215 ;
        RECT 83.520 38.720 83.595 38.865 ;
        RECT 83.520 37.370 83.595 37.515 ;
        RECT 83.520 36.020 83.595 36.165 ;
        RECT 83.520 34.670 83.595 34.815 ;
        RECT 83.520 33.320 83.595 33.465 ;
        RECT 83.520 31.970 83.595 32.115 ;
        RECT 83.520 30.620 83.595 30.765 ;
        RECT 83.520 29.270 83.595 29.415 ;
        RECT 83.520 27.920 83.595 28.065 ;
        RECT 83.520 26.570 83.595 26.715 ;
        RECT 83.520 25.220 83.595 25.365 ;
        RECT 83.520 23.870 83.595 24.015 ;
        RECT 83.520 22.520 83.595 22.665 ;
        RECT 83.520 21.170 83.595 21.315 ;
        RECT 83.520 19.820 83.595 19.965 ;
        RECT 83.520 18.470 83.595 18.615 ;
        RECT 83.520 17.120 83.595 17.265 ;
        RECT 83.520 15.770 83.595 15.915 ;
        RECT 83.520 14.420 83.595 14.565 ;
        RECT 83.520 13.070 83.595 13.215 ;
        RECT 83.520 11.720 83.595 11.865 ;
        RECT 83.520 10.370 83.595 10.515 ;
        RECT 83.520 9.020 83.595 9.165 ;
        RECT 83.520 7.670 83.595 7.815 ;
        RECT 83.520 6.320 83.595 6.465 ;
        RECT 83.520 4.970 83.595 5.115 ;
        RECT 83.520 3.620 83.595 3.765 ;
        RECT 83.520 2.275 83.595 2.420 ;
        RECT 83.520 0.925 83.595 1.070 ;
    END
  END WBL_12
  PIN WBLb_12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.739575 ;
    PORT
      LAYER li1 ;
        RECT 35.170 42.770 35.245 42.910 ;
        RECT 35.170 41.420 35.245 41.560 ;
        RECT 35.170 40.070 35.245 40.210 ;
        RECT 35.170 38.720 35.245 38.860 ;
        RECT 35.170 37.370 35.245 37.510 ;
        RECT 35.170 36.020 35.245 36.160 ;
        RECT 35.170 34.670 35.245 34.810 ;
        RECT 35.170 33.320 35.245 33.460 ;
        RECT 35.170 31.970 35.245 32.110 ;
        RECT 35.170 30.620 35.245 30.760 ;
        RECT 35.170 29.270 35.245 29.410 ;
        RECT 35.170 27.920 35.245 28.060 ;
        RECT 35.170 26.570 35.245 26.710 ;
        RECT 35.170 25.220 35.245 25.360 ;
        RECT 35.170 23.870 35.245 24.010 ;
        RECT 35.170 22.520 35.245 22.660 ;
        RECT 35.170 21.170 35.245 21.310 ;
        RECT 35.170 19.820 35.245 19.960 ;
        RECT 35.170 18.470 35.245 18.610 ;
        RECT 35.170 17.120 35.245 17.260 ;
        RECT 35.170 15.770 35.245 15.910 ;
        RECT 35.170 14.420 35.245 14.560 ;
        RECT 35.170 13.070 35.245 13.210 ;
        RECT 35.170 11.720 35.245 11.860 ;
        RECT 35.170 10.370 35.245 10.510 ;
        RECT 35.170 9.020 35.245 9.160 ;
        RECT 35.170 7.670 35.245 7.810 ;
        RECT 35.170 6.320 35.245 6.460 ;
        RECT 35.170 4.970 35.245 5.110 ;
        RECT 35.170 3.620 35.245 3.760 ;
        RECT 35.170 2.275 35.245 2.415 ;
        RECT 35.170 0.920 35.245 1.065 ;
    END
    PORT
      LAYER li1 ;
        RECT 81.570 42.770 81.645 42.910 ;
        RECT 81.570 41.420 81.645 41.560 ;
        RECT 81.570 40.070 81.645 40.210 ;
        RECT 81.570 38.720 81.645 38.860 ;
        RECT 81.570 37.370 81.645 37.510 ;
        RECT 81.570 36.020 81.645 36.160 ;
        RECT 81.570 34.670 81.645 34.810 ;
        RECT 81.570 33.320 81.645 33.460 ;
        RECT 81.570 31.970 81.645 32.110 ;
        RECT 81.570 30.620 81.645 30.760 ;
        RECT 81.570 29.270 81.645 29.410 ;
        RECT 81.570 27.920 81.645 28.060 ;
        RECT 81.570 26.570 81.645 26.710 ;
        RECT 81.570 25.220 81.645 25.360 ;
        RECT 81.570 23.870 81.645 24.010 ;
        RECT 81.570 22.520 81.645 22.660 ;
        RECT 81.570 21.170 81.645 21.310 ;
        RECT 81.570 19.820 81.645 19.960 ;
        RECT 81.570 18.470 81.645 18.610 ;
        RECT 81.570 17.120 81.645 17.260 ;
        RECT 81.570 15.770 81.645 15.910 ;
        RECT 81.570 14.420 81.645 14.560 ;
        RECT 81.570 13.070 81.645 13.210 ;
        RECT 81.570 11.720 81.645 11.860 ;
        RECT 81.570 10.370 81.645 10.510 ;
        RECT 81.570 9.020 81.645 9.160 ;
        RECT 81.570 7.670 81.645 7.810 ;
        RECT 81.570 6.320 81.645 6.460 ;
        RECT 81.570 4.970 81.645 5.110 ;
        RECT 81.570 3.620 81.645 3.760 ;
        RECT 81.570 2.275 81.645 2.415 ;
        RECT 81.570 0.925 81.645 1.065 ;
    END
  END WBLb_12
  PIN WBL_13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.773975 ;
    PORT
      LAYER li1 ;
        RECT 40.020 42.770 40.095 42.915 ;
        RECT 40.020 41.420 40.095 41.565 ;
        RECT 40.020 40.070 40.095 40.215 ;
        RECT 40.020 38.720 40.095 38.865 ;
        RECT 40.020 37.370 40.095 37.515 ;
        RECT 40.020 36.020 40.095 36.165 ;
        RECT 40.020 34.670 40.095 34.815 ;
        RECT 40.020 33.320 40.095 33.465 ;
        RECT 40.020 31.970 40.095 32.115 ;
        RECT 40.020 30.620 40.095 30.765 ;
        RECT 40.020 29.270 40.095 29.415 ;
        RECT 40.020 27.920 40.095 28.065 ;
        RECT 40.020 26.570 40.095 26.715 ;
        RECT 40.020 25.220 40.095 25.365 ;
        RECT 40.020 23.870 40.095 24.015 ;
        RECT 40.020 22.520 40.095 22.665 ;
        RECT 40.020 21.170 40.095 21.315 ;
        RECT 40.020 19.820 40.095 19.965 ;
        RECT 40.020 18.470 40.095 18.615 ;
        RECT 40.020 17.120 40.095 17.265 ;
        RECT 40.020 15.770 40.095 15.915 ;
        RECT 40.020 14.420 40.095 14.565 ;
        RECT 40.020 13.070 40.095 13.215 ;
        RECT 40.020 11.720 40.095 11.865 ;
        RECT 40.020 10.370 40.095 10.515 ;
        RECT 40.020 9.020 40.095 9.165 ;
        RECT 40.020 7.670 40.095 7.815 ;
        RECT 40.020 6.320 40.095 6.465 ;
        RECT 40.020 4.970 40.095 5.115 ;
        RECT 40.020 3.620 40.095 3.765 ;
        RECT 40.020 2.275 40.095 2.420 ;
        RECT 40.020 0.920 40.095 1.070 ;
    END
    PORT
      LAYER li1 ;
        RECT 86.420 42.770 86.495 42.915 ;
        RECT 86.420 41.420 86.495 41.565 ;
        RECT 86.420 40.070 86.495 40.215 ;
        RECT 86.420 38.720 86.495 38.865 ;
        RECT 86.420 37.370 86.495 37.515 ;
        RECT 86.420 36.020 86.495 36.165 ;
        RECT 86.420 34.670 86.495 34.815 ;
        RECT 86.420 33.320 86.495 33.465 ;
        RECT 86.420 31.970 86.495 32.115 ;
        RECT 86.420 30.620 86.495 30.765 ;
        RECT 86.420 29.270 86.495 29.415 ;
        RECT 86.420 27.920 86.495 28.065 ;
        RECT 86.420 26.570 86.495 26.715 ;
        RECT 86.420 25.220 86.495 25.365 ;
        RECT 86.420 23.870 86.495 24.015 ;
        RECT 86.420 22.520 86.495 22.665 ;
        RECT 86.420 21.170 86.495 21.315 ;
        RECT 86.420 19.820 86.495 19.965 ;
        RECT 86.420 18.470 86.495 18.615 ;
        RECT 86.420 17.120 86.495 17.265 ;
        RECT 86.420 15.770 86.495 15.915 ;
        RECT 86.420 14.420 86.495 14.565 ;
        RECT 86.420 13.070 86.495 13.215 ;
        RECT 86.420 11.720 86.495 11.865 ;
        RECT 86.420 10.370 86.495 10.515 ;
        RECT 86.420 9.020 86.495 9.165 ;
        RECT 86.420 7.670 86.495 7.815 ;
        RECT 86.420 6.320 86.495 6.465 ;
        RECT 86.420 4.970 86.495 5.115 ;
        RECT 86.420 3.620 86.495 3.765 ;
        RECT 86.420 2.275 86.495 2.420 ;
        RECT 86.420 0.925 86.495 1.070 ;
    END
  END WBL_13
  PIN WBLb_13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.739575 ;
    PORT
      LAYER li1 ;
        RECT 38.070 42.770 38.145 42.910 ;
        RECT 38.070 41.420 38.145 41.560 ;
        RECT 38.070 40.070 38.145 40.210 ;
        RECT 38.070 38.720 38.145 38.860 ;
        RECT 38.070 37.370 38.145 37.510 ;
        RECT 38.070 36.020 38.145 36.160 ;
        RECT 38.070 34.670 38.145 34.810 ;
        RECT 38.070 33.320 38.145 33.460 ;
        RECT 38.070 31.970 38.145 32.110 ;
        RECT 38.070 30.620 38.145 30.760 ;
        RECT 38.070 29.270 38.145 29.410 ;
        RECT 38.070 27.920 38.145 28.060 ;
        RECT 38.070 26.570 38.145 26.710 ;
        RECT 38.070 25.220 38.145 25.360 ;
        RECT 38.070 23.870 38.145 24.010 ;
        RECT 38.070 22.520 38.145 22.660 ;
        RECT 38.070 21.170 38.145 21.310 ;
        RECT 38.070 19.820 38.145 19.960 ;
        RECT 38.070 18.470 38.145 18.610 ;
        RECT 38.070 17.120 38.145 17.260 ;
        RECT 38.070 15.770 38.145 15.910 ;
        RECT 38.070 14.420 38.145 14.560 ;
        RECT 38.070 13.070 38.145 13.210 ;
        RECT 38.070 11.720 38.145 11.860 ;
        RECT 38.070 10.370 38.145 10.510 ;
        RECT 38.070 9.020 38.145 9.160 ;
        RECT 38.070 7.670 38.145 7.810 ;
        RECT 38.070 6.320 38.145 6.460 ;
        RECT 38.070 4.970 38.145 5.110 ;
        RECT 38.070 3.620 38.145 3.760 ;
        RECT 38.070 2.275 38.145 2.415 ;
        RECT 38.070 0.920 38.145 1.065 ;
    END
    PORT
      LAYER li1 ;
        RECT 84.470 42.770 84.545 42.910 ;
        RECT 84.470 41.420 84.545 41.560 ;
        RECT 84.470 40.070 84.545 40.210 ;
        RECT 84.470 38.720 84.545 38.860 ;
        RECT 84.470 37.370 84.545 37.510 ;
        RECT 84.470 36.020 84.545 36.160 ;
        RECT 84.470 34.670 84.545 34.810 ;
        RECT 84.470 33.320 84.545 33.460 ;
        RECT 84.470 31.970 84.545 32.110 ;
        RECT 84.470 30.620 84.545 30.760 ;
        RECT 84.470 29.270 84.545 29.410 ;
        RECT 84.470 27.920 84.545 28.060 ;
        RECT 84.470 26.570 84.545 26.710 ;
        RECT 84.470 25.220 84.545 25.360 ;
        RECT 84.470 23.870 84.545 24.010 ;
        RECT 84.470 22.520 84.545 22.660 ;
        RECT 84.470 21.170 84.545 21.310 ;
        RECT 84.470 19.820 84.545 19.960 ;
        RECT 84.470 18.470 84.545 18.610 ;
        RECT 84.470 17.120 84.545 17.260 ;
        RECT 84.470 15.770 84.545 15.910 ;
        RECT 84.470 14.420 84.545 14.560 ;
        RECT 84.470 13.070 84.545 13.210 ;
        RECT 84.470 11.720 84.545 11.860 ;
        RECT 84.470 10.370 84.545 10.510 ;
        RECT 84.470 9.020 84.545 9.160 ;
        RECT 84.470 7.670 84.545 7.810 ;
        RECT 84.470 6.320 84.545 6.460 ;
        RECT 84.470 4.970 84.545 5.110 ;
        RECT 84.470 3.620 84.545 3.760 ;
        RECT 84.470 2.275 84.545 2.415 ;
        RECT 84.470 0.925 84.545 1.065 ;
    END
  END WBLb_13
  PIN WBL_14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.773975 ;
    PORT
      LAYER li1 ;
        RECT 42.920 42.770 42.995 42.915 ;
        RECT 42.920 41.420 42.995 41.565 ;
        RECT 42.920 40.070 42.995 40.215 ;
        RECT 42.920 38.720 42.995 38.865 ;
        RECT 42.920 37.370 42.995 37.515 ;
        RECT 42.920 36.020 42.995 36.165 ;
        RECT 42.920 34.670 42.995 34.815 ;
        RECT 42.920 33.320 42.995 33.465 ;
        RECT 42.920 31.970 42.995 32.115 ;
        RECT 42.920 30.620 42.995 30.765 ;
        RECT 42.920 29.270 42.995 29.415 ;
        RECT 42.920 27.920 42.995 28.065 ;
        RECT 42.920 26.570 42.995 26.715 ;
        RECT 42.920 25.220 42.995 25.365 ;
        RECT 42.920 23.870 42.995 24.015 ;
        RECT 42.920 22.520 42.995 22.665 ;
        RECT 42.920 21.170 42.995 21.315 ;
        RECT 42.920 19.820 42.995 19.965 ;
        RECT 42.920 18.470 42.995 18.615 ;
        RECT 42.920 17.120 42.995 17.265 ;
        RECT 42.920 15.770 42.995 15.915 ;
        RECT 42.920 14.420 42.995 14.565 ;
        RECT 42.920 13.070 42.995 13.215 ;
        RECT 42.920 11.720 42.995 11.865 ;
        RECT 42.920 10.370 42.995 10.515 ;
        RECT 42.920 9.020 42.995 9.165 ;
        RECT 42.920 7.670 42.995 7.815 ;
        RECT 42.920 6.320 42.995 6.465 ;
        RECT 42.920 4.970 42.995 5.115 ;
        RECT 42.920 3.620 42.995 3.765 ;
        RECT 42.920 2.275 42.995 2.420 ;
        RECT 42.920 0.920 42.995 1.070 ;
    END
    PORT
      LAYER li1 ;
        RECT 89.320 42.770 89.395 42.915 ;
        RECT 89.320 41.420 89.395 41.565 ;
        RECT 89.320 40.070 89.395 40.215 ;
        RECT 89.320 38.720 89.395 38.865 ;
        RECT 89.320 37.370 89.395 37.515 ;
        RECT 89.320 36.020 89.395 36.165 ;
        RECT 89.320 34.670 89.395 34.815 ;
        RECT 89.320 33.320 89.395 33.465 ;
        RECT 89.320 31.970 89.395 32.115 ;
        RECT 89.320 30.620 89.395 30.765 ;
        RECT 89.320 29.270 89.395 29.415 ;
        RECT 89.320 27.920 89.395 28.065 ;
        RECT 89.320 26.570 89.395 26.715 ;
        RECT 89.320 25.220 89.395 25.365 ;
        RECT 89.320 23.870 89.395 24.015 ;
        RECT 89.320 22.520 89.395 22.665 ;
        RECT 89.320 21.170 89.395 21.315 ;
        RECT 89.320 19.820 89.395 19.965 ;
        RECT 89.320 18.470 89.395 18.615 ;
        RECT 89.320 17.120 89.395 17.265 ;
        RECT 89.320 15.770 89.395 15.915 ;
        RECT 89.320 14.420 89.395 14.565 ;
        RECT 89.320 13.070 89.395 13.215 ;
        RECT 89.320 11.720 89.395 11.865 ;
        RECT 89.320 10.370 89.395 10.515 ;
        RECT 89.320 9.020 89.395 9.165 ;
        RECT 89.320 7.670 89.395 7.815 ;
        RECT 89.320 6.320 89.395 6.465 ;
        RECT 89.320 4.970 89.395 5.115 ;
        RECT 89.320 3.620 89.395 3.765 ;
        RECT 89.320 2.275 89.395 2.420 ;
        RECT 89.320 0.925 89.395 1.070 ;
    END
  END WBL_14
  PIN WBLb_14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.739575 ;
    PORT
      LAYER li1 ;
        RECT 40.970 42.770 41.045 42.910 ;
        RECT 40.970 41.420 41.045 41.560 ;
        RECT 40.970 40.070 41.045 40.210 ;
        RECT 40.970 38.720 41.045 38.860 ;
        RECT 40.970 37.370 41.045 37.510 ;
        RECT 40.970 36.020 41.045 36.160 ;
        RECT 40.970 34.670 41.045 34.810 ;
        RECT 40.970 33.320 41.045 33.460 ;
        RECT 40.970 31.970 41.045 32.110 ;
        RECT 40.970 30.620 41.045 30.760 ;
        RECT 40.970 29.270 41.045 29.410 ;
        RECT 40.970 27.920 41.045 28.060 ;
        RECT 40.970 26.570 41.045 26.710 ;
        RECT 40.970 25.220 41.045 25.360 ;
        RECT 40.970 23.870 41.045 24.010 ;
        RECT 40.970 22.520 41.045 22.660 ;
        RECT 40.970 21.170 41.045 21.310 ;
        RECT 40.970 19.820 41.045 19.960 ;
        RECT 40.970 18.470 41.045 18.610 ;
        RECT 40.970 17.120 41.045 17.260 ;
        RECT 40.970 15.770 41.045 15.910 ;
        RECT 40.970 14.420 41.045 14.560 ;
        RECT 40.970 13.070 41.045 13.210 ;
        RECT 40.970 11.720 41.045 11.860 ;
        RECT 40.970 10.370 41.045 10.510 ;
        RECT 40.970 9.020 41.045 9.160 ;
        RECT 40.970 7.670 41.045 7.810 ;
        RECT 40.970 6.320 41.045 6.460 ;
        RECT 40.970 4.970 41.045 5.110 ;
        RECT 40.970 3.620 41.045 3.760 ;
        RECT 40.970 2.275 41.045 2.415 ;
        RECT 40.970 0.920 41.045 1.065 ;
    END
    PORT
      LAYER li1 ;
        RECT 87.370 42.770 87.445 42.910 ;
        RECT 87.370 41.420 87.445 41.560 ;
        RECT 87.370 40.070 87.445 40.210 ;
        RECT 87.370 38.720 87.445 38.860 ;
        RECT 87.370 37.370 87.445 37.510 ;
        RECT 87.370 36.020 87.445 36.160 ;
        RECT 87.370 34.670 87.445 34.810 ;
        RECT 87.370 33.320 87.445 33.460 ;
        RECT 87.370 31.970 87.445 32.110 ;
        RECT 87.370 30.620 87.445 30.760 ;
        RECT 87.370 29.270 87.445 29.410 ;
        RECT 87.370 27.920 87.445 28.060 ;
        RECT 87.370 26.570 87.445 26.710 ;
        RECT 87.370 25.220 87.445 25.360 ;
        RECT 87.370 23.870 87.445 24.010 ;
        RECT 87.370 22.520 87.445 22.660 ;
        RECT 87.370 21.170 87.445 21.310 ;
        RECT 87.370 19.820 87.445 19.960 ;
        RECT 87.370 18.470 87.445 18.610 ;
        RECT 87.370 17.120 87.445 17.260 ;
        RECT 87.370 15.770 87.445 15.910 ;
        RECT 87.370 14.420 87.445 14.560 ;
        RECT 87.370 13.070 87.445 13.210 ;
        RECT 87.370 11.720 87.445 11.860 ;
        RECT 87.370 10.370 87.445 10.510 ;
        RECT 87.370 9.020 87.445 9.160 ;
        RECT 87.370 7.670 87.445 7.810 ;
        RECT 87.370 6.320 87.445 6.460 ;
        RECT 87.370 4.970 87.445 5.110 ;
        RECT 87.370 3.620 87.445 3.760 ;
        RECT 87.370 2.275 87.445 2.415 ;
        RECT 87.370 0.925 87.445 1.065 ;
    END
  END WBLb_14
  PIN WBL_15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.773975 ;
    PORT
      LAYER li1 ;
        RECT 45.820 42.770 45.895 42.915 ;
        RECT 45.820 41.420 45.895 41.565 ;
        RECT 45.820 40.070 45.895 40.215 ;
        RECT 45.820 38.720 45.895 38.865 ;
        RECT 45.820 37.370 45.895 37.515 ;
        RECT 45.820 36.020 45.895 36.165 ;
        RECT 45.820 34.670 45.895 34.815 ;
        RECT 45.820 33.320 45.895 33.465 ;
        RECT 45.820 31.970 45.895 32.115 ;
        RECT 45.820 30.620 45.895 30.765 ;
        RECT 45.820 29.270 45.895 29.415 ;
        RECT 45.820 27.920 45.895 28.065 ;
        RECT 45.820 26.570 45.895 26.715 ;
        RECT 45.820 25.220 45.895 25.365 ;
        RECT 45.820 23.870 45.895 24.015 ;
        RECT 45.820 22.520 45.895 22.665 ;
        RECT 45.820 21.170 45.895 21.315 ;
        RECT 45.820 19.820 45.895 19.965 ;
        RECT 45.820 18.470 45.895 18.615 ;
        RECT 45.820 17.120 45.895 17.265 ;
        RECT 45.820 15.770 45.895 15.915 ;
        RECT 45.820 14.420 45.895 14.565 ;
        RECT 45.820 13.070 45.895 13.215 ;
        RECT 45.820 11.720 45.895 11.865 ;
        RECT 45.820 10.370 45.895 10.515 ;
        RECT 45.820 9.020 45.895 9.165 ;
        RECT 45.820 7.670 45.895 7.815 ;
        RECT 45.820 6.320 45.895 6.465 ;
        RECT 45.820 4.970 45.895 5.115 ;
        RECT 45.820 3.620 45.895 3.765 ;
        RECT 45.820 2.275 45.895 2.420 ;
        RECT 45.820 0.920 45.895 1.070 ;
    END
    PORT
      LAYER li1 ;
        RECT 92.220 42.770 92.295 42.915 ;
        RECT 92.220 41.420 92.295 41.565 ;
        RECT 92.220 40.070 92.295 40.215 ;
        RECT 92.220 38.720 92.295 38.865 ;
        RECT 92.220 37.370 92.295 37.515 ;
        RECT 92.220 36.020 92.295 36.165 ;
        RECT 92.220 34.670 92.295 34.815 ;
        RECT 92.220 33.320 92.295 33.465 ;
        RECT 92.220 31.970 92.295 32.115 ;
        RECT 92.220 30.620 92.295 30.765 ;
        RECT 92.220 29.270 92.295 29.415 ;
        RECT 92.220 27.920 92.295 28.065 ;
        RECT 92.220 26.570 92.295 26.715 ;
        RECT 92.220 25.220 92.295 25.365 ;
        RECT 92.220 23.870 92.295 24.015 ;
        RECT 92.220 22.520 92.295 22.665 ;
        RECT 92.220 21.170 92.295 21.315 ;
        RECT 92.220 19.820 92.295 19.965 ;
        RECT 92.220 18.470 92.295 18.615 ;
        RECT 92.220 17.120 92.295 17.265 ;
        RECT 92.220 15.770 92.295 15.915 ;
        RECT 92.220 14.420 92.295 14.565 ;
        RECT 92.220 13.070 92.295 13.215 ;
        RECT 92.220 11.720 92.295 11.865 ;
        RECT 92.220 10.370 92.295 10.515 ;
        RECT 92.220 9.020 92.295 9.165 ;
        RECT 92.220 7.670 92.295 7.815 ;
        RECT 92.220 6.320 92.295 6.465 ;
        RECT 92.220 4.970 92.295 5.115 ;
        RECT 92.220 3.620 92.295 3.765 ;
        RECT 92.220 2.275 92.295 2.420 ;
        RECT 92.220 0.925 92.295 1.070 ;
    END
  END WBL_15
  PIN WBLb_15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.739575 ;
    PORT
      LAYER li1 ;
        RECT 43.870 42.770 43.945 42.910 ;
        RECT 43.870 41.420 43.945 41.560 ;
        RECT 43.870 40.070 43.945 40.210 ;
        RECT 43.870 38.720 43.945 38.860 ;
        RECT 43.870 37.370 43.945 37.510 ;
        RECT 43.870 36.020 43.945 36.160 ;
        RECT 43.870 34.670 43.945 34.810 ;
        RECT 43.870 33.320 43.945 33.460 ;
        RECT 43.870 31.970 43.945 32.110 ;
        RECT 43.870 30.620 43.945 30.760 ;
        RECT 43.870 29.270 43.945 29.410 ;
        RECT 43.870 27.920 43.945 28.060 ;
        RECT 43.870 26.570 43.945 26.710 ;
        RECT 43.870 25.220 43.945 25.360 ;
        RECT 43.870 23.870 43.945 24.010 ;
        RECT 43.870 22.520 43.945 22.660 ;
        RECT 43.870 21.170 43.945 21.310 ;
        RECT 43.870 19.820 43.945 19.960 ;
        RECT 43.870 18.470 43.945 18.610 ;
        RECT 43.870 17.120 43.945 17.260 ;
        RECT 43.870 15.770 43.945 15.910 ;
        RECT 43.870 14.420 43.945 14.560 ;
        RECT 43.870 13.070 43.945 13.210 ;
        RECT 43.870 11.720 43.945 11.860 ;
        RECT 43.870 10.370 43.945 10.510 ;
        RECT 43.870 9.020 43.945 9.160 ;
        RECT 43.870 7.670 43.945 7.810 ;
        RECT 43.870 6.320 43.945 6.460 ;
        RECT 43.870 4.970 43.945 5.110 ;
        RECT 43.870 3.620 43.945 3.760 ;
        RECT 43.870 2.275 43.945 2.415 ;
        RECT 43.870 0.920 43.945 1.065 ;
    END
    PORT
      LAYER li1 ;
        RECT 90.270 42.770 90.345 42.910 ;
        RECT 90.270 41.420 90.345 41.560 ;
        RECT 90.270 40.070 90.345 40.210 ;
        RECT 90.270 38.720 90.345 38.860 ;
        RECT 90.270 37.370 90.345 37.510 ;
        RECT 90.270 36.020 90.345 36.160 ;
        RECT 90.270 34.670 90.345 34.810 ;
        RECT 90.270 33.320 90.345 33.460 ;
        RECT 90.270 31.970 90.345 32.110 ;
        RECT 90.270 30.620 90.345 30.760 ;
        RECT 90.270 29.270 90.345 29.410 ;
        RECT 90.270 27.920 90.345 28.060 ;
        RECT 90.270 26.570 90.345 26.710 ;
        RECT 90.270 25.220 90.345 25.360 ;
        RECT 90.270 23.870 90.345 24.010 ;
        RECT 90.270 22.520 90.345 22.660 ;
        RECT 90.270 21.170 90.345 21.310 ;
        RECT 90.270 19.820 90.345 19.960 ;
        RECT 90.270 18.470 90.345 18.610 ;
        RECT 90.270 17.120 90.345 17.260 ;
        RECT 90.270 15.770 90.345 15.910 ;
        RECT 90.270 14.420 90.345 14.560 ;
        RECT 90.270 13.070 90.345 13.210 ;
        RECT 90.270 11.720 90.345 11.860 ;
        RECT 90.270 10.370 90.345 10.510 ;
        RECT 90.270 9.020 90.345 9.160 ;
        RECT 90.270 7.670 90.345 7.810 ;
        RECT 90.270 6.320 90.345 6.460 ;
        RECT 90.270 4.970 90.345 5.110 ;
        RECT 90.270 3.620 90.345 3.760 ;
        RECT 90.270 2.275 90.345 2.415 ;
        RECT 90.270 0.925 90.345 1.065 ;
    END
  END WBLb_15
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER nwell ;
        RECT 0.990 42.570 1.755 43.050 ;
        RECT 3.890 42.570 4.655 43.050 ;
        RECT 6.790 42.570 7.555 43.050 ;
        RECT 9.690 42.570 10.455 43.050 ;
        RECT 12.590 42.570 13.355 43.050 ;
        RECT 15.490 42.570 16.255 43.050 ;
        RECT 18.390 42.570 19.155 43.050 ;
        RECT 21.290 42.570 22.055 43.050 ;
        RECT 24.190 42.570 24.955 43.050 ;
        RECT 27.090 42.570 27.855 43.050 ;
        RECT 29.990 42.570 30.755 43.050 ;
        RECT 32.890 42.570 33.655 43.050 ;
        RECT 35.790 42.570 36.555 43.050 ;
        RECT 38.690 42.570 39.455 43.050 ;
        RECT 41.590 42.570 42.355 43.050 ;
        RECT 44.490 42.570 45.255 43.050 ;
        RECT 47.390 42.570 48.155 43.050 ;
        RECT 50.290 42.570 51.055 43.050 ;
        RECT 53.190 42.570 53.955 43.050 ;
        RECT 56.090 42.570 56.855 43.050 ;
        RECT 58.990 42.570 59.755 43.050 ;
        RECT 61.890 42.570 62.655 43.050 ;
        RECT 64.790 42.570 65.555 43.050 ;
        RECT 67.690 42.570 68.455 43.050 ;
        RECT 70.590 42.570 71.355 43.050 ;
        RECT 73.490 42.570 74.255 43.050 ;
        RECT 76.390 42.570 77.155 43.050 ;
        RECT 79.290 42.570 80.055 43.050 ;
        RECT 82.190 42.570 82.955 43.050 ;
        RECT 85.090 42.570 85.855 43.050 ;
        RECT 87.990 42.570 88.755 43.050 ;
        RECT 90.890 42.570 91.655 43.050 ;
      LAYER li1 ;
        RECT 1.300 42.980 1.460 43.050 ;
        RECT 4.200 42.980 4.360 43.050 ;
        RECT 7.100 42.980 7.260 43.050 ;
        RECT 10.000 42.980 10.160 43.050 ;
        RECT 12.900 42.980 13.060 43.050 ;
        RECT 15.800 42.980 15.960 43.050 ;
        RECT 18.700 42.980 18.860 43.050 ;
        RECT 21.600 42.980 21.760 43.050 ;
        RECT 24.500 42.980 24.660 43.050 ;
        RECT 27.400 42.980 27.560 43.050 ;
        RECT 30.300 42.980 30.460 43.050 ;
        RECT 33.200 42.980 33.360 43.050 ;
        RECT 36.100 42.980 36.260 43.050 ;
        RECT 39.000 42.980 39.160 43.050 ;
        RECT 41.900 42.980 42.060 43.050 ;
        RECT 44.800 42.980 44.960 43.050 ;
        RECT 47.700 42.980 47.860 43.050 ;
        RECT 50.600 42.980 50.760 43.050 ;
        RECT 53.500 42.980 53.660 43.050 ;
        RECT 56.400 42.980 56.560 43.050 ;
        RECT 59.300 42.980 59.460 43.050 ;
        RECT 62.200 42.980 62.360 43.050 ;
        RECT 65.100 42.980 65.260 43.050 ;
        RECT 68.000 42.980 68.160 43.050 ;
        RECT 70.900 42.980 71.060 43.050 ;
        RECT 73.800 42.980 73.960 43.050 ;
        RECT 76.700 42.980 76.860 43.050 ;
        RECT 79.600 42.980 79.760 43.050 ;
        RECT 82.500 42.980 82.660 43.050 ;
        RECT 85.400 42.980 85.560 43.050 ;
        RECT 88.300 42.980 88.460 43.050 ;
        RECT 91.200 42.980 91.360 43.050 ;
        RECT 1.310 42.970 1.450 42.980 ;
        RECT 4.210 42.970 4.350 42.980 ;
        RECT 7.110 42.970 7.250 42.980 ;
        RECT 10.010 42.970 10.150 42.980 ;
        RECT 12.910 42.970 13.050 42.980 ;
        RECT 15.810 42.970 15.950 42.980 ;
        RECT 18.710 42.970 18.850 42.980 ;
        RECT 21.610 42.970 21.750 42.980 ;
        RECT 24.510 42.970 24.650 42.980 ;
        RECT 27.410 42.970 27.550 42.980 ;
        RECT 30.310 42.970 30.450 42.980 ;
        RECT 33.210 42.970 33.350 42.980 ;
        RECT 36.110 42.970 36.250 42.980 ;
        RECT 39.010 42.970 39.150 42.980 ;
        RECT 41.910 42.970 42.050 42.980 ;
        RECT 44.810 42.970 44.950 42.980 ;
        RECT 47.710 42.970 47.850 42.980 ;
        RECT 50.610 42.970 50.750 42.980 ;
        RECT 53.510 42.970 53.650 42.980 ;
        RECT 56.410 42.970 56.550 42.980 ;
        RECT 59.310 42.970 59.450 42.980 ;
        RECT 62.210 42.970 62.350 42.980 ;
        RECT 65.110 42.970 65.250 42.980 ;
        RECT 68.010 42.970 68.150 42.980 ;
        RECT 70.910 42.970 71.050 42.980 ;
        RECT 73.810 42.970 73.950 42.980 ;
        RECT 76.710 42.970 76.850 42.980 ;
        RECT 79.610 42.970 79.750 42.980 ;
        RECT 82.510 42.970 82.650 42.980 ;
        RECT 85.410 42.970 85.550 42.980 ;
        RECT 88.310 42.970 88.450 42.980 ;
        RECT 91.210 42.970 91.350 42.980 ;
      LAYER met1 ;
        RECT 0.000 42.980 92.660 43.050 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.990 41.220 1.755 41.700 ;
        RECT 3.890 41.220 4.655 41.700 ;
        RECT 6.790 41.220 7.555 41.700 ;
        RECT 9.690 41.220 10.455 41.700 ;
        RECT 12.590 41.220 13.355 41.700 ;
        RECT 15.490 41.220 16.255 41.700 ;
        RECT 18.390 41.220 19.155 41.700 ;
        RECT 21.290 41.220 22.055 41.700 ;
        RECT 24.190 41.220 24.955 41.700 ;
        RECT 27.090 41.220 27.855 41.700 ;
        RECT 29.990 41.220 30.755 41.700 ;
        RECT 32.890 41.220 33.655 41.700 ;
        RECT 35.790 41.220 36.555 41.700 ;
        RECT 38.690 41.220 39.455 41.700 ;
        RECT 41.590 41.220 42.355 41.700 ;
        RECT 44.490 41.220 45.255 41.700 ;
        RECT 47.390 41.220 48.155 41.700 ;
        RECT 50.290 41.220 51.055 41.700 ;
        RECT 53.190 41.220 53.955 41.700 ;
        RECT 56.090 41.220 56.855 41.700 ;
        RECT 58.990 41.220 59.755 41.700 ;
        RECT 61.890 41.220 62.655 41.700 ;
        RECT 64.790 41.220 65.555 41.700 ;
        RECT 67.690 41.220 68.455 41.700 ;
        RECT 70.590 41.220 71.355 41.700 ;
        RECT 73.490 41.220 74.255 41.700 ;
        RECT 76.390 41.220 77.155 41.700 ;
        RECT 79.290 41.220 80.055 41.700 ;
        RECT 82.190 41.220 82.955 41.700 ;
        RECT 85.090 41.220 85.855 41.700 ;
        RECT 87.990 41.220 88.755 41.700 ;
        RECT 90.890 41.220 91.655 41.700 ;
      LAYER li1 ;
        RECT 1.300 41.630 1.460 41.700 ;
        RECT 4.200 41.630 4.360 41.700 ;
        RECT 7.100 41.630 7.260 41.700 ;
        RECT 10.000 41.630 10.160 41.700 ;
        RECT 12.900 41.630 13.060 41.700 ;
        RECT 15.800 41.630 15.960 41.700 ;
        RECT 18.700 41.630 18.860 41.700 ;
        RECT 21.600 41.630 21.760 41.700 ;
        RECT 24.500 41.630 24.660 41.700 ;
        RECT 27.400 41.630 27.560 41.700 ;
        RECT 30.300 41.630 30.460 41.700 ;
        RECT 33.200 41.630 33.360 41.700 ;
        RECT 36.100 41.630 36.260 41.700 ;
        RECT 39.000 41.630 39.160 41.700 ;
        RECT 41.900 41.630 42.060 41.700 ;
        RECT 44.800 41.630 44.960 41.700 ;
        RECT 47.700 41.630 47.860 41.700 ;
        RECT 50.600 41.630 50.760 41.700 ;
        RECT 53.500 41.630 53.660 41.700 ;
        RECT 56.400 41.630 56.560 41.700 ;
        RECT 59.300 41.630 59.460 41.700 ;
        RECT 62.200 41.630 62.360 41.700 ;
        RECT 65.100 41.630 65.260 41.700 ;
        RECT 68.000 41.630 68.160 41.700 ;
        RECT 70.900 41.630 71.060 41.700 ;
        RECT 73.800 41.630 73.960 41.700 ;
        RECT 76.700 41.630 76.860 41.700 ;
        RECT 79.600 41.630 79.760 41.700 ;
        RECT 82.500 41.630 82.660 41.700 ;
        RECT 85.400 41.630 85.560 41.700 ;
        RECT 88.300 41.630 88.460 41.700 ;
        RECT 91.200 41.630 91.360 41.700 ;
        RECT 1.310 41.620 1.450 41.630 ;
        RECT 4.210 41.620 4.350 41.630 ;
        RECT 7.110 41.620 7.250 41.630 ;
        RECT 10.010 41.620 10.150 41.630 ;
        RECT 12.910 41.620 13.050 41.630 ;
        RECT 15.810 41.620 15.950 41.630 ;
        RECT 18.710 41.620 18.850 41.630 ;
        RECT 21.610 41.620 21.750 41.630 ;
        RECT 24.510 41.620 24.650 41.630 ;
        RECT 27.410 41.620 27.550 41.630 ;
        RECT 30.310 41.620 30.450 41.630 ;
        RECT 33.210 41.620 33.350 41.630 ;
        RECT 36.110 41.620 36.250 41.630 ;
        RECT 39.010 41.620 39.150 41.630 ;
        RECT 41.910 41.620 42.050 41.630 ;
        RECT 44.810 41.620 44.950 41.630 ;
        RECT 47.710 41.620 47.850 41.630 ;
        RECT 50.610 41.620 50.750 41.630 ;
        RECT 53.510 41.620 53.650 41.630 ;
        RECT 56.410 41.620 56.550 41.630 ;
        RECT 59.310 41.620 59.450 41.630 ;
        RECT 62.210 41.620 62.350 41.630 ;
        RECT 65.110 41.620 65.250 41.630 ;
        RECT 68.010 41.620 68.150 41.630 ;
        RECT 70.910 41.620 71.050 41.630 ;
        RECT 73.810 41.620 73.950 41.630 ;
        RECT 76.710 41.620 76.850 41.630 ;
        RECT 79.610 41.620 79.750 41.630 ;
        RECT 82.510 41.620 82.650 41.630 ;
        RECT 85.410 41.620 85.550 41.630 ;
        RECT 88.310 41.620 88.450 41.630 ;
        RECT 91.210 41.620 91.350 41.630 ;
      LAYER met1 ;
        RECT 0.000 41.630 92.660 41.700 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.990 39.870 1.755 40.350 ;
        RECT 3.890 39.870 4.655 40.350 ;
        RECT 6.790 39.870 7.555 40.350 ;
        RECT 9.690 39.870 10.455 40.350 ;
        RECT 12.590 39.870 13.355 40.350 ;
        RECT 15.490 39.870 16.255 40.350 ;
        RECT 18.390 39.870 19.155 40.350 ;
        RECT 21.290 39.870 22.055 40.350 ;
        RECT 24.190 39.870 24.955 40.350 ;
        RECT 27.090 39.870 27.855 40.350 ;
        RECT 29.990 39.870 30.755 40.350 ;
        RECT 32.890 39.870 33.655 40.350 ;
        RECT 35.790 39.870 36.555 40.350 ;
        RECT 38.690 39.870 39.455 40.350 ;
        RECT 41.590 39.870 42.355 40.350 ;
        RECT 44.490 39.870 45.255 40.350 ;
        RECT 47.390 39.870 48.155 40.350 ;
        RECT 50.290 39.870 51.055 40.350 ;
        RECT 53.190 39.870 53.955 40.350 ;
        RECT 56.090 39.870 56.855 40.350 ;
        RECT 58.990 39.870 59.755 40.350 ;
        RECT 61.890 39.870 62.655 40.350 ;
        RECT 64.790 39.870 65.555 40.350 ;
        RECT 67.690 39.870 68.455 40.350 ;
        RECT 70.590 39.870 71.355 40.350 ;
        RECT 73.490 39.870 74.255 40.350 ;
        RECT 76.390 39.870 77.155 40.350 ;
        RECT 79.290 39.870 80.055 40.350 ;
        RECT 82.190 39.870 82.955 40.350 ;
        RECT 85.090 39.870 85.855 40.350 ;
        RECT 87.990 39.870 88.755 40.350 ;
        RECT 90.890 39.870 91.655 40.350 ;
      LAYER li1 ;
        RECT 1.300 40.280 1.460 40.350 ;
        RECT 4.200 40.280 4.360 40.350 ;
        RECT 7.100 40.280 7.260 40.350 ;
        RECT 10.000 40.280 10.160 40.350 ;
        RECT 12.900 40.280 13.060 40.350 ;
        RECT 15.800 40.280 15.960 40.350 ;
        RECT 18.700 40.280 18.860 40.350 ;
        RECT 21.600 40.280 21.760 40.350 ;
        RECT 24.500 40.280 24.660 40.350 ;
        RECT 27.400 40.280 27.560 40.350 ;
        RECT 30.300 40.280 30.460 40.350 ;
        RECT 33.200 40.280 33.360 40.350 ;
        RECT 36.100 40.280 36.260 40.350 ;
        RECT 39.000 40.280 39.160 40.350 ;
        RECT 41.900 40.280 42.060 40.350 ;
        RECT 44.800 40.280 44.960 40.350 ;
        RECT 47.700 40.280 47.860 40.350 ;
        RECT 50.600 40.280 50.760 40.350 ;
        RECT 53.500 40.280 53.660 40.350 ;
        RECT 56.400 40.280 56.560 40.350 ;
        RECT 59.300 40.280 59.460 40.350 ;
        RECT 62.200 40.280 62.360 40.350 ;
        RECT 65.100 40.280 65.260 40.350 ;
        RECT 68.000 40.280 68.160 40.350 ;
        RECT 70.900 40.280 71.060 40.350 ;
        RECT 73.800 40.280 73.960 40.350 ;
        RECT 76.700 40.280 76.860 40.350 ;
        RECT 79.600 40.280 79.760 40.350 ;
        RECT 82.500 40.280 82.660 40.350 ;
        RECT 85.400 40.280 85.560 40.350 ;
        RECT 88.300 40.280 88.460 40.350 ;
        RECT 91.200 40.280 91.360 40.350 ;
        RECT 1.310 40.270 1.450 40.280 ;
        RECT 4.210 40.270 4.350 40.280 ;
        RECT 7.110 40.270 7.250 40.280 ;
        RECT 10.010 40.270 10.150 40.280 ;
        RECT 12.910 40.270 13.050 40.280 ;
        RECT 15.810 40.270 15.950 40.280 ;
        RECT 18.710 40.270 18.850 40.280 ;
        RECT 21.610 40.270 21.750 40.280 ;
        RECT 24.510 40.270 24.650 40.280 ;
        RECT 27.410 40.270 27.550 40.280 ;
        RECT 30.310 40.270 30.450 40.280 ;
        RECT 33.210 40.270 33.350 40.280 ;
        RECT 36.110 40.270 36.250 40.280 ;
        RECT 39.010 40.270 39.150 40.280 ;
        RECT 41.910 40.270 42.050 40.280 ;
        RECT 44.810 40.270 44.950 40.280 ;
        RECT 47.710 40.270 47.850 40.280 ;
        RECT 50.610 40.270 50.750 40.280 ;
        RECT 53.510 40.270 53.650 40.280 ;
        RECT 56.410 40.270 56.550 40.280 ;
        RECT 59.310 40.270 59.450 40.280 ;
        RECT 62.210 40.270 62.350 40.280 ;
        RECT 65.110 40.270 65.250 40.280 ;
        RECT 68.010 40.270 68.150 40.280 ;
        RECT 70.910 40.270 71.050 40.280 ;
        RECT 73.810 40.270 73.950 40.280 ;
        RECT 76.710 40.270 76.850 40.280 ;
        RECT 79.610 40.270 79.750 40.280 ;
        RECT 82.510 40.270 82.650 40.280 ;
        RECT 85.410 40.270 85.550 40.280 ;
        RECT 88.310 40.270 88.450 40.280 ;
        RECT 91.210 40.270 91.350 40.280 ;
      LAYER met1 ;
        RECT 0.000 40.280 92.660 40.350 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.990 38.520 1.755 39.000 ;
        RECT 3.890 38.520 4.655 39.000 ;
        RECT 6.790 38.520 7.555 39.000 ;
        RECT 9.690 38.520 10.455 39.000 ;
        RECT 12.590 38.520 13.355 39.000 ;
        RECT 15.490 38.520 16.255 39.000 ;
        RECT 18.390 38.520 19.155 39.000 ;
        RECT 21.290 38.520 22.055 39.000 ;
        RECT 24.190 38.520 24.955 39.000 ;
        RECT 27.090 38.520 27.855 39.000 ;
        RECT 29.990 38.520 30.755 39.000 ;
        RECT 32.890 38.520 33.655 39.000 ;
        RECT 35.790 38.520 36.555 39.000 ;
        RECT 38.690 38.520 39.455 39.000 ;
        RECT 41.590 38.520 42.355 39.000 ;
        RECT 44.490 38.520 45.255 39.000 ;
        RECT 47.390 38.520 48.155 39.000 ;
        RECT 50.290 38.520 51.055 39.000 ;
        RECT 53.190 38.520 53.955 39.000 ;
        RECT 56.090 38.520 56.855 39.000 ;
        RECT 58.990 38.520 59.755 39.000 ;
        RECT 61.890 38.520 62.655 39.000 ;
        RECT 64.790 38.520 65.555 39.000 ;
        RECT 67.690 38.520 68.455 39.000 ;
        RECT 70.590 38.520 71.355 39.000 ;
        RECT 73.490 38.520 74.255 39.000 ;
        RECT 76.390 38.520 77.155 39.000 ;
        RECT 79.290 38.520 80.055 39.000 ;
        RECT 82.190 38.520 82.955 39.000 ;
        RECT 85.090 38.520 85.855 39.000 ;
        RECT 87.990 38.520 88.755 39.000 ;
        RECT 90.890 38.520 91.655 39.000 ;
      LAYER li1 ;
        RECT 1.300 38.930 1.460 39.000 ;
        RECT 4.200 38.930 4.360 39.000 ;
        RECT 7.100 38.930 7.260 39.000 ;
        RECT 10.000 38.930 10.160 39.000 ;
        RECT 12.900 38.930 13.060 39.000 ;
        RECT 15.800 38.930 15.960 39.000 ;
        RECT 18.700 38.930 18.860 39.000 ;
        RECT 21.600 38.930 21.760 39.000 ;
        RECT 24.500 38.930 24.660 39.000 ;
        RECT 27.400 38.930 27.560 39.000 ;
        RECT 30.300 38.930 30.460 39.000 ;
        RECT 33.200 38.930 33.360 39.000 ;
        RECT 36.100 38.930 36.260 39.000 ;
        RECT 39.000 38.930 39.160 39.000 ;
        RECT 41.900 38.930 42.060 39.000 ;
        RECT 44.800 38.930 44.960 39.000 ;
        RECT 47.700 38.930 47.860 39.000 ;
        RECT 50.600 38.930 50.760 39.000 ;
        RECT 53.500 38.930 53.660 39.000 ;
        RECT 56.400 38.930 56.560 39.000 ;
        RECT 59.300 38.930 59.460 39.000 ;
        RECT 62.200 38.930 62.360 39.000 ;
        RECT 65.100 38.930 65.260 39.000 ;
        RECT 68.000 38.930 68.160 39.000 ;
        RECT 70.900 38.930 71.060 39.000 ;
        RECT 73.800 38.930 73.960 39.000 ;
        RECT 76.700 38.930 76.860 39.000 ;
        RECT 79.600 38.930 79.760 39.000 ;
        RECT 82.500 38.930 82.660 39.000 ;
        RECT 85.400 38.930 85.560 39.000 ;
        RECT 88.300 38.930 88.460 39.000 ;
        RECT 91.200 38.930 91.360 39.000 ;
        RECT 1.310 38.920 1.450 38.930 ;
        RECT 4.210 38.920 4.350 38.930 ;
        RECT 7.110 38.920 7.250 38.930 ;
        RECT 10.010 38.920 10.150 38.930 ;
        RECT 12.910 38.920 13.050 38.930 ;
        RECT 15.810 38.920 15.950 38.930 ;
        RECT 18.710 38.920 18.850 38.930 ;
        RECT 21.610 38.920 21.750 38.930 ;
        RECT 24.510 38.920 24.650 38.930 ;
        RECT 27.410 38.920 27.550 38.930 ;
        RECT 30.310 38.920 30.450 38.930 ;
        RECT 33.210 38.920 33.350 38.930 ;
        RECT 36.110 38.920 36.250 38.930 ;
        RECT 39.010 38.920 39.150 38.930 ;
        RECT 41.910 38.920 42.050 38.930 ;
        RECT 44.810 38.920 44.950 38.930 ;
        RECT 47.710 38.920 47.850 38.930 ;
        RECT 50.610 38.920 50.750 38.930 ;
        RECT 53.510 38.920 53.650 38.930 ;
        RECT 56.410 38.920 56.550 38.930 ;
        RECT 59.310 38.920 59.450 38.930 ;
        RECT 62.210 38.920 62.350 38.930 ;
        RECT 65.110 38.920 65.250 38.930 ;
        RECT 68.010 38.920 68.150 38.930 ;
        RECT 70.910 38.920 71.050 38.930 ;
        RECT 73.810 38.920 73.950 38.930 ;
        RECT 76.710 38.920 76.850 38.930 ;
        RECT 79.610 38.920 79.750 38.930 ;
        RECT 82.510 38.920 82.650 38.930 ;
        RECT 85.410 38.920 85.550 38.930 ;
        RECT 88.310 38.920 88.450 38.930 ;
        RECT 91.210 38.920 91.350 38.930 ;
      LAYER met1 ;
        RECT 0.000 38.930 92.660 39.000 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.990 37.170 1.755 37.650 ;
        RECT 3.890 37.170 4.655 37.650 ;
        RECT 6.790 37.170 7.555 37.650 ;
        RECT 9.690 37.170 10.455 37.650 ;
        RECT 12.590 37.170 13.355 37.650 ;
        RECT 15.490 37.170 16.255 37.650 ;
        RECT 18.390 37.170 19.155 37.650 ;
        RECT 21.290 37.170 22.055 37.650 ;
        RECT 24.190 37.170 24.955 37.650 ;
        RECT 27.090 37.170 27.855 37.650 ;
        RECT 29.990 37.170 30.755 37.650 ;
        RECT 32.890 37.170 33.655 37.650 ;
        RECT 35.790 37.170 36.555 37.650 ;
        RECT 38.690 37.170 39.455 37.650 ;
        RECT 41.590 37.170 42.355 37.650 ;
        RECT 44.490 37.170 45.255 37.650 ;
        RECT 47.390 37.170 48.155 37.650 ;
        RECT 50.290 37.170 51.055 37.650 ;
        RECT 53.190 37.170 53.955 37.650 ;
        RECT 56.090 37.170 56.855 37.650 ;
        RECT 58.990 37.170 59.755 37.650 ;
        RECT 61.890 37.170 62.655 37.650 ;
        RECT 64.790 37.170 65.555 37.650 ;
        RECT 67.690 37.170 68.455 37.650 ;
        RECT 70.590 37.170 71.355 37.650 ;
        RECT 73.490 37.170 74.255 37.650 ;
        RECT 76.390 37.170 77.155 37.650 ;
        RECT 79.290 37.170 80.055 37.650 ;
        RECT 82.190 37.170 82.955 37.650 ;
        RECT 85.090 37.170 85.855 37.650 ;
        RECT 87.990 37.170 88.755 37.650 ;
        RECT 90.890 37.170 91.655 37.650 ;
      LAYER li1 ;
        RECT 1.300 37.580 1.460 37.650 ;
        RECT 4.200 37.580 4.360 37.650 ;
        RECT 7.100 37.580 7.260 37.650 ;
        RECT 10.000 37.580 10.160 37.650 ;
        RECT 12.900 37.580 13.060 37.650 ;
        RECT 15.800 37.580 15.960 37.650 ;
        RECT 18.700 37.580 18.860 37.650 ;
        RECT 21.600 37.580 21.760 37.650 ;
        RECT 24.500 37.580 24.660 37.650 ;
        RECT 27.400 37.580 27.560 37.650 ;
        RECT 30.300 37.580 30.460 37.650 ;
        RECT 33.200 37.580 33.360 37.650 ;
        RECT 36.100 37.580 36.260 37.650 ;
        RECT 39.000 37.580 39.160 37.650 ;
        RECT 41.900 37.580 42.060 37.650 ;
        RECT 44.800 37.580 44.960 37.650 ;
        RECT 47.700 37.580 47.860 37.650 ;
        RECT 50.600 37.580 50.760 37.650 ;
        RECT 53.500 37.580 53.660 37.650 ;
        RECT 56.400 37.580 56.560 37.650 ;
        RECT 59.300 37.580 59.460 37.650 ;
        RECT 62.200 37.580 62.360 37.650 ;
        RECT 65.100 37.580 65.260 37.650 ;
        RECT 68.000 37.580 68.160 37.650 ;
        RECT 70.900 37.580 71.060 37.650 ;
        RECT 73.800 37.580 73.960 37.650 ;
        RECT 76.700 37.580 76.860 37.650 ;
        RECT 79.600 37.580 79.760 37.650 ;
        RECT 82.500 37.580 82.660 37.650 ;
        RECT 85.400 37.580 85.560 37.650 ;
        RECT 88.300 37.580 88.460 37.650 ;
        RECT 91.200 37.580 91.360 37.650 ;
        RECT 1.310 37.570 1.450 37.580 ;
        RECT 4.210 37.570 4.350 37.580 ;
        RECT 7.110 37.570 7.250 37.580 ;
        RECT 10.010 37.570 10.150 37.580 ;
        RECT 12.910 37.570 13.050 37.580 ;
        RECT 15.810 37.570 15.950 37.580 ;
        RECT 18.710 37.570 18.850 37.580 ;
        RECT 21.610 37.570 21.750 37.580 ;
        RECT 24.510 37.570 24.650 37.580 ;
        RECT 27.410 37.570 27.550 37.580 ;
        RECT 30.310 37.570 30.450 37.580 ;
        RECT 33.210 37.570 33.350 37.580 ;
        RECT 36.110 37.570 36.250 37.580 ;
        RECT 39.010 37.570 39.150 37.580 ;
        RECT 41.910 37.570 42.050 37.580 ;
        RECT 44.810 37.570 44.950 37.580 ;
        RECT 47.710 37.570 47.850 37.580 ;
        RECT 50.610 37.570 50.750 37.580 ;
        RECT 53.510 37.570 53.650 37.580 ;
        RECT 56.410 37.570 56.550 37.580 ;
        RECT 59.310 37.570 59.450 37.580 ;
        RECT 62.210 37.570 62.350 37.580 ;
        RECT 65.110 37.570 65.250 37.580 ;
        RECT 68.010 37.570 68.150 37.580 ;
        RECT 70.910 37.570 71.050 37.580 ;
        RECT 73.810 37.570 73.950 37.580 ;
        RECT 76.710 37.570 76.850 37.580 ;
        RECT 79.610 37.570 79.750 37.580 ;
        RECT 82.510 37.570 82.650 37.580 ;
        RECT 85.410 37.570 85.550 37.580 ;
        RECT 88.310 37.570 88.450 37.580 ;
        RECT 91.210 37.570 91.350 37.580 ;
      LAYER met1 ;
        RECT 0.000 37.580 92.660 37.650 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.990 35.820 1.755 36.300 ;
        RECT 3.890 35.820 4.655 36.300 ;
        RECT 6.790 35.820 7.555 36.300 ;
        RECT 9.690 35.820 10.455 36.300 ;
        RECT 12.590 35.820 13.355 36.300 ;
        RECT 15.490 35.820 16.255 36.300 ;
        RECT 18.390 35.820 19.155 36.300 ;
        RECT 21.290 35.820 22.055 36.300 ;
        RECT 24.190 35.820 24.955 36.300 ;
        RECT 27.090 35.820 27.855 36.300 ;
        RECT 29.990 35.820 30.755 36.300 ;
        RECT 32.890 35.820 33.655 36.300 ;
        RECT 35.790 35.820 36.555 36.300 ;
        RECT 38.690 35.820 39.455 36.300 ;
        RECT 41.590 35.820 42.355 36.300 ;
        RECT 44.490 35.820 45.255 36.300 ;
        RECT 47.390 35.820 48.155 36.300 ;
        RECT 50.290 35.820 51.055 36.300 ;
        RECT 53.190 35.820 53.955 36.300 ;
        RECT 56.090 35.820 56.855 36.300 ;
        RECT 58.990 35.820 59.755 36.300 ;
        RECT 61.890 35.820 62.655 36.300 ;
        RECT 64.790 35.820 65.555 36.300 ;
        RECT 67.690 35.820 68.455 36.300 ;
        RECT 70.590 35.820 71.355 36.300 ;
        RECT 73.490 35.820 74.255 36.300 ;
        RECT 76.390 35.820 77.155 36.300 ;
        RECT 79.290 35.820 80.055 36.300 ;
        RECT 82.190 35.820 82.955 36.300 ;
        RECT 85.090 35.820 85.855 36.300 ;
        RECT 87.990 35.820 88.755 36.300 ;
        RECT 90.890 35.820 91.655 36.300 ;
      LAYER li1 ;
        RECT 1.300 36.230 1.460 36.300 ;
        RECT 4.200 36.230 4.360 36.300 ;
        RECT 7.100 36.230 7.260 36.300 ;
        RECT 10.000 36.230 10.160 36.300 ;
        RECT 12.900 36.230 13.060 36.300 ;
        RECT 15.800 36.230 15.960 36.300 ;
        RECT 18.700 36.230 18.860 36.300 ;
        RECT 21.600 36.230 21.760 36.300 ;
        RECT 24.500 36.230 24.660 36.300 ;
        RECT 27.400 36.230 27.560 36.300 ;
        RECT 30.300 36.230 30.460 36.300 ;
        RECT 33.200 36.230 33.360 36.300 ;
        RECT 36.100 36.230 36.260 36.300 ;
        RECT 39.000 36.230 39.160 36.300 ;
        RECT 41.900 36.230 42.060 36.300 ;
        RECT 44.800 36.230 44.960 36.300 ;
        RECT 47.700 36.230 47.860 36.300 ;
        RECT 50.600 36.230 50.760 36.300 ;
        RECT 53.500 36.230 53.660 36.300 ;
        RECT 56.400 36.230 56.560 36.300 ;
        RECT 59.300 36.230 59.460 36.300 ;
        RECT 62.200 36.230 62.360 36.300 ;
        RECT 65.100 36.230 65.260 36.300 ;
        RECT 68.000 36.230 68.160 36.300 ;
        RECT 70.900 36.230 71.060 36.300 ;
        RECT 73.800 36.230 73.960 36.300 ;
        RECT 76.700 36.230 76.860 36.300 ;
        RECT 79.600 36.230 79.760 36.300 ;
        RECT 82.500 36.230 82.660 36.300 ;
        RECT 85.400 36.230 85.560 36.300 ;
        RECT 88.300 36.230 88.460 36.300 ;
        RECT 91.200 36.230 91.360 36.300 ;
        RECT 1.310 36.220 1.450 36.230 ;
        RECT 4.210 36.220 4.350 36.230 ;
        RECT 7.110 36.220 7.250 36.230 ;
        RECT 10.010 36.220 10.150 36.230 ;
        RECT 12.910 36.220 13.050 36.230 ;
        RECT 15.810 36.220 15.950 36.230 ;
        RECT 18.710 36.220 18.850 36.230 ;
        RECT 21.610 36.220 21.750 36.230 ;
        RECT 24.510 36.220 24.650 36.230 ;
        RECT 27.410 36.220 27.550 36.230 ;
        RECT 30.310 36.220 30.450 36.230 ;
        RECT 33.210 36.220 33.350 36.230 ;
        RECT 36.110 36.220 36.250 36.230 ;
        RECT 39.010 36.220 39.150 36.230 ;
        RECT 41.910 36.220 42.050 36.230 ;
        RECT 44.810 36.220 44.950 36.230 ;
        RECT 47.710 36.220 47.850 36.230 ;
        RECT 50.610 36.220 50.750 36.230 ;
        RECT 53.510 36.220 53.650 36.230 ;
        RECT 56.410 36.220 56.550 36.230 ;
        RECT 59.310 36.220 59.450 36.230 ;
        RECT 62.210 36.220 62.350 36.230 ;
        RECT 65.110 36.220 65.250 36.230 ;
        RECT 68.010 36.220 68.150 36.230 ;
        RECT 70.910 36.220 71.050 36.230 ;
        RECT 73.810 36.220 73.950 36.230 ;
        RECT 76.710 36.220 76.850 36.230 ;
        RECT 79.610 36.220 79.750 36.230 ;
        RECT 82.510 36.220 82.650 36.230 ;
        RECT 85.410 36.220 85.550 36.230 ;
        RECT 88.310 36.220 88.450 36.230 ;
        RECT 91.210 36.220 91.350 36.230 ;
      LAYER met1 ;
        RECT 0.000 36.230 92.660 36.300 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.990 34.470 1.755 34.950 ;
        RECT 3.890 34.470 4.655 34.950 ;
        RECT 6.790 34.470 7.555 34.950 ;
        RECT 9.690 34.470 10.455 34.950 ;
        RECT 12.590 34.470 13.355 34.950 ;
        RECT 15.490 34.470 16.255 34.950 ;
        RECT 18.390 34.470 19.155 34.950 ;
        RECT 21.290 34.470 22.055 34.950 ;
        RECT 24.190 34.470 24.955 34.950 ;
        RECT 27.090 34.470 27.855 34.950 ;
        RECT 29.990 34.470 30.755 34.950 ;
        RECT 32.890 34.470 33.655 34.950 ;
        RECT 35.790 34.470 36.555 34.950 ;
        RECT 38.690 34.470 39.455 34.950 ;
        RECT 41.590 34.470 42.355 34.950 ;
        RECT 44.490 34.470 45.255 34.950 ;
        RECT 47.390 34.470 48.155 34.950 ;
        RECT 50.290 34.470 51.055 34.950 ;
        RECT 53.190 34.470 53.955 34.950 ;
        RECT 56.090 34.470 56.855 34.950 ;
        RECT 58.990 34.470 59.755 34.950 ;
        RECT 61.890 34.470 62.655 34.950 ;
        RECT 64.790 34.470 65.555 34.950 ;
        RECT 67.690 34.470 68.455 34.950 ;
        RECT 70.590 34.470 71.355 34.950 ;
        RECT 73.490 34.470 74.255 34.950 ;
        RECT 76.390 34.470 77.155 34.950 ;
        RECT 79.290 34.470 80.055 34.950 ;
        RECT 82.190 34.470 82.955 34.950 ;
        RECT 85.090 34.470 85.855 34.950 ;
        RECT 87.990 34.470 88.755 34.950 ;
        RECT 90.890 34.470 91.655 34.950 ;
      LAYER li1 ;
        RECT 1.300 34.880 1.460 34.950 ;
        RECT 4.200 34.880 4.360 34.950 ;
        RECT 7.100 34.880 7.260 34.950 ;
        RECT 10.000 34.880 10.160 34.950 ;
        RECT 12.900 34.880 13.060 34.950 ;
        RECT 15.800 34.880 15.960 34.950 ;
        RECT 18.700 34.880 18.860 34.950 ;
        RECT 21.600 34.880 21.760 34.950 ;
        RECT 24.500 34.880 24.660 34.950 ;
        RECT 27.400 34.880 27.560 34.950 ;
        RECT 30.300 34.880 30.460 34.950 ;
        RECT 33.200 34.880 33.360 34.950 ;
        RECT 36.100 34.880 36.260 34.950 ;
        RECT 39.000 34.880 39.160 34.950 ;
        RECT 41.900 34.880 42.060 34.950 ;
        RECT 44.800 34.880 44.960 34.950 ;
        RECT 47.700 34.880 47.860 34.950 ;
        RECT 50.600 34.880 50.760 34.950 ;
        RECT 53.500 34.880 53.660 34.950 ;
        RECT 56.400 34.880 56.560 34.950 ;
        RECT 59.300 34.880 59.460 34.950 ;
        RECT 62.200 34.880 62.360 34.950 ;
        RECT 65.100 34.880 65.260 34.950 ;
        RECT 68.000 34.880 68.160 34.950 ;
        RECT 70.900 34.880 71.060 34.950 ;
        RECT 73.800 34.880 73.960 34.950 ;
        RECT 76.700 34.880 76.860 34.950 ;
        RECT 79.600 34.880 79.760 34.950 ;
        RECT 82.500 34.880 82.660 34.950 ;
        RECT 85.400 34.880 85.560 34.950 ;
        RECT 88.300 34.880 88.460 34.950 ;
        RECT 91.200 34.880 91.360 34.950 ;
        RECT 1.310 34.870 1.450 34.880 ;
        RECT 4.210 34.870 4.350 34.880 ;
        RECT 7.110 34.870 7.250 34.880 ;
        RECT 10.010 34.870 10.150 34.880 ;
        RECT 12.910 34.870 13.050 34.880 ;
        RECT 15.810 34.870 15.950 34.880 ;
        RECT 18.710 34.870 18.850 34.880 ;
        RECT 21.610 34.870 21.750 34.880 ;
        RECT 24.510 34.870 24.650 34.880 ;
        RECT 27.410 34.870 27.550 34.880 ;
        RECT 30.310 34.870 30.450 34.880 ;
        RECT 33.210 34.870 33.350 34.880 ;
        RECT 36.110 34.870 36.250 34.880 ;
        RECT 39.010 34.870 39.150 34.880 ;
        RECT 41.910 34.870 42.050 34.880 ;
        RECT 44.810 34.870 44.950 34.880 ;
        RECT 47.710 34.870 47.850 34.880 ;
        RECT 50.610 34.870 50.750 34.880 ;
        RECT 53.510 34.870 53.650 34.880 ;
        RECT 56.410 34.870 56.550 34.880 ;
        RECT 59.310 34.870 59.450 34.880 ;
        RECT 62.210 34.870 62.350 34.880 ;
        RECT 65.110 34.870 65.250 34.880 ;
        RECT 68.010 34.870 68.150 34.880 ;
        RECT 70.910 34.870 71.050 34.880 ;
        RECT 73.810 34.870 73.950 34.880 ;
        RECT 76.710 34.870 76.850 34.880 ;
        RECT 79.610 34.870 79.750 34.880 ;
        RECT 82.510 34.870 82.650 34.880 ;
        RECT 85.410 34.870 85.550 34.880 ;
        RECT 88.310 34.870 88.450 34.880 ;
        RECT 91.210 34.870 91.350 34.880 ;
      LAYER met1 ;
        RECT 0.000 34.880 92.660 34.950 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.990 33.120 1.755 33.600 ;
        RECT 3.890 33.120 4.655 33.600 ;
        RECT 6.790 33.120 7.555 33.600 ;
        RECT 9.690 33.120 10.455 33.600 ;
        RECT 12.590 33.120 13.355 33.600 ;
        RECT 15.490 33.120 16.255 33.600 ;
        RECT 18.390 33.120 19.155 33.600 ;
        RECT 21.290 33.120 22.055 33.600 ;
        RECT 24.190 33.120 24.955 33.600 ;
        RECT 27.090 33.120 27.855 33.600 ;
        RECT 29.990 33.120 30.755 33.600 ;
        RECT 32.890 33.120 33.655 33.600 ;
        RECT 35.790 33.120 36.555 33.600 ;
        RECT 38.690 33.120 39.455 33.600 ;
        RECT 41.590 33.120 42.355 33.600 ;
        RECT 44.490 33.120 45.255 33.600 ;
        RECT 47.390 33.120 48.155 33.600 ;
        RECT 50.290 33.120 51.055 33.600 ;
        RECT 53.190 33.120 53.955 33.600 ;
        RECT 56.090 33.120 56.855 33.600 ;
        RECT 58.990 33.120 59.755 33.600 ;
        RECT 61.890 33.120 62.655 33.600 ;
        RECT 64.790 33.120 65.555 33.600 ;
        RECT 67.690 33.120 68.455 33.600 ;
        RECT 70.590 33.120 71.355 33.600 ;
        RECT 73.490 33.120 74.255 33.600 ;
        RECT 76.390 33.120 77.155 33.600 ;
        RECT 79.290 33.120 80.055 33.600 ;
        RECT 82.190 33.120 82.955 33.600 ;
        RECT 85.090 33.120 85.855 33.600 ;
        RECT 87.990 33.120 88.755 33.600 ;
        RECT 90.890 33.120 91.655 33.600 ;
      LAYER li1 ;
        RECT 1.300 33.530 1.460 33.600 ;
        RECT 4.200 33.530 4.360 33.600 ;
        RECT 7.100 33.530 7.260 33.600 ;
        RECT 10.000 33.530 10.160 33.600 ;
        RECT 12.900 33.530 13.060 33.600 ;
        RECT 15.800 33.530 15.960 33.600 ;
        RECT 18.700 33.530 18.860 33.600 ;
        RECT 21.600 33.530 21.760 33.600 ;
        RECT 24.500 33.530 24.660 33.600 ;
        RECT 27.400 33.530 27.560 33.600 ;
        RECT 30.300 33.530 30.460 33.600 ;
        RECT 33.200 33.530 33.360 33.600 ;
        RECT 36.100 33.530 36.260 33.600 ;
        RECT 39.000 33.530 39.160 33.600 ;
        RECT 41.900 33.530 42.060 33.600 ;
        RECT 44.800 33.530 44.960 33.600 ;
        RECT 47.700 33.530 47.860 33.600 ;
        RECT 50.600 33.530 50.760 33.600 ;
        RECT 53.500 33.530 53.660 33.600 ;
        RECT 56.400 33.530 56.560 33.600 ;
        RECT 59.300 33.530 59.460 33.600 ;
        RECT 62.200 33.530 62.360 33.600 ;
        RECT 65.100 33.530 65.260 33.600 ;
        RECT 68.000 33.530 68.160 33.600 ;
        RECT 70.900 33.530 71.060 33.600 ;
        RECT 73.800 33.530 73.960 33.600 ;
        RECT 76.700 33.530 76.860 33.600 ;
        RECT 79.600 33.530 79.760 33.600 ;
        RECT 82.500 33.530 82.660 33.600 ;
        RECT 85.400 33.530 85.560 33.600 ;
        RECT 88.300 33.530 88.460 33.600 ;
        RECT 91.200 33.530 91.360 33.600 ;
        RECT 1.310 33.520 1.450 33.530 ;
        RECT 4.210 33.520 4.350 33.530 ;
        RECT 7.110 33.520 7.250 33.530 ;
        RECT 10.010 33.520 10.150 33.530 ;
        RECT 12.910 33.520 13.050 33.530 ;
        RECT 15.810 33.520 15.950 33.530 ;
        RECT 18.710 33.520 18.850 33.530 ;
        RECT 21.610 33.520 21.750 33.530 ;
        RECT 24.510 33.520 24.650 33.530 ;
        RECT 27.410 33.520 27.550 33.530 ;
        RECT 30.310 33.520 30.450 33.530 ;
        RECT 33.210 33.520 33.350 33.530 ;
        RECT 36.110 33.520 36.250 33.530 ;
        RECT 39.010 33.520 39.150 33.530 ;
        RECT 41.910 33.520 42.050 33.530 ;
        RECT 44.810 33.520 44.950 33.530 ;
        RECT 47.710 33.520 47.850 33.530 ;
        RECT 50.610 33.520 50.750 33.530 ;
        RECT 53.510 33.520 53.650 33.530 ;
        RECT 56.410 33.520 56.550 33.530 ;
        RECT 59.310 33.520 59.450 33.530 ;
        RECT 62.210 33.520 62.350 33.530 ;
        RECT 65.110 33.520 65.250 33.530 ;
        RECT 68.010 33.520 68.150 33.530 ;
        RECT 70.910 33.520 71.050 33.530 ;
        RECT 73.810 33.520 73.950 33.530 ;
        RECT 76.710 33.520 76.850 33.530 ;
        RECT 79.610 33.520 79.750 33.530 ;
        RECT 82.510 33.520 82.650 33.530 ;
        RECT 85.410 33.520 85.550 33.530 ;
        RECT 88.310 33.520 88.450 33.530 ;
        RECT 91.210 33.520 91.350 33.530 ;
      LAYER met1 ;
        RECT 0.000 33.530 92.660 33.600 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.990 31.770 1.755 32.250 ;
        RECT 3.890 31.770 4.655 32.250 ;
        RECT 6.790 31.770 7.555 32.250 ;
        RECT 9.690 31.770 10.455 32.250 ;
        RECT 12.590 31.770 13.355 32.250 ;
        RECT 15.490 31.770 16.255 32.250 ;
        RECT 18.390 31.770 19.155 32.250 ;
        RECT 21.290 31.770 22.055 32.250 ;
        RECT 24.190 31.770 24.955 32.250 ;
        RECT 27.090 31.770 27.855 32.250 ;
        RECT 29.990 31.770 30.755 32.250 ;
        RECT 32.890 31.770 33.655 32.250 ;
        RECT 35.790 31.770 36.555 32.250 ;
        RECT 38.690 31.770 39.455 32.250 ;
        RECT 41.590 31.770 42.355 32.250 ;
        RECT 44.490 31.770 45.255 32.250 ;
        RECT 47.390 31.770 48.155 32.250 ;
        RECT 50.290 31.770 51.055 32.250 ;
        RECT 53.190 31.770 53.955 32.250 ;
        RECT 56.090 31.770 56.855 32.250 ;
        RECT 58.990 31.770 59.755 32.250 ;
        RECT 61.890 31.770 62.655 32.250 ;
        RECT 64.790 31.770 65.555 32.250 ;
        RECT 67.690 31.770 68.455 32.250 ;
        RECT 70.590 31.770 71.355 32.250 ;
        RECT 73.490 31.770 74.255 32.250 ;
        RECT 76.390 31.770 77.155 32.250 ;
        RECT 79.290 31.770 80.055 32.250 ;
        RECT 82.190 31.770 82.955 32.250 ;
        RECT 85.090 31.770 85.855 32.250 ;
        RECT 87.990 31.770 88.755 32.250 ;
        RECT 90.890 31.770 91.655 32.250 ;
      LAYER li1 ;
        RECT 1.300 32.180 1.460 32.250 ;
        RECT 4.200 32.180 4.360 32.250 ;
        RECT 7.100 32.180 7.260 32.250 ;
        RECT 10.000 32.180 10.160 32.250 ;
        RECT 12.900 32.180 13.060 32.250 ;
        RECT 15.800 32.180 15.960 32.250 ;
        RECT 18.700 32.180 18.860 32.250 ;
        RECT 21.600 32.180 21.760 32.250 ;
        RECT 24.500 32.180 24.660 32.250 ;
        RECT 27.400 32.180 27.560 32.250 ;
        RECT 30.300 32.180 30.460 32.250 ;
        RECT 33.200 32.180 33.360 32.250 ;
        RECT 36.100 32.180 36.260 32.250 ;
        RECT 39.000 32.180 39.160 32.250 ;
        RECT 41.900 32.180 42.060 32.250 ;
        RECT 44.800 32.180 44.960 32.250 ;
        RECT 47.700 32.180 47.860 32.250 ;
        RECT 50.600 32.180 50.760 32.250 ;
        RECT 53.500 32.180 53.660 32.250 ;
        RECT 56.400 32.180 56.560 32.250 ;
        RECT 59.300 32.180 59.460 32.250 ;
        RECT 62.200 32.180 62.360 32.250 ;
        RECT 65.100 32.180 65.260 32.250 ;
        RECT 68.000 32.180 68.160 32.250 ;
        RECT 70.900 32.180 71.060 32.250 ;
        RECT 73.800 32.180 73.960 32.250 ;
        RECT 76.700 32.180 76.860 32.250 ;
        RECT 79.600 32.180 79.760 32.250 ;
        RECT 82.500 32.180 82.660 32.250 ;
        RECT 85.400 32.180 85.560 32.250 ;
        RECT 88.300 32.180 88.460 32.250 ;
        RECT 91.200 32.180 91.360 32.250 ;
        RECT 1.310 32.170 1.450 32.180 ;
        RECT 4.210 32.170 4.350 32.180 ;
        RECT 7.110 32.170 7.250 32.180 ;
        RECT 10.010 32.170 10.150 32.180 ;
        RECT 12.910 32.170 13.050 32.180 ;
        RECT 15.810 32.170 15.950 32.180 ;
        RECT 18.710 32.170 18.850 32.180 ;
        RECT 21.610 32.170 21.750 32.180 ;
        RECT 24.510 32.170 24.650 32.180 ;
        RECT 27.410 32.170 27.550 32.180 ;
        RECT 30.310 32.170 30.450 32.180 ;
        RECT 33.210 32.170 33.350 32.180 ;
        RECT 36.110 32.170 36.250 32.180 ;
        RECT 39.010 32.170 39.150 32.180 ;
        RECT 41.910 32.170 42.050 32.180 ;
        RECT 44.810 32.170 44.950 32.180 ;
        RECT 47.710 32.170 47.850 32.180 ;
        RECT 50.610 32.170 50.750 32.180 ;
        RECT 53.510 32.170 53.650 32.180 ;
        RECT 56.410 32.170 56.550 32.180 ;
        RECT 59.310 32.170 59.450 32.180 ;
        RECT 62.210 32.170 62.350 32.180 ;
        RECT 65.110 32.170 65.250 32.180 ;
        RECT 68.010 32.170 68.150 32.180 ;
        RECT 70.910 32.170 71.050 32.180 ;
        RECT 73.810 32.170 73.950 32.180 ;
        RECT 76.710 32.170 76.850 32.180 ;
        RECT 79.610 32.170 79.750 32.180 ;
        RECT 82.510 32.170 82.650 32.180 ;
        RECT 85.410 32.170 85.550 32.180 ;
        RECT 88.310 32.170 88.450 32.180 ;
        RECT 91.210 32.170 91.350 32.180 ;
      LAYER met1 ;
        RECT 0.000 32.180 92.660 32.250 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.990 30.420 1.755 30.900 ;
        RECT 3.890 30.420 4.655 30.900 ;
        RECT 6.790 30.420 7.555 30.900 ;
        RECT 9.690 30.420 10.455 30.900 ;
        RECT 12.590 30.420 13.355 30.900 ;
        RECT 15.490 30.420 16.255 30.900 ;
        RECT 18.390 30.420 19.155 30.900 ;
        RECT 21.290 30.420 22.055 30.900 ;
        RECT 24.190 30.420 24.955 30.900 ;
        RECT 27.090 30.420 27.855 30.900 ;
        RECT 29.990 30.420 30.755 30.900 ;
        RECT 32.890 30.420 33.655 30.900 ;
        RECT 35.790 30.420 36.555 30.900 ;
        RECT 38.690 30.420 39.455 30.900 ;
        RECT 41.590 30.420 42.355 30.900 ;
        RECT 44.490 30.420 45.255 30.900 ;
        RECT 47.390 30.420 48.155 30.900 ;
        RECT 50.290 30.420 51.055 30.900 ;
        RECT 53.190 30.420 53.955 30.900 ;
        RECT 56.090 30.420 56.855 30.900 ;
        RECT 58.990 30.420 59.755 30.900 ;
        RECT 61.890 30.420 62.655 30.900 ;
        RECT 64.790 30.420 65.555 30.900 ;
        RECT 67.690 30.420 68.455 30.900 ;
        RECT 70.590 30.420 71.355 30.900 ;
        RECT 73.490 30.420 74.255 30.900 ;
        RECT 76.390 30.420 77.155 30.900 ;
        RECT 79.290 30.420 80.055 30.900 ;
        RECT 82.190 30.420 82.955 30.900 ;
        RECT 85.090 30.420 85.855 30.900 ;
        RECT 87.990 30.420 88.755 30.900 ;
        RECT 90.890 30.420 91.655 30.900 ;
      LAYER li1 ;
        RECT 1.300 30.830 1.460 30.900 ;
        RECT 4.200 30.830 4.360 30.900 ;
        RECT 7.100 30.830 7.260 30.900 ;
        RECT 10.000 30.830 10.160 30.900 ;
        RECT 12.900 30.830 13.060 30.900 ;
        RECT 15.800 30.830 15.960 30.900 ;
        RECT 18.700 30.830 18.860 30.900 ;
        RECT 21.600 30.830 21.760 30.900 ;
        RECT 24.500 30.830 24.660 30.900 ;
        RECT 27.400 30.830 27.560 30.900 ;
        RECT 30.300 30.830 30.460 30.900 ;
        RECT 33.200 30.830 33.360 30.900 ;
        RECT 36.100 30.830 36.260 30.900 ;
        RECT 39.000 30.830 39.160 30.900 ;
        RECT 41.900 30.830 42.060 30.900 ;
        RECT 44.800 30.830 44.960 30.900 ;
        RECT 47.700 30.830 47.860 30.900 ;
        RECT 50.600 30.830 50.760 30.900 ;
        RECT 53.500 30.830 53.660 30.900 ;
        RECT 56.400 30.830 56.560 30.900 ;
        RECT 59.300 30.830 59.460 30.900 ;
        RECT 62.200 30.830 62.360 30.900 ;
        RECT 65.100 30.830 65.260 30.900 ;
        RECT 68.000 30.830 68.160 30.900 ;
        RECT 70.900 30.830 71.060 30.900 ;
        RECT 73.800 30.830 73.960 30.900 ;
        RECT 76.700 30.830 76.860 30.900 ;
        RECT 79.600 30.830 79.760 30.900 ;
        RECT 82.500 30.830 82.660 30.900 ;
        RECT 85.400 30.830 85.560 30.900 ;
        RECT 88.300 30.830 88.460 30.900 ;
        RECT 91.200 30.830 91.360 30.900 ;
        RECT 1.310 30.820 1.450 30.830 ;
        RECT 4.210 30.820 4.350 30.830 ;
        RECT 7.110 30.820 7.250 30.830 ;
        RECT 10.010 30.820 10.150 30.830 ;
        RECT 12.910 30.820 13.050 30.830 ;
        RECT 15.810 30.820 15.950 30.830 ;
        RECT 18.710 30.820 18.850 30.830 ;
        RECT 21.610 30.820 21.750 30.830 ;
        RECT 24.510 30.820 24.650 30.830 ;
        RECT 27.410 30.820 27.550 30.830 ;
        RECT 30.310 30.820 30.450 30.830 ;
        RECT 33.210 30.820 33.350 30.830 ;
        RECT 36.110 30.820 36.250 30.830 ;
        RECT 39.010 30.820 39.150 30.830 ;
        RECT 41.910 30.820 42.050 30.830 ;
        RECT 44.810 30.820 44.950 30.830 ;
        RECT 47.710 30.820 47.850 30.830 ;
        RECT 50.610 30.820 50.750 30.830 ;
        RECT 53.510 30.820 53.650 30.830 ;
        RECT 56.410 30.820 56.550 30.830 ;
        RECT 59.310 30.820 59.450 30.830 ;
        RECT 62.210 30.820 62.350 30.830 ;
        RECT 65.110 30.820 65.250 30.830 ;
        RECT 68.010 30.820 68.150 30.830 ;
        RECT 70.910 30.820 71.050 30.830 ;
        RECT 73.810 30.820 73.950 30.830 ;
        RECT 76.710 30.820 76.850 30.830 ;
        RECT 79.610 30.820 79.750 30.830 ;
        RECT 82.510 30.820 82.650 30.830 ;
        RECT 85.410 30.820 85.550 30.830 ;
        RECT 88.310 30.820 88.450 30.830 ;
        RECT 91.210 30.820 91.350 30.830 ;
      LAYER met1 ;
        RECT 0.000 30.830 92.660 30.900 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.990 29.070 1.755 29.550 ;
        RECT 3.890 29.070 4.655 29.550 ;
        RECT 6.790 29.070 7.555 29.550 ;
        RECT 9.690 29.070 10.455 29.550 ;
        RECT 12.590 29.070 13.355 29.550 ;
        RECT 15.490 29.070 16.255 29.550 ;
        RECT 18.390 29.070 19.155 29.550 ;
        RECT 21.290 29.070 22.055 29.550 ;
        RECT 24.190 29.070 24.955 29.550 ;
        RECT 27.090 29.070 27.855 29.550 ;
        RECT 29.990 29.070 30.755 29.550 ;
        RECT 32.890 29.070 33.655 29.550 ;
        RECT 35.790 29.070 36.555 29.550 ;
        RECT 38.690 29.070 39.455 29.550 ;
        RECT 41.590 29.070 42.355 29.550 ;
        RECT 44.490 29.070 45.255 29.550 ;
        RECT 47.390 29.070 48.155 29.550 ;
        RECT 50.290 29.070 51.055 29.550 ;
        RECT 53.190 29.070 53.955 29.550 ;
        RECT 56.090 29.070 56.855 29.550 ;
        RECT 58.990 29.070 59.755 29.550 ;
        RECT 61.890 29.070 62.655 29.550 ;
        RECT 64.790 29.070 65.555 29.550 ;
        RECT 67.690 29.070 68.455 29.550 ;
        RECT 70.590 29.070 71.355 29.550 ;
        RECT 73.490 29.070 74.255 29.550 ;
        RECT 76.390 29.070 77.155 29.550 ;
        RECT 79.290 29.070 80.055 29.550 ;
        RECT 82.190 29.070 82.955 29.550 ;
        RECT 85.090 29.070 85.855 29.550 ;
        RECT 87.990 29.070 88.755 29.550 ;
        RECT 90.890 29.070 91.655 29.550 ;
      LAYER li1 ;
        RECT 1.300 29.480 1.460 29.550 ;
        RECT 4.200 29.480 4.360 29.550 ;
        RECT 7.100 29.480 7.260 29.550 ;
        RECT 10.000 29.480 10.160 29.550 ;
        RECT 12.900 29.480 13.060 29.550 ;
        RECT 15.800 29.480 15.960 29.550 ;
        RECT 18.700 29.480 18.860 29.550 ;
        RECT 21.600 29.480 21.760 29.550 ;
        RECT 24.500 29.480 24.660 29.550 ;
        RECT 27.400 29.480 27.560 29.550 ;
        RECT 30.300 29.480 30.460 29.550 ;
        RECT 33.200 29.480 33.360 29.550 ;
        RECT 36.100 29.480 36.260 29.550 ;
        RECT 39.000 29.480 39.160 29.550 ;
        RECT 41.900 29.480 42.060 29.550 ;
        RECT 44.800 29.480 44.960 29.550 ;
        RECT 47.700 29.480 47.860 29.550 ;
        RECT 50.600 29.480 50.760 29.550 ;
        RECT 53.500 29.480 53.660 29.550 ;
        RECT 56.400 29.480 56.560 29.550 ;
        RECT 59.300 29.480 59.460 29.550 ;
        RECT 62.200 29.480 62.360 29.550 ;
        RECT 65.100 29.480 65.260 29.550 ;
        RECT 68.000 29.480 68.160 29.550 ;
        RECT 70.900 29.480 71.060 29.550 ;
        RECT 73.800 29.480 73.960 29.550 ;
        RECT 76.700 29.480 76.860 29.550 ;
        RECT 79.600 29.480 79.760 29.550 ;
        RECT 82.500 29.480 82.660 29.550 ;
        RECT 85.400 29.480 85.560 29.550 ;
        RECT 88.300 29.480 88.460 29.550 ;
        RECT 91.200 29.480 91.360 29.550 ;
        RECT 1.310 29.470 1.450 29.480 ;
        RECT 4.210 29.470 4.350 29.480 ;
        RECT 7.110 29.470 7.250 29.480 ;
        RECT 10.010 29.470 10.150 29.480 ;
        RECT 12.910 29.470 13.050 29.480 ;
        RECT 15.810 29.470 15.950 29.480 ;
        RECT 18.710 29.470 18.850 29.480 ;
        RECT 21.610 29.470 21.750 29.480 ;
        RECT 24.510 29.470 24.650 29.480 ;
        RECT 27.410 29.470 27.550 29.480 ;
        RECT 30.310 29.470 30.450 29.480 ;
        RECT 33.210 29.470 33.350 29.480 ;
        RECT 36.110 29.470 36.250 29.480 ;
        RECT 39.010 29.470 39.150 29.480 ;
        RECT 41.910 29.470 42.050 29.480 ;
        RECT 44.810 29.470 44.950 29.480 ;
        RECT 47.710 29.470 47.850 29.480 ;
        RECT 50.610 29.470 50.750 29.480 ;
        RECT 53.510 29.470 53.650 29.480 ;
        RECT 56.410 29.470 56.550 29.480 ;
        RECT 59.310 29.470 59.450 29.480 ;
        RECT 62.210 29.470 62.350 29.480 ;
        RECT 65.110 29.470 65.250 29.480 ;
        RECT 68.010 29.470 68.150 29.480 ;
        RECT 70.910 29.470 71.050 29.480 ;
        RECT 73.810 29.470 73.950 29.480 ;
        RECT 76.710 29.470 76.850 29.480 ;
        RECT 79.610 29.470 79.750 29.480 ;
        RECT 82.510 29.470 82.650 29.480 ;
        RECT 85.410 29.470 85.550 29.480 ;
        RECT 88.310 29.470 88.450 29.480 ;
        RECT 91.210 29.470 91.350 29.480 ;
      LAYER met1 ;
        RECT 0.000 29.480 92.660 29.550 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.990 27.720 1.755 28.200 ;
        RECT 3.890 27.720 4.655 28.200 ;
        RECT 6.790 27.720 7.555 28.200 ;
        RECT 9.690 27.720 10.455 28.200 ;
        RECT 12.590 27.720 13.355 28.200 ;
        RECT 15.490 27.720 16.255 28.200 ;
        RECT 18.390 27.720 19.155 28.200 ;
        RECT 21.290 27.720 22.055 28.200 ;
        RECT 24.190 27.720 24.955 28.200 ;
        RECT 27.090 27.720 27.855 28.200 ;
        RECT 29.990 27.720 30.755 28.200 ;
        RECT 32.890 27.720 33.655 28.200 ;
        RECT 35.790 27.720 36.555 28.200 ;
        RECT 38.690 27.720 39.455 28.200 ;
        RECT 41.590 27.720 42.355 28.200 ;
        RECT 44.490 27.720 45.255 28.200 ;
        RECT 47.390 27.720 48.155 28.200 ;
        RECT 50.290 27.720 51.055 28.200 ;
        RECT 53.190 27.720 53.955 28.200 ;
        RECT 56.090 27.720 56.855 28.200 ;
        RECT 58.990 27.720 59.755 28.200 ;
        RECT 61.890 27.720 62.655 28.200 ;
        RECT 64.790 27.720 65.555 28.200 ;
        RECT 67.690 27.720 68.455 28.200 ;
        RECT 70.590 27.720 71.355 28.200 ;
        RECT 73.490 27.720 74.255 28.200 ;
        RECT 76.390 27.720 77.155 28.200 ;
        RECT 79.290 27.720 80.055 28.200 ;
        RECT 82.190 27.720 82.955 28.200 ;
        RECT 85.090 27.720 85.855 28.200 ;
        RECT 87.990 27.720 88.755 28.200 ;
        RECT 90.890 27.720 91.655 28.200 ;
      LAYER li1 ;
        RECT 1.300 28.130 1.460 28.200 ;
        RECT 4.200 28.130 4.360 28.200 ;
        RECT 7.100 28.130 7.260 28.200 ;
        RECT 10.000 28.130 10.160 28.200 ;
        RECT 12.900 28.130 13.060 28.200 ;
        RECT 15.800 28.130 15.960 28.200 ;
        RECT 18.700 28.130 18.860 28.200 ;
        RECT 21.600 28.130 21.760 28.200 ;
        RECT 24.500 28.130 24.660 28.200 ;
        RECT 27.400 28.130 27.560 28.200 ;
        RECT 30.300 28.130 30.460 28.200 ;
        RECT 33.200 28.130 33.360 28.200 ;
        RECT 36.100 28.130 36.260 28.200 ;
        RECT 39.000 28.130 39.160 28.200 ;
        RECT 41.900 28.130 42.060 28.200 ;
        RECT 44.800 28.130 44.960 28.200 ;
        RECT 47.700 28.130 47.860 28.200 ;
        RECT 50.600 28.130 50.760 28.200 ;
        RECT 53.500 28.130 53.660 28.200 ;
        RECT 56.400 28.130 56.560 28.200 ;
        RECT 59.300 28.130 59.460 28.200 ;
        RECT 62.200 28.130 62.360 28.200 ;
        RECT 65.100 28.130 65.260 28.200 ;
        RECT 68.000 28.130 68.160 28.200 ;
        RECT 70.900 28.130 71.060 28.200 ;
        RECT 73.800 28.130 73.960 28.200 ;
        RECT 76.700 28.130 76.860 28.200 ;
        RECT 79.600 28.130 79.760 28.200 ;
        RECT 82.500 28.130 82.660 28.200 ;
        RECT 85.400 28.130 85.560 28.200 ;
        RECT 88.300 28.130 88.460 28.200 ;
        RECT 91.200 28.130 91.360 28.200 ;
        RECT 1.310 28.120 1.450 28.130 ;
        RECT 4.210 28.120 4.350 28.130 ;
        RECT 7.110 28.120 7.250 28.130 ;
        RECT 10.010 28.120 10.150 28.130 ;
        RECT 12.910 28.120 13.050 28.130 ;
        RECT 15.810 28.120 15.950 28.130 ;
        RECT 18.710 28.120 18.850 28.130 ;
        RECT 21.610 28.120 21.750 28.130 ;
        RECT 24.510 28.120 24.650 28.130 ;
        RECT 27.410 28.120 27.550 28.130 ;
        RECT 30.310 28.120 30.450 28.130 ;
        RECT 33.210 28.120 33.350 28.130 ;
        RECT 36.110 28.120 36.250 28.130 ;
        RECT 39.010 28.120 39.150 28.130 ;
        RECT 41.910 28.120 42.050 28.130 ;
        RECT 44.810 28.120 44.950 28.130 ;
        RECT 47.710 28.120 47.850 28.130 ;
        RECT 50.610 28.120 50.750 28.130 ;
        RECT 53.510 28.120 53.650 28.130 ;
        RECT 56.410 28.120 56.550 28.130 ;
        RECT 59.310 28.120 59.450 28.130 ;
        RECT 62.210 28.120 62.350 28.130 ;
        RECT 65.110 28.120 65.250 28.130 ;
        RECT 68.010 28.120 68.150 28.130 ;
        RECT 70.910 28.120 71.050 28.130 ;
        RECT 73.810 28.120 73.950 28.130 ;
        RECT 76.710 28.120 76.850 28.130 ;
        RECT 79.610 28.120 79.750 28.130 ;
        RECT 82.510 28.120 82.650 28.130 ;
        RECT 85.410 28.120 85.550 28.130 ;
        RECT 88.310 28.120 88.450 28.130 ;
        RECT 91.210 28.120 91.350 28.130 ;
      LAYER met1 ;
        RECT 0.000 28.130 92.660 28.200 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.990 26.370 1.755 26.850 ;
        RECT 3.890 26.370 4.655 26.850 ;
        RECT 6.790 26.370 7.555 26.850 ;
        RECT 9.690 26.370 10.455 26.850 ;
        RECT 12.590 26.370 13.355 26.850 ;
        RECT 15.490 26.370 16.255 26.850 ;
        RECT 18.390 26.370 19.155 26.850 ;
        RECT 21.290 26.370 22.055 26.850 ;
        RECT 24.190 26.370 24.955 26.850 ;
        RECT 27.090 26.370 27.855 26.850 ;
        RECT 29.990 26.370 30.755 26.850 ;
        RECT 32.890 26.370 33.655 26.850 ;
        RECT 35.790 26.370 36.555 26.850 ;
        RECT 38.690 26.370 39.455 26.850 ;
        RECT 41.590 26.370 42.355 26.850 ;
        RECT 44.490 26.370 45.255 26.850 ;
        RECT 47.390 26.370 48.155 26.850 ;
        RECT 50.290 26.370 51.055 26.850 ;
        RECT 53.190 26.370 53.955 26.850 ;
        RECT 56.090 26.370 56.855 26.850 ;
        RECT 58.990 26.370 59.755 26.850 ;
        RECT 61.890 26.370 62.655 26.850 ;
        RECT 64.790 26.370 65.555 26.850 ;
        RECT 67.690 26.370 68.455 26.850 ;
        RECT 70.590 26.370 71.355 26.850 ;
        RECT 73.490 26.370 74.255 26.850 ;
        RECT 76.390 26.370 77.155 26.850 ;
        RECT 79.290 26.370 80.055 26.850 ;
        RECT 82.190 26.370 82.955 26.850 ;
        RECT 85.090 26.370 85.855 26.850 ;
        RECT 87.990 26.370 88.755 26.850 ;
        RECT 90.890 26.370 91.655 26.850 ;
      LAYER li1 ;
        RECT 1.300 26.780 1.460 26.850 ;
        RECT 4.200 26.780 4.360 26.850 ;
        RECT 7.100 26.780 7.260 26.850 ;
        RECT 10.000 26.780 10.160 26.850 ;
        RECT 12.900 26.780 13.060 26.850 ;
        RECT 15.800 26.780 15.960 26.850 ;
        RECT 18.700 26.780 18.860 26.850 ;
        RECT 21.600 26.780 21.760 26.850 ;
        RECT 24.500 26.780 24.660 26.850 ;
        RECT 27.400 26.780 27.560 26.850 ;
        RECT 30.300 26.780 30.460 26.850 ;
        RECT 33.200 26.780 33.360 26.850 ;
        RECT 36.100 26.780 36.260 26.850 ;
        RECT 39.000 26.780 39.160 26.850 ;
        RECT 41.900 26.780 42.060 26.850 ;
        RECT 44.800 26.780 44.960 26.850 ;
        RECT 47.700 26.780 47.860 26.850 ;
        RECT 50.600 26.780 50.760 26.850 ;
        RECT 53.500 26.780 53.660 26.850 ;
        RECT 56.400 26.780 56.560 26.850 ;
        RECT 59.300 26.780 59.460 26.850 ;
        RECT 62.200 26.780 62.360 26.850 ;
        RECT 65.100 26.780 65.260 26.850 ;
        RECT 68.000 26.780 68.160 26.850 ;
        RECT 70.900 26.780 71.060 26.850 ;
        RECT 73.800 26.780 73.960 26.850 ;
        RECT 76.700 26.780 76.860 26.850 ;
        RECT 79.600 26.780 79.760 26.850 ;
        RECT 82.500 26.780 82.660 26.850 ;
        RECT 85.400 26.780 85.560 26.850 ;
        RECT 88.300 26.780 88.460 26.850 ;
        RECT 91.200 26.780 91.360 26.850 ;
        RECT 1.310 26.770 1.450 26.780 ;
        RECT 4.210 26.770 4.350 26.780 ;
        RECT 7.110 26.770 7.250 26.780 ;
        RECT 10.010 26.770 10.150 26.780 ;
        RECT 12.910 26.770 13.050 26.780 ;
        RECT 15.810 26.770 15.950 26.780 ;
        RECT 18.710 26.770 18.850 26.780 ;
        RECT 21.610 26.770 21.750 26.780 ;
        RECT 24.510 26.770 24.650 26.780 ;
        RECT 27.410 26.770 27.550 26.780 ;
        RECT 30.310 26.770 30.450 26.780 ;
        RECT 33.210 26.770 33.350 26.780 ;
        RECT 36.110 26.770 36.250 26.780 ;
        RECT 39.010 26.770 39.150 26.780 ;
        RECT 41.910 26.770 42.050 26.780 ;
        RECT 44.810 26.770 44.950 26.780 ;
        RECT 47.710 26.770 47.850 26.780 ;
        RECT 50.610 26.770 50.750 26.780 ;
        RECT 53.510 26.770 53.650 26.780 ;
        RECT 56.410 26.770 56.550 26.780 ;
        RECT 59.310 26.770 59.450 26.780 ;
        RECT 62.210 26.770 62.350 26.780 ;
        RECT 65.110 26.770 65.250 26.780 ;
        RECT 68.010 26.770 68.150 26.780 ;
        RECT 70.910 26.770 71.050 26.780 ;
        RECT 73.810 26.770 73.950 26.780 ;
        RECT 76.710 26.770 76.850 26.780 ;
        RECT 79.610 26.770 79.750 26.780 ;
        RECT 82.510 26.770 82.650 26.780 ;
        RECT 85.410 26.770 85.550 26.780 ;
        RECT 88.310 26.770 88.450 26.780 ;
        RECT 91.210 26.770 91.350 26.780 ;
      LAYER met1 ;
        RECT 0.000 26.780 92.660 26.850 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.990 25.020 1.755 25.500 ;
        RECT 3.890 25.020 4.655 25.500 ;
        RECT 6.790 25.020 7.555 25.500 ;
        RECT 9.690 25.020 10.455 25.500 ;
        RECT 12.590 25.020 13.355 25.500 ;
        RECT 15.490 25.020 16.255 25.500 ;
        RECT 18.390 25.020 19.155 25.500 ;
        RECT 21.290 25.020 22.055 25.500 ;
        RECT 24.190 25.020 24.955 25.500 ;
        RECT 27.090 25.020 27.855 25.500 ;
        RECT 29.990 25.020 30.755 25.500 ;
        RECT 32.890 25.020 33.655 25.500 ;
        RECT 35.790 25.020 36.555 25.500 ;
        RECT 38.690 25.020 39.455 25.500 ;
        RECT 41.590 25.020 42.355 25.500 ;
        RECT 44.490 25.020 45.255 25.500 ;
        RECT 47.390 25.020 48.155 25.500 ;
        RECT 50.290 25.020 51.055 25.500 ;
        RECT 53.190 25.020 53.955 25.500 ;
        RECT 56.090 25.020 56.855 25.500 ;
        RECT 58.990 25.020 59.755 25.500 ;
        RECT 61.890 25.020 62.655 25.500 ;
        RECT 64.790 25.020 65.555 25.500 ;
        RECT 67.690 25.020 68.455 25.500 ;
        RECT 70.590 25.020 71.355 25.500 ;
        RECT 73.490 25.020 74.255 25.500 ;
        RECT 76.390 25.020 77.155 25.500 ;
        RECT 79.290 25.020 80.055 25.500 ;
        RECT 82.190 25.020 82.955 25.500 ;
        RECT 85.090 25.020 85.855 25.500 ;
        RECT 87.990 25.020 88.755 25.500 ;
        RECT 90.890 25.020 91.655 25.500 ;
      LAYER li1 ;
        RECT 1.300 25.430 1.460 25.500 ;
        RECT 4.200 25.430 4.360 25.500 ;
        RECT 7.100 25.430 7.260 25.500 ;
        RECT 10.000 25.430 10.160 25.500 ;
        RECT 12.900 25.430 13.060 25.500 ;
        RECT 15.800 25.430 15.960 25.500 ;
        RECT 18.700 25.430 18.860 25.500 ;
        RECT 21.600 25.430 21.760 25.500 ;
        RECT 24.500 25.430 24.660 25.500 ;
        RECT 27.400 25.430 27.560 25.500 ;
        RECT 30.300 25.430 30.460 25.500 ;
        RECT 33.200 25.430 33.360 25.500 ;
        RECT 36.100 25.430 36.260 25.500 ;
        RECT 39.000 25.430 39.160 25.500 ;
        RECT 41.900 25.430 42.060 25.500 ;
        RECT 44.800 25.430 44.960 25.500 ;
        RECT 47.700 25.430 47.860 25.500 ;
        RECT 50.600 25.430 50.760 25.500 ;
        RECT 53.500 25.430 53.660 25.500 ;
        RECT 56.400 25.430 56.560 25.500 ;
        RECT 59.300 25.430 59.460 25.500 ;
        RECT 62.200 25.430 62.360 25.500 ;
        RECT 65.100 25.430 65.260 25.500 ;
        RECT 68.000 25.430 68.160 25.500 ;
        RECT 70.900 25.430 71.060 25.500 ;
        RECT 73.800 25.430 73.960 25.500 ;
        RECT 76.700 25.430 76.860 25.500 ;
        RECT 79.600 25.430 79.760 25.500 ;
        RECT 82.500 25.430 82.660 25.500 ;
        RECT 85.400 25.430 85.560 25.500 ;
        RECT 88.300 25.430 88.460 25.500 ;
        RECT 91.200 25.430 91.360 25.500 ;
        RECT 1.310 25.420 1.450 25.430 ;
        RECT 4.210 25.420 4.350 25.430 ;
        RECT 7.110 25.420 7.250 25.430 ;
        RECT 10.010 25.420 10.150 25.430 ;
        RECT 12.910 25.420 13.050 25.430 ;
        RECT 15.810 25.420 15.950 25.430 ;
        RECT 18.710 25.420 18.850 25.430 ;
        RECT 21.610 25.420 21.750 25.430 ;
        RECT 24.510 25.420 24.650 25.430 ;
        RECT 27.410 25.420 27.550 25.430 ;
        RECT 30.310 25.420 30.450 25.430 ;
        RECT 33.210 25.420 33.350 25.430 ;
        RECT 36.110 25.420 36.250 25.430 ;
        RECT 39.010 25.420 39.150 25.430 ;
        RECT 41.910 25.420 42.050 25.430 ;
        RECT 44.810 25.420 44.950 25.430 ;
        RECT 47.710 25.420 47.850 25.430 ;
        RECT 50.610 25.420 50.750 25.430 ;
        RECT 53.510 25.420 53.650 25.430 ;
        RECT 56.410 25.420 56.550 25.430 ;
        RECT 59.310 25.420 59.450 25.430 ;
        RECT 62.210 25.420 62.350 25.430 ;
        RECT 65.110 25.420 65.250 25.430 ;
        RECT 68.010 25.420 68.150 25.430 ;
        RECT 70.910 25.420 71.050 25.430 ;
        RECT 73.810 25.420 73.950 25.430 ;
        RECT 76.710 25.420 76.850 25.430 ;
        RECT 79.610 25.420 79.750 25.430 ;
        RECT 82.510 25.420 82.650 25.430 ;
        RECT 85.410 25.420 85.550 25.430 ;
        RECT 88.310 25.420 88.450 25.430 ;
        RECT 91.210 25.420 91.350 25.430 ;
      LAYER met1 ;
        RECT 0.000 25.430 92.660 25.500 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.990 23.670 1.755 24.150 ;
        RECT 3.890 23.670 4.655 24.150 ;
        RECT 6.790 23.670 7.555 24.150 ;
        RECT 9.690 23.670 10.455 24.150 ;
        RECT 12.590 23.670 13.355 24.150 ;
        RECT 15.490 23.670 16.255 24.150 ;
        RECT 18.390 23.670 19.155 24.150 ;
        RECT 21.290 23.670 22.055 24.150 ;
        RECT 24.190 23.670 24.955 24.150 ;
        RECT 27.090 23.670 27.855 24.150 ;
        RECT 29.990 23.670 30.755 24.150 ;
        RECT 32.890 23.670 33.655 24.150 ;
        RECT 35.790 23.670 36.555 24.150 ;
        RECT 38.690 23.670 39.455 24.150 ;
        RECT 41.590 23.670 42.355 24.150 ;
        RECT 44.490 23.670 45.255 24.150 ;
        RECT 47.390 23.670 48.155 24.150 ;
        RECT 50.290 23.670 51.055 24.150 ;
        RECT 53.190 23.670 53.955 24.150 ;
        RECT 56.090 23.670 56.855 24.150 ;
        RECT 58.990 23.670 59.755 24.150 ;
        RECT 61.890 23.670 62.655 24.150 ;
        RECT 64.790 23.670 65.555 24.150 ;
        RECT 67.690 23.670 68.455 24.150 ;
        RECT 70.590 23.670 71.355 24.150 ;
        RECT 73.490 23.670 74.255 24.150 ;
        RECT 76.390 23.670 77.155 24.150 ;
        RECT 79.290 23.670 80.055 24.150 ;
        RECT 82.190 23.670 82.955 24.150 ;
        RECT 85.090 23.670 85.855 24.150 ;
        RECT 87.990 23.670 88.755 24.150 ;
        RECT 90.890 23.670 91.655 24.150 ;
      LAYER li1 ;
        RECT 1.300 24.080 1.460 24.150 ;
        RECT 4.200 24.080 4.360 24.150 ;
        RECT 7.100 24.080 7.260 24.150 ;
        RECT 10.000 24.080 10.160 24.150 ;
        RECT 12.900 24.080 13.060 24.150 ;
        RECT 15.800 24.080 15.960 24.150 ;
        RECT 18.700 24.080 18.860 24.150 ;
        RECT 21.600 24.080 21.760 24.150 ;
        RECT 24.500 24.080 24.660 24.150 ;
        RECT 27.400 24.080 27.560 24.150 ;
        RECT 30.300 24.080 30.460 24.150 ;
        RECT 33.200 24.080 33.360 24.150 ;
        RECT 36.100 24.080 36.260 24.150 ;
        RECT 39.000 24.080 39.160 24.150 ;
        RECT 41.900 24.080 42.060 24.150 ;
        RECT 44.800 24.080 44.960 24.150 ;
        RECT 47.700 24.080 47.860 24.150 ;
        RECT 50.600 24.080 50.760 24.150 ;
        RECT 53.500 24.080 53.660 24.150 ;
        RECT 56.400 24.080 56.560 24.150 ;
        RECT 59.300 24.080 59.460 24.150 ;
        RECT 62.200 24.080 62.360 24.150 ;
        RECT 65.100 24.080 65.260 24.150 ;
        RECT 68.000 24.080 68.160 24.150 ;
        RECT 70.900 24.080 71.060 24.150 ;
        RECT 73.800 24.080 73.960 24.150 ;
        RECT 76.700 24.080 76.860 24.150 ;
        RECT 79.600 24.080 79.760 24.150 ;
        RECT 82.500 24.080 82.660 24.150 ;
        RECT 85.400 24.080 85.560 24.150 ;
        RECT 88.300 24.080 88.460 24.150 ;
        RECT 91.200 24.080 91.360 24.150 ;
        RECT 1.310 24.070 1.450 24.080 ;
        RECT 4.210 24.070 4.350 24.080 ;
        RECT 7.110 24.070 7.250 24.080 ;
        RECT 10.010 24.070 10.150 24.080 ;
        RECT 12.910 24.070 13.050 24.080 ;
        RECT 15.810 24.070 15.950 24.080 ;
        RECT 18.710 24.070 18.850 24.080 ;
        RECT 21.610 24.070 21.750 24.080 ;
        RECT 24.510 24.070 24.650 24.080 ;
        RECT 27.410 24.070 27.550 24.080 ;
        RECT 30.310 24.070 30.450 24.080 ;
        RECT 33.210 24.070 33.350 24.080 ;
        RECT 36.110 24.070 36.250 24.080 ;
        RECT 39.010 24.070 39.150 24.080 ;
        RECT 41.910 24.070 42.050 24.080 ;
        RECT 44.810 24.070 44.950 24.080 ;
        RECT 47.710 24.070 47.850 24.080 ;
        RECT 50.610 24.070 50.750 24.080 ;
        RECT 53.510 24.070 53.650 24.080 ;
        RECT 56.410 24.070 56.550 24.080 ;
        RECT 59.310 24.070 59.450 24.080 ;
        RECT 62.210 24.070 62.350 24.080 ;
        RECT 65.110 24.070 65.250 24.080 ;
        RECT 68.010 24.070 68.150 24.080 ;
        RECT 70.910 24.070 71.050 24.080 ;
        RECT 73.810 24.070 73.950 24.080 ;
        RECT 76.710 24.070 76.850 24.080 ;
        RECT 79.610 24.070 79.750 24.080 ;
        RECT 82.510 24.070 82.650 24.080 ;
        RECT 85.410 24.070 85.550 24.080 ;
        RECT 88.310 24.070 88.450 24.080 ;
        RECT 91.210 24.070 91.350 24.080 ;
      LAYER met1 ;
        RECT 0.000 24.080 92.660 24.150 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.990 22.320 1.755 22.800 ;
        RECT 3.890 22.320 4.655 22.800 ;
        RECT 6.790 22.320 7.555 22.800 ;
        RECT 9.690 22.320 10.455 22.800 ;
        RECT 12.590 22.320 13.355 22.800 ;
        RECT 15.490 22.320 16.255 22.800 ;
        RECT 18.390 22.320 19.155 22.800 ;
        RECT 21.290 22.320 22.055 22.800 ;
        RECT 24.190 22.320 24.955 22.800 ;
        RECT 27.090 22.320 27.855 22.800 ;
        RECT 29.990 22.320 30.755 22.800 ;
        RECT 32.890 22.320 33.655 22.800 ;
        RECT 35.790 22.320 36.555 22.800 ;
        RECT 38.690 22.320 39.455 22.800 ;
        RECT 41.590 22.320 42.355 22.800 ;
        RECT 44.490 22.320 45.255 22.800 ;
        RECT 47.390 22.320 48.155 22.800 ;
        RECT 50.290 22.320 51.055 22.800 ;
        RECT 53.190 22.320 53.955 22.800 ;
        RECT 56.090 22.320 56.855 22.800 ;
        RECT 58.990 22.320 59.755 22.800 ;
        RECT 61.890 22.320 62.655 22.800 ;
        RECT 64.790 22.320 65.555 22.800 ;
        RECT 67.690 22.320 68.455 22.800 ;
        RECT 70.590 22.320 71.355 22.800 ;
        RECT 73.490 22.320 74.255 22.800 ;
        RECT 76.390 22.320 77.155 22.800 ;
        RECT 79.290 22.320 80.055 22.800 ;
        RECT 82.190 22.320 82.955 22.800 ;
        RECT 85.090 22.320 85.855 22.800 ;
        RECT 87.990 22.320 88.755 22.800 ;
        RECT 90.890 22.320 91.655 22.800 ;
      LAYER li1 ;
        RECT 1.300 22.730 1.460 22.800 ;
        RECT 4.200 22.730 4.360 22.800 ;
        RECT 7.100 22.730 7.260 22.800 ;
        RECT 10.000 22.730 10.160 22.800 ;
        RECT 12.900 22.730 13.060 22.800 ;
        RECT 15.800 22.730 15.960 22.800 ;
        RECT 18.700 22.730 18.860 22.800 ;
        RECT 21.600 22.730 21.760 22.800 ;
        RECT 24.500 22.730 24.660 22.800 ;
        RECT 27.400 22.730 27.560 22.800 ;
        RECT 30.300 22.730 30.460 22.800 ;
        RECT 33.200 22.730 33.360 22.800 ;
        RECT 36.100 22.730 36.260 22.800 ;
        RECT 39.000 22.730 39.160 22.800 ;
        RECT 41.900 22.730 42.060 22.800 ;
        RECT 44.800 22.730 44.960 22.800 ;
        RECT 47.700 22.730 47.860 22.800 ;
        RECT 50.600 22.730 50.760 22.800 ;
        RECT 53.500 22.730 53.660 22.800 ;
        RECT 56.400 22.730 56.560 22.800 ;
        RECT 59.300 22.730 59.460 22.800 ;
        RECT 62.200 22.730 62.360 22.800 ;
        RECT 65.100 22.730 65.260 22.800 ;
        RECT 68.000 22.730 68.160 22.800 ;
        RECT 70.900 22.730 71.060 22.800 ;
        RECT 73.800 22.730 73.960 22.800 ;
        RECT 76.700 22.730 76.860 22.800 ;
        RECT 79.600 22.730 79.760 22.800 ;
        RECT 82.500 22.730 82.660 22.800 ;
        RECT 85.400 22.730 85.560 22.800 ;
        RECT 88.300 22.730 88.460 22.800 ;
        RECT 91.200 22.730 91.360 22.800 ;
        RECT 1.310 22.720 1.450 22.730 ;
        RECT 4.210 22.720 4.350 22.730 ;
        RECT 7.110 22.720 7.250 22.730 ;
        RECT 10.010 22.720 10.150 22.730 ;
        RECT 12.910 22.720 13.050 22.730 ;
        RECT 15.810 22.720 15.950 22.730 ;
        RECT 18.710 22.720 18.850 22.730 ;
        RECT 21.610 22.720 21.750 22.730 ;
        RECT 24.510 22.720 24.650 22.730 ;
        RECT 27.410 22.720 27.550 22.730 ;
        RECT 30.310 22.720 30.450 22.730 ;
        RECT 33.210 22.720 33.350 22.730 ;
        RECT 36.110 22.720 36.250 22.730 ;
        RECT 39.010 22.720 39.150 22.730 ;
        RECT 41.910 22.720 42.050 22.730 ;
        RECT 44.810 22.720 44.950 22.730 ;
        RECT 47.710 22.720 47.850 22.730 ;
        RECT 50.610 22.720 50.750 22.730 ;
        RECT 53.510 22.720 53.650 22.730 ;
        RECT 56.410 22.720 56.550 22.730 ;
        RECT 59.310 22.720 59.450 22.730 ;
        RECT 62.210 22.720 62.350 22.730 ;
        RECT 65.110 22.720 65.250 22.730 ;
        RECT 68.010 22.720 68.150 22.730 ;
        RECT 70.910 22.720 71.050 22.730 ;
        RECT 73.810 22.720 73.950 22.730 ;
        RECT 76.710 22.720 76.850 22.730 ;
        RECT 79.610 22.720 79.750 22.730 ;
        RECT 82.510 22.720 82.650 22.730 ;
        RECT 85.410 22.720 85.550 22.730 ;
        RECT 88.310 22.720 88.450 22.730 ;
        RECT 91.210 22.720 91.350 22.730 ;
      LAYER met1 ;
        RECT 0.000 22.730 92.660 22.800 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.990 20.970 1.755 21.450 ;
        RECT 3.890 20.970 4.655 21.450 ;
        RECT 6.790 20.970 7.555 21.450 ;
        RECT 9.690 20.970 10.455 21.450 ;
        RECT 12.590 20.970 13.355 21.450 ;
        RECT 15.490 20.970 16.255 21.450 ;
        RECT 18.390 20.970 19.155 21.450 ;
        RECT 21.290 20.970 22.055 21.450 ;
        RECT 24.190 20.970 24.955 21.450 ;
        RECT 27.090 20.970 27.855 21.450 ;
        RECT 29.990 20.970 30.755 21.450 ;
        RECT 32.890 20.970 33.655 21.450 ;
        RECT 35.790 20.970 36.555 21.450 ;
        RECT 38.690 20.970 39.455 21.450 ;
        RECT 41.590 20.970 42.355 21.450 ;
        RECT 44.490 20.970 45.255 21.450 ;
        RECT 47.390 20.970 48.155 21.450 ;
        RECT 50.290 20.970 51.055 21.450 ;
        RECT 53.190 20.970 53.955 21.450 ;
        RECT 56.090 20.970 56.855 21.450 ;
        RECT 58.990 20.970 59.755 21.450 ;
        RECT 61.890 20.970 62.655 21.450 ;
        RECT 64.790 20.970 65.555 21.450 ;
        RECT 67.690 20.970 68.455 21.450 ;
        RECT 70.590 20.970 71.355 21.450 ;
        RECT 73.490 20.970 74.255 21.450 ;
        RECT 76.390 20.970 77.155 21.450 ;
        RECT 79.290 20.970 80.055 21.450 ;
        RECT 82.190 20.970 82.955 21.450 ;
        RECT 85.090 20.970 85.855 21.450 ;
        RECT 87.990 20.970 88.755 21.450 ;
        RECT 90.890 20.970 91.655 21.450 ;
      LAYER li1 ;
        RECT 1.300 21.380 1.460 21.450 ;
        RECT 4.200 21.380 4.360 21.450 ;
        RECT 7.100 21.380 7.260 21.450 ;
        RECT 10.000 21.380 10.160 21.450 ;
        RECT 12.900 21.380 13.060 21.450 ;
        RECT 15.800 21.380 15.960 21.450 ;
        RECT 18.700 21.380 18.860 21.450 ;
        RECT 21.600 21.380 21.760 21.450 ;
        RECT 24.500 21.380 24.660 21.450 ;
        RECT 27.400 21.380 27.560 21.450 ;
        RECT 30.300 21.380 30.460 21.450 ;
        RECT 33.200 21.380 33.360 21.450 ;
        RECT 36.100 21.380 36.260 21.450 ;
        RECT 39.000 21.380 39.160 21.450 ;
        RECT 41.900 21.380 42.060 21.450 ;
        RECT 44.800 21.380 44.960 21.450 ;
        RECT 47.700 21.380 47.860 21.450 ;
        RECT 50.600 21.380 50.760 21.450 ;
        RECT 53.500 21.380 53.660 21.450 ;
        RECT 56.400 21.380 56.560 21.450 ;
        RECT 59.300 21.380 59.460 21.450 ;
        RECT 62.200 21.380 62.360 21.450 ;
        RECT 65.100 21.380 65.260 21.450 ;
        RECT 68.000 21.380 68.160 21.450 ;
        RECT 70.900 21.380 71.060 21.450 ;
        RECT 73.800 21.380 73.960 21.450 ;
        RECT 76.700 21.380 76.860 21.450 ;
        RECT 79.600 21.380 79.760 21.450 ;
        RECT 82.500 21.380 82.660 21.450 ;
        RECT 85.400 21.380 85.560 21.450 ;
        RECT 88.300 21.380 88.460 21.450 ;
        RECT 91.200 21.380 91.360 21.450 ;
        RECT 1.310 21.370 1.450 21.380 ;
        RECT 4.210 21.370 4.350 21.380 ;
        RECT 7.110 21.370 7.250 21.380 ;
        RECT 10.010 21.370 10.150 21.380 ;
        RECT 12.910 21.370 13.050 21.380 ;
        RECT 15.810 21.370 15.950 21.380 ;
        RECT 18.710 21.370 18.850 21.380 ;
        RECT 21.610 21.370 21.750 21.380 ;
        RECT 24.510 21.370 24.650 21.380 ;
        RECT 27.410 21.370 27.550 21.380 ;
        RECT 30.310 21.370 30.450 21.380 ;
        RECT 33.210 21.370 33.350 21.380 ;
        RECT 36.110 21.370 36.250 21.380 ;
        RECT 39.010 21.370 39.150 21.380 ;
        RECT 41.910 21.370 42.050 21.380 ;
        RECT 44.810 21.370 44.950 21.380 ;
        RECT 47.710 21.370 47.850 21.380 ;
        RECT 50.610 21.370 50.750 21.380 ;
        RECT 53.510 21.370 53.650 21.380 ;
        RECT 56.410 21.370 56.550 21.380 ;
        RECT 59.310 21.370 59.450 21.380 ;
        RECT 62.210 21.370 62.350 21.380 ;
        RECT 65.110 21.370 65.250 21.380 ;
        RECT 68.010 21.370 68.150 21.380 ;
        RECT 70.910 21.370 71.050 21.380 ;
        RECT 73.810 21.370 73.950 21.380 ;
        RECT 76.710 21.370 76.850 21.380 ;
        RECT 79.610 21.370 79.750 21.380 ;
        RECT 82.510 21.370 82.650 21.380 ;
        RECT 85.410 21.370 85.550 21.380 ;
        RECT 88.310 21.370 88.450 21.380 ;
        RECT 91.210 21.370 91.350 21.380 ;
      LAYER met1 ;
        RECT 0.000 21.380 92.660 21.450 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.990 19.620 1.755 20.100 ;
        RECT 3.890 19.620 4.655 20.100 ;
        RECT 6.790 19.620 7.555 20.100 ;
        RECT 9.690 19.620 10.455 20.100 ;
        RECT 12.590 19.620 13.355 20.100 ;
        RECT 15.490 19.620 16.255 20.100 ;
        RECT 18.390 19.620 19.155 20.100 ;
        RECT 21.290 19.620 22.055 20.100 ;
        RECT 24.190 19.620 24.955 20.100 ;
        RECT 27.090 19.620 27.855 20.100 ;
        RECT 29.990 19.620 30.755 20.100 ;
        RECT 32.890 19.620 33.655 20.100 ;
        RECT 35.790 19.620 36.555 20.100 ;
        RECT 38.690 19.620 39.455 20.100 ;
        RECT 41.590 19.620 42.355 20.100 ;
        RECT 44.490 19.620 45.255 20.100 ;
        RECT 47.390 19.620 48.155 20.100 ;
        RECT 50.290 19.620 51.055 20.100 ;
        RECT 53.190 19.620 53.955 20.100 ;
        RECT 56.090 19.620 56.855 20.100 ;
        RECT 58.990 19.620 59.755 20.100 ;
        RECT 61.890 19.620 62.655 20.100 ;
        RECT 64.790 19.620 65.555 20.100 ;
        RECT 67.690 19.620 68.455 20.100 ;
        RECT 70.590 19.620 71.355 20.100 ;
        RECT 73.490 19.620 74.255 20.100 ;
        RECT 76.390 19.620 77.155 20.100 ;
        RECT 79.290 19.620 80.055 20.100 ;
        RECT 82.190 19.620 82.955 20.100 ;
        RECT 85.090 19.620 85.855 20.100 ;
        RECT 87.990 19.620 88.755 20.100 ;
        RECT 90.890 19.620 91.655 20.100 ;
      LAYER li1 ;
        RECT 1.300 20.030 1.460 20.100 ;
        RECT 4.200 20.030 4.360 20.100 ;
        RECT 7.100 20.030 7.260 20.100 ;
        RECT 10.000 20.030 10.160 20.100 ;
        RECT 12.900 20.030 13.060 20.100 ;
        RECT 15.800 20.030 15.960 20.100 ;
        RECT 18.700 20.030 18.860 20.100 ;
        RECT 21.600 20.030 21.760 20.100 ;
        RECT 24.500 20.030 24.660 20.100 ;
        RECT 27.400 20.030 27.560 20.100 ;
        RECT 30.300 20.030 30.460 20.100 ;
        RECT 33.200 20.030 33.360 20.100 ;
        RECT 36.100 20.030 36.260 20.100 ;
        RECT 39.000 20.030 39.160 20.100 ;
        RECT 41.900 20.030 42.060 20.100 ;
        RECT 44.800 20.030 44.960 20.100 ;
        RECT 47.700 20.030 47.860 20.100 ;
        RECT 50.600 20.030 50.760 20.100 ;
        RECT 53.500 20.030 53.660 20.100 ;
        RECT 56.400 20.030 56.560 20.100 ;
        RECT 59.300 20.030 59.460 20.100 ;
        RECT 62.200 20.030 62.360 20.100 ;
        RECT 65.100 20.030 65.260 20.100 ;
        RECT 68.000 20.030 68.160 20.100 ;
        RECT 70.900 20.030 71.060 20.100 ;
        RECT 73.800 20.030 73.960 20.100 ;
        RECT 76.700 20.030 76.860 20.100 ;
        RECT 79.600 20.030 79.760 20.100 ;
        RECT 82.500 20.030 82.660 20.100 ;
        RECT 85.400 20.030 85.560 20.100 ;
        RECT 88.300 20.030 88.460 20.100 ;
        RECT 91.200 20.030 91.360 20.100 ;
        RECT 1.310 20.020 1.450 20.030 ;
        RECT 4.210 20.020 4.350 20.030 ;
        RECT 7.110 20.020 7.250 20.030 ;
        RECT 10.010 20.020 10.150 20.030 ;
        RECT 12.910 20.020 13.050 20.030 ;
        RECT 15.810 20.020 15.950 20.030 ;
        RECT 18.710 20.020 18.850 20.030 ;
        RECT 21.610 20.020 21.750 20.030 ;
        RECT 24.510 20.020 24.650 20.030 ;
        RECT 27.410 20.020 27.550 20.030 ;
        RECT 30.310 20.020 30.450 20.030 ;
        RECT 33.210 20.020 33.350 20.030 ;
        RECT 36.110 20.020 36.250 20.030 ;
        RECT 39.010 20.020 39.150 20.030 ;
        RECT 41.910 20.020 42.050 20.030 ;
        RECT 44.810 20.020 44.950 20.030 ;
        RECT 47.710 20.020 47.850 20.030 ;
        RECT 50.610 20.020 50.750 20.030 ;
        RECT 53.510 20.020 53.650 20.030 ;
        RECT 56.410 20.020 56.550 20.030 ;
        RECT 59.310 20.020 59.450 20.030 ;
        RECT 62.210 20.020 62.350 20.030 ;
        RECT 65.110 20.020 65.250 20.030 ;
        RECT 68.010 20.020 68.150 20.030 ;
        RECT 70.910 20.020 71.050 20.030 ;
        RECT 73.810 20.020 73.950 20.030 ;
        RECT 76.710 20.020 76.850 20.030 ;
        RECT 79.610 20.020 79.750 20.030 ;
        RECT 82.510 20.020 82.650 20.030 ;
        RECT 85.410 20.020 85.550 20.030 ;
        RECT 88.310 20.020 88.450 20.030 ;
        RECT 91.210 20.020 91.350 20.030 ;
      LAYER met1 ;
        RECT 0.000 20.030 92.660 20.100 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.990 18.270 1.755 18.750 ;
        RECT 3.890 18.270 4.655 18.750 ;
        RECT 6.790 18.270 7.555 18.750 ;
        RECT 9.690 18.270 10.455 18.750 ;
        RECT 12.590 18.270 13.355 18.750 ;
        RECT 15.490 18.270 16.255 18.750 ;
        RECT 18.390 18.270 19.155 18.750 ;
        RECT 21.290 18.270 22.055 18.750 ;
        RECT 24.190 18.270 24.955 18.750 ;
        RECT 27.090 18.270 27.855 18.750 ;
        RECT 29.990 18.270 30.755 18.750 ;
        RECT 32.890 18.270 33.655 18.750 ;
        RECT 35.790 18.270 36.555 18.750 ;
        RECT 38.690 18.270 39.455 18.750 ;
        RECT 41.590 18.270 42.355 18.750 ;
        RECT 44.490 18.270 45.255 18.750 ;
        RECT 47.390 18.270 48.155 18.750 ;
        RECT 50.290 18.270 51.055 18.750 ;
        RECT 53.190 18.270 53.955 18.750 ;
        RECT 56.090 18.270 56.855 18.750 ;
        RECT 58.990 18.270 59.755 18.750 ;
        RECT 61.890 18.270 62.655 18.750 ;
        RECT 64.790 18.270 65.555 18.750 ;
        RECT 67.690 18.270 68.455 18.750 ;
        RECT 70.590 18.270 71.355 18.750 ;
        RECT 73.490 18.270 74.255 18.750 ;
        RECT 76.390 18.270 77.155 18.750 ;
        RECT 79.290 18.270 80.055 18.750 ;
        RECT 82.190 18.270 82.955 18.750 ;
        RECT 85.090 18.270 85.855 18.750 ;
        RECT 87.990 18.270 88.755 18.750 ;
        RECT 90.890 18.270 91.655 18.750 ;
      LAYER li1 ;
        RECT 1.300 18.680 1.460 18.750 ;
        RECT 4.200 18.680 4.360 18.750 ;
        RECT 7.100 18.680 7.260 18.750 ;
        RECT 10.000 18.680 10.160 18.750 ;
        RECT 12.900 18.680 13.060 18.750 ;
        RECT 15.800 18.680 15.960 18.750 ;
        RECT 18.700 18.680 18.860 18.750 ;
        RECT 21.600 18.680 21.760 18.750 ;
        RECT 24.500 18.680 24.660 18.750 ;
        RECT 27.400 18.680 27.560 18.750 ;
        RECT 30.300 18.680 30.460 18.750 ;
        RECT 33.200 18.680 33.360 18.750 ;
        RECT 36.100 18.680 36.260 18.750 ;
        RECT 39.000 18.680 39.160 18.750 ;
        RECT 41.900 18.680 42.060 18.750 ;
        RECT 44.800 18.680 44.960 18.750 ;
        RECT 47.700 18.680 47.860 18.750 ;
        RECT 50.600 18.680 50.760 18.750 ;
        RECT 53.500 18.680 53.660 18.750 ;
        RECT 56.400 18.680 56.560 18.750 ;
        RECT 59.300 18.680 59.460 18.750 ;
        RECT 62.200 18.680 62.360 18.750 ;
        RECT 65.100 18.680 65.260 18.750 ;
        RECT 68.000 18.680 68.160 18.750 ;
        RECT 70.900 18.680 71.060 18.750 ;
        RECT 73.800 18.680 73.960 18.750 ;
        RECT 76.700 18.680 76.860 18.750 ;
        RECT 79.600 18.680 79.760 18.750 ;
        RECT 82.500 18.680 82.660 18.750 ;
        RECT 85.400 18.680 85.560 18.750 ;
        RECT 88.300 18.680 88.460 18.750 ;
        RECT 91.200 18.680 91.360 18.750 ;
        RECT 1.310 18.670 1.450 18.680 ;
        RECT 4.210 18.670 4.350 18.680 ;
        RECT 7.110 18.670 7.250 18.680 ;
        RECT 10.010 18.670 10.150 18.680 ;
        RECT 12.910 18.670 13.050 18.680 ;
        RECT 15.810 18.670 15.950 18.680 ;
        RECT 18.710 18.670 18.850 18.680 ;
        RECT 21.610 18.670 21.750 18.680 ;
        RECT 24.510 18.670 24.650 18.680 ;
        RECT 27.410 18.670 27.550 18.680 ;
        RECT 30.310 18.670 30.450 18.680 ;
        RECT 33.210 18.670 33.350 18.680 ;
        RECT 36.110 18.670 36.250 18.680 ;
        RECT 39.010 18.670 39.150 18.680 ;
        RECT 41.910 18.670 42.050 18.680 ;
        RECT 44.810 18.670 44.950 18.680 ;
        RECT 47.710 18.670 47.850 18.680 ;
        RECT 50.610 18.670 50.750 18.680 ;
        RECT 53.510 18.670 53.650 18.680 ;
        RECT 56.410 18.670 56.550 18.680 ;
        RECT 59.310 18.670 59.450 18.680 ;
        RECT 62.210 18.670 62.350 18.680 ;
        RECT 65.110 18.670 65.250 18.680 ;
        RECT 68.010 18.670 68.150 18.680 ;
        RECT 70.910 18.670 71.050 18.680 ;
        RECT 73.810 18.670 73.950 18.680 ;
        RECT 76.710 18.670 76.850 18.680 ;
        RECT 79.610 18.670 79.750 18.680 ;
        RECT 82.510 18.670 82.650 18.680 ;
        RECT 85.410 18.670 85.550 18.680 ;
        RECT 88.310 18.670 88.450 18.680 ;
        RECT 91.210 18.670 91.350 18.680 ;
      LAYER met1 ;
        RECT 0.000 18.680 92.660 18.750 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.990 16.920 1.755 17.400 ;
        RECT 3.890 16.920 4.655 17.400 ;
        RECT 6.790 16.920 7.555 17.400 ;
        RECT 9.690 16.920 10.455 17.400 ;
        RECT 12.590 16.920 13.355 17.400 ;
        RECT 15.490 16.920 16.255 17.400 ;
        RECT 18.390 16.920 19.155 17.400 ;
        RECT 21.290 16.920 22.055 17.400 ;
        RECT 24.190 16.920 24.955 17.400 ;
        RECT 27.090 16.920 27.855 17.400 ;
        RECT 29.990 16.920 30.755 17.400 ;
        RECT 32.890 16.920 33.655 17.400 ;
        RECT 35.790 16.920 36.555 17.400 ;
        RECT 38.690 16.920 39.455 17.400 ;
        RECT 41.590 16.920 42.355 17.400 ;
        RECT 44.490 16.920 45.255 17.400 ;
        RECT 47.390 16.920 48.155 17.400 ;
        RECT 50.290 16.920 51.055 17.400 ;
        RECT 53.190 16.920 53.955 17.400 ;
        RECT 56.090 16.920 56.855 17.400 ;
        RECT 58.990 16.920 59.755 17.400 ;
        RECT 61.890 16.920 62.655 17.400 ;
        RECT 64.790 16.920 65.555 17.400 ;
        RECT 67.690 16.920 68.455 17.400 ;
        RECT 70.590 16.920 71.355 17.400 ;
        RECT 73.490 16.920 74.255 17.400 ;
        RECT 76.390 16.920 77.155 17.400 ;
        RECT 79.290 16.920 80.055 17.400 ;
        RECT 82.190 16.920 82.955 17.400 ;
        RECT 85.090 16.920 85.855 17.400 ;
        RECT 87.990 16.920 88.755 17.400 ;
        RECT 90.890 16.920 91.655 17.400 ;
      LAYER li1 ;
        RECT 1.300 17.330 1.460 17.400 ;
        RECT 4.200 17.330 4.360 17.400 ;
        RECT 7.100 17.330 7.260 17.400 ;
        RECT 10.000 17.330 10.160 17.400 ;
        RECT 12.900 17.330 13.060 17.400 ;
        RECT 15.800 17.330 15.960 17.400 ;
        RECT 18.700 17.330 18.860 17.400 ;
        RECT 21.600 17.330 21.760 17.400 ;
        RECT 24.500 17.330 24.660 17.400 ;
        RECT 27.400 17.330 27.560 17.400 ;
        RECT 30.300 17.330 30.460 17.400 ;
        RECT 33.200 17.330 33.360 17.400 ;
        RECT 36.100 17.330 36.260 17.400 ;
        RECT 39.000 17.330 39.160 17.400 ;
        RECT 41.900 17.330 42.060 17.400 ;
        RECT 44.800 17.330 44.960 17.400 ;
        RECT 47.700 17.330 47.860 17.400 ;
        RECT 50.600 17.330 50.760 17.400 ;
        RECT 53.500 17.330 53.660 17.400 ;
        RECT 56.400 17.330 56.560 17.400 ;
        RECT 59.300 17.330 59.460 17.400 ;
        RECT 62.200 17.330 62.360 17.400 ;
        RECT 65.100 17.330 65.260 17.400 ;
        RECT 68.000 17.330 68.160 17.400 ;
        RECT 70.900 17.330 71.060 17.400 ;
        RECT 73.800 17.330 73.960 17.400 ;
        RECT 76.700 17.330 76.860 17.400 ;
        RECT 79.600 17.330 79.760 17.400 ;
        RECT 82.500 17.330 82.660 17.400 ;
        RECT 85.400 17.330 85.560 17.400 ;
        RECT 88.300 17.330 88.460 17.400 ;
        RECT 91.200 17.330 91.360 17.400 ;
        RECT 1.310 17.320 1.450 17.330 ;
        RECT 4.210 17.320 4.350 17.330 ;
        RECT 7.110 17.320 7.250 17.330 ;
        RECT 10.010 17.320 10.150 17.330 ;
        RECT 12.910 17.320 13.050 17.330 ;
        RECT 15.810 17.320 15.950 17.330 ;
        RECT 18.710 17.320 18.850 17.330 ;
        RECT 21.610 17.320 21.750 17.330 ;
        RECT 24.510 17.320 24.650 17.330 ;
        RECT 27.410 17.320 27.550 17.330 ;
        RECT 30.310 17.320 30.450 17.330 ;
        RECT 33.210 17.320 33.350 17.330 ;
        RECT 36.110 17.320 36.250 17.330 ;
        RECT 39.010 17.320 39.150 17.330 ;
        RECT 41.910 17.320 42.050 17.330 ;
        RECT 44.810 17.320 44.950 17.330 ;
        RECT 47.710 17.320 47.850 17.330 ;
        RECT 50.610 17.320 50.750 17.330 ;
        RECT 53.510 17.320 53.650 17.330 ;
        RECT 56.410 17.320 56.550 17.330 ;
        RECT 59.310 17.320 59.450 17.330 ;
        RECT 62.210 17.320 62.350 17.330 ;
        RECT 65.110 17.320 65.250 17.330 ;
        RECT 68.010 17.320 68.150 17.330 ;
        RECT 70.910 17.320 71.050 17.330 ;
        RECT 73.810 17.320 73.950 17.330 ;
        RECT 76.710 17.320 76.850 17.330 ;
        RECT 79.610 17.320 79.750 17.330 ;
        RECT 82.510 17.320 82.650 17.330 ;
        RECT 85.410 17.320 85.550 17.330 ;
        RECT 88.310 17.320 88.450 17.330 ;
        RECT 91.210 17.320 91.350 17.330 ;
      LAYER met1 ;
        RECT 0.000 17.330 92.660 17.400 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.990 15.570 1.755 16.050 ;
        RECT 3.890 15.570 4.655 16.050 ;
        RECT 6.790 15.570 7.555 16.050 ;
        RECT 9.690 15.570 10.455 16.050 ;
        RECT 12.590 15.570 13.355 16.050 ;
        RECT 15.490 15.570 16.255 16.050 ;
        RECT 18.390 15.570 19.155 16.050 ;
        RECT 21.290 15.570 22.055 16.050 ;
        RECT 24.190 15.570 24.955 16.050 ;
        RECT 27.090 15.570 27.855 16.050 ;
        RECT 29.990 15.570 30.755 16.050 ;
        RECT 32.890 15.570 33.655 16.050 ;
        RECT 35.790 15.570 36.555 16.050 ;
        RECT 38.690 15.570 39.455 16.050 ;
        RECT 41.590 15.570 42.355 16.050 ;
        RECT 44.490 15.570 45.255 16.050 ;
        RECT 47.390 15.570 48.155 16.050 ;
        RECT 50.290 15.570 51.055 16.050 ;
        RECT 53.190 15.570 53.955 16.050 ;
        RECT 56.090 15.570 56.855 16.050 ;
        RECT 58.990 15.570 59.755 16.050 ;
        RECT 61.890 15.570 62.655 16.050 ;
        RECT 64.790 15.570 65.555 16.050 ;
        RECT 67.690 15.570 68.455 16.050 ;
        RECT 70.590 15.570 71.355 16.050 ;
        RECT 73.490 15.570 74.255 16.050 ;
        RECT 76.390 15.570 77.155 16.050 ;
        RECT 79.290 15.570 80.055 16.050 ;
        RECT 82.190 15.570 82.955 16.050 ;
        RECT 85.090 15.570 85.855 16.050 ;
        RECT 87.990 15.570 88.755 16.050 ;
        RECT 90.890 15.570 91.655 16.050 ;
      LAYER li1 ;
        RECT 1.300 15.980 1.460 16.050 ;
        RECT 4.200 15.980 4.360 16.050 ;
        RECT 7.100 15.980 7.260 16.050 ;
        RECT 10.000 15.980 10.160 16.050 ;
        RECT 12.900 15.980 13.060 16.050 ;
        RECT 15.800 15.980 15.960 16.050 ;
        RECT 18.700 15.980 18.860 16.050 ;
        RECT 21.600 15.980 21.760 16.050 ;
        RECT 24.500 15.980 24.660 16.050 ;
        RECT 27.400 15.980 27.560 16.050 ;
        RECT 30.300 15.980 30.460 16.050 ;
        RECT 33.200 15.980 33.360 16.050 ;
        RECT 36.100 15.980 36.260 16.050 ;
        RECT 39.000 15.980 39.160 16.050 ;
        RECT 41.900 15.980 42.060 16.050 ;
        RECT 44.800 15.980 44.960 16.050 ;
        RECT 47.700 15.980 47.860 16.050 ;
        RECT 50.600 15.980 50.760 16.050 ;
        RECT 53.500 15.980 53.660 16.050 ;
        RECT 56.400 15.980 56.560 16.050 ;
        RECT 59.300 15.980 59.460 16.050 ;
        RECT 62.200 15.980 62.360 16.050 ;
        RECT 65.100 15.980 65.260 16.050 ;
        RECT 68.000 15.980 68.160 16.050 ;
        RECT 70.900 15.980 71.060 16.050 ;
        RECT 73.800 15.980 73.960 16.050 ;
        RECT 76.700 15.980 76.860 16.050 ;
        RECT 79.600 15.980 79.760 16.050 ;
        RECT 82.500 15.980 82.660 16.050 ;
        RECT 85.400 15.980 85.560 16.050 ;
        RECT 88.300 15.980 88.460 16.050 ;
        RECT 91.200 15.980 91.360 16.050 ;
        RECT 1.310 15.970 1.450 15.980 ;
        RECT 4.210 15.970 4.350 15.980 ;
        RECT 7.110 15.970 7.250 15.980 ;
        RECT 10.010 15.970 10.150 15.980 ;
        RECT 12.910 15.970 13.050 15.980 ;
        RECT 15.810 15.970 15.950 15.980 ;
        RECT 18.710 15.970 18.850 15.980 ;
        RECT 21.610 15.970 21.750 15.980 ;
        RECT 24.510 15.970 24.650 15.980 ;
        RECT 27.410 15.970 27.550 15.980 ;
        RECT 30.310 15.970 30.450 15.980 ;
        RECT 33.210 15.970 33.350 15.980 ;
        RECT 36.110 15.970 36.250 15.980 ;
        RECT 39.010 15.970 39.150 15.980 ;
        RECT 41.910 15.970 42.050 15.980 ;
        RECT 44.810 15.970 44.950 15.980 ;
        RECT 47.710 15.970 47.850 15.980 ;
        RECT 50.610 15.970 50.750 15.980 ;
        RECT 53.510 15.970 53.650 15.980 ;
        RECT 56.410 15.970 56.550 15.980 ;
        RECT 59.310 15.970 59.450 15.980 ;
        RECT 62.210 15.970 62.350 15.980 ;
        RECT 65.110 15.970 65.250 15.980 ;
        RECT 68.010 15.970 68.150 15.980 ;
        RECT 70.910 15.970 71.050 15.980 ;
        RECT 73.810 15.970 73.950 15.980 ;
        RECT 76.710 15.970 76.850 15.980 ;
        RECT 79.610 15.970 79.750 15.980 ;
        RECT 82.510 15.970 82.650 15.980 ;
        RECT 85.410 15.970 85.550 15.980 ;
        RECT 88.310 15.970 88.450 15.980 ;
        RECT 91.210 15.970 91.350 15.980 ;
      LAYER met1 ;
        RECT 0.000 15.980 92.660 16.050 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.990 14.220 1.755 14.700 ;
        RECT 3.890 14.220 4.655 14.700 ;
        RECT 6.790 14.220 7.555 14.700 ;
        RECT 9.690 14.220 10.455 14.700 ;
        RECT 12.590 14.220 13.355 14.700 ;
        RECT 15.490 14.220 16.255 14.700 ;
        RECT 18.390 14.220 19.155 14.700 ;
        RECT 21.290 14.220 22.055 14.700 ;
        RECT 24.190 14.220 24.955 14.700 ;
        RECT 27.090 14.220 27.855 14.700 ;
        RECT 29.990 14.220 30.755 14.700 ;
        RECT 32.890 14.220 33.655 14.700 ;
        RECT 35.790 14.220 36.555 14.700 ;
        RECT 38.690 14.220 39.455 14.700 ;
        RECT 41.590 14.220 42.355 14.700 ;
        RECT 44.490 14.220 45.255 14.700 ;
        RECT 47.390 14.220 48.155 14.700 ;
        RECT 50.290 14.220 51.055 14.700 ;
        RECT 53.190 14.220 53.955 14.700 ;
        RECT 56.090 14.220 56.855 14.700 ;
        RECT 58.990 14.220 59.755 14.700 ;
        RECT 61.890 14.220 62.655 14.700 ;
        RECT 64.790 14.220 65.555 14.700 ;
        RECT 67.690 14.220 68.455 14.700 ;
        RECT 70.590 14.220 71.355 14.700 ;
        RECT 73.490 14.220 74.255 14.700 ;
        RECT 76.390 14.220 77.155 14.700 ;
        RECT 79.290 14.220 80.055 14.700 ;
        RECT 82.190 14.220 82.955 14.700 ;
        RECT 85.090 14.220 85.855 14.700 ;
        RECT 87.990 14.220 88.755 14.700 ;
        RECT 90.890 14.220 91.655 14.700 ;
      LAYER li1 ;
        RECT 1.300 14.630 1.460 14.700 ;
        RECT 4.200 14.630 4.360 14.700 ;
        RECT 7.100 14.630 7.260 14.700 ;
        RECT 10.000 14.630 10.160 14.700 ;
        RECT 12.900 14.630 13.060 14.700 ;
        RECT 15.800 14.630 15.960 14.700 ;
        RECT 18.700 14.630 18.860 14.700 ;
        RECT 21.600 14.630 21.760 14.700 ;
        RECT 24.500 14.630 24.660 14.700 ;
        RECT 27.400 14.630 27.560 14.700 ;
        RECT 30.300 14.630 30.460 14.700 ;
        RECT 33.200 14.630 33.360 14.700 ;
        RECT 36.100 14.630 36.260 14.700 ;
        RECT 39.000 14.630 39.160 14.700 ;
        RECT 41.900 14.630 42.060 14.700 ;
        RECT 44.800 14.630 44.960 14.700 ;
        RECT 47.700 14.630 47.860 14.700 ;
        RECT 50.600 14.630 50.760 14.700 ;
        RECT 53.500 14.630 53.660 14.700 ;
        RECT 56.400 14.630 56.560 14.700 ;
        RECT 59.300 14.630 59.460 14.700 ;
        RECT 62.200 14.630 62.360 14.700 ;
        RECT 65.100 14.630 65.260 14.700 ;
        RECT 68.000 14.630 68.160 14.700 ;
        RECT 70.900 14.630 71.060 14.700 ;
        RECT 73.800 14.630 73.960 14.700 ;
        RECT 76.700 14.630 76.860 14.700 ;
        RECT 79.600 14.630 79.760 14.700 ;
        RECT 82.500 14.630 82.660 14.700 ;
        RECT 85.400 14.630 85.560 14.700 ;
        RECT 88.300 14.630 88.460 14.700 ;
        RECT 91.200 14.630 91.360 14.700 ;
        RECT 1.310 14.620 1.450 14.630 ;
        RECT 4.210 14.620 4.350 14.630 ;
        RECT 7.110 14.620 7.250 14.630 ;
        RECT 10.010 14.620 10.150 14.630 ;
        RECT 12.910 14.620 13.050 14.630 ;
        RECT 15.810 14.620 15.950 14.630 ;
        RECT 18.710 14.620 18.850 14.630 ;
        RECT 21.610 14.620 21.750 14.630 ;
        RECT 24.510 14.620 24.650 14.630 ;
        RECT 27.410 14.620 27.550 14.630 ;
        RECT 30.310 14.620 30.450 14.630 ;
        RECT 33.210 14.620 33.350 14.630 ;
        RECT 36.110 14.620 36.250 14.630 ;
        RECT 39.010 14.620 39.150 14.630 ;
        RECT 41.910 14.620 42.050 14.630 ;
        RECT 44.810 14.620 44.950 14.630 ;
        RECT 47.710 14.620 47.850 14.630 ;
        RECT 50.610 14.620 50.750 14.630 ;
        RECT 53.510 14.620 53.650 14.630 ;
        RECT 56.410 14.620 56.550 14.630 ;
        RECT 59.310 14.620 59.450 14.630 ;
        RECT 62.210 14.620 62.350 14.630 ;
        RECT 65.110 14.620 65.250 14.630 ;
        RECT 68.010 14.620 68.150 14.630 ;
        RECT 70.910 14.620 71.050 14.630 ;
        RECT 73.810 14.620 73.950 14.630 ;
        RECT 76.710 14.620 76.850 14.630 ;
        RECT 79.610 14.620 79.750 14.630 ;
        RECT 82.510 14.620 82.650 14.630 ;
        RECT 85.410 14.620 85.550 14.630 ;
        RECT 88.310 14.620 88.450 14.630 ;
        RECT 91.210 14.620 91.350 14.630 ;
      LAYER met1 ;
        RECT 0.000 14.630 92.660 14.700 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.990 12.870 1.755 13.350 ;
        RECT 3.890 12.870 4.655 13.350 ;
        RECT 6.790 12.870 7.555 13.350 ;
        RECT 9.690 12.870 10.455 13.350 ;
        RECT 12.590 12.870 13.355 13.350 ;
        RECT 15.490 12.870 16.255 13.350 ;
        RECT 18.390 12.870 19.155 13.350 ;
        RECT 21.290 12.870 22.055 13.350 ;
        RECT 24.190 12.870 24.955 13.350 ;
        RECT 27.090 12.870 27.855 13.350 ;
        RECT 29.990 12.870 30.755 13.350 ;
        RECT 32.890 12.870 33.655 13.350 ;
        RECT 35.790 12.870 36.555 13.350 ;
        RECT 38.690 12.870 39.455 13.350 ;
        RECT 41.590 12.870 42.355 13.350 ;
        RECT 44.490 12.870 45.255 13.350 ;
        RECT 47.390 12.870 48.155 13.350 ;
        RECT 50.290 12.870 51.055 13.350 ;
        RECT 53.190 12.870 53.955 13.350 ;
        RECT 56.090 12.870 56.855 13.350 ;
        RECT 58.990 12.870 59.755 13.350 ;
        RECT 61.890 12.870 62.655 13.350 ;
        RECT 64.790 12.870 65.555 13.350 ;
        RECT 67.690 12.870 68.455 13.350 ;
        RECT 70.590 12.870 71.355 13.350 ;
        RECT 73.490 12.870 74.255 13.350 ;
        RECT 76.390 12.870 77.155 13.350 ;
        RECT 79.290 12.870 80.055 13.350 ;
        RECT 82.190 12.870 82.955 13.350 ;
        RECT 85.090 12.870 85.855 13.350 ;
        RECT 87.990 12.870 88.755 13.350 ;
        RECT 90.890 12.870 91.655 13.350 ;
      LAYER li1 ;
        RECT 1.300 13.280 1.460 13.350 ;
        RECT 4.200 13.280 4.360 13.350 ;
        RECT 7.100 13.280 7.260 13.350 ;
        RECT 10.000 13.280 10.160 13.350 ;
        RECT 12.900 13.280 13.060 13.350 ;
        RECT 15.800 13.280 15.960 13.350 ;
        RECT 18.700 13.280 18.860 13.350 ;
        RECT 21.600 13.280 21.760 13.350 ;
        RECT 24.500 13.280 24.660 13.350 ;
        RECT 27.400 13.280 27.560 13.350 ;
        RECT 30.300 13.280 30.460 13.350 ;
        RECT 33.200 13.280 33.360 13.350 ;
        RECT 36.100 13.280 36.260 13.350 ;
        RECT 39.000 13.280 39.160 13.350 ;
        RECT 41.900 13.280 42.060 13.350 ;
        RECT 44.800 13.280 44.960 13.350 ;
        RECT 47.700 13.280 47.860 13.350 ;
        RECT 50.600 13.280 50.760 13.350 ;
        RECT 53.500 13.280 53.660 13.350 ;
        RECT 56.400 13.280 56.560 13.350 ;
        RECT 59.300 13.280 59.460 13.350 ;
        RECT 62.200 13.280 62.360 13.350 ;
        RECT 65.100 13.280 65.260 13.350 ;
        RECT 68.000 13.280 68.160 13.350 ;
        RECT 70.900 13.280 71.060 13.350 ;
        RECT 73.800 13.280 73.960 13.350 ;
        RECT 76.700 13.280 76.860 13.350 ;
        RECT 79.600 13.280 79.760 13.350 ;
        RECT 82.500 13.280 82.660 13.350 ;
        RECT 85.400 13.280 85.560 13.350 ;
        RECT 88.300 13.280 88.460 13.350 ;
        RECT 91.200 13.280 91.360 13.350 ;
        RECT 1.310 13.270 1.450 13.280 ;
        RECT 4.210 13.270 4.350 13.280 ;
        RECT 7.110 13.270 7.250 13.280 ;
        RECT 10.010 13.270 10.150 13.280 ;
        RECT 12.910 13.270 13.050 13.280 ;
        RECT 15.810 13.270 15.950 13.280 ;
        RECT 18.710 13.270 18.850 13.280 ;
        RECT 21.610 13.270 21.750 13.280 ;
        RECT 24.510 13.270 24.650 13.280 ;
        RECT 27.410 13.270 27.550 13.280 ;
        RECT 30.310 13.270 30.450 13.280 ;
        RECT 33.210 13.270 33.350 13.280 ;
        RECT 36.110 13.270 36.250 13.280 ;
        RECT 39.010 13.270 39.150 13.280 ;
        RECT 41.910 13.270 42.050 13.280 ;
        RECT 44.810 13.270 44.950 13.280 ;
        RECT 47.710 13.270 47.850 13.280 ;
        RECT 50.610 13.270 50.750 13.280 ;
        RECT 53.510 13.270 53.650 13.280 ;
        RECT 56.410 13.270 56.550 13.280 ;
        RECT 59.310 13.270 59.450 13.280 ;
        RECT 62.210 13.270 62.350 13.280 ;
        RECT 65.110 13.270 65.250 13.280 ;
        RECT 68.010 13.270 68.150 13.280 ;
        RECT 70.910 13.270 71.050 13.280 ;
        RECT 73.810 13.270 73.950 13.280 ;
        RECT 76.710 13.270 76.850 13.280 ;
        RECT 79.610 13.270 79.750 13.280 ;
        RECT 82.510 13.270 82.650 13.280 ;
        RECT 85.410 13.270 85.550 13.280 ;
        RECT 88.310 13.270 88.450 13.280 ;
        RECT 91.210 13.270 91.350 13.280 ;
      LAYER met1 ;
        RECT 0.000 13.280 92.660 13.350 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.990 11.520 1.755 12.000 ;
        RECT 3.890 11.520 4.655 12.000 ;
        RECT 6.790 11.520 7.555 12.000 ;
        RECT 9.690 11.520 10.455 12.000 ;
        RECT 12.590 11.520 13.355 12.000 ;
        RECT 15.490 11.520 16.255 12.000 ;
        RECT 18.390 11.520 19.155 12.000 ;
        RECT 21.290 11.520 22.055 12.000 ;
        RECT 24.190 11.520 24.955 12.000 ;
        RECT 27.090 11.520 27.855 12.000 ;
        RECT 29.990 11.520 30.755 12.000 ;
        RECT 32.890 11.520 33.655 12.000 ;
        RECT 35.790 11.520 36.555 12.000 ;
        RECT 38.690 11.520 39.455 12.000 ;
        RECT 41.590 11.520 42.355 12.000 ;
        RECT 44.490 11.520 45.255 12.000 ;
        RECT 47.390 11.520 48.155 12.000 ;
        RECT 50.290 11.520 51.055 12.000 ;
        RECT 53.190 11.520 53.955 12.000 ;
        RECT 56.090 11.520 56.855 12.000 ;
        RECT 58.990 11.520 59.755 12.000 ;
        RECT 61.890 11.520 62.655 12.000 ;
        RECT 64.790 11.520 65.555 12.000 ;
        RECT 67.690 11.520 68.455 12.000 ;
        RECT 70.590 11.520 71.355 12.000 ;
        RECT 73.490 11.520 74.255 12.000 ;
        RECT 76.390 11.520 77.155 12.000 ;
        RECT 79.290 11.520 80.055 12.000 ;
        RECT 82.190 11.520 82.955 12.000 ;
        RECT 85.090 11.520 85.855 12.000 ;
        RECT 87.990 11.520 88.755 12.000 ;
        RECT 90.890 11.520 91.655 12.000 ;
      LAYER li1 ;
        RECT 1.300 11.930 1.460 12.000 ;
        RECT 4.200 11.930 4.360 12.000 ;
        RECT 7.100 11.930 7.260 12.000 ;
        RECT 10.000 11.930 10.160 12.000 ;
        RECT 12.900 11.930 13.060 12.000 ;
        RECT 15.800 11.930 15.960 12.000 ;
        RECT 18.700 11.930 18.860 12.000 ;
        RECT 21.600 11.930 21.760 12.000 ;
        RECT 24.500 11.930 24.660 12.000 ;
        RECT 27.400 11.930 27.560 12.000 ;
        RECT 30.300 11.930 30.460 12.000 ;
        RECT 33.200 11.930 33.360 12.000 ;
        RECT 36.100 11.930 36.260 12.000 ;
        RECT 39.000 11.930 39.160 12.000 ;
        RECT 41.900 11.930 42.060 12.000 ;
        RECT 44.800 11.930 44.960 12.000 ;
        RECT 47.700 11.930 47.860 12.000 ;
        RECT 50.600 11.930 50.760 12.000 ;
        RECT 53.500 11.930 53.660 12.000 ;
        RECT 56.400 11.930 56.560 12.000 ;
        RECT 59.300 11.930 59.460 12.000 ;
        RECT 62.200 11.930 62.360 12.000 ;
        RECT 65.100 11.930 65.260 12.000 ;
        RECT 68.000 11.930 68.160 12.000 ;
        RECT 70.900 11.930 71.060 12.000 ;
        RECT 73.800 11.930 73.960 12.000 ;
        RECT 76.700 11.930 76.860 12.000 ;
        RECT 79.600 11.930 79.760 12.000 ;
        RECT 82.500 11.930 82.660 12.000 ;
        RECT 85.400 11.930 85.560 12.000 ;
        RECT 88.300 11.930 88.460 12.000 ;
        RECT 91.200 11.930 91.360 12.000 ;
        RECT 1.310 11.920 1.450 11.930 ;
        RECT 4.210 11.920 4.350 11.930 ;
        RECT 7.110 11.920 7.250 11.930 ;
        RECT 10.010 11.920 10.150 11.930 ;
        RECT 12.910 11.920 13.050 11.930 ;
        RECT 15.810 11.920 15.950 11.930 ;
        RECT 18.710 11.920 18.850 11.930 ;
        RECT 21.610 11.920 21.750 11.930 ;
        RECT 24.510 11.920 24.650 11.930 ;
        RECT 27.410 11.920 27.550 11.930 ;
        RECT 30.310 11.920 30.450 11.930 ;
        RECT 33.210 11.920 33.350 11.930 ;
        RECT 36.110 11.920 36.250 11.930 ;
        RECT 39.010 11.920 39.150 11.930 ;
        RECT 41.910 11.920 42.050 11.930 ;
        RECT 44.810 11.920 44.950 11.930 ;
        RECT 47.710 11.920 47.850 11.930 ;
        RECT 50.610 11.920 50.750 11.930 ;
        RECT 53.510 11.920 53.650 11.930 ;
        RECT 56.410 11.920 56.550 11.930 ;
        RECT 59.310 11.920 59.450 11.930 ;
        RECT 62.210 11.920 62.350 11.930 ;
        RECT 65.110 11.920 65.250 11.930 ;
        RECT 68.010 11.920 68.150 11.930 ;
        RECT 70.910 11.920 71.050 11.930 ;
        RECT 73.810 11.920 73.950 11.930 ;
        RECT 76.710 11.920 76.850 11.930 ;
        RECT 79.610 11.920 79.750 11.930 ;
        RECT 82.510 11.920 82.650 11.930 ;
        RECT 85.410 11.920 85.550 11.930 ;
        RECT 88.310 11.920 88.450 11.930 ;
        RECT 91.210 11.920 91.350 11.930 ;
      LAYER met1 ;
        RECT 0.000 11.930 92.660 12.000 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.990 10.170 1.755 10.650 ;
        RECT 3.890 10.170 4.655 10.650 ;
        RECT 6.790 10.170 7.555 10.650 ;
        RECT 9.690 10.170 10.455 10.650 ;
        RECT 12.590 10.170 13.355 10.650 ;
        RECT 15.490 10.170 16.255 10.650 ;
        RECT 18.390 10.170 19.155 10.650 ;
        RECT 21.290 10.170 22.055 10.650 ;
        RECT 24.190 10.170 24.955 10.650 ;
        RECT 27.090 10.170 27.855 10.650 ;
        RECT 29.990 10.170 30.755 10.650 ;
        RECT 32.890 10.170 33.655 10.650 ;
        RECT 35.790 10.170 36.555 10.650 ;
        RECT 38.690 10.170 39.455 10.650 ;
        RECT 41.590 10.170 42.355 10.650 ;
        RECT 44.490 10.170 45.255 10.650 ;
        RECT 47.390 10.170 48.155 10.650 ;
        RECT 50.290 10.170 51.055 10.650 ;
        RECT 53.190 10.170 53.955 10.650 ;
        RECT 56.090 10.170 56.855 10.650 ;
        RECT 58.990 10.170 59.755 10.650 ;
        RECT 61.890 10.170 62.655 10.650 ;
        RECT 64.790 10.170 65.555 10.650 ;
        RECT 67.690 10.170 68.455 10.650 ;
        RECT 70.590 10.170 71.355 10.650 ;
        RECT 73.490 10.170 74.255 10.650 ;
        RECT 76.390 10.170 77.155 10.650 ;
        RECT 79.290 10.170 80.055 10.650 ;
        RECT 82.190 10.170 82.955 10.650 ;
        RECT 85.090 10.170 85.855 10.650 ;
        RECT 87.990 10.170 88.755 10.650 ;
        RECT 90.890 10.170 91.655 10.650 ;
      LAYER li1 ;
        RECT 1.300 10.580 1.460 10.650 ;
        RECT 4.200 10.580 4.360 10.650 ;
        RECT 7.100 10.580 7.260 10.650 ;
        RECT 10.000 10.580 10.160 10.650 ;
        RECT 12.900 10.580 13.060 10.650 ;
        RECT 15.800 10.580 15.960 10.650 ;
        RECT 18.700 10.580 18.860 10.650 ;
        RECT 21.600 10.580 21.760 10.650 ;
        RECT 24.500 10.580 24.660 10.650 ;
        RECT 27.400 10.580 27.560 10.650 ;
        RECT 30.300 10.580 30.460 10.650 ;
        RECT 33.200 10.580 33.360 10.650 ;
        RECT 36.100 10.580 36.260 10.650 ;
        RECT 39.000 10.580 39.160 10.650 ;
        RECT 41.900 10.580 42.060 10.650 ;
        RECT 44.800 10.580 44.960 10.650 ;
        RECT 47.700 10.580 47.860 10.650 ;
        RECT 50.600 10.580 50.760 10.650 ;
        RECT 53.500 10.580 53.660 10.650 ;
        RECT 56.400 10.580 56.560 10.650 ;
        RECT 59.300 10.580 59.460 10.650 ;
        RECT 62.200 10.580 62.360 10.650 ;
        RECT 65.100 10.580 65.260 10.650 ;
        RECT 68.000 10.580 68.160 10.650 ;
        RECT 70.900 10.580 71.060 10.650 ;
        RECT 73.800 10.580 73.960 10.650 ;
        RECT 76.700 10.580 76.860 10.650 ;
        RECT 79.600 10.580 79.760 10.650 ;
        RECT 82.500 10.580 82.660 10.650 ;
        RECT 85.400 10.580 85.560 10.650 ;
        RECT 88.300 10.580 88.460 10.650 ;
        RECT 91.200 10.580 91.360 10.650 ;
        RECT 1.310 10.570 1.450 10.580 ;
        RECT 4.210 10.570 4.350 10.580 ;
        RECT 7.110 10.570 7.250 10.580 ;
        RECT 10.010 10.570 10.150 10.580 ;
        RECT 12.910 10.570 13.050 10.580 ;
        RECT 15.810 10.570 15.950 10.580 ;
        RECT 18.710 10.570 18.850 10.580 ;
        RECT 21.610 10.570 21.750 10.580 ;
        RECT 24.510 10.570 24.650 10.580 ;
        RECT 27.410 10.570 27.550 10.580 ;
        RECT 30.310 10.570 30.450 10.580 ;
        RECT 33.210 10.570 33.350 10.580 ;
        RECT 36.110 10.570 36.250 10.580 ;
        RECT 39.010 10.570 39.150 10.580 ;
        RECT 41.910 10.570 42.050 10.580 ;
        RECT 44.810 10.570 44.950 10.580 ;
        RECT 47.710 10.570 47.850 10.580 ;
        RECT 50.610 10.570 50.750 10.580 ;
        RECT 53.510 10.570 53.650 10.580 ;
        RECT 56.410 10.570 56.550 10.580 ;
        RECT 59.310 10.570 59.450 10.580 ;
        RECT 62.210 10.570 62.350 10.580 ;
        RECT 65.110 10.570 65.250 10.580 ;
        RECT 68.010 10.570 68.150 10.580 ;
        RECT 70.910 10.570 71.050 10.580 ;
        RECT 73.810 10.570 73.950 10.580 ;
        RECT 76.710 10.570 76.850 10.580 ;
        RECT 79.610 10.570 79.750 10.580 ;
        RECT 82.510 10.570 82.650 10.580 ;
        RECT 85.410 10.570 85.550 10.580 ;
        RECT 88.310 10.570 88.450 10.580 ;
        RECT 91.210 10.570 91.350 10.580 ;
      LAYER met1 ;
        RECT 0.000 10.580 92.660 10.650 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.990 8.820 1.755 9.300 ;
        RECT 3.890 8.820 4.655 9.300 ;
        RECT 6.790 8.820 7.555 9.300 ;
        RECT 9.690 8.820 10.455 9.300 ;
        RECT 12.590 8.820 13.355 9.300 ;
        RECT 15.490 8.820 16.255 9.300 ;
        RECT 18.390 8.820 19.155 9.300 ;
        RECT 21.290 8.820 22.055 9.300 ;
        RECT 24.190 8.820 24.955 9.300 ;
        RECT 27.090 8.820 27.855 9.300 ;
        RECT 29.990 8.820 30.755 9.300 ;
        RECT 32.890 8.820 33.655 9.300 ;
        RECT 35.790 8.820 36.555 9.300 ;
        RECT 38.690 8.820 39.455 9.300 ;
        RECT 41.590 8.820 42.355 9.300 ;
        RECT 44.490 8.820 45.255 9.300 ;
        RECT 47.390 8.820 48.155 9.300 ;
        RECT 50.290 8.820 51.055 9.300 ;
        RECT 53.190 8.820 53.955 9.300 ;
        RECT 56.090 8.820 56.855 9.300 ;
        RECT 58.990 8.820 59.755 9.300 ;
        RECT 61.890 8.820 62.655 9.300 ;
        RECT 64.790 8.820 65.555 9.300 ;
        RECT 67.690 8.820 68.455 9.300 ;
        RECT 70.590 8.820 71.355 9.300 ;
        RECT 73.490 8.820 74.255 9.300 ;
        RECT 76.390 8.820 77.155 9.300 ;
        RECT 79.290 8.820 80.055 9.300 ;
        RECT 82.190 8.820 82.955 9.300 ;
        RECT 85.090 8.820 85.855 9.300 ;
        RECT 87.990 8.820 88.755 9.300 ;
        RECT 90.890 8.820 91.655 9.300 ;
      LAYER li1 ;
        RECT 1.300 9.230 1.460 9.300 ;
        RECT 4.200 9.230 4.360 9.300 ;
        RECT 7.100 9.230 7.260 9.300 ;
        RECT 10.000 9.230 10.160 9.300 ;
        RECT 12.900 9.230 13.060 9.300 ;
        RECT 15.800 9.230 15.960 9.300 ;
        RECT 18.700 9.230 18.860 9.300 ;
        RECT 21.600 9.230 21.760 9.300 ;
        RECT 24.500 9.230 24.660 9.300 ;
        RECT 27.400 9.230 27.560 9.300 ;
        RECT 30.300 9.230 30.460 9.300 ;
        RECT 33.200 9.230 33.360 9.300 ;
        RECT 36.100 9.230 36.260 9.300 ;
        RECT 39.000 9.230 39.160 9.300 ;
        RECT 41.900 9.230 42.060 9.300 ;
        RECT 44.800 9.230 44.960 9.300 ;
        RECT 47.700 9.230 47.860 9.300 ;
        RECT 50.600 9.230 50.760 9.300 ;
        RECT 53.500 9.230 53.660 9.300 ;
        RECT 56.400 9.230 56.560 9.300 ;
        RECT 59.300 9.230 59.460 9.300 ;
        RECT 62.200 9.230 62.360 9.300 ;
        RECT 65.100 9.230 65.260 9.300 ;
        RECT 68.000 9.230 68.160 9.300 ;
        RECT 70.900 9.230 71.060 9.300 ;
        RECT 73.800 9.230 73.960 9.300 ;
        RECT 76.700 9.230 76.860 9.300 ;
        RECT 79.600 9.230 79.760 9.300 ;
        RECT 82.500 9.230 82.660 9.300 ;
        RECT 85.400 9.230 85.560 9.300 ;
        RECT 88.300 9.230 88.460 9.300 ;
        RECT 91.200 9.230 91.360 9.300 ;
        RECT 1.310 9.220 1.450 9.230 ;
        RECT 4.210 9.220 4.350 9.230 ;
        RECT 7.110 9.220 7.250 9.230 ;
        RECT 10.010 9.220 10.150 9.230 ;
        RECT 12.910 9.220 13.050 9.230 ;
        RECT 15.810 9.220 15.950 9.230 ;
        RECT 18.710 9.220 18.850 9.230 ;
        RECT 21.610 9.220 21.750 9.230 ;
        RECT 24.510 9.220 24.650 9.230 ;
        RECT 27.410 9.220 27.550 9.230 ;
        RECT 30.310 9.220 30.450 9.230 ;
        RECT 33.210 9.220 33.350 9.230 ;
        RECT 36.110 9.220 36.250 9.230 ;
        RECT 39.010 9.220 39.150 9.230 ;
        RECT 41.910 9.220 42.050 9.230 ;
        RECT 44.810 9.220 44.950 9.230 ;
        RECT 47.710 9.220 47.850 9.230 ;
        RECT 50.610 9.220 50.750 9.230 ;
        RECT 53.510 9.220 53.650 9.230 ;
        RECT 56.410 9.220 56.550 9.230 ;
        RECT 59.310 9.220 59.450 9.230 ;
        RECT 62.210 9.220 62.350 9.230 ;
        RECT 65.110 9.220 65.250 9.230 ;
        RECT 68.010 9.220 68.150 9.230 ;
        RECT 70.910 9.220 71.050 9.230 ;
        RECT 73.810 9.220 73.950 9.230 ;
        RECT 76.710 9.220 76.850 9.230 ;
        RECT 79.610 9.220 79.750 9.230 ;
        RECT 82.510 9.220 82.650 9.230 ;
        RECT 85.410 9.220 85.550 9.230 ;
        RECT 88.310 9.220 88.450 9.230 ;
        RECT 91.210 9.220 91.350 9.230 ;
      LAYER met1 ;
        RECT 0.000 9.230 92.660 9.300 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.990 7.470 1.755 7.950 ;
        RECT 3.890 7.470 4.655 7.950 ;
        RECT 6.790 7.470 7.555 7.950 ;
        RECT 9.690 7.470 10.455 7.950 ;
        RECT 12.590 7.470 13.355 7.950 ;
        RECT 15.490 7.470 16.255 7.950 ;
        RECT 18.390 7.470 19.155 7.950 ;
        RECT 21.290 7.470 22.055 7.950 ;
        RECT 24.190 7.470 24.955 7.950 ;
        RECT 27.090 7.470 27.855 7.950 ;
        RECT 29.990 7.470 30.755 7.950 ;
        RECT 32.890 7.470 33.655 7.950 ;
        RECT 35.790 7.470 36.555 7.950 ;
        RECT 38.690 7.470 39.455 7.950 ;
        RECT 41.590 7.470 42.355 7.950 ;
        RECT 44.490 7.470 45.255 7.950 ;
        RECT 47.390 7.470 48.155 7.950 ;
        RECT 50.290 7.470 51.055 7.950 ;
        RECT 53.190 7.470 53.955 7.950 ;
        RECT 56.090 7.470 56.855 7.950 ;
        RECT 58.990 7.470 59.755 7.950 ;
        RECT 61.890 7.470 62.655 7.950 ;
        RECT 64.790 7.470 65.555 7.950 ;
        RECT 67.690 7.470 68.455 7.950 ;
        RECT 70.590 7.470 71.355 7.950 ;
        RECT 73.490 7.470 74.255 7.950 ;
        RECT 76.390 7.470 77.155 7.950 ;
        RECT 79.290 7.470 80.055 7.950 ;
        RECT 82.190 7.470 82.955 7.950 ;
        RECT 85.090 7.470 85.855 7.950 ;
        RECT 87.990 7.470 88.755 7.950 ;
        RECT 90.890 7.470 91.655 7.950 ;
      LAYER li1 ;
        RECT 1.300 7.880 1.460 7.950 ;
        RECT 4.200 7.880 4.360 7.950 ;
        RECT 7.100 7.880 7.260 7.950 ;
        RECT 10.000 7.880 10.160 7.950 ;
        RECT 12.900 7.880 13.060 7.950 ;
        RECT 15.800 7.880 15.960 7.950 ;
        RECT 18.700 7.880 18.860 7.950 ;
        RECT 21.600 7.880 21.760 7.950 ;
        RECT 24.500 7.880 24.660 7.950 ;
        RECT 27.400 7.880 27.560 7.950 ;
        RECT 30.300 7.880 30.460 7.950 ;
        RECT 33.200 7.880 33.360 7.950 ;
        RECT 36.100 7.880 36.260 7.950 ;
        RECT 39.000 7.880 39.160 7.950 ;
        RECT 41.900 7.880 42.060 7.950 ;
        RECT 44.800 7.880 44.960 7.950 ;
        RECT 47.700 7.880 47.860 7.950 ;
        RECT 50.600 7.880 50.760 7.950 ;
        RECT 53.500 7.880 53.660 7.950 ;
        RECT 56.400 7.880 56.560 7.950 ;
        RECT 59.300 7.880 59.460 7.950 ;
        RECT 62.200 7.880 62.360 7.950 ;
        RECT 65.100 7.880 65.260 7.950 ;
        RECT 68.000 7.880 68.160 7.950 ;
        RECT 70.900 7.880 71.060 7.950 ;
        RECT 73.800 7.880 73.960 7.950 ;
        RECT 76.700 7.880 76.860 7.950 ;
        RECT 79.600 7.880 79.760 7.950 ;
        RECT 82.500 7.880 82.660 7.950 ;
        RECT 85.400 7.880 85.560 7.950 ;
        RECT 88.300 7.880 88.460 7.950 ;
        RECT 91.200 7.880 91.360 7.950 ;
        RECT 1.310 7.870 1.450 7.880 ;
        RECT 4.210 7.870 4.350 7.880 ;
        RECT 7.110 7.870 7.250 7.880 ;
        RECT 10.010 7.870 10.150 7.880 ;
        RECT 12.910 7.870 13.050 7.880 ;
        RECT 15.810 7.870 15.950 7.880 ;
        RECT 18.710 7.870 18.850 7.880 ;
        RECT 21.610 7.870 21.750 7.880 ;
        RECT 24.510 7.870 24.650 7.880 ;
        RECT 27.410 7.870 27.550 7.880 ;
        RECT 30.310 7.870 30.450 7.880 ;
        RECT 33.210 7.870 33.350 7.880 ;
        RECT 36.110 7.870 36.250 7.880 ;
        RECT 39.010 7.870 39.150 7.880 ;
        RECT 41.910 7.870 42.050 7.880 ;
        RECT 44.810 7.870 44.950 7.880 ;
        RECT 47.710 7.870 47.850 7.880 ;
        RECT 50.610 7.870 50.750 7.880 ;
        RECT 53.510 7.870 53.650 7.880 ;
        RECT 56.410 7.870 56.550 7.880 ;
        RECT 59.310 7.870 59.450 7.880 ;
        RECT 62.210 7.870 62.350 7.880 ;
        RECT 65.110 7.870 65.250 7.880 ;
        RECT 68.010 7.870 68.150 7.880 ;
        RECT 70.910 7.870 71.050 7.880 ;
        RECT 73.810 7.870 73.950 7.880 ;
        RECT 76.710 7.870 76.850 7.880 ;
        RECT 79.610 7.870 79.750 7.880 ;
        RECT 82.510 7.870 82.650 7.880 ;
        RECT 85.410 7.870 85.550 7.880 ;
        RECT 88.310 7.870 88.450 7.880 ;
        RECT 91.210 7.870 91.350 7.880 ;
      LAYER met1 ;
        RECT 0.000 7.880 92.660 7.950 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.990 6.120 1.755 6.600 ;
        RECT 3.890 6.120 4.655 6.600 ;
        RECT 6.790 6.120 7.555 6.600 ;
        RECT 9.690 6.120 10.455 6.600 ;
        RECT 12.590 6.120 13.355 6.600 ;
        RECT 15.490 6.120 16.255 6.600 ;
        RECT 18.390 6.120 19.155 6.600 ;
        RECT 21.290 6.120 22.055 6.600 ;
        RECT 24.190 6.120 24.955 6.600 ;
        RECT 27.090 6.120 27.855 6.600 ;
        RECT 29.990 6.120 30.755 6.600 ;
        RECT 32.890 6.120 33.655 6.600 ;
        RECT 35.790 6.120 36.555 6.600 ;
        RECT 38.690 6.120 39.455 6.600 ;
        RECT 41.590 6.120 42.355 6.600 ;
        RECT 44.490 6.120 45.255 6.600 ;
        RECT 47.390 6.120 48.155 6.600 ;
        RECT 50.290 6.120 51.055 6.600 ;
        RECT 53.190 6.120 53.955 6.600 ;
        RECT 56.090 6.120 56.855 6.600 ;
        RECT 58.990 6.120 59.755 6.600 ;
        RECT 61.890 6.120 62.655 6.600 ;
        RECT 64.790 6.120 65.555 6.600 ;
        RECT 67.690 6.120 68.455 6.600 ;
        RECT 70.590 6.120 71.355 6.600 ;
        RECT 73.490 6.120 74.255 6.600 ;
        RECT 76.390 6.120 77.155 6.600 ;
        RECT 79.290 6.120 80.055 6.600 ;
        RECT 82.190 6.120 82.955 6.600 ;
        RECT 85.090 6.120 85.855 6.600 ;
        RECT 87.990 6.120 88.755 6.600 ;
        RECT 90.890 6.120 91.655 6.600 ;
      LAYER li1 ;
        RECT 1.300 6.530 1.460 6.600 ;
        RECT 4.200 6.530 4.360 6.600 ;
        RECT 7.100 6.530 7.260 6.600 ;
        RECT 10.000 6.530 10.160 6.600 ;
        RECT 12.900 6.530 13.060 6.600 ;
        RECT 15.800 6.530 15.960 6.600 ;
        RECT 18.700 6.530 18.860 6.600 ;
        RECT 21.600 6.530 21.760 6.600 ;
        RECT 24.500 6.530 24.660 6.600 ;
        RECT 27.400 6.530 27.560 6.600 ;
        RECT 30.300 6.530 30.460 6.600 ;
        RECT 33.200 6.530 33.360 6.600 ;
        RECT 36.100 6.530 36.260 6.600 ;
        RECT 39.000 6.530 39.160 6.600 ;
        RECT 41.900 6.530 42.060 6.600 ;
        RECT 44.800 6.530 44.960 6.600 ;
        RECT 47.700 6.530 47.860 6.600 ;
        RECT 50.600 6.530 50.760 6.600 ;
        RECT 53.500 6.530 53.660 6.600 ;
        RECT 56.400 6.530 56.560 6.600 ;
        RECT 59.300 6.530 59.460 6.600 ;
        RECT 62.200 6.530 62.360 6.600 ;
        RECT 65.100 6.530 65.260 6.600 ;
        RECT 68.000 6.530 68.160 6.600 ;
        RECT 70.900 6.530 71.060 6.600 ;
        RECT 73.800 6.530 73.960 6.600 ;
        RECT 76.700 6.530 76.860 6.600 ;
        RECT 79.600 6.530 79.760 6.600 ;
        RECT 82.500 6.530 82.660 6.600 ;
        RECT 85.400 6.530 85.560 6.600 ;
        RECT 88.300 6.530 88.460 6.600 ;
        RECT 91.200 6.530 91.360 6.600 ;
        RECT 1.310 6.520 1.450 6.530 ;
        RECT 4.210 6.520 4.350 6.530 ;
        RECT 7.110 6.520 7.250 6.530 ;
        RECT 10.010 6.520 10.150 6.530 ;
        RECT 12.910 6.520 13.050 6.530 ;
        RECT 15.810 6.520 15.950 6.530 ;
        RECT 18.710 6.520 18.850 6.530 ;
        RECT 21.610 6.520 21.750 6.530 ;
        RECT 24.510 6.520 24.650 6.530 ;
        RECT 27.410 6.520 27.550 6.530 ;
        RECT 30.310 6.520 30.450 6.530 ;
        RECT 33.210 6.520 33.350 6.530 ;
        RECT 36.110 6.520 36.250 6.530 ;
        RECT 39.010 6.520 39.150 6.530 ;
        RECT 41.910 6.520 42.050 6.530 ;
        RECT 44.810 6.520 44.950 6.530 ;
        RECT 47.710 6.520 47.850 6.530 ;
        RECT 50.610 6.520 50.750 6.530 ;
        RECT 53.510 6.520 53.650 6.530 ;
        RECT 56.410 6.520 56.550 6.530 ;
        RECT 59.310 6.520 59.450 6.530 ;
        RECT 62.210 6.520 62.350 6.530 ;
        RECT 65.110 6.520 65.250 6.530 ;
        RECT 68.010 6.520 68.150 6.530 ;
        RECT 70.910 6.520 71.050 6.530 ;
        RECT 73.810 6.520 73.950 6.530 ;
        RECT 76.710 6.520 76.850 6.530 ;
        RECT 79.610 6.520 79.750 6.530 ;
        RECT 82.510 6.520 82.650 6.530 ;
        RECT 85.410 6.520 85.550 6.530 ;
        RECT 88.310 6.520 88.450 6.530 ;
        RECT 91.210 6.520 91.350 6.530 ;
      LAYER met1 ;
        RECT 0.000 6.530 92.660 6.600 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.990 4.770 1.755 5.250 ;
        RECT 3.890 4.770 4.655 5.250 ;
        RECT 6.790 4.770 7.555 5.250 ;
        RECT 9.690 4.770 10.455 5.250 ;
        RECT 12.590 4.770 13.355 5.250 ;
        RECT 15.490 4.770 16.255 5.250 ;
        RECT 18.390 4.770 19.155 5.250 ;
        RECT 21.290 4.770 22.055 5.250 ;
        RECT 24.190 4.770 24.955 5.250 ;
        RECT 27.090 4.770 27.855 5.250 ;
        RECT 29.990 4.770 30.755 5.250 ;
        RECT 32.890 4.770 33.655 5.250 ;
        RECT 35.790 4.770 36.555 5.250 ;
        RECT 38.690 4.770 39.455 5.250 ;
        RECT 41.590 4.770 42.355 5.250 ;
        RECT 44.490 4.770 45.255 5.250 ;
        RECT 47.390 4.770 48.155 5.250 ;
        RECT 50.290 4.770 51.055 5.250 ;
        RECT 53.190 4.770 53.955 5.250 ;
        RECT 56.090 4.770 56.855 5.250 ;
        RECT 58.990 4.770 59.755 5.250 ;
        RECT 61.890 4.770 62.655 5.250 ;
        RECT 64.790 4.770 65.555 5.250 ;
        RECT 67.690 4.770 68.455 5.250 ;
        RECT 70.590 4.770 71.355 5.250 ;
        RECT 73.490 4.770 74.255 5.250 ;
        RECT 76.390 4.770 77.155 5.250 ;
        RECT 79.290 4.770 80.055 5.250 ;
        RECT 82.190 4.770 82.955 5.250 ;
        RECT 85.090 4.770 85.855 5.250 ;
        RECT 87.990 4.770 88.755 5.250 ;
        RECT 90.890 4.770 91.655 5.250 ;
      LAYER li1 ;
        RECT 1.300 5.180 1.460 5.250 ;
        RECT 4.200 5.180 4.360 5.250 ;
        RECT 7.100 5.180 7.260 5.250 ;
        RECT 10.000 5.180 10.160 5.250 ;
        RECT 12.900 5.180 13.060 5.250 ;
        RECT 15.800 5.180 15.960 5.250 ;
        RECT 18.700 5.180 18.860 5.250 ;
        RECT 21.600 5.180 21.760 5.250 ;
        RECT 24.500 5.180 24.660 5.250 ;
        RECT 27.400 5.180 27.560 5.250 ;
        RECT 30.300 5.180 30.460 5.250 ;
        RECT 33.200 5.180 33.360 5.250 ;
        RECT 36.100 5.180 36.260 5.250 ;
        RECT 39.000 5.180 39.160 5.250 ;
        RECT 41.900 5.180 42.060 5.250 ;
        RECT 44.800 5.180 44.960 5.250 ;
        RECT 47.700 5.180 47.860 5.250 ;
        RECT 50.600 5.180 50.760 5.250 ;
        RECT 53.500 5.180 53.660 5.250 ;
        RECT 56.400 5.180 56.560 5.250 ;
        RECT 59.300 5.180 59.460 5.250 ;
        RECT 62.200 5.180 62.360 5.250 ;
        RECT 65.100 5.180 65.260 5.250 ;
        RECT 68.000 5.180 68.160 5.250 ;
        RECT 70.900 5.180 71.060 5.250 ;
        RECT 73.800 5.180 73.960 5.250 ;
        RECT 76.700 5.180 76.860 5.250 ;
        RECT 79.600 5.180 79.760 5.250 ;
        RECT 82.500 5.180 82.660 5.250 ;
        RECT 85.400 5.180 85.560 5.250 ;
        RECT 88.300 5.180 88.460 5.250 ;
        RECT 91.200 5.180 91.360 5.250 ;
        RECT 1.310 5.170 1.450 5.180 ;
        RECT 4.210 5.170 4.350 5.180 ;
        RECT 7.110 5.170 7.250 5.180 ;
        RECT 10.010 5.170 10.150 5.180 ;
        RECT 12.910 5.170 13.050 5.180 ;
        RECT 15.810 5.170 15.950 5.180 ;
        RECT 18.710 5.170 18.850 5.180 ;
        RECT 21.610 5.170 21.750 5.180 ;
        RECT 24.510 5.170 24.650 5.180 ;
        RECT 27.410 5.170 27.550 5.180 ;
        RECT 30.310 5.170 30.450 5.180 ;
        RECT 33.210 5.170 33.350 5.180 ;
        RECT 36.110 5.170 36.250 5.180 ;
        RECT 39.010 5.170 39.150 5.180 ;
        RECT 41.910 5.170 42.050 5.180 ;
        RECT 44.810 5.170 44.950 5.180 ;
        RECT 47.710 5.170 47.850 5.180 ;
        RECT 50.610 5.170 50.750 5.180 ;
        RECT 53.510 5.170 53.650 5.180 ;
        RECT 56.410 5.170 56.550 5.180 ;
        RECT 59.310 5.170 59.450 5.180 ;
        RECT 62.210 5.170 62.350 5.180 ;
        RECT 65.110 5.170 65.250 5.180 ;
        RECT 68.010 5.170 68.150 5.180 ;
        RECT 70.910 5.170 71.050 5.180 ;
        RECT 73.810 5.170 73.950 5.180 ;
        RECT 76.710 5.170 76.850 5.180 ;
        RECT 79.610 5.170 79.750 5.180 ;
        RECT 82.510 5.170 82.650 5.180 ;
        RECT 85.410 5.170 85.550 5.180 ;
        RECT 88.310 5.170 88.450 5.180 ;
        RECT 91.210 5.170 91.350 5.180 ;
      LAYER met1 ;
        RECT 0.000 5.180 92.660 5.250 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.990 3.420 1.755 3.900 ;
        RECT 3.890 3.420 4.655 3.900 ;
        RECT 6.790 3.420 7.555 3.900 ;
        RECT 9.690 3.420 10.455 3.900 ;
        RECT 12.590 3.420 13.355 3.900 ;
        RECT 15.490 3.420 16.255 3.900 ;
        RECT 18.390 3.420 19.155 3.900 ;
        RECT 21.290 3.420 22.055 3.900 ;
        RECT 24.190 3.420 24.955 3.900 ;
        RECT 27.090 3.420 27.855 3.900 ;
        RECT 29.990 3.420 30.755 3.900 ;
        RECT 32.890 3.420 33.655 3.900 ;
        RECT 35.790 3.420 36.555 3.900 ;
        RECT 38.690 3.420 39.455 3.900 ;
        RECT 41.590 3.420 42.355 3.900 ;
        RECT 44.490 3.420 45.255 3.900 ;
        RECT 47.390 3.420 48.155 3.900 ;
        RECT 50.290 3.420 51.055 3.900 ;
        RECT 53.190 3.420 53.955 3.900 ;
        RECT 56.090 3.420 56.855 3.900 ;
        RECT 58.990 3.420 59.755 3.900 ;
        RECT 61.890 3.420 62.655 3.900 ;
        RECT 64.790 3.420 65.555 3.900 ;
        RECT 67.690 3.420 68.455 3.900 ;
        RECT 70.590 3.420 71.355 3.900 ;
        RECT 73.490 3.420 74.255 3.900 ;
        RECT 76.390 3.420 77.155 3.900 ;
        RECT 79.290 3.420 80.055 3.900 ;
        RECT 82.190 3.420 82.955 3.900 ;
        RECT 85.090 3.420 85.855 3.900 ;
        RECT 87.990 3.420 88.755 3.900 ;
        RECT 90.890 3.420 91.655 3.900 ;
      LAYER li1 ;
        RECT 1.300 3.830 1.460 3.900 ;
        RECT 4.200 3.830 4.360 3.900 ;
        RECT 7.100 3.830 7.260 3.900 ;
        RECT 10.000 3.830 10.160 3.900 ;
        RECT 12.900 3.830 13.060 3.900 ;
        RECT 15.800 3.830 15.960 3.900 ;
        RECT 18.700 3.830 18.860 3.900 ;
        RECT 21.600 3.830 21.760 3.900 ;
        RECT 24.500 3.830 24.660 3.900 ;
        RECT 27.400 3.830 27.560 3.900 ;
        RECT 30.300 3.830 30.460 3.900 ;
        RECT 33.200 3.830 33.360 3.900 ;
        RECT 36.100 3.830 36.260 3.900 ;
        RECT 39.000 3.830 39.160 3.900 ;
        RECT 41.900 3.830 42.060 3.900 ;
        RECT 44.800 3.830 44.960 3.900 ;
        RECT 47.700 3.830 47.860 3.900 ;
        RECT 50.600 3.830 50.760 3.900 ;
        RECT 53.500 3.830 53.660 3.900 ;
        RECT 56.400 3.830 56.560 3.900 ;
        RECT 59.300 3.830 59.460 3.900 ;
        RECT 62.200 3.830 62.360 3.900 ;
        RECT 65.100 3.830 65.260 3.900 ;
        RECT 68.000 3.830 68.160 3.900 ;
        RECT 70.900 3.830 71.060 3.900 ;
        RECT 73.800 3.830 73.960 3.900 ;
        RECT 76.700 3.830 76.860 3.900 ;
        RECT 79.600 3.830 79.760 3.900 ;
        RECT 82.500 3.830 82.660 3.900 ;
        RECT 85.400 3.830 85.560 3.900 ;
        RECT 88.300 3.830 88.460 3.900 ;
        RECT 91.200 3.830 91.360 3.900 ;
        RECT 1.310 3.820 1.450 3.830 ;
        RECT 4.210 3.820 4.350 3.830 ;
        RECT 7.110 3.820 7.250 3.830 ;
        RECT 10.010 3.820 10.150 3.830 ;
        RECT 12.910 3.820 13.050 3.830 ;
        RECT 15.810 3.820 15.950 3.830 ;
        RECT 18.710 3.820 18.850 3.830 ;
        RECT 21.610 3.820 21.750 3.830 ;
        RECT 24.510 3.820 24.650 3.830 ;
        RECT 27.410 3.820 27.550 3.830 ;
        RECT 30.310 3.820 30.450 3.830 ;
        RECT 33.210 3.820 33.350 3.830 ;
        RECT 36.110 3.820 36.250 3.830 ;
        RECT 39.010 3.820 39.150 3.830 ;
        RECT 41.910 3.820 42.050 3.830 ;
        RECT 44.810 3.820 44.950 3.830 ;
        RECT 47.710 3.820 47.850 3.830 ;
        RECT 50.610 3.820 50.750 3.830 ;
        RECT 53.510 3.820 53.650 3.830 ;
        RECT 56.410 3.820 56.550 3.830 ;
        RECT 59.310 3.820 59.450 3.830 ;
        RECT 62.210 3.820 62.350 3.830 ;
        RECT 65.110 3.820 65.250 3.830 ;
        RECT 68.010 3.820 68.150 3.830 ;
        RECT 70.910 3.820 71.050 3.830 ;
        RECT 73.810 3.820 73.950 3.830 ;
        RECT 76.710 3.820 76.850 3.830 ;
        RECT 79.610 3.820 79.750 3.830 ;
        RECT 82.510 3.820 82.650 3.830 ;
        RECT 85.410 3.820 85.550 3.830 ;
        RECT 88.310 3.820 88.450 3.830 ;
        RECT 91.210 3.820 91.350 3.830 ;
      LAYER met1 ;
        RECT 0.000 3.830 92.660 3.900 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.990 0.720 1.755 1.200 ;
        RECT 3.890 0.720 4.655 1.200 ;
        RECT 6.790 0.720 7.555 1.200 ;
        RECT 9.690 0.720 10.455 1.200 ;
        RECT 12.590 0.720 13.355 1.200 ;
        RECT 15.490 0.720 16.255 1.200 ;
        RECT 18.390 0.720 19.155 1.200 ;
        RECT 21.290 0.720 22.055 1.200 ;
        RECT 24.190 0.725 24.955 1.205 ;
        RECT 27.090 0.725 27.855 1.205 ;
        RECT 29.990 0.725 30.755 1.205 ;
        RECT 32.890 0.725 33.655 1.205 ;
        RECT 35.790 0.725 36.555 1.205 ;
        RECT 38.690 0.725 39.455 1.205 ;
        RECT 41.590 0.725 42.355 1.205 ;
        RECT 44.490 0.725 45.255 1.205 ;
        RECT 47.390 0.725 48.155 1.205 ;
        RECT 50.290 0.725 51.055 1.205 ;
        RECT 53.190 0.725 53.955 1.205 ;
        RECT 56.090 0.725 56.855 1.205 ;
        RECT 58.990 0.725 59.755 1.205 ;
        RECT 61.890 0.725 62.655 1.205 ;
        RECT 64.790 0.725 65.555 1.205 ;
        RECT 67.690 0.725 68.455 1.205 ;
        RECT 70.590 0.725 71.355 1.205 ;
        RECT 73.490 0.725 74.255 1.205 ;
        RECT 76.390 0.725 77.155 1.205 ;
        RECT 79.290 0.725 80.055 1.205 ;
        RECT 82.190 0.725 82.955 1.205 ;
        RECT 85.090 0.725 85.855 1.205 ;
        RECT 87.990 0.725 88.755 1.205 ;
        RECT 90.890 0.725 91.655 1.205 ;
      LAYER li1 ;
        RECT 1.300 1.130 1.460 1.200 ;
        RECT 4.200 1.130 4.360 1.200 ;
        RECT 7.100 1.130 7.260 1.200 ;
        RECT 10.000 1.130 10.160 1.200 ;
        RECT 12.900 1.130 13.060 1.200 ;
        RECT 15.800 1.130 15.960 1.200 ;
        RECT 18.700 1.130 18.860 1.200 ;
        RECT 21.600 1.130 21.760 1.200 ;
        RECT 24.500 1.135 24.660 1.205 ;
        RECT 27.400 1.135 27.560 1.205 ;
        RECT 30.300 1.135 30.460 1.205 ;
        RECT 33.200 1.135 33.360 1.205 ;
        RECT 36.100 1.135 36.260 1.205 ;
        RECT 39.000 1.135 39.160 1.205 ;
        RECT 41.900 1.135 42.060 1.205 ;
        RECT 44.800 1.135 44.960 1.205 ;
        RECT 47.700 1.135 47.860 1.205 ;
        RECT 50.600 1.135 50.760 1.205 ;
        RECT 53.500 1.135 53.660 1.205 ;
        RECT 56.400 1.135 56.560 1.205 ;
        RECT 59.300 1.135 59.460 1.205 ;
        RECT 62.200 1.135 62.360 1.205 ;
        RECT 65.100 1.135 65.260 1.205 ;
        RECT 68.000 1.135 68.160 1.205 ;
        RECT 70.900 1.135 71.060 1.205 ;
        RECT 73.800 1.135 73.960 1.205 ;
        RECT 76.700 1.135 76.860 1.205 ;
        RECT 79.600 1.135 79.760 1.205 ;
        RECT 82.500 1.135 82.660 1.205 ;
        RECT 85.400 1.135 85.560 1.205 ;
        RECT 88.300 1.135 88.460 1.205 ;
        RECT 91.200 1.135 91.360 1.205 ;
        RECT 1.310 1.120 1.450 1.130 ;
        RECT 4.210 1.120 4.350 1.130 ;
        RECT 7.110 1.120 7.250 1.130 ;
        RECT 10.010 1.120 10.150 1.130 ;
        RECT 12.910 1.120 13.050 1.130 ;
        RECT 15.810 1.120 15.950 1.130 ;
        RECT 18.710 1.120 18.850 1.130 ;
        RECT 21.610 1.120 21.750 1.130 ;
        RECT 24.510 1.125 24.650 1.135 ;
        RECT 27.410 1.125 27.550 1.135 ;
        RECT 30.310 1.125 30.450 1.135 ;
        RECT 33.210 1.125 33.350 1.135 ;
        RECT 36.110 1.125 36.250 1.135 ;
        RECT 39.010 1.125 39.150 1.135 ;
        RECT 41.910 1.125 42.050 1.135 ;
        RECT 44.810 1.125 44.950 1.135 ;
        RECT 47.710 1.125 47.850 1.135 ;
        RECT 50.610 1.125 50.750 1.135 ;
        RECT 53.510 1.125 53.650 1.135 ;
        RECT 56.410 1.125 56.550 1.135 ;
        RECT 59.310 1.125 59.450 1.135 ;
        RECT 62.210 1.125 62.350 1.135 ;
        RECT 65.110 1.125 65.250 1.135 ;
        RECT 68.010 1.125 68.150 1.135 ;
        RECT 70.910 1.125 71.050 1.135 ;
        RECT 73.810 1.125 73.950 1.135 ;
        RECT 76.710 1.125 76.850 1.135 ;
        RECT 79.610 1.125 79.750 1.135 ;
        RECT 82.510 1.125 82.650 1.135 ;
        RECT 85.410 1.125 85.550 1.135 ;
        RECT 88.310 1.125 88.450 1.135 ;
        RECT 91.210 1.125 91.350 1.135 ;
      LAYER met1 ;
        RECT 23.155 1.200 92.660 1.205 ;
        RECT 0.000 1.135 92.660 1.200 ;
        RECT 0.000 1.130 23.155 1.135 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.990 2.070 1.755 2.550 ;
        RECT 3.890 2.070 4.655 2.550 ;
        RECT 6.790 2.070 7.555 2.550 ;
        RECT 9.690 2.070 10.455 2.550 ;
        RECT 12.590 2.070 13.355 2.550 ;
        RECT 15.490 2.070 16.255 2.550 ;
        RECT 18.390 2.070 19.155 2.550 ;
        RECT 21.290 2.070 22.055 2.550 ;
        RECT 24.190 2.075 24.955 2.555 ;
        RECT 27.090 2.075 27.855 2.555 ;
        RECT 29.990 2.075 30.755 2.555 ;
        RECT 32.890 2.075 33.655 2.555 ;
        RECT 35.790 2.075 36.555 2.555 ;
        RECT 38.690 2.075 39.455 2.555 ;
        RECT 41.590 2.075 42.355 2.555 ;
        RECT 44.490 2.075 45.255 2.555 ;
        RECT 47.390 2.075 48.155 2.555 ;
        RECT 50.290 2.075 51.055 2.555 ;
        RECT 53.190 2.075 53.955 2.555 ;
        RECT 56.090 2.075 56.855 2.555 ;
        RECT 58.990 2.075 59.755 2.555 ;
        RECT 61.890 2.075 62.655 2.555 ;
        RECT 64.790 2.075 65.555 2.555 ;
        RECT 67.690 2.075 68.455 2.555 ;
        RECT 70.590 2.075 71.355 2.555 ;
        RECT 73.490 2.075 74.255 2.555 ;
        RECT 76.390 2.075 77.155 2.555 ;
        RECT 79.290 2.075 80.055 2.555 ;
        RECT 82.190 2.075 82.955 2.555 ;
        RECT 85.090 2.075 85.855 2.555 ;
        RECT 87.990 2.075 88.755 2.555 ;
        RECT 90.890 2.075 91.655 2.555 ;
      LAYER li1 ;
        RECT 1.300 2.480 1.460 2.550 ;
        RECT 4.200 2.480 4.360 2.550 ;
        RECT 7.100 2.480 7.260 2.550 ;
        RECT 10.000 2.480 10.160 2.550 ;
        RECT 12.900 2.480 13.060 2.550 ;
        RECT 15.800 2.480 15.960 2.550 ;
        RECT 18.700 2.480 18.860 2.550 ;
        RECT 21.600 2.480 21.760 2.550 ;
        RECT 24.500 2.485 24.660 2.555 ;
        RECT 27.400 2.485 27.560 2.555 ;
        RECT 30.300 2.485 30.460 2.555 ;
        RECT 33.200 2.485 33.360 2.555 ;
        RECT 36.100 2.485 36.260 2.555 ;
        RECT 39.000 2.485 39.160 2.555 ;
        RECT 41.900 2.485 42.060 2.555 ;
        RECT 44.800 2.485 44.960 2.555 ;
        RECT 47.700 2.485 47.860 2.555 ;
        RECT 50.600 2.485 50.760 2.555 ;
        RECT 53.500 2.485 53.660 2.555 ;
        RECT 56.400 2.485 56.560 2.555 ;
        RECT 59.300 2.485 59.460 2.555 ;
        RECT 62.200 2.485 62.360 2.555 ;
        RECT 65.100 2.485 65.260 2.555 ;
        RECT 68.000 2.485 68.160 2.555 ;
        RECT 70.900 2.485 71.060 2.555 ;
        RECT 73.800 2.485 73.960 2.555 ;
        RECT 76.700 2.485 76.860 2.555 ;
        RECT 79.600 2.485 79.760 2.555 ;
        RECT 82.500 2.485 82.660 2.555 ;
        RECT 85.400 2.485 85.560 2.555 ;
        RECT 88.300 2.485 88.460 2.555 ;
        RECT 91.200 2.485 91.360 2.555 ;
        RECT 1.310 2.470 1.450 2.480 ;
        RECT 4.210 2.470 4.350 2.480 ;
        RECT 7.110 2.470 7.250 2.480 ;
        RECT 10.010 2.470 10.150 2.480 ;
        RECT 12.910 2.470 13.050 2.480 ;
        RECT 15.810 2.470 15.950 2.480 ;
        RECT 18.710 2.470 18.850 2.480 ;
        RECT 21.610 2.470 21.750 2.480 ;
        RECT 24.510 2.475 24.650 2.485 ;
        RECT 27.410 2.475 27.550 2.485 ;
        RECT 30.310 2.475 30.450 2.485 ;
        RECT 33.210 2.475 33.350 2.485 ;
        RECT 36.110 2.475 36.250 2.485 ;
        RECT 39.010 2.475 39.150 2.485 ;
        RECT 41.910 2.475 42.050 2.485 ;
        RECT 44.810 2.475 44.950 2.485 ;
        RECT 47.710 2.475 47.850 2.485 ;
        RECT 50.610 2.475 50.750 2.485 ;
        RECT 53.510 2.475 53.650 2.485 ;
        RECT 56.410 2.475 56.550 2.485 ;
        RECT 59.310 2.475 59.450 2.485 ;
        RECT 62.210 2.475 62.350 2.485 ;
        RECT 65.110 2.475 65.250 2.485 ;
        RECT 68.010 2.475 68.150 2.485 ;
        RECT 70.910 2.475 71.050 2.485 ;
        RECT 73.810 2.475 73.950 2.485 ;
        RECT 76.710 2.475 76.850 2.485 ;
        RECT 79.610 2.475 79.750 2.485 ;
        RECT 82.510 2.475 82.650 2.485 ;
        RECT 85.410 2.475 85.550 2.485 ;
        RECT 88.310 2.475 88.450 2.485 ;
        RECT 91.210 2.475 91.350 2.485 ;
      LAYER met1 ;
        RECT 23.200 2.550 69.460 2.555 ;
        RECT 69.600 2.550 92.660 2.555 ;
        RECT 0.000 2.485 92.660 2.550 ;
        RECT 0.000 2.480 23.275 2.485 ;
        RECT 69.460 2.480 69.675 2.485 ;
        RECT 0.000 2.475 0.075 2.480 ;
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER pwell ;
        RECT 0.000 42.340 0.850 43.200 ;
        RECT 1.910 42.340 3.750 43.200 ;
        RECT 4.810 42.340 6.650 43.200 ;
        RECT 7.710 42.340 9.550 43.200 ;
        RECT 10.610 42.340 12.450 43.200 ;
        RECT 13.510 42.340 15.350 43.200 ;
        RECT 16.410 42.340 18.250 43.200 ;
        RECT 19.310 42.340 21.150 43.200 ;
        RECT 22.210 42.340 23.060 43.200 ;
        RECT 0.000 41.850 23.060 42.340 ;
        RECT 0.000 40.990 0.850 41.850 ;
        RECT 1.910 40.990 3.750 41.850 ;
        RECT 4.810 40.990 6.650 41.850 ;
        RECT 7.710 40.990 9.550 41.850 ;
        RECT 10.610 40.990 12.450 41.850 ;
        RECT 13.510 40.990 15.350 41.850 ;
        RECT 16.410 40.990 18.250 41.850 ;
        RECT 19.310 40.990 21.150 41.850 ;
        RECT 22.210 40.990 23.060 41.850 ;
        RECT 0.000 40.500 23.060 40.990 ;
        RECT 0.000 39.640 0.850 40.500 ;
        RECT 1.910 39.640 3.750 40.500 ;
        RECT 4.810 39.640 6.650 40.500 ;
        RECT 7.710 39.640 9.550 40.500 ;
        RECT 10.610 39.640 12.450 40.500 ;
        RECT 13.510 39.640 15.350 40.500 ;
        RECT 16.410 39.640 18.250 40.500 ;
        RECT 19.310 39.640 21.150 40.500 ;
        RECT 22.210 39.640 23.060 40.500 ;
        RECT 0.000 39.150 23.060 39.640 ;
        RECT 0.000 38.290 0.850 39.150 ;
        RECT 1.910 38.290 3.750 39.150 ;
        RECT 4.810 38.290 6.650 39.150 ;
        RECT 7.710 38.290 9.550 39.150 ;
        RECT 10.610 38.290 12.450 39.150 ;
        RECT 13.510 38.290 15.350 39.150 ;
        RECT 16.410 38.290 18.250 39.150 ;
        RECT 19.310 38.290 21.150 39.150 ;
        RECT 22.210 38.290 23.060 39.150 ;
        RECT 0.000 37.870 23.060 38.290 ;
        RECT 23.200 42.340 24.050 43.200 ;
        RECT 25.110 42.340 26.950 43.200 ;
        RECT 28.010 42.340 29.850 43.200 ;
        RECT 30.910 42.340 32.750 43.200 ;
        RECT 33.810 42.340 35.650 43.200 ;
        RECT 36.710 42.340 38.550 43.200 ;
        RECT 39.610 42.340 41.450 43.200 ;
        RECT 42.510 42.340 44.350 43.200 ;
        RECT 45.410 42.340 46.260 43.200 ;
        RECT 23.200 41.850 46.260 42.340 ;
        RECT 23.200 40.990 24.050 41.850 ;
        RECT 25.110 40.990 26.950 41.850 ;
        RECT 28.010 40.990 29.850 41.850 ;
        RECT 30.910 40.990 32.750 41.850 ;
        RECT 33.810 40.990 35.650 41.850 ;
        RECT 36.710 40.990 38.550 41.850 ;
        RECT 39.610 40.990 41.450 41.850 ;
        RECT 42.510 40.990 44.350 41.850 ;
        RECT 45.410 40.990 46.260 41.850 ;
        RECT 23.200 40.500 46.260 40.990 ;
        RECT 23.200 39.640 24.050 40.500 ;
        RECT 25.110 39.640 26.950 40.500 ;
        RECT 28.010 39.640 29.850 40.500 ;
        RECT 30.910 39.640 32.750 40.500 ;
        RECT 33.810 39.640 35.650 40.500 ;
        RECT 36.710 39.640 38.550 40.500 ;
        RECT 39.610 39.640 41.450 40.500 ;
        RECT 42.510 39.640 44.350 40.500 ;
        RECT 45.410 39.640 46.260 40.500 ;
        RECT 23.200 39.150 46.260 39.640 ;
        RECT 23.200 38.290 24.050 39.150 ;
        RECT 25.110 38.290 26.950 39.150 ;
        RECT 28.010 38.290 29.850 39.150 ;
        RECT 30.910 38.290 32.750 39.150 ;
        RECT 33.810 38.290 35.650 39.150 ;
        RECT 36.710 38.290 38.550 39.150 ;
        RECT 39.610 38.290 41.450 39.150 ;
        RECT 42.510 38.290 44.350 39.150 ;
        RECT 45.410 38.290 46.260 39.150 ;
        RECT 23.200 37.870 46.260 38.290 ;
        RECT 0.000 37.800 46.260 37.870 ;
        RECT 0.000 36.940 0.850 37.800 ;
        RECT 1.910 36.940 3.750 37.800 ;
        RECT 4.810 36.940 6.650 37.800 ;
        RECT 7.710 36.940 9.550 37.800 ;
        RECT 10.610 36.940 12.450 37.800 ;
        RECT 13.510 36.940 15.350 37.800 ;
        RECT 16.410 36.940 18.250 37.800 ;
        RECT 19.310 36.940 21.150 37.800 ;
        RECT 22.210 37.650 23.060 37.800 ;
        RECT 23.200 37.650 24.050 37.800 ;
        RECT 22.210 37.580 24.050 37.650 ;
        RECT 22.210 36.940 23.060 37.580 ;
        RECT 0.000 36.520 23.060 36.940 ;
        RECT 23.200 36.940 24.050 37.580 ;
        RECT 25.110 36.940 26.950 37.800 ;
        RECT 28.010 36.940 29.850 37.800 ;
        RECT 30.910 36.940 32.750 37.800 ;
        RECT 33.810 36.940 35.650 37.800 ;
        RECT 36.710 36.940 38.550 37.800 ;
        RECT 39.610 36.940 41.450 37.800 ;
        RECT 42.510 36.940 44.350 37.800 ;
        RECT 45.410 36.940 46.260 37.800 ;
        RECT 23.200 36.520 46.260 36.940 ;
        RECT 0.000 36.450 46.260 36.520 ;
        RECT 0.000 35.590 0.850 36.450 ;
        RECT 1.910 35.590 3.750 36.450 ;
        RECT 4.810 35.590 6.650 36.450 ;
        RECT 7.710 35.590 9.550 36.450 ;
        RECT 10.610 35.590 12.450 36.450 ;
        RECT 13.510 35.590 15.350 36.450 ;
        RECT 16.410 35.590 18.250 36.450 ;
        RECT 19.310 35.590 21.150 36.450 ;
        RECT 22.210 36.300 23.060 36.450 ;
        RECT 23.200 36.300 24.050 36.450 ;
        RECT 22.210 36.230 24.050 36.300 ;
        RECT 22.210 35.590 23.060 36.230 ;
        RECT 0.000 35.170 23.060 35.590 ;
        RECT 23.200 35.590 24.050 36.230 ;
        RECT 25.110 35.590 26.950 36.450 ;
        RECT 28.010 35.590 29.850 36.450 ;
        RECT 30.910 35.590 32.750 36.450 ;
        RECT 33.810 35.590 35.650 36.450 ;
        RECT 36.710 35.590 38.550 36.450 ;
        RECT 39.610 35.590 41.450 36.450 ;
        RECT 42.510 35.590 44.350 36.450 ;
        RECT 45.410 35.590 46.260 36.450 ;
        RECT 23.200 35.170 46.260 35.590 ;
        RECT 0.000 35.100 46.260 35.170 ;
        RECT 0.000 34.240 0.850 35.100 ;
        RECT 1.910 34.240 3.750 35.100 ;
        RECT 4.810 34.240 6.650 35.100 ;
        RECT 7.710 34.240 9.550 35.100 ;
        RECT 10.610 34.240 12.450 35.100 ;
        RECT 13.510 34.240 15.350 35.100 ;
        RECT 16.410 34.240 18.250 35.100 ;
        RECT 19.310 34.240 21.150 35.100 ;
        RECT 22.210 34.950 23.060 35.100 ;
        RECT 23.200 34.950 24.050 35.100 ;
        RECT 22.210 34.880 24.050 34.950 ;
        RECT 22.210 34.240 23.060 34.880 ;
        RECT 0.000 33.820 23.060 34.240 ;
        RECT 23.200 34.240 24.050 34.880 ;
        RECT 25.110 34.240 26.950 35.100 ;
        RECT 28.010 34.240 29.850 35.100 ;
        RECT 30.910 34.240 32.750 35.100 ;
        RECT 33.810 34.240 35.650 35.100 ;
        RECT 36.710 34.240 38.550 35.100 ;
        RECT 39.610 34.240 41.450 35.100 ;
        RECT 42.510 34.240 44.350 35.100 ;
        RECT 45.410 34.240 46.260 35.100 ;
        RECT 23.200 33.820 46.260 34.240 ;
        RECT 0.000 33.750 46.260 33.820 ;
        RECT 0.000 32.890 0.850 33.750 ;
        RECT 1.910 32.890 3.750 33.750 ;
        RECT 4.810 32.890 6.650 33.750 ;
        RECT 7.710 32.890 9.550 33.750 ;
        RECT 10.610 32.890 12.450 33.750 ;
        RECT 13.510 32.890 15.350 33.750 ;
        RECT 16.410 32.890 18.250 33.750 ;
        RECT 19.310 32.890 21.150 33.750 ;
        RECT 22.210 33.600 23.060 33.750 ;
        RECT 23.200 33.600 24.050 33.750 ;
        RECT 22.210 33.530 24.050 33.600 ;
        RECT 22.210 32.890 23.060 33.530 ;
        RECT 0.000 32.470 23.060 32.890 ;
        RECT 23.200 32.890 24.050 33.530 ;
        RECT 25.110 32.890 26.950 33.750 ;
        RECT 28.010 32.890 29.850 33.750 ;
        RECT 30.910 32.890 32.750 33.750 ;
        RECT 33.810 32.890 35.650 33.750 ;
        RECT 36.710 32.890 38.550 33.750 ;
        RECT 39.610 32.890 41.450 33.750 ;
        RECT 42.510 32.890 44.350 33.750 ;
        RECT 45.410 32.890 46.260 33.750 ;
        RECT 23.200 32.470 46.260 32.890 ;
        RECT 0.000 32.400 46.260 32.470 ;
        RECT 0.000 31.540 0.850 32.400 ;
        RECT 1.910 31.540 3.750 32.400 ;
        RECT 4.810 31.540 6.650 32.400 ;
        RECT 7.710 31.540 9.550 32.400 ;
        RECT 10.610 31.540 12.450 32.400 ;
        RECT 13.510 31.540 15.350 32.400 ;
        RECT 16.410 31.540 18.250 32.400 ;
        RECT 19.310 31.540 21.150 32.400 ;
        RECT 22.210 32.250 23.060 32.400 ;
        RECT 23.200 32.250 24.050 32.400 ;
        RECT 22.210 32.180 24.050 32.250 ;
        RECT 22.210 31.540 23.060 32.180 ;
        RECT 0.000 31.120 23.060 31.540 ;
        RECT 23.200 31.540 24.050 32.180 ;
        RECT 25.110 31.540 26.950 32.400 ;
        RECT 28.010 31.540 29.850 32.400 ;
        RECT 30.910 31.540 32.750 32.400 ;
        RECT 33.810 31.540 35.650 32.400 ;
        RECT 36.710 31.540 38.550 32.400 ;
        RECT 39.610 31.540 41.450 32.400 ;
        RECT 42.510 31.540 44.350 32.400 ;
        RECT 45.410 31.540 46.260 32.400 ;
        RECT 23.200 31.120 46.260 31.540 ;
        RECT 0.000 31.050 46.260 31.120 ;
        RECT 0.000 30.190 0.850 31.050 ;
        RECT 1.910 30.190 3.750 31.050 ;
        RECT 4.810 30.190 6.650 31.050 ;
        RECT 7.710 30.190 9.550 31.050 ;
        RECT 10.610 30.190 12.450 31.050 ;
        RECT 13.510 30.190 15.350 31.050 ;
        RECT 16.410 30.190 18.250 31.050 ;
        RECT 19.310 30.190 21.150 31.050 ;
        RECT 22.210 30.900 23.060 31.050 ;
        RECT 23.200 30.900 24.050 31.050 ;
        RECT 22.210 30.830 24.050 30.900 ;
        RECT 22.210 30.190 23.060 30.830 ;
        RECT 0.000 29.770 23.060 30.190 ;
        RECT 23.200 30.190 24.050 30.830 ;
        RECT 25.110 30.190 26.950 31.050 ;
        RECT 28.010 30.190 29.850 31.050 ;
        RECT 30.910 30.190 32.750 31.050 ;
        RECT 33.810 30.190 35.650 31.050 ;
        RECT 36.710 30.190 38.550 31.050 ;
        RECT 39.610 30.190 41.450 31.050 ;
        RECT 42.510 30.190 44.350 31.050 ;
        RECT 45.410 30.190 46.260 31.050 ;
        RECT 23.200 29.770 46.260 30.190 ;
        RECT 0.000 29.700 46.260 29.770 ;
        RECT 0.000 28.840 0.850 29.700 ;
        RECT 1.910 28.840 3.750 29.700 ;
        RECT 4.810 28.840 6.650 29.700 ;
        RECT 7.710 28.840 9.550 29.700 ;
        RECT 10.610 28.840 12.450 29.700 ;
        RECT 13.510 28.840 15.350 29.700 ;
        RECT 16.410 28.840 18.250 29.700 ;
        RECT 19.310 28.840 21.150 29.700 ;
        RECT 22.210 29.550 23.060 29.700 ;
        RECT 23.200 29.550 24.050 29.700 ;
        RECT 22.210 29.480 24.050 29.550 ;
        RECT 22.210 28.840 23.060 29.480 ;
        RECT 0.000 28.420 23.060 28.840 ;
        RECT 23.200 28.840 24.050 29.480 ;
        RECT 25.110 28.840 26.950 29.700 ;
        RECT 28.010 28.840 29.850 29.700 ;
        RECT 30.910 28.840 32.750 29.700 ;
        RECT 33.810 28.840 35.650 29.700 ;
        RECT 36.710 28.840 38.550 29.700 ;
        RECT 39.610 28.840 41.450 29.700 ;
        RECT 42.510 28.840 44.350 29.700 ;
        RECT 45.410 28.840 46.260 29.700 ;
        RECT 23.200 28.420 46.260 28.840 ;
        RECT 0.000 28.350 46.260 28.420 ;
        RECT 0.000 27.490 0.850 28.350 ;
        RECT 1.910 27.490 3.750 28.350 ;
        RECT 4.810 27.490 6.650 28.350 ;
        RECT 7.710 27.490 9.550 28.350 ;
        RECT 10.610 27.490 12.450 28.350 ;
        RECT 13.510 27.490 15.350 28.350 ;
        RECT 16.410 27.490 18.250 28.350 ;
        RECT 19.310 27.490 21.150 28.350 ;
        RECT 22.210 28.200 23.060 28.350 ;
        RECT 23.200 28.200 24.050 28.350 ;
        RECT 22.210 28.130 24.050 28.200 ;
        RECT 22.210 27.490 23.060 28.130 ;
        RECT 0.000 27.070 23.060 27.490 ;
        RECT 23.200 27.490 24.050 28.130 ;
        RECT 25.110 27.490 26.950 28.350 ;
        RECT 28.010 27.490 29.850 28.350 ;
        RECT 30.910 27.490 32.750 28.350 ;
        RECT 33.810 27.490 35.650 28.350 ;
        RECT 36.710 27.490 38.550 28.350 ;
        RECT 39.610 27.490 41.450 28.350 ;
        RECT 42.510 27.490 44.350 28.350 ;
        RECT 45.410 27.490 46.260 28.350 ;
        RECT 23.200 27.070 46.260 27.490 ;
        RECT 0.000 27.000 46.260 27.070 ;
        RECT 0.000 26.140 0.850 27.000 ;
        RECT 1.910 26.140 3.750 27.000 ;
        RECT 4.810 26.140 6.650 27.000 ;
        RECT 7.710 26.140 9.550 27.000 ;
        RECT 10.610 26.140 12.450 27.000 ;
        RECT 13.510 26.140 15.350 27.000 ;
        RECT 16.410 26.140 18.250 27.000 ;
        RECT 19.310 26.140 21.150 27.000 ;
        RECT 22.210 26.850 23.060 27.000 ;
        RECT 23.200 26.850 24.050 27.000 ;
        RECT 22.210 26.780 24.050 26.850 ;
        RECT 22.210 26.140 23.060 26.780 ;
        RECT 0.000 25.720 23.060 26.140 ;
        RECT 23.200 26.140 24.050 26.780 ;
        RECT 25.110 26.140 26.950 27.000 ;
        RECT 28.010 26.140 29.850 27.000 ;
        RECT 30.910 26.140 32.750 27.000 ;
        RECT 33.810 26.140 35.650 27.000 ;
        RECT 36.710 26.140 38.550 27.000 ;
        RECT 39.610 26.140 41.450 27.000 ;
        RECT 42.510 26.140 44.350 27.000 ;
        RECT 45.410 26.140 46.260 27.000 ;
        RECT 23.200 25.720 46.260 26.140 ;
        RECT 0.000 25.650 46.260 25.720 ;
        RECT 0.000 24.790 0.850 25.650 ;
        RECT 1.910 24.790 3.750 25.650 ;
        RECT 4.810 24.790 6.650 25.650 ;
        RECT 7.710 24.790 9.550 25.650 ;
        RECT 10.610 24.790 12.450 25.650 ;
        RECT 13.510 24.790 15.350 25.650 ;
        RECT 16.410 24.790 18.250 25.650 ;
        RECT 19.310 24.790 21.150 25.650 ;
        RECT 22.210 25.500 23.060 25.650 ;
        RECT 23.200 25.500 24.050 25.650 ;
        RECT 22.210 25.430 24.050 25.500 ;
        RECT 22.210 24.790 23.060 25.430 ;
        RECT 0.000 24.370 23.060 24.790 ;
        RECT 23.200 24.790 24.050 25.430 ;
        RECT 25.110 24.790 26.950 25.650 ;
        RECT 28.010 24.790 29.850 25.650 ;
        RECT 30.910 24.790 32.750 25.650 ;
        RECT 33.810 24.790 35.650 25.650 ;
        RECT 36.710 24.790 38.550 25.650 ;
        RECT 39.610 24.790 41.450 25.650 ;
        RECT 42.510 24.790 44.350 25.650 ;
        RECT 45.410 24.790 46.260 25.650 ;
        RECT 23.200 24.370 46.260 24.790 ;
        RECT 0.000 24.300 46.260 24.370 ;
        RECT 0.000 23.440 0.850 24.300 ;
        RECT 1.910 23.440 3.750 24.300 ;
        RECT 4.810 23.440 6.650 24.300 ;
        RECT 7.710 23.440 9.550 24.300 ;
        RECT 10.610 23.440 12.450 24.300 ;
        RECT 13.510 23.440 15.350 24.300 ;
        RECT 16.410 23.440 18.250 24.300 ;
        RECT 19.310 23.440 21.150 24.300 ;
        RECT 22.210 24.150 23.060 24.300 ;
        RECT 23.200 24.150 24.050 24.300 ;
        RECT 22.210 24.080 24.050 24.150 ;
        RECT 22.210 23.440 23.060 24.080 ;
        RECT 0.000 23.020 23.060 23.440 ;
        RECT 23.200 23.440 24.050 24.080 ;
        RECT 25.110 23.440 26.950 24.300 ;
        RECT 28.010 23.440 29.850 24.300 ;
        RECT 30.910 23.440 32.750 24.300 ;
        RECT 33.810 23.440 35.650 24.300 ;
        RECT 36.710 23.440 38.550 24.300 ;
        RECT 39.610 23.440 41.450 24.300 ;
        RECT 42.510 23.440 44.350 24.300 ;
        RECT 45.410 23.440 46.260 24.300 ;
        RECT 23.200 23.020 46.260 23.440 ;
        RECT 0.000 22.950 46.260 23.020 ;
        RECT 0.000 22.090 0.850 22.950 ;
        RECT 1.910 22.090 3.750 22.950 ;
        RECT 4.810 22.090 6.650 22.950 ;
        RECT 7.710 22.090 9.550 22.950 ;
        RECT 10.610 22.090 12.450 22.950 ;
        RECT 13.510 22.090 15.350 22.950 ;
        RECT 16.410 22.090 18.250 22.950 ;
        RECT 19.310 22.090 21.150 22.950 ;
        RECT 22.210 22.800 23.060 22.950 ;
        RECT 23.200 22.800 24.050 22.950 ;
        RECT 22.210 22.730 24.050 22.800 ;
        RECT 22.210 22.090 23.060 22.730 ;
        RECT 0.000 21.670 23.060 22.090 ;
        RECT 23.200 22.090 24.050 22.730 ;
        RECT 25.110 22.090 26.950 22.950 ;
        RECT 28.010 22.090 29.850 22.950 ;
        RECT 30.910 22.090 32.750 22.950 ;
        RECT 33.810 22.090 35.650 22.950 ;
        RECT 36.710 22.090 38.550 22.950 ;
        RECT 39.610 22.090 41.450 22.950 ;
        RECT 42.510 22.090 44.350 22.950 ;
        RECT 45.410 22.090 46.260 22.950 ;
        RECT 23.200 21.670 46.260 22.090 ;
        RECT 0.000 21.600 46.260 21.670 ;
        RECT 0.000 20.740 0.850 21.600 ;
        RECT 1.910 20.740 3.750 21.600 ;
        RECT 4.810 20.740 6.650 21.600 ;
        RECT 7.710 20.740 9.550 21.600 ;
        RECT 10.610 20.740 12.450 21.600 ;
        RECT 13.510 20.740 15.350 21.600 ;
        RECT 16.410 20.740 18.250 21.600 ;
        RECT 19.310 20.740 21.150 21.600 ;
        RECT 22.210 21.450 23.060 21.600 ;
        RECT 23.200 21.450 24.050 21.600 ;
        RECT 22.210 21.380 24.050 21.450 ;
        RECT 22.210 20.740 23.060 21.380 ;
        RECT 0.000 20.320 23.060 20.740 ;
        RECT 23.200 20.740 24.050 21.380 ;
        RECT 25.110 20.740 26.950 21.600 ;
        RECT 28.010 20.740 29.850 21.600 ;
        RECT 30.910 20.740 32.750 21.600 ;
        RECT 33.810 20.740 35.650 21.600 ;
        RECT 36.710 20.740 38.550 21.600 ;
        RECT 39.610 20.740 41.450 21.600 ;
        RECT 42.510 20.740 44.350 21.600 ;
        RECT 45.410 20.740 46.260 21.600 ;
        RECT 23.200 20.320 46.260 20.740 ;
        RECT 0.000 20.250 46.260 20.320 ;
        RECT 0.000 19.390 0.850 20.250 ;
        RECT 1.910 19.390 3.750 20.250 ;
        RECT 4.810 19.390 6.650 20.250 ;
        RECT 7.710 19.390 9.550 20.250 ;
        RECT 10.610 19.390 12.450 20.250 ;
        RECT 13.510 19.390 15.350 20.250 ;
        RECT 16.410 19.390 18.250 20.250 ;
        RECT 19.310 19.390 21.150 20.250 ;
        RECT 22.210 20.100 23.060 20.250 ;
        RECT 23.200 20.100 24.050 20.250 ;
        RECT 22.210 20.030 24.050 20.100 ;
        RECT 22.210 19.390 23.060 20.030 ;
        RECT 0.000 18.970 23.060 19.390 ;
        RECT 23.200 19.390 24.050 20.030 ;
        RECT 25.110 19.390 26.950 20.250 ;
        RECT 28.010 19.390 29.850 20.250 ;
        RECT 30.910 19.390 32.750 20.250 ;
        RECT 33.810 19.390 35.650 20.250 ;
        RECT 36.710 19.390 38.550 20.250 ;
        RECT 39.610 19.390 41.450 20.250 ;
        RECT 42.510 19.390 44.350 20.250 ;
        RECT 45.410 19.390 46.260 20.250 ;
        RECT 23.200 18.970 46.260 19.390 ;
        RECT 0.000 18.900 46.260 18.970 ;
        RECT 0.000 18.040 0.850 18.900 ;
        RECT 1.910 18.040 3.750 18.900 ;
        RECT 4.810 18.040 6.650 18.900 ;
        RECT 7.710 18.040 9.550 18.900 ;
        RECT 10.610 18.040 12.450 18.900 ;
        RECT 13.510 18.040 15.350 18.900 ;
        RECT 16.410 18.040 18.250 18.900 ;
        RECT 19.310 18.040 21.150 18.900 ;
        RECT 22.210 18.750 23.060 18.900 ;
        RECT 23.200 18.750 24.050 18.900 ;
        RECT 22.210 18.680 24.050 18.750 ;
        RECT 22.210 18.040 23.060 18.680 ;
        RECT 0.000 17.620 23.060 18.040 ;
        RECT 23.200 18.040 24.050 18.680 ;
        RECT 25.110 18.040 26.950 18.900 ;
        RECT 28.010 18.040 29.850 18.900 ;
        RECT 30.910 18.040 32.750 18.900 ;
        RECT 33.810 18.040 35.650 18.900 ;
        RECT 36.710 18.040 38.550 18.900 ;
        RECT 39.610 18.040 41.450 18.900 ;
        RECT 42.510 18.040 44.350 18.900 ;
        RECT 45.410 18.040 46.260 18.900 ;
        RECT 23.200 17.620 46.260 18.040 ;
        RECT 0.000 17.550 46.260 17.620 ;
        RECT 0.000 16.690 0.850 17.550 ;
        RECT 1.910 16.690 3.750 17.550 ;
        RECT 4.810 16.690 6.650 17.550 ;
        RECT 7.710 16.690 9.550 17.550 ;
        RECT 10.610 16.690 12.450 17.550 ;
        RECT 13.510 16.690 15.350 17.550 ;
        RECT 16.410 16.690 18.250 17.550 ;
        RECT 19.310 16.690 21.150 17.550 ;
        RECT 22.210 17.400 23.060 17.550 ;
        RECT 23.200 17.400 24.050 17.550 ;
        RECT 22.210 17.330 24.050 17.400 ;
        RECT 22.210 16.690 23.060 17.330 ;
        RECT 0.000 16.270 23.060 16.690 ;
        RECT 23.200 16.690 24.050 17.330 ;
        RECT 25.110 16.690 26.950 17.550 ;
        RECT 28.010 16.690 29.850 17.550 ;
        RECT 30.910 16.690 32.750 17.550 ;
        RECT 33.810 16.690 35.650 17.550 ;
        RECT 36.710 16.690 38.550 17.550 ;
        RECT 39.610 16.690 41.450 17.550 ;
        RECT 42.510 16.690 44.350 17.550 ;
        RECT 45.410 16.690 46.260 17.550 ;
        RECT 23.200 16.270 46.260 16.690 ;
        RECT 0.000 16.200 46.260 16.270 ;
        RECT 0.000 15.340 0.850 16.200 ;
        RECT 1.910 15.340 3.750 16.200 ;
        RECT 4.810 15.340 6.650 16.200 ;
        RECT 7.710 15.340 9.550 16.200 ;
        RECT 10.610 15.340 12.450 16.200 ;
        RECT 13.510 15.340 15.350 16.200 ;
        RECT 16.410 15.340 18.250 16.200 ;
        RECT 19.310 15.340 21.150 16.200 ;
        RECT 22.210 16.050 23.060 16.200 ;
        RECT 23.200 16.050 24.050 16.200 ;
        RECT 22.210 15.980 24.050 16.050 ;
        RECT 22.210 15.340 23.060 15.980 ;
        RECT 0.000 14.920 23.060 15.340 ;
        RECT 23.200 15.340 24.050 15.980 ;
        RECT 25.110 15.340 26.950 16.200 ;
        RECT 28.010 15.340 29.850 16.200 ;
        RECT 30.910 15.340 32.750 16.200 ;
        RECT 33.810 15.340 35.650 16.200 ;
        RECT 36.710 15.340 38.550 16.200 ;
        RECT 39.610 15.340 41.450 16.200 ;
        RECT 42.510 15.340 44.350 16.200 ;
        RECT 45.410 15.340 46.260 16.200 ;
        RECT 23.200 14.920 46.260 15.340 ;
        RECT 0.000 14.850 46.260 14.920 ;
        RECT 0.000 13.990 0.850 14.850 ;
        RECT 1.910 13.990 3.750 14.850 ;
        RECT 4.810 13.990 6.650 14.850 ;
        RECT 7.710 13.990 9.550 14.850 ;
        RECT 10.610 13.990 12.450 14.850 ;
        RECT 13.510 13.990 15.350 14.850 ;
        RECT 16.410 13.990 18.250 14.850 ;
        RECT 19.310 13.990 21.150 14.850 ;
        RECT 22.210 14.700 23.060 14.850 ;
        RECT 23.200 14.700 24.050 14.850 ;
        RECT 22.210 14.630 24.050 14.700 ;
        RECT 22.210 13.990 23.060 14.630 ;
        RECT 0.000 13.570 23.060 13.990 ;
        RECT 23.200 13.990 24.050 14.630 ;
        RECT 25.110 13.990 26.950 14.850 ;
        RECT 28.010 13.990 29.850 14.850 ;
        RECT 30.910 13.990 32.750 14.850 ;
        RECT 33.810 13.990 35.650 14.850 ;
        RECT 36.710 13.990 38.550 14.850 ;
        RECT 39.610 13.990 41.450 14.850 ;
        RECT 42.510 13.990 44.350 14.850 ;
        RECT 45.410 13.990 46.260 14.850 ;
        RECT 23.200 13.570 46.260 13.990 ;
        RECT 0.000 13.500 46.260 13.570 ;
        RECT 0.000 12.640 0.850 13.500 ;
        RECT 1.910 12.640 3.750 13.500 ;
        RECT 4.810 12.640 6.650 13.500 ;
        RECT 7.710 12.640 9.550 13.500 ;
        RECT 10.610 12.640 12.450 13.500 ;
        RECT 13.510 12.640 15.350 13.500 ;
        RECT 16.410 12.640 18.250 13.500 ;
        RECT 19.310 12.640 21.150 13.500 ;
        RECT 22.210 13.350 23.060 13.500 ;
        RECT 23.200 13.350 24.050 13.500 ;
        RECT 22.210 13.280 24.050 13.350 ;
        RECT 22.210 12.640 23.060 13.280 ;
        RECT 0.000 12.220 23.060 12.640 ;
        RECT 23.200 12.640 24.050 13.280 ;
        RECT 25.110 12.640 26.950 13.500 ;
        RECT 28.010 12.640 29.850 13.500 ;
        RECT 30.910 12.640 32.750 13.500 ;
        RECT 33.810 12.640 35.650 13.500 ;
        RECT 36.710 12.640 38.550 13.500 ;
        RECT 39.610 12.640 41.450 13.500 ;
        RECT 42.510 12.640 44.350 13.500 ;
        RECT 45.410 12.640 46.260 13.500 ;
        RECT 23.200 12.220 46.260 12.640 ;
        RECT 0.000 12.150 46.260 12.220 ;
        RECT 0.000 11.290 0.850 12.150 ;
        RECT 1.910 11.290 3.750 12.150 ;
        RECT 4.810 11.290 6.650 12.150 ;
        RECT 7.710 11.290 9.550 12.150 ;
        RECT 10.610 11.290 12.450 12.150 ;
        RECT 13.510 11.290 15.350 12.150 ;
        RECT 16.410 11.290 18.250 12.150 ;
        RECT 19.310 11.290 21.150 12.150 ;
        RECT 22.210 12.000 23.060 12.150 ;
        RECT 23.200 12.000 24.050 12.150 ;
        RECT 22.210 11.930 24.050 12.000 ;
        RECT 22.210 11.290 23.060 11.930 ;
        RECT 0.000 10.870 23.060 11.290 ;
        RECT 23.200 11.290 24.050 11.930 ;
        RECT 25.110 11.290 26.950 12.150 ;
        RECT 28.010 11.290 29.850 12.150 ;
        RECT 30.910 11.290 32.750 12.150 ;
        RECT 33.810 11.290 35.650 12.150 ;
        RECT 36.710 11.290 38.550 12.150 ;
        RECT 39.610 11.290 41.450 12.150 ;
        RECT 42.510 11.290 44.350 12.150 ;
        RECT 45.410 11.290 46.260 12.150 ;
        RECT 23.200 10.870 46.260 11.290 ;
        RECT 0.000 10.800 46.260 10.870 ;
        RECT 0.000 9.940 0.850 10.800 ;
        RECT 1.910 9.940 3.750 10.800 ;
        RECT 4.810 9.940 6.650 10.800 ;
        RECT 7.710 9.940 9.550 10.800 ;
        RECT 10.610 9.940 12.450 10.800 ;
        RECT 13.510 9.940 15.350 10.800 ;
        RECT 16.410 9.940 18.250 10.800 ;
        RECT 19.310 9.940 21.150 10.800 ;
        RECT 22.210 10.650 23.060 10.800 ;
        RECT 23.200 10.650 24.050 10.800 ;
        RECT 22.210 10.580 24.050 10.650 ;
        RECT 22.210 9.940 23.060 10.580 ;
        RECT 0.000 9.520 23.060 9.940 ;
        RECT 23.200 9.940 24.050 10.580 ;
        RECT 25.110 9.940 26.950 10.800 ;
        RECT 28.010 9.940 29.850 10.800 ;
        RECT 30.910 9.940 32.750 10.800 ;
        RECT 33.810 9.940 35.650 10.800 ;
        RECT 36.710 9.940 38.550 10.800 ;
        RECT 39.610 9.940 41.450 10.800 ;
        RECT 42.510 9.940 44.350 10.800 ;
        RECT 45.410 9.940 46.260 10.800 ;
        RECT 23.200 9.520 46.260 9.940 ;
        RECT 0.000 9.450 46.260 9.520 ;
        RECT 0.000 8.590 0.850 9.450 ;
        RECT 1.910 8.590 3.750 9.450 ;
        RECT 4.810 8.590 6.650 9.450 ;
        RECT 7.710 8.590 9.550 9.450 ;
        RECT 10.610 8.590 12.450 9.450 ;
        RECT 13.510 8.590 15.350 9.450 ;
        RECT 16.410 8.590 18.250 9.450 ;
        RECT 19.310 8.590 21.150 9.450 ;
        RECT 22.210 9.300 23.060 9.450 ;
        RECT 23.200 9.300 24.050 9.450 ;
        RECT 22.210 9.230 24.050 9.300 ;
        RECT 22.210 8.590 23.060 9.230 ;
        RECT 0.000 8.170 23.060 8.590 ;
        RECT 23.200 8.590 24.050 9.230 ;
        RECT 25.110 8.590 26.950 9.450 ;
        RECT 28.010 8.590 29.850 9.450 ;
        RECT 30.910 8.590 32.750 9.450 ;
        RECT 33.810 8.590 35.650 9.450 ;
        RECT 36.710 8.590 38.550 9.450 ;
        RECT 39.610 8.590 41.450 9.450 ;
        RECT 42.510 8.590 44.350 9.450 ;
        RECT 45.410 8.590 46.260 9.450 ;
        RECT 23.200 8.170 46.260 8.590 ;
        RECT 0.000 8.100 46.260 8.170 ;
        RECT 0.000 7.240 0.850 8.100 ;
        RECT 1.910 7.240 3.750 8.100 ;
        RECT 4.810 7.240 6.650 8.100 ;
        RECT 7.710 7.240 9.550 8.100 ;
        RECT 10.610 7.240 12.450 8.100 ;
        RECT 13.510 7.240 15.350 8.100 ;
        RECT 16.410 7.240 18.250 8.100 ;
        RECT 19.310 7.240 21.150 8.100 ;
        RECT 22.210 7.950 23.060 8.100 ;
        RECT 23.200 7.950 24.050 8.100 ;
        RECT 22.210 7.880 24.050 7.950 ;
        RECT 22.210 7.240 23.060 7.880 ;
        RECT 0.000 6.820 23.060 7.240 ;
        RECT 23.200 7.240 24.050 7.880 ;
        RECT 25.110 7.240 26.950 8.100 ;
        RECT 28.010 7.240 29.850 8.100 ;
        RECT 30.910 7.240 32.750 8.100 ;
        RECT 33.810 7.240 35.650 8.100 ;
        RECT 36.710 7.240 38.550 8.100 ;
        RECT 39.610 7.240 41.450 8.100 ;
        RECT 42.510 7.240 44.350 8.100 ;
        RECT 45.410 7.240 46.260 8.100 ;
        RECT 23.200 6.820 46.260 7.240 ;
        RECT 0.000 6.750 46.260 6.820 ;
        RECT 0.000 5.890 0.850 6.750 ;
        RECT 1.910 5.890 3.750 6.750 ;
        RECT 4.810 5.890 6.650 6.750 ;
        RECT 7.710 5.890 9.550 6.750 ;
        RECT 10.610 5.890 12.450 6.750 ;
        RECT 13.510 5.890 15.350 6.750 ;
        RECT 16.410 5.890 18.250 6.750 ;
        RECT 19.310 5.890 21.150 6.750 ;
        RECT 22.210 6.600 23.060 6.750 ;
        RECT 23.200 6.600 24.050 6.750 ;
        RECT 22.210 6.530 24.050 6.600 ;
        RECT 22.210 5.890 23.060 6.530 ;
        RECT 0.000 5.470 23.060 5.890 ;
        RECT 23.200 5.890 24.050 6.530 ;
        RECT 25.110 5.890 26.950 6.750 ;
        RECT 28.010 5.890 29.850 6.750 ;
        RECT 30.910 5.890 32.750 6.750 ;
        RECT 33.810 5.890 35.650 6.750 ;
        RECT 36.710 5.890 38.550 6.750 ;
        RECT 39.610 5.890 41.450 6.750 ;
        RECT 42.510 5.890 44.350 6.750 ;
        RECT 45.410 5.890 46.260 6.750 ;
        RECT 23.200 5.470 46.260 5.890 ;
        RECT 0.000 5.400 46.260 5.470 ;
        RECT 0.000 4.540 0.850 5.400 ;
        RECT 1.910 4.540 3.750 5.400 ;
        RECT 4.810 4.540 6.650 5.400 ;
        RECT 7.710 4.540 9.550 5.400 ;
        RECT 10.610 4.540 12.450 5.400 ;
        RECT 13.510 4.540 15.350 5.400 ;
        RECT 16.410 4.540 18.250 5.400 ;
        RECT 19.310 4.540 21.150 5.400 ;
        RECT 22.210 5.250 23.060 5.400 ;
        RECT 23.200 5.250 24.050 5.400 ;
        RECT 22.210 5.180 24.050 5.250 ;
        RECT 22.210 4.540 23.060 5.180 ;
        RECT 0.000 4.120 23.060 4.540 ;
        RECT 23.200 4.540 24.050 5.180 ;
        RECT 25.110 4.540 26.950 5.400 ;
        RECT 28.010 4.540 29.850 5.400 ;
        RECT 30.910 4.540 32.750 5.400 ;
        RECT 33.810 4.540 35.650 5.400 ;
        RECT 36.710 4.540 38.550 5.400 ;
        RECT 39.610 4.540 41.450 5.400 ;
        RECT 42.510 4.540 44.350 5.400 ;
        RECT 45.410 4.540 46.260 5.400 ;
        RECT 23.200 4.120 46.260 4.540 ;
        RECT 0.000 4.050 46.260 4.120 ;
        RECT 0.000 3.190 0.850 4.050 ;
        RECT 1.910 3.190 3.750 4.050 ;
        RECT 4.810 3.190 6.650 4.050 ;
        RECT 7.710 3.190 9.550 4.050 ;
        RECT 10.610 3.190 12.450 4.050 ;
        RECT 13.510 3.190 15.350 4.050 ;
        RECT 16.410 3.190 18.250 4.050 ;
        RECT 19.310 3.190 21.150 4.050 ;
        RECT 22.210 3.900 23.060 4.050 ;
        RECT 23.200 3.900 24.050 4.050 ;
        RECT 22.210 3.830 24.050 3.900 ;
        RECT 22.210 3.190 23.060 3.830 ;
        RECT 0.000 2.770 23.060 3.190 ;
        RECT 23.200 3.190 24.050 3.830 ;
        RECT 25.110 3.190 26.950 4.050 ;
        RECT 28.010 3.190 29.850 4.050 ;
        RECT 30.910 3.190 32.750 4.050 ;
        RECT 33.810 3.190 35.650 4.050 ;
        RECT 36.710 3.190 38.550 4.050 ;
        RECT 39.610 3.190 41.450 4.050 ;
        RECT 42.510 3.190 44.350 4.050 ;
        RECT 45.410 3.190 46.260 4.050 ;
        RECT 23.200 2.770 46.260 3.190 ;
        RECT 0.000 2.700 46.260 2.770 ;
        RECT 0.000 1.840 0.850 2.700 ;
        RECT 1.910 1.840 3.750 2.700 ;
        RECT 4.810 1.840 6.650 2.700 ;
        RECT 7.710 1.840 9.550 2.700 ;
        RECT 10.610 1.840 12.450 2.700 ;
        RECT 13.510 1.840 15.350 2.700 ;
        RECT 16.410 1.840 18.250 2.700 ;
        RECT 19.310 1.840 21.150 2.700 ;
        RECT 22.210 2.550 23.060 2.700 ;
        RECT 23.200 2.550 24.050 2.700 ;
        RECT 22.210 2.480 24.050 2.550 ;
        RECT 22.210 1.840 23.060 2.480 ;
        RECT 0.000 1.420 23.060 1.840 ;
        RECT 23.200 1.845 24.050 2.480 ;
        RECT 25.110 1.845 26.950 2.700 ;
        RECT 28.010 1.845 29.850 2.700 ;
        RECT 30.910 1.845 32.750 2.700 ;
        RECT 33.810 1.845 35.650 2.700 ;
        RECT 36.710 1.845 38.550 2.700 ;
        RECT 39.610 1.845 41.450 2.700 ;
        RECT 42.510 1.845 44.350 2.700 ;
        RECT 45.410 1.845 46.260 2.700 ;
        RECT 23.200 1.420 46.260 1.845 ;
        RECT 0.000 1.355 46.260 1.420 ;
        RECT 0.000 1.350 24.050 1.355 ;
        RECT 0.000 0.490 0.850 1.350 ;
        RECT 1.910 0.490 3.750 1.350 ;
        RECT 4.810 0.490 6.650 1.350 ;
        RECT 7.710 0.490 9.550 1.350 ;
        RECT 10.610 0.490 12.450 1.350 ;
        RECT 13.510 0.490 15.350 1.350 ;
        RECT 16.410 0.490 18.250 1.350 ;
        RECT 19.310 0.490 21.150 1.350 ;
        RECT 22.210 1.200 23.060 1.350 ;
        RECT 23.200 1.200 24.050 1.350 ;
        RECT 22.210 1.130 24.050 1.200 ;
        RECT 22.210 0.490 23.060 1.130 ;
        RECT 0.000 0.070 23.060 0.490 ;
        RECT 23.200 0.495 24.050 1.130 ;
        RECT 25.110 0.495 26.950 1.355 ;
        RECT 28.010 0.495 29.850 1.355 ;
        RECT 30.910 0.495 32.750 1.355 ;
        RECT 33.810 0.495 35.650 1.355 ;
        RECT 36.710 0.495 38.550 1.355 ;
        RECT 39.610 0.495 41.450 1.355 ;
        RECT 42.510 0.495 44.350 1.355 ;
        RECT 45.410 0.495 46.260 1.355 ;
        RECT 23.200 0.070 46.260 0.495 ;
        RECT 0.000 0.005 46.260 0.070 ;
        RECT 46.400 42.340 47.250 43.200 ;
        RECT 48.310 42.340 50.150 43.200 ;
        RECT 51.210 42.340 53.050 43.200 ;
        RECT 54.110 42.340 55.950 43.200 ;
        RECT 57.010 42.340 58.850 43.200 ;
        RECT 59.910 42.340 61.750 43.200 ;
        RECT 62.810 42.340 64.650 43.200 ;
        RECT 65.710 42.340 67.550 43.200 ;
        RECT 68.610 42.340 69.460 43.200 ;
        RECT 46.400 41.850 69.460 42.340 ;
        RECT 46.400 40.990 47.250 41.850 ;
        RECT 48.310 40.990 50.150 41.850 ;
        RECT 51.210 40.990 53.050 41.850 ;
        RECT 54.110 40.990 55.950 41.850 ;
        RECT 57.010 40.990 58.850 41.850 ;
        RECT 59.910 40.990 61.750 41.850 ;
        RECT 62.810 40.990 64.650 41.850 ;
        RECT 65.710 40.990 67.550 41.850 ;
        RECT 68.610 40.990 69.460 41.850 ;
        RECT 46.400 40.500 69.460 40.990 ;
        RECT 46.400 39.640 47.250 40.500 ;
        RECT 48.310 39.640 50.150 40.500 ;
        RECT 51.210 39.640 53.050 40.500 ;
        RECT 54.110 39.640 55.950 40.500 ;
        RECT 57.010 39.640 58.850 40.500 ;
        RECT 59.910 39.640 61.750 40.500 ;
        RECT 62.810 39.640 64.650 40.500 ;
        RECT 65.710 39.640 67.550 40.500 ;
        RECT 68.610 39.640 69.460 40.500 ;
        RECT 46.400 39.150 69.460 39.640 ;
        RECT 46.400 38.290 47.250 39.150 ;
        RECT 48.310 38.290 50.150 39.150 ;
        RECT 51.210 38.290 53.050 39.150 ;
        RECT 54.110 38.290 55.950 39.150 ;
        RECT 57.010 38.290 58.850 39.150 ;
        RECT 59.910 38.290 61.750 39.150 ;
        RECT 62.810 38.290 64.650 39.150 ;
        RECT 65.710 38.290 67.550 39.150 ;
        RECT 68.610 38.290 69.460 39.150 ;
        RECT 46.400 37.800 69.460 38.290 ;
        RECT 46.400 36.940 47.250 37.800 ;
        RECT 48.310 36.940 50.150 37.800 ;
        RECT 51.210 36.940 53.050 37.800 ;
        RECT 54.110 36.940 55.950 37.800 ;
        RECT 57.010 36.940 58.850 37.800 ;
        RECT 59.910 36.940 61.750 37.800 ;
        RECT 62.810 36.940 64.650 37.800 ;
        RECT 65.710 36.940 67.550 37.800 ;
        RECT 68.610 36.940 69.460 37.800 ;
        RECT 46.400 36.450 69.460 36.940 ;
        RECT 46.400 35.590 47.250 36.450 ;
        RECT 48.310 35.590 50.150 36.450 ;
        RECT 51.210 35.590 53.050 36.450 ;
        RECT 54.110 35.590 55.950 36.450 ;
        RECT 57.010 35.590 58.850 36.450 ;
        RECT 59.910 35.590 61.750 36.450 ;
        RECT 62.810 35.590 64.650 36.450 ;
        RECT 65.710 35.590 67.550 36.450 ;
        RECT 68.610 35.590 69.460 36.450 ;
        RECT 46.400 35.100 69.460 35.590 ;
        RECT 46.400 34.240 47.250 35.100 ;
        RECT 48.310 34.240 50.150 35.100 ;
        RECT 51.210 34.240 53.050 35.100 ;
        RECT 54.110 34.240 55.950 35.100 ;
        RECT 57.010 34.240 58.850 35.100 ;
        RECT 59.910 34.240 61.750 35.100 ;
        RECT 62.810 34.240 64.650 35.100 ;
        RECT 65.710 34.240 67.550 35.100 ;
        RECT 68.610 34.240 69.460 35.100 ;
        RECT 46.400 33.750 69.460 34.240 ;
        RECT 46.400 32.890 47.250 33.750 ;
        RECT 48.310 32.890 50.150 33.750 ;
        RECT 51.210 32.890 53.050 33.750 ;
        RECT 54.110 32.890 55.950 33.750 ;
        RECT 57.010 32.890 58.850 33.750 ;
        RECT 59.910 32.890 61.750 33.750 ;
        RECT 62.810 32.890 64.650 33.750 ;
        RECT 65.710 32.890 67.550 33.750 ;
        RECT 68.610 32.890 69.460 33.750 ;
        RECT 46.400 32.400 69.460 32.890 ;
        RECT 46.400 31.540 47.250 32.400 ;
        RECT 48.310 31.540 50.150 32.400 ;
        RECT 51.210 31.540 53.050 32.400 ;
        RECT 54.110 31.540 55.950 32.400 ;
        RECT 57.010 31.540 58.850 32.400 ;
        RECT 59.910 31.540 61.750 32.400 ;
        RECT 62.810 31.540 64.650 32.400 ;
        RECT 65.710 31.540 67.550 32.400 ;
        RECT 68.610 31.540 69.460 32.400 ;
        RECT 46.400 31.050 69.460 31.540 ;
        RECT 46.400 30.190 47.250 31.050 ;
        RECT 48.310 30.190 50.150 31.050 ;
        RECT 51.210 30.190 53.050 31.050 ;
        RECT 54.110 30.190 55.950 31.050 ;
        RECT 57.010 30.190 58.850 31.050 ;
        RECT 59.910 30.190 61.750 31.050 ;
        RECT 62.810 30.190 64.650 31.050 ;
        RECT 65.710 30.190 67.550 31.050 ;
        RECT 68.610 30.190 69.460 31.050 ;
        RECT 46.400 29.700 69.460 30.190 ;
        RECT 46.400 28.840 47.250 29.700 ;
        RECT 48.310 28.840 50.150 29.700 ;
        RECT 51.210 28.840 53.050 29.700 ;
        RECT 54.110 28.840 55.950 29.700 ;
        RECT 57.010 28.840 58.850 29.700 ;
        RECT 59.910 28.840 61.750 29.700 ;
        RECT 62.810 28.840 64.650 29.700 ;
        RECT 65.710 28.840 67.550 29.700 ;
        RECT 68.610 28.840 69.460 29.700 ;
        RECT 46.400 28.350 69.460 28.840 ;
        RECT 46.400 27.490 47.250 28.350 ;
        RECT 48.310 27.490 50.150 28.350 ;
        RECT 51.210 27.490 53.050 28.350 ;
        RECT 54.110 27.490 55.950 28.350 ;
        RECT 57.010 27.490 58.850 28.350 ;
        RECT 59.910 27.490 61.750 28.350 ;
        RECT 62.810 27.490 64.650 28.350 ;
        RECT 65.710 27.490 67.550 28.350 ;
        RECT 68.610 27.490 69.460 28.350 ;
        RECT 46.400 27.000 69.460 27.490 ;
        RECT 46.400 26.140 47.250 27.000 ;
        RECT 48.310 26.140 50.150 27.000 ;
        RECT 51.210 26.140 53.050 27.000 ;
        RECT 54.110 26.140 55.950 27.000 ;
        RECT 57.010 26.140 58.850 27.000 ;
        RECT 59.910 26.140 61.750 27.000 ;
        RECT 62.810 26.140 64.650 27.000 ;
        RECT 65.710 26.140 67.550 27.000 ;
        RECT 68.610 26.140 69.460 27.000 ;
        RECT 46.400 25.650 69.460 26.140 ;
        RECT 46.400 24.790 47.250 25.650 ;
        RECT 48.310 24.790 50.150 25.650 ;
        RECT 51.210 24.790 53.050 25.650 ;
        RECT 54.110 24.790 55.950 25.650 ;
        RECT 57.010 24.790 58.850 25.650 ;
        RECT 59.910 24.790 61.750 25.650 ;
        RECT 62.810 24.790 64.650 25.650 ;
        RECT 65.710 24.790 67.550 25.650 ;
        RECT 68.610 24.790 69.460 25.650 ;
        RECT 46.400 24.300 69.460 24.790 ;
        RECT 46.400 23.440 47.250 24.300 ;
        RECT 48.310 23.440 50.150 24.300 ;
        RECT 51.210 23.440 53.050 24.300 ;
        RECT 54.110 23.440 55.950 24.300 ;
        RECT 57.010 23.440 58.850 24.300 ;
        RECT 59.910 23.440 61.750 24.300 ;
        RECT 62.810 23.440 64.650 24.300 ;
        RECT 65.710 23.440 67.550 24.300 ;
        RECT 68.610 23.440 69.460 24.300 ;
        RECT 46.400 22.950 69.460 23.440 ;
        RECT 46.400 22.090 47.250 22.950 ;
        RECT 48.310 22.090 50.150 22.950 ;
        RECT 51.210 22.090 53.050 22.950 ;
        RECT 54.110 22.090 55.950 22.950 ;
        RECT 57.010 22.090 58.850 22.950 ;
        RECT 59.910 22.090 61.750 22.950 ;
        RECT 62.810 22.090 64.650 22.950 ;
        RECT 65.710 22.090 67.550 22.950 ;
        RECT 68.610 22.090 69.460 22.950 ;
        RECT 46.400 21.600 69.460 22.090 ;
        RECT 46.400 20.740 47.250 21.600 ;
        RECT 48.310 20.740 50.150 21.600 ;
        RECT 51.210 20.740 53.050 21.600 ;
        RECT 54.110 20.740 55.950 21.600 ;
        RECT 57.010 20.740 58.850 21.600 ;
        RECT 59.910 20.740 61.750 21.600 ;
        RECT 62.810 20.740 64.650 21.600 ;
        RECT 65.710 20.740 67.550 21.600 ;
        RECT 68.610 20.740 69.460 21.600 ;
        RECT 46.400 20.250 69.460 20.740 ;
        RECT 46.400 19.390 47.250 20.250 ;
        RECT 48.310 19.390 50.150 20.250 ;
        RECT 51.210 19.390 53.050 20.250 ;
        RECT 54.110 19.390 55.950 20.250 ;
        RECT 57.010 19.390 58.850 20.250 ;
        RECT 59.910 19.390 61.750 20.250 ;
        RECT 62.810 19.390 64.650 20.250 ;
        RECT 65.710 19.390 67.550 20.250 ;
        RECT 68.610 19.390 69.460 20.250 ;
        RECT 46.400 18.900 69.460 19.390 ;
        RECT 46.400 18.040 47.250 18.900 ;
        RECT 48.310 18.040 50.150 18.900 ;
        RECT 51.210 18.040 53.050 18.900 ;
        RECT 54.110 18.040 55.950 18.900 ;
        RECT 57.010 18.040 58.850 18.900 ;
        RECT 59.910 18.040 61.750 18.900 ;
        RECT 62.810 18.040 64.650 18.900 ;
        RECT 65.710 18.040 67.550 18.900 ;
        RECT 68.610 18.040 69.460 18.900 ;
        RECT 46.400 17.550 69.460 18.040 ;
        RECT 46.400 16.690 47.250 17.550 ;
        RECT 48.310 16.690 50.150 17.550 ;
        RECT 51.210 16.690 53.050 17.550 ;
        RECT 54.110 16.690 55.950 17.550 ;
        RECT 57.010 16.690 58.850 17.550 ;
        RECT 59.910 16.690 61.750 17.550 ;
        RECT 62.810 16.690 64.650 17.550 ;
        RECT 65.710 16.690 67.550 17.550 ;
        RECT 68.610 16.690 69.460 17.550 ;
        RECT 46.400 16.200 69.460 16.690 ;
        RECT 46.400 15.340 47.250 16.200 ;
        RECT 48.310 15.340 50.150 16.200 ;
        RECT 51.210 15.340 53.050 16.200 ;
        RECT 54.110 15.340 55.950 16.200 ;
        RECT 57.010 15.340 58.850 16.200 ;
        RECT 59.910 15.340 61.750 16.200 ;
        RECT 62.810 15.340 64.650 16.200 ;
        RECT 65.710 15.340 67.550 16.200 ;
        RECT 68.610 15.340 69.460 16.200 ;
        RECT 46.400 14.850 69.460 15.340 ;
        RECT 46.400 13.990 47.250 14.850 ;
        RECT 48.310 13.990 50.150 14.850 ;
        RECT 51.210 13.990 53.050 14.850 ;
        RECT 54.110 13.990 55.950 14.850 ;
        RECT 57.010 13.990 58.850 14.850 ;
        RECT 59.910 13.990 61.750 14.850 ;
        RECT 62.810 13.990 64.650 14.850 ;
        RECT 65.710 13.990 67.550 14.850 ;
        RECT 68.610 13.990 69.460 14.850 ;
        RECT 46.400 13.500 69.460 13.990 ;
        RECT 46.400 12.640 47.250 13.500 ;
        RECT 48.310 12.640 50.150 13.500 ;
        RECT 51.210 12.640 53.050 13.500 ;
        RECT 54.110 12.640 55.950 13.500 ;
        RECT 57.010 12.640 58.850 13.500 ;
        RECT 59.910 12.640 61.750 13.500 ;
        RECT 62.810 12.640 64.650 13.500 ;
        RECT 65.710 12.640 67.550 13.500 ;
        RECT 68.610 12.640 69.460 13.500 ;
        RECT 46.400 12.150 69.460 12.640 ;
        RECT 46.400 11.290 47.250 12.150 ;
        RECT 48.310 11.290 50.150 12.150 ;
        RECT 51.210 11.290 53.050 12.150 ;
        RECT 54.110 11.290 55.950 12.150 ;
        RECT 57.010 11.290 58.850 12.150 ;
        RECT 59.910 11.290 61.750 12.150 ;
        RECT 62.810 11.290 64.650 12.150 ;
        RECT 65.710 11.290 67.550 12.150 ;
        RECT 68.610 11.290 69.460 12.150 ;
        RECT 46.400 10.800 69.460 11.290 ;
        RECT 46.400 9.940 47.250 10.800 ;
        RECT 48.310 9.940 50.150 10.800 ;
        RECT 51.210 9.940 53.050 10.800 ;
        RECT 54.110 9.940 55.950 10.800 ;
        RECT 57.010 9.940 58.850 10.800 ;
        RECT 59.910 9.940 61.750 10.800 ;
        RECT 62.810 9.940 64.650 10.800 ;
        RECT 65.710 9.940 67.550 10.800 ;
        RECT 68.610 9.940 69.460 10.800 ;
        RECT 46.400 9.450 69.460 9.940 ;
        RECT 46.400 8.590 47.250 9.450 ;
        RECT 48.310 8.590 50.150 9.450 ;
        RECT 51.210 8.590 53.050 9.450 ;
        RECT 54.110 8.590 55.950 9.450 ;
        RECT 57.010 8.590 58.850 9.450 ;
        RECT 59.910 8.590 61.750 9.450 ;
        RECT 62.810 8.590 64.650 9.450 ;
        RECT 65.710 8.590 67.550 9.450 ;
        RECT 68.610 8.590 69.460 9.450 ;
        RECT 46.400 8.100 69.460 8.590 ;
        RECT 46.400 7.240 47.250 8.100 ;
        RECT 48.310 7.240 50.150 8.100 ;
        RECT 51.210 7.240 53.050 8.100 ;
        RECT 54.110 7.240 55.950 8.100 ;
        RECT 57.010 7.240 58.850 8.100 ;
        RECT 59.910 7.240 61.750 8.100 ;
        RECT 62.810 7.240 64.650 8.100 ;
        RECT 65.710 7.240 67.550 8.100 ;
        RECT 68.610 7.240 69.460 8.100 ;
        RECT 46.400 6.750 69.460 7.240 ;
        RECT 46.400 5.890 47.250 6.750 ;
        RECT 48.310 5.890 50.150 6.750 ;
        RECT 51.210 5.890 53.050 6.750 ;
        RECT 54.110 5.890 55.950 6.750 ;
        RECT 57.010 5.890 58.850 6.750 ;
        RECT 59.910 5.890 61.750 6.750 ;
        RECT 62.810 5.890 64.650 6.750 ;
        RECT 65.710 5.890 67.550 6.750 ;
        RECT 68.610 5.890 69.460 6.750 ;
        RECT 46.400 5.400 69.460 5.890 ;
        RECT 46.400 4.540 47.250 5.400 ;
        RECT 48.310 4.540 50.150 5.400 ;
        RECT 51.210 4.540 53.050 5.400 ;
        RECT 54.110 4.540 55.950 5.400 ;
        RECT 57.010 4.540 58.850 5.400 ;
        RECT 59.910 4.540 61.750 5.400 ;
        RECT 62.810 4.540 64.650 5.400 ;
        RECT 65.710 4.540 67.550 5.400 ;
        RECT 68.610 4.540 69.460 5.400 ;
        RECT 46.400 4.050 69.460 4.540 ;
        RECT 46.400 3.190 47.250 4.050 ;
        RECT 48.310 3.190 50.150 4.050 ;
        RECT 51.210 3.190 53.050 4.050 ;
        RECT 54.110 3.190 55.950 4.050 ;
        RECT 57.010 3.190 58.850 4.050 ;
        RECT 59.910 3.190 61.750 4.050 ;
        RECT 62.810 3.190 64.650 4.050 ;
        RECT 65.710 3.190 67.550 4.050 ;
        RECT 68.610 3.190 69.460 4.050 ;
        RECT 46.400 2.700 69.460 3.190 ;
        RECT 46.400 1.845 47.250 2.700 ;
        RECT 48.310 1.845 50.150 2.700 ;
        RECT 51.210 1.845 53.050 2.700 ;
        RECT 54.110 1.845 55.950 2.700 ;
        RECT 57.010 1.845 58.850 2.700 ;
        RECT 59.910 1.845 61.750 2.700 ;
        RECT 62.810 1.845 64.650 2.700 ;
        RECT 65.710 1.845 67.550 2.700 ;
        RECT 68.610 1.845 69.460 2.700 ;
        RECT 46.400 1.355 69.460 1.845 ;
        RECT 46.400 0.495 47.250 1.355 ;
        RECT 48.310 0.495 50.150 1.355 ;
        RECT 51.210 0.495 53.050 1.355 ;
        RECT 54.110 0.495 55.950 1.355 ;
        RECT 57.010 0.495 58.850 1.355 ;
        RECT 59.910 0.495 61.750 1.355 ;
        RECT 62.810 0.495 64.650 1.355 ;
        RECT 65.710 0.495 67.550 1.355 ;
        RECT 68.610 0.495 69.460 1.355 ;
        RECT 46.400 0.005 69.460 0.495 ;
        RECT 69.600 42.340 70.450 43.200 ;
        RECT 71.510 42.340 73.350 43.200 ;
        RECT 74.410 42.340 76.250 43.200 ;
        RECT 77.310 42.340 79.150 43.200 ;
        RECT 80.210 42.340 82.050 43.200 ;
        RECT 83.110 42.340 84.950 43.200 ;
        RECT 86.010 42.340 87.850 43.200 ;
        RECT 88.910 42.340 90.750 43.200 ;
        RECT 91.810 42.340 92.660 43.200 ;
        RECT 69.600 41.850 92.660 42.340 ;
        RECT 69.600 40.990 70.450 41.850 ;
        RECT 71.510 40.990 73.350 41.850 ;
        RECT 74.410 40.990 76.250 41.850 ;
        RECT 77.310 40.990 79.150 41.850 ;
        RECT 80.210 40.990 82.050 41.850 ;
        RECT 83.110 40.990 84.950 41.850 ;
        RECT 86.010 40.990 87.850 41.850 ;
        RECT 88.910 40.990 90.750 41.850 ;
        RECT 91.810 40.990 92.660 41.850 ;
        RECT 69.600 40.500 92.660 40.990 ;
        RECT 69.600 39.640 70.450 40.500 ;
        RECT 71.510 39.640 73.350 40.500 ;
        RECT 74.410 39.640 76.250 40.500 ;
        RECT 77.310 39.640 79.150 40.500 ;
        RECT 80.210 39.640 82.050 40.500 ;
        RECT 83.110 39.640 84.950 40.500 ;
        RECT 86.010 39.640 87.850 40.500 ;
        RECT 88.910 39.640 90.750 40.500 ;
        RECT 91.810 39.640 92.660 40.500 ;
        RECT 69.600 39.150 92.660 39.640 ;
        RECT 69.600 38.290 70.450 39.150 ;
        RECT 71.510 38.290 73.350 39.150 ;
        RECT 74.410 38.290 76.250 39.150 ;
        RECT 77.310 38.290 79.150 39.150 ;
        RECT 80.210 38.290 82.050 39.150 ;
        RECT 83.110 38.290 84.950 39.150 ;
        RECT 86.010 38.290 87.850 39.150 ;
        RECT 88.910 38.290 90.750 39.150 ;
        RECT 91.810 38.290 92.660 39.150 ;
        RECT 69.600 37.800 92.660 38.290 ;
        RECT 69.600 36.940 70.450 37.800 ;
        RECT 71.510 36.940 73.350 37.800 ;
        RECT 74.410 36.940 76.250 37.800 ;
        RECT 77.310 36.940 79.150 37.800 ;
        RECT 80.210 36.940 82.050 37.800 ;
        RECT 83.110 36.940 84.950 37.800 ;
        RECT 86.010 36.940 87.850 37.800 ;
        RECT 88.910 36.940 90.750 37.800 ;
        RECT 91.810 36.940 92.660 37.800 ;
        RECT 69.600 36.450 92.660 36.940 ;
        RECT 69.600 35.590 70.450 36.450 ;
        RECT 71.510 35.590 73.350 36.450 ;
        RECT 74.410 35.590 76.250 36.450 ;
        RECT 77.310 35.590 79.150 36.450 ;
        RECT 80.210 35.590 82.050 36.450 ;
        RECT 83.110 35.590 84.950 36.450 ;
        RECT 86.010 35.590 87.850 36.450 ;
        RECT 88.910 35.590 90.750 36.450 ;
        RECT 91.810 35.590 92.660 36.450 ;
        RECT 69.600 35.100 92.660 35.590 ;
        RECT 69.600 34.240 70.450 35.100 ;
        RECT 71.510 34.240 73.350 35.100 ;
        RECT 74.410 34.240 76.250 35.100 ;
        RECT 77.310 34.240 79.150 35.100 ;
        RECT 80.210 34.240 82.050 35.100 ;
        RECT 83.110 34.240 84.950 35.100 ;
        RECT 86.010 34.240 87.850 35.100 ;
        RECT 88.910 34.240 90.750 35.100 ;
        RECT 91.810 34.240 92.660 35.100 ;
        RECT 69.600 33.750 92.660 34.240 ;
        RECT 69.600 32.890 70.450 33.750 ;
        RECT 71.510 32.890 73.350 33.750 ;
        RECT 74.410 32.890 76.250 33.750 ;
        RECT 77.310 32.890 79.150 33.750 ;
        RECT 80.210 32.890 82.050 33.750 ;
        RECT 83.110 32.890 84.950 33.750 ;
        RECT 86.010 32.890 87.850 33.750 ;
        RECT 88.910 32.890 90.750 33.750 ;
        RECT 91.810 32.890 92.660 33.750 ;
        RECT 69.600 32.400 92.660 32.890 ;
        RECT 69.600 31.540 70.450 32.400 ;
        RECT 71.510 31.540 73.350 32.400 ;
        RECT 74.410 31.540 76.250 32.400 ;
        RECT 77.310 31.540 79.150 32.400 ;
        RECT 80.210 31.540 82.050 32.400 ;
        RECT 83.110 31.540 84.950 32.400 ;
        RECT 86.010 31.540 87.850 32.400 ;
        RECT 88.910 31.540 90.750 32.400 ;
        RECT 91.810 31.540 92.660 32.400 ;
        RECT 69.600 31.050 92.660 31.540 ;
        RECT 69.600 30.190 70.450 31.050 ;
        RECT 71.510 30.190 73.350 31.050 ;
        RECT 74.410 30.190 76.250 31.050 ;
        RECT 77.310 30.190 79.150 31.050 ;
        RECT 80.210 30.190 82.050 31.050 ;
        RECT 83.110 30.190 84.950 31.050 ;
        RECT 86.010 30.190 87.850 31.050 ;
        RECT 88.910 30.190 90.750 31.050 ;
        RECT 91.810 30.190 92.660 31.050 ;
        RECT 69.600 29.700 92.660 30.190 ;
        RECT 69.600 28.840 70.450 29.700 ;
        RECT 71.510 28.840 73.350 29.700 ;
        RECT 74.410 28.840 76.250 29.700 ;
        RECT 77.310 28.840 79.150 29.700 ;
        RECT 80.210 28.840 82.050 29.700 ;
        RECT 83.110 28.840 84.950 29.700 ;
        RECT 86.010 28.840 87.850 29.700 ;
        RECT 88.910 28.840 90.750 29.700 ;
        RECT 91.810 28.840 92.660 29.700 ;
        RECT 69.600 28.350 92.660 28.840 ;
        RECT 69.600 27.490 70.450 28.350 ;
        RECT 71.510 27.490 73.350 28.350 ;
        RECT 74.410 27.490 76.250 28.350 ;
        RECT 77.310 27.490 79.150 28.350 ;
        RECT 80.210 27.490 82.050 28.350 ;
        RECT 83.110 27.490 84.950 28.350 ;
        RECT 86.010 27.490 87.850 28.350 ;
        RECT 88.910 27.490 90.750 28.350 ;
        RECT 91.810 27.490 92.660 28.350 ;
        RECT 69.600 27.000 92.660 27.490 ;
        RECT 69.600 26.140 70.450 27.000 ;
        RECT 71.510 26.140 73.350 27.000 ;
        RECT 74.410 26.140 76.250 27.000 ;
        RECT 77.310 26.140 79.150 27.000 ;
        RECT 80.210 26.140 82.050 27.000 ;
        RECT 83.110 26.140 84.950 27.000 ;
        RECT 86.010 26.140 87.850 27.000 ;
        RECT 88.910 26.140 90.750 27.000 ;
        RECT 91.810 26.140 92.660 27.000 ;
        RECT 69.600 25.650 92.660 26.140 ;
        RECT 69.600 24.790 70.450 25.650 ;
        RECT 71.510 24.790 73.350 25.650 ;
        RECT 74.410 24.790 76.250 25.650 ;
        RECT 77.310 24.790 79.150 25.650 ;
        RECT 80.210 24.790 82.050 25.650 ;
        RECT 83.110 24.790 84.950 25.650 ;
        RECT 86.010 24.790 87.850 25.650 ;
        RECT 88.910 24.790 90.750 25.650 ;
        RECT 91.810 24.790 92.660 25.650 ;
        RECT 69.600 24.300 92.660 24.790 ;
        RECT 69.600 23.440 70.450 24.300 ;
        RECT 71.510 23.440 73.350 24.300 ;
        RECT 74.410 23.440 76.250 24.300 ;
        RECT 77.310 23.440 79.150 24.300 ;
        RECT 80.210 23.440 82.050 24.300 ;
        RECT 83.110 23.440 84.950 24.300 ;
        RECT 86.010 23.440 87.850 24.300 ;
        RECT 88.910 23.440 90.750 24.300 ;
        RECT 91.810 23.440 92.660 24.300 ;
        RECT 69.600 22.950 92.660 23.440 ;
        RECT 69.600 22.090 70.450 22.950 ;
        RECT 71.510 22.090 73.350 22.950 ;
        RECT 74.410 22.090 76.250 22.950 ;
        RECT 77.310 22.090 79.150 22.950 ;
        RECT 80.210 22.090 82.050 22.950 ;
        RECT 83.110 22.090 84.950 22.950 ;
        RECT 86.010 22.090 87.850 22.950 ;
        RECT 88.910 22.090 90.750 22.950 ;
        RECT 91.810 22.090 92.660 22.950 ;
        RECT 69.600 21.600 92.660 22.090 ;
        RECT 69.600 20.740 70.450 21.600 ;
        RECT 71.510 20.740 73.350 21.600 ;
        RECT 74.410 20.740 76.250 21.600 ;
        RECT 77.310 20.740 79.150 21.600 ;
        RECT 80.210 20.740 82.050 21.600 ;
        RECT 83.110 20.740 84.950 21.600 ;
        RECT 86.010 20.740 87.850 21.600 ;
        RECT 88.910 20.740 90.750 21.600 ;
        RECT 91.810 20.740 92.660 21.600 ;
        RECT 69.600 20.250 92.660 20.740 ;
        RECT 69.600 19.390 70.450 20.250 ;
        RECT 71.510 19.390 73.350 20.250 ;
        RECT 74.410 19.390 76.250 20.250 ;
        RECT 77.310 19.390 79.150 20.250 ;
        RECT 80.210 19.390 82.050 20.250 ;
        RECT 83.110 19.390 84.950 20.250 ;
        RECT 86.010 19.390 87.850 20.250 ;
        RECT 88.910 19.390 90.750 20.250 ;
        RECT 91.810 19.390 92.660 20.250 ;
        RECT 69.600 18.900 92.660 19.390 ;
        RECT 69.600 18.040 70.450 18.900 ;
        RECT 71.510 18.040 73.350 18.900 ;
        RECT 74.410 18.040 76.250 18.900 ;
        RECT 77.310 18.040 79.150 18.900 ;
        RECT 80.210 18.040 82.050 18.900 ;
        RECT 83.110 18.040 84.950 18.900 ;
        RECT 86.010 18.040 87.850 18.900 ;
        RECT 88.910 18.040 90.750 18.900 ;
        RECT 91.810 18.040 92.660 18.900 ;
        RECT 69.600 17.550 92.660 18.040 ;
        RECT 69.600 16.690 70.450 17.550 ;
        RECT 71.510 16.690 73.350 17.550 ;
        RECT 74.410 16.690 76.250 17.550 ;
        RECT 77.310 16.690 79.150 17.550 ;
        RECT 80.210 16.690 82.050 17.550 ;
        RECT 83.110 16.690 84.950 17.550 ;
        RECT 86.010 16.690 87.850 17.550 ;
        RECT 88.910 16.690 90.750 17.550 ;
        RECT 91.810 16.690 92.660 17.550 ;
        RECT 69.600 16.200 92.660 16.690 ;
        RECT 69.600 15.340 70.450 16.200 ;
        RECT 71.510 15.340 73.350 16.200 ;
        RECT 74.410 15.340 76.250 16.200 ;
        RECT 77.310 15.340 79.150 16.200 ;
        RECT 80.210 15.340 82.050 16.200 ;
        RECT 83.110 15.340 84.950 16.200 ;
        RECT 86.010 15.340 87.850 16.200 ;
        RECT 88.910 15.340 90.750 16.200 ;
        RECT 91.810 15.340 92.660 16.200 ;
        RECT 69.600 14.850 92.660 15.340 ;
        RECT 69.600 13.990 70.450 14.850 ;
        RECT 71.510 13.990 73.350 14.850 ;
        RECT 74.410 13.990 76.250 14.850 ;
        RECT 77.310 13.990 79.150 14.850 ;
        RECT 80.210 13.990 82.050 14.850 ;
        RECT 83.110 13.990 84.950 14.850 ;
        RECT 86.010 13.990 87.850 14.850 ;
        RECT 88.910 13.990 90.750 14.850 ;
        RECT 91.810 13.990 92.660 14.850 ;
        RECT 69.600 13.500 92.660 13.990 ;
        RECT 69.600 12.640 70.450 13.500 ;
        RECT 71.510 12.640 73.350 13.500 ;
        RECT 74.410 12.640 76.250 13.500 ;
        RECT 77.310 12.640 79.150 13.500 ;
        RECT 80.210 12.640 82.050 13.500 ;
        RECT 83.110 12.640 84.950 13.500 ;
        RECT 86.010 12.640 87.850 13.500 ;
        RECT 88.910 12.640 90.750 13.500 ;
        RECT 91.810 12.640 92.660 13.500 ;
        RECT 69.600 12.150 92.660 12.640 ;
        RECT 69.600 11.290 70.450 12.150 ;
        RECT 71.510 11.290 73.350 12.150 ;
        RECT 74.410 11.290 76.250 12.150 ;
        RECT 77.310 11.290 79.150 12.150 ;
        RECT 80.210 11.290 82.050 12.150 ;
        RECT 83.110 11.290 84.950 12.150 ;
        RECT 86.010 11.290 87.850 12.150 ;
        RECT 88.910 11.290 90.750 12.150 ;
        RECT 91.810 11.290 92.660 12.150 ;
        RECT 69.600 10.800 92.660 11.290 ;
        RECT 69.600 9.940 70.450 10.800 ;
        RECT 71.510 9.940 73.350 10.800 ;
        RECT 74.410 9.940 76.250 10.800 ;
        RECT 77.310 9.940 79.150 10.800 ;
        RECT 80.210 9.940 82.050 10.800 ;
        RECT 83.110 9.940 84.950 10.800 ;
        RECT 86.010 9.940 87.850 10.800 ;
        RECT 88.910 9.940 90.750 10.800 ;
        RECT 91.810 9.940 92.660 10.800 ;
        RECT 69.600 9.450 92.660 9.940 ;
        RECT 69.600 8.590 70.450 9.450 ;
        RECT 71.510 8.590 73.350 9.450 ;
        RECT 74.410 8.590 76.250 9.450 ;
        RECT 77.310 8.590 79.150 9.450 ;
        RECT 80.210 8.590 82.050 9.450 ;
        RECT 83.110 8.590 84.950 9.450 ;
        RECT 86.010 8.590 87.850 9.450 ;
        RECT 88.910 8.590 90.750 9.450 ;
        RECT 91.810 8.590 92.660 9.450 ;
        RECT 69.600 8.100 92.660 8.590 ;
        RECT 69.600 7.240 70.450 8.100 ;
        RECT 71.510 7.240 73.350 8.100 ;
        RECT 74.410 7.240 76.250 8.100 ;
        RECT 77.310 7.240 79.150 8.100 ;
        RECT 80.210 7.240 82.050 8.100 ;
        RECT 83.110 7.240 84.950 8.100 ;
        RECT 86.010 7.240 87.850 8.100 ;
        RECT 88.910 7.240 90.750 8.100 ;
        RECT 91.810 7.240 92.660 8.100 ;
        RECT 69.600 6.750 92.660 7.240 ;
        RECT 69.600 5.890 70.450 6.750 ;
        RECT 71.510 5.890 73.350 6.750 ;
        RECT 74.410 5.890 76.250 6.750 ;
        RECT 77.310 5.890 79.150 6.750 ;
        RECT 80.210 5.890 82.050 6.750 ;
        RECT 83.110 5.890 84.950 6.750 ;
        RECT 86.010 5.890 87.850 6.750 ;
        RECT 88.910 5.890 90.750 6.750 ;
        RECT 91.810 5.890 92.660 6.750 ;
        RECT 69.600 5.400 92.660 5.890 ;
        RECT 69.600 4.540 70.450 5.400 ;
        RECT 71.510 4.540 73.350 5.400 ;
        RECT 74.410 4.540 76.250 5.400 ;
        RECT 77.310 4.540 79.150 5.400 ;
        RECT 80.210 4.540 82.050 5.400 ;
        RECT 83.110 4.540 84.950 5.400 ;
        RECT 86.010 4.540 87.850 5.400 ;
        RECT 88.910 4.540 90.750 5.400 ;
        RECT 91.810 4.540 92.660 5.400 ;
        RECT 69.600 4.050 92.660 4.540 ;
        RECT 69.600 3.190 70.450 4.050 ;
        RECT 71.510 3.190 73.350 4.050 ;
        RECT 74.410 3.190 76.250 4.050 ;
        RECT 77.310 3.190 79.150 4.050 ;
        RECT 80.210 3.190 82.050 4.050 ;
        RECT 83.110 3.190 84.950 4.050 ;
        RECT 86.010 3.190 87.850 4.050 ;
        RECT 88.910 3.190 90.750 4.050 ;
        RECT 91.810 3.190 92.660 4.050 ;
        RECT 69.600 2.700 92.660 3.190 ;
        RECT 69.600 1.845 70.450 2.700 ;
        RECT 71.510 1.845 73.350 2.700 ;
        RECT 74.410 1.845 76.250 2.700 ;
        RECT 77.310 1.845 79.150 2.700 ;
        RECT 80.210 1.845 82.050 2.700 ;
        RECT 83.110 1.845 84.950 2.700 ;
        RECT 86.010 1.845 87.850 2.700 ;
        RECT 88.910 1.845 90.750 2.700 ;
        RECT 91.810 1.845 92.660 2.700 ;
        RECT 69.600 1.355 92.660 1.845 ;
        RECT 69.600 0.495 70.450 1.355 ;
        RECT 71.510 0.495 73.350 1.355 ;
        RECT 74.410 0.495 76.250 1.355 ;
        RECT 77.310 0.495 79.150 1.355 ;
        RECT 80.210 0.495 82.050 1.355 ;
        RECT 83.110 0.495 84.950 1.355 ;
        RECT 86.010 0.495 87.850 1.355 ;
        RECT 88.910 0.495 90.750 1.355 ;
        RECT 91.810 0.495 92.660 1.355 ;
        RECT 69.600 0.005 92.660 0.495 ;
        RECT 0.000 0.000 23.200 0.005 ;
      LAYER li1 ;
        RECT 1.310 41.920 1.450 41.930 ;
        RECT 4.210 41.920 4.350 41.930 ;
        RECT 7.110 41.920 7.250 41.930 ;
        RECT 10.010 41.920 10.150 41.930 ;
        RECT 12.910 41.920 13.050 41.930 ;
        RECT 15.810 41.920 15.950 41.930 ;
        RECT 18.710 41.920 18.850 41.930 ;
        RECT 21.610 41.920 21.750 41.930 ;
        RECT 24.510 41.920 24.650 41.930 ;
        RECT 27.410 41.920 27.550 41.930 ;
        RECT 30.310 41.920 30.450 41.930 ;
        RECT 33.210 41.920 33.350 41.930 ;
        RECT 36.110 41.920 36.250 41.930 ;
        RECT 39.010 41.920 39.150 41.930 ;
        RECT 41.910 41.920 42.050 41.930 ;
        RECT 44.810 41.920 44.950 41.930 ;
        RECT 47.710 41.920 47.850 41.930 ;
        RECT 50.610 41.920 50.750 41.930 ;
        RECT 53.510 41.920 53.650 41.930 ;
        RECT 56.410 41.920 56.550 41.930 ;
        RECT 59.310 41.920 59.450 41.930 ;
        RECT 62.210 41.920 62.350 41.930 ;
        RECT 65.110 41.920 65.250 41.930 ;
        RECT 68.010 41.920 68.150 41.930 ;
        RECT 70.910 41.920 71.050 41.930 ;
        RECT 73.810 41.920 73.950 41.930 ;
        RECT 76.710 41.920 76.850 41.930 ;
        RECT 79.610 41.920 79.750 41.930 ;
        RECT 82.510 41.920 82.650 41.930 ;
        RECT 85.410 41.920 85.550 41.930 ;
        RECT 88.310 41.920 88.450 41.930 ;
        RECT 91.210 41.920 91.350 41.930 ;
        RECT 1.300 41.850 1.460 41.920 ;
        RECT 4.200 41.850 4.360 41.920 ;
        RECT 7.100 41.850 7.260 41.920 ;
        RECT 10.000 41.850 10.160 41.920 ;
        RECT 12.900 41.850 13.060 41.920 ;
        RECT 15.800 41.850 15.960 41.920 ;
        RECT 18.700 41.850 18.860 41.920 ;
        RECT 21.600 41.850 21.760 41.920 ;
        RECT 24.500 41.850 24.660 41.920 ;
        RECT 27.400 41.850 27.560 41.920 ;
        RECT 30.300 41.850 30.460 41.920 ;
        RECT 33.200 41.850 33.360 41.920 ;
        RECT 36.100 41.850 36.260 41.920 ;
        RECT 39.000 41.850 39.160 41.920 ;
        RECT 41.900 41.850 42.060 41.920 ;
        RECT 44.800 41.850 44.960 41.920 ;
        RECT 47.700 41.850 47.860 41.920 ;
        RECT 50.600 41.850 50.760 41.920 ;
        RECT 53.500 41.850 53.660 41.920 ;
        RECT 56.400 41.850 56.560 41.920 ;
        RECT 59.300 41.850 59.460 41.920 ;
        RECT 62.200 41.850 62.360 41.920 ;
        RECT 65.100 41.850 65.260 41.920 ;
        RECT 68.000 41.850 68.160 41.920 ;
        RECT 70.900 41.850 71.060 41.920 ;
        RECT 73.800 41.850 73.960 41.920 ;
        RECT 76.700 41.850 76.860 41.920 ;
        RECT 79.600 41.850 79.760 41.920 ;
        RECT 82.500 41.850 82.660 41.920 ;
        RECT 85.400 41.850 85.560 41.920 ;
        RECT 88.300 41.850 88.460 41.920 ;
        RECT 91.200 41.850 91.360 41.920 ;
        RECT 1.310 40.570 1.450 40.580 ;
        RECT 4.210 40.570 4.350 40.580 ;
        RECT 7.110 40.570 7.250 40.580 ;
        RECT 10.010 40.570 10.150 40.580 ;
        RECT 12.910 40.570 13.050 40.580 ;
        RECT 15.810 40.570 15.950 40.580 ;
        RECT 18.710 40.570 18.850 40.580 ;
        RECT 21.610 40.570 21.750 40.580 ;
        RECT 24.510 40.570 24.650 40.580 ;
        RECT 27.410 40.570 27.550 40.580 ;
        RECT 30.310 40.570 30.450 40.580 ;
        RECT 33.210 40.570 33.350 40.580 ;
        RECT 36.110 40.570 36.250 40.580 ;
        RECT 39.010 40.570 39.150 40.580 ;
        RECT 41.910 40.570 42.050 40.580 ;
        RECT 44.810 40.570 44.950 40.580 ;
        RECT 47.710 40.570 47.850 40.580 ;
        RECT 50.610 40.570 50.750 40.580 ;
        RECT 53.510 40.570 53.650 40.580 ;
        RECT 56.410 40.570 56.550 40.580 ;
        RECT 59.310 40.570 59.450 40.580 ;
        RECT 62.210 40.570 62.350 40.580 ;
        RECT 65.110 40.570 65.250 40.580 ;
        RECT 68.010 40.570 68.150 40.580 ;
        RECT 70.910 40.570 71.050 40.580 ;
        RECT 73.810 40.570 73.950 40.580 ;
        RECT 76.710 40.570 76.850 40.580 ;
        RECT 79.610 40.570 79.750 40.580 ;
        RECT 82.510 40.570 82.650 40.580 ;
        RECT 85.410 40.570 85.550 40.580 ;
        RECT 88.310 40.570 88.450 40.580 ;
        RECT 91.210 40.570 91.350 40.580 ;
        RECT 1.300 40.500 1.460 40.570 ;
        RECT 4.200 40.500 4.360 40.570 ;
        RECT 7.100 40.500 7.260 40.570 ;
        RECT 10.000 40.500 10.160 40.570 ;
        RECT 12.900 40.500 13.060 40.570 ;
        RECT 15.800 40.500 15.960 40.570 ;
        RECT 18.700 40.500 18.860 40.570 ;
        RECT 21.600 40.500 21.760 40.570 ;
        RECT 24.500 40.500 24.660 40.570 ;
        RECT 27.400 40.500 27.560 40.570 ;
        RECT 30.300 40.500 30.460 40.570 ;
        RECT 33.200 40.500 33.360 40.570 ;
        RECT 36.100 40.500 36.260 40.570 ;
        RECT 39.000 40.500 39.160 40.570 ;
        RECT 41.900 40.500 42.060 40.570 ;
        RECT 44.800 40.500 44.960 40.570 ;
        RECT 47.700 40.500 47.860 40.570 ;
        RECT 50.600 40.500 50.760 40.570 ;
        RECT 53.500 40.500 53.660 40.570 ;
        RECT 56.400 40.500 56.560 40.570 ;
        RECT 59.300 40.500 59.460 40.570 ;
        RECT 62.200 40.500 62.360 40.570 ;
        RECT 65.100 40.500 65.260 40.570 ;
        RECT 68.000 40.500 68.160 40.570 ;
        RECT 70.900 40.500 71.060 40.570 ;
        RECT 73.800 40.500 73.960 40.570 ;
        RECT 76.700 40.500 76.860 40.570 ;
        RECT 79.600 40.500 79.760 40.570 ;
        RECT 82.500 40.500 82.660 40.570 ;
        RECT 85.400 40.500 85.560 40.570 ;
        RECT 88.300 40.500 88.460 40.570 ;
        RECT 91.200 40.500 91.360 40.570 ;
        RECT 1.310 39.220 1.450 39.230 ;
        RECT 4.210 39.220 4.350 39.230 ;
        RECT 7.110 39.220 7.250 39.230 ;
        RECT 10.010 39.220 10.150 39.230 ;
        RECT 12.910 39.220 13.050 39.230 ;
        RECT 15.810 39.220 15.950 39.230 ;
        RECT 18.710 39.220 18.850 39.230 ;
        RECT 21.610 39.220 21.750 39.230 ;
        RECT 24.510 39.220 24.650 39.230 ;
        RECT 27.410 39.220 27.550 39.230 ;
        RECT 30.310 39.220 30.450 39.230 ;
        RECT 33.210 39.220 33.350 39.230 ;
        RECT 36.110 39.220 36.250 39.230 ;
        RECT 39.010 39.220 39.150 39.230 ;
        RECT 41.910 39.220 42.050 39.230 ;
        RECT 44.810 39.220 44.950 39.230 ;
        RECT 47.710 39.220 47.850 39.230 ;
        RECT 50.610 39.220 50.750 39.230 ;
        RECT 53.510 39.220 53.650 39.230 ;
        RECT 56.410 39.220 56.550 39.230 ;
        RECT 59.310 39.220 59.450 39.230 ;
        RECT 62.210 39.220 62.350 39.230 ;
        RECT 65.110 39.220 65.250 39.230 ;
        RECT 68.010 39.220 68.150 39.230 ;
        RECT 70.910 39.220 71.050 39.230 ;
        RECT 73.810 39.220 73.950 39.230 ;
        RECT 76.710 39.220 76.850 39.230 ;
        RECT 79.610 39.220 79.750 39.230 ;
        RECT 82.510 39.220 82.650 39.230 ;
        RECT 85.410 39.220 85.550 39.230 ;
        RECT 88.310 39.220 88.450 39.230 ;
        RECT 91.210 39.220 91.350 39.230 ;
        RECT 1.300 39.150 1.460 39.220 ;
        RECT 4.200 39.150 4.360 39.220 ;
        RECT 7.100 39.150 7.260 39.220 ;
        RECT 10.000 39.150 10.160 39.220 ;
        RECT 12.900 39.150 13.060 39.220 ;
        RECT 15.800 39.150 15.960 39.220 ;
        RECT 18.700 39.150 18.860 39.220 ;
        RECT 21.600 39.150 21.760 39.220 ;
        RECT 24.500 39.150 24.660 39.220 ;
        RECT 27.400 39.150 27.560 39.220 ;
        RECT 30.300 39.150 30.460 39.220 ;
        RECT 33.200 39.150 33.360 39.220 ;
        RECT 36.100 39.150 36.260 39.220 ;
        RECT 39.000 39.150 39.160 39.220 ;
        RECT 41.900 39.150 42.060 39.220 ;
        RECT 44.800 39.150 44.960 39.220 ;
        RECT 47.700 39.150 47.860 39.220 ;
        RECT 50.600 39.150 50.760 39.220 ;
        RECT 53.500 39.150 53.660 39.220 ;
        RECT 56.400 39.150 56.560 39.220 ;
        RECT 59.300 39.150 59.460 39.220 ;
        RECT 62.200 39.150 62.360 39.220 ;
        RECT 65.100 39.150 65.260 39.220 ;
        RECT 68.000 39.150 68.160 39.220 ;
        RECT 70.900 39.150 71.060 39.220 ;
        RECT 73.800 39.150 73.960 39.220 ;
        RECT 76.700 39.150 76.860 39.220 ;
        RECT 79.600 39.150 79.760 39.220 ;
        RECT 82.500 39.150 82.660 39.220 ;
        RECT 85.400 39.150 85.560 39.220 ;
        RECT 88.300 39.150 88.460 39.220 ;
        RECT 91.200 39.150 91.360 39.220 ;
        RECT 1.310 37.870 1.450 37.880 ;
        RECT 4.210 37.870 4.350 37.880 ;
        RECT 7.110 37.870 7.250 37.880 ;
        RECT 10.010 37.870 10.150 37.880 ;
        RECT 12.910 37.870 13.050 37.880 ;
        RECT 15.810 37.870 15.950 37.880 ;
        RECT 18.710 37.870 18.850 37.880 ;
        RECT 21.610 37.870 21.750 37.880 ;
        RECT 24.510 37.870 24.650 37.880 ;
        RECT 27.410 37.870 27.550 37.880 ;
        RECT 30.310 37.870 30.450 37.880 ;
        RECT 33.210 37.870 33.350 37.880 ;
        RECT 36.110 37.870 36.250 37.880 ;
        RECT 39.010 37.870 39.150 37.880 ;
        RECT 41.910 37.870 42.050 37.880 ;
        RECT 44.810 37.870 44.950 37.880 ;
        RECT 47.710 37.870 47.850 37.880 ;
        RECT 50.610 37.870 50.750 37.880 ;
        RECT 53.510 37.870 53.650 37.880 ;
        RECT 56.410 37.870 56.550 37.880 ;
        RECT 59.310 37.870 59.450 37.880 ;
        RECT 62.210 37.870 62.350 37.880 ;
        RECT 65.110 37.870 65.250 37.880 ;
        RECT 68.010 37.870 68.150 37.880 ;
        RECT 70.910 37.870 71.050 37.880 ;
        RECT 73.810 37.870 73.950 37.880 ;
        RECT 76.710 37.870 76.850 37.880 ;
        RECT 79.610 37.870 79.750 37.880 ;
        RECT 82.510 37.870 82.650 37.880 ;
        RECT 85.410 37.870 85.550 37.880 ;
        RECT 88.310 37.870 88.450 37.880 ;
        RECT 91.210 37.870 91.350 37.880 ;
        RECT 1.300 37.800 1.460 37.870 ;
        RECT 4.200 37.800 4.360 37.870 ;
        RECT 7.100 37.800 7.260 37.870 ;
        RECT 10.000 37.800 10.160 37.870 ;
        RECT 12.900 37.800 13.060 37.870 ;
        RECT 15.800 37.800 15.960 37.870 ;
        RECT 18.700 37.800 18.860 37.870 ;
        RECT 21.600 37.800 21.760 37.870 ;
        RECT 24.500 37.800 24.660 37.870 ;
        RECT 27.400 37.800 27.560 37.870 ;
        RECT 30.300 37.800 30.460 37.870 ;
        RECT 33.200 37.800 33.360 37.870 ;
        RECT 36.100 37.800 36.260 37.870 ;
        RECT 39.000 37.800 39.160 37.870 ;
        RECT 41.900 37.800 42.060 37.870 ;
        RECT 44.800 37.800 44.960 37.870 ;
        RECT 47.700 37.800 47.860 37.870 ;
        RECT 50.600 37.800 50.760 37.870 ;
        RECT 53.500 37.800 53.660 37.870 ;
        RECT 56.400 37.800 56.560 37.870 ;
        RECT 59.300 37.800 59.460 37.870 ;
        RECT 62.200 37.800 62.360 37.870 ;
        RECT 65.100 37.800 65.260 37.870 ;
        RECT 68.000 37.800 68.160 37.870 ;
        RECT 70.900 37.800 71.060 37.870 ;
        RECT 73.800 37.800 73.960 37.870 ;
        RECT 76.700 37.800 76.860 37.870 ;
        RECT 79.600 37.800 79.760 37.870 ;
        RECT 82.500 37.800 82.660 37.870 ;
        RECT 85.400 37.800 85.560 37.870 ;
        RECT 88.300 37.800 88.460 37.870 ;
        RECT 91.200 37.800 91.360 37.870 ;
        RECT 1.310 36.520 1.450 36.530 ;
        RECT 4.210 36.520 4.350 36.530 ;
        RECT 7.110 36.520 7.250 36.530 ;
        RECT 10.010 36.520 10.150 36.530 ;
        RECT 12.910 36.520 13.050 36.530 ;
        RECT 15.810 36.520 15.950 36.530 ;
        RECT 18.710 36.520 18.850 36.530 ;
        RECT 21.610 36.520 21.750 36.530 ;
        RECT 24.510 36.520 24.650 36.530 ;
        RECT 27.410 36.520 27.550 36.530 ;
        RECT 30.310 36.520 30.450 36.530 ;
        RECT 33.210 36.520 33.350 36.530 ;
        RECT 36.110 36.520 36.250 36.530 ;
        RECT 39.010 36.520 39.150 36.530 ;
        RECT 41.910 36.520 42.050 36.530 ;
        RECT 44.810 36.520 44.950 36.530 ;
        RECT 47.710 36.520 47.850 36.530 ;
        RECT 50.610 36.520 50.750 36.530 ;
        RECT 53.510 36.520 53.650 36.530 ;
        RECT 56.410 36.520 56.550 36.530 ;
        RECT 59.310 36.520 59.450 36.530 ;
        RECT 62.210 36.520 62.350 36.530 ;
        RECT 65.110 36.520 65.250 36.530 ;
        RECT 68.010 36.520 68.150 36.530 ;
        RECT 70.910 36.520 71.050 36.530 ;
        RECT 73.810 36.520 73.950 36.530 ;
        RECT 76.710 36.520 76.850 36.530 ;
        RECT 79.610 36.520 79.750 36.530 ;
        RECT 82.510 36.520 82.650 36.530 ;
        RECT 85.410 36.520 85.550 36.530 ;
        RECT 88.310 36.520 88.450 36.530 ;
        RECT 91.210 36.520 91.350 36.530 ;
        RECT 1.300 36.450 1.460 36.520 ;
        RECT 4.200 36.450 4.360 36.520 ;
        RECT 7.100 36.450 7.260 36.520 ;
        RECT 10.000 36.450 10.160 36.520 ;
        RECT 12.900 36.450 13.060 36.520 ;
        RECT 15.800 36.450 15.960 36.520 ;
        RECT 18.700 36.450 18.860 36.520 ;
        RECT 21.600 36.450 21.760 36.520 ;
        RECT 24.500 36.450 24.660 36.520 ;
        RECT 27.400 36.450 27.560 36.520 ;
        RECT 30.300 36.450 30.460 36.520 ;
        RECT 33.200 36.450 33.360 36.520 ;
        RECT 36.100 36.450 36.260 36.520 ;
        RECT 39.000 36.450 39.160 36.520 ;
        RECT 41.900 36.450 42.060 36.520 ;
        RECT 44.800 36.450 44.960 36.520 ;
        RECT 47.700 36.450 47.860 36.520 ;
        RECT 50.600 36.450 50.760 36.520 ;
        RECT 53.500 36.450 53.660 36.520 ;
        RECT 56.400 36.450 56.560 36.520 ;
        RECT 59.300 36.450 59.460 36.520 ;
        RECT 62.200 36.450 62.360 36.520 ;
        RECT 65.100 36.450 65.260 36.520 ;
        RECT 68.000 36.450 68.160 36.520 ;
        RECT 70.900 36.450 71.060 36.520 ;
        RECT 73.800 36.450 73.960 36.520 ;
        RECT 76.700 36.450 76.860 36.520 ;
        RECT 79.600 36.450 79.760 36.520 ;
        RECT 82.500 36.450 82.660 36.520 ;
        RECT 85.400 36.450 85.560 36.520 ;
        RECT 88.300 36.450 88.460 36.520 ;
        RECT 91.200 36.450 91.360 36.520 ;
        RECT 1.310 35.170 1.450 35.180 ;
        RECT 4.210 35.170 4.350 35.180 ;
        RECT 7.110 35.170 7.250 35.180 ;
        RECT 10.010 35.170 10.150 35.180 ;
        RECT 12.910 35.170 13.050 35.180 ;
        RECT 15.810 35.170 15.950 35.180 ;
        RECT 18.710 35.170 18.850 35.180 ;
        RECT 21.610 35.170 21.750 35.180 ;
        RECT 24.510 35.170 24.650 35.180 ;
        RECT 27.410 35.170 27.550 35.180 ;
        RECT 30.310 35.170 30.450 35.180 ;
        RECT 33.210 35.170 33.350 35.180 ;
        RECT 36.110 35.170 36.250 35.180 ;
        RECT 39.010 35.170 39.150 35.180 ;
        RECT 41.910 35.170 42.050 35.180 ;
        RECT 44.810 35.170 44.950 35.180 ;
        RECT 47.710 35.170 47.850 35.180 ;
        RECT 50.610 35.170 50.750 35.180 ;
        RECT 53.510 35.170 53.650 35.180 ;
        RECT 56.410 35.170 56.550 35.180 ;
        RECT 59.310 35.170 59.450 35.180 ;
        RECT 62.210 35.170 62.350 35.180 ;
        RECT 65.110 35.170 65.250 35.180 ;
        RECT 68.010 35.170 68.150 35.180 ;
        RECT 70.910 35.170 71.050 35.180 ;
        RECT 73.810 35.170 73.950 35.180 ;
        RECT 76.710 35.170 76.850 35.180 ;
        RECT 79.610 35.170 79.750 35.180 ;
        RECT 82.510 35.170 82.650 35.180 ;
        RECT 85.410 35.170 85.550 35.180 ;
        RECT 88.310 35.170 88.450 35.180 ;
        RECT 91.210 35.170 91.350 35.180 ;
        RECT 1.300 35.100 1.460 35.170 ;
        RECT 4.200 35.100 4.360 35.170 ;
        RECT 7.100 35.100 7.260 35.170 ;
        RECT 10.000 35.100 10.160 35.170 ;
        RECT 12.900 35.100 13.060 35.170 ;
        RECT 15.800 35.100 15.960 35.170 ;
        RECT 18.700 35.100 18.860 35.170 ;
        RECT 21.600 35.100 21.760 35.170 ;
        RECT 24.500 35.100 24.660 35.170 ;
        RECT 27.400 35.100 27.560 35.170 ;
        RECT 30.300 35.100 30.460 35.170 ;
        RECT 33.200 35.100 33.360 35.170 ;
        RECT 36.100 35.100 36.260 35.170 ;
        RECT 39.000 35.100 39.160 35.170 ;
        RECT 41.900 35.100 42.060 35.170 ;
        RECT 44.800 35.100 44.960 35.170 ;
        RECT 47.700 35.100 47.860 35.170 ;
        RECT 50.600 35.100 50.760 35.170 ;
        RECT 53.500 35.100 53.660 35.170 ;
        RECT 56.400 35.100 56.560 35.170 ;
        RECT 59.300 35.100 59.460 35.170 ;
        RECT 62.200 35.100 62.360 35.170 ;
        RECT 65.100 35.100 65.260 35.170 ;
        RECT 68.000 35.100 68.160 35.170 ;
        RECT 70.900 35.100 71.060 35.170 ;
        RECT 73.800 35.100 73.960 35.170 ;
        RECT 76.700 35.100 76.860 35.170 ;
        RECT 79.600 35.100 79.760 35.170 ;
        RECT 82.500 35.100 82.660 35.170 ;
        RECT 85.400 35.100 85.560 35.170 ;
        RECT 88.300 35.100 88.460 35.170 ;
        RECT 91.200 35.100 91.360 35.170 ;
        RECT 1.310 33.820 1.450 33.830 ;
        RECT 4.210 33.820 4.350 33.830 ;
        RECT 7.110 33.820 7.250 33.830 ;
        RECT 10.010 33.820 10.150 33.830 ;
        RECT 12.910 33.820 13.050 33.830 ;
        RECT 15.810 33.820 15.950 33.830 ;
        RECT 18.710 33.820 18.850 33.830 ;
        RECT 21.610 33.820 21.750 33.830 ;
        RECT 24.510 33.820 24.650 33.830 ;
        RECT 27.410 33.820 27.550 33.830 ;
        RECT 30.310 33.820 30.450 33.830 ;
        RECT 33.210 33.820 33.350 33.830 ;
        RECT 36.110 33.820 36.250 33.830 ;
        RECT 39.010 33.820 39.150 33.830 ;
        RECT 41.910 33.820 42.050 33.830 ;
        RECT 44.810 33.820 44.950 33.830 ;
        RECT 47.710 33.820 47.850 33.830 ;
        RECT 50.610 33.820 50.750 33.830 ;
        RECT 53.510 33.820 53.650 33.830 ;
        RECT 56.410 33.820 56.550 33.830 ;
        RECT 59.310 33.820 59.450 33.830 ;
        RECT 62.210 33.820 62.350 33.830 ;
        RECT 65.110 33.820 65.250 33.830 ;
        RECT 68.010 33.820 68.150 33.830 ;
        RECT 70.910 33.820 71.050 33.830 ;
        RECT 73.810 33.820 73.950 33.830 ;
        RECT 76.710 33.820 76.850 33.830 ;
        RECT 79.610 33.820 79.750 33.830 ;
        RECT 82.510 33.820 82.650 33.830 ;
        RECT 85.410 33.820 85.550 33.830 ;
        RECT 88.310 33.820 88.450 33.830 ;
        RECT 91.210 33.820 91.350 33.830 ;
        RECT 1.300 33.750 1.460 33.820 ;
        RECT 4.200 33.750 4.360 33.820 ;
        RECT 7.100 33.750 7.260 33.820 ;
        RECT 10.000 33.750 10.160 33.820 ;
        RECT 12.900 33.750 13.060 33.820 ;
        RECT 15.800 33.750 15.960 33.820 ;
        RECT 18.700 33.750 18.860 33.820 ;
        RECT 21.600 33.750 21.760 33.820 ;
        RECT 24.500 33.750 24.660 33.820 ;
        RECT 27.400 33.750 27.560 33.820 ;
        RECT 30.300 33.750 30.460 33.820 ;
        RECT 33.200 33.750 33.360 33.820 ;
        RECT 36.100 33.750 36.260 33.820 ;
        RECT 39.000 33.750 39.160 33.820 ;
        RECT 41.900 33.750 42.060 33.820 ;
        RECT 44.800 33.750 44.960 33.820 ;
        RECT 47.700 33.750 47.860 33.820 ;
        RECT 50.600 33.750 50.760 33.820 ;
        RECT 53.500 33.750 53.660 33.820 ;
        RECT 56.400 33.750 56.560 33.820 ;
        RECT 59.300 33.750 59.460 33.820 ;
        RECT 62.200 33.750 62.360 33.820 ;
        RECT 65.100 33.750 65.260 33.820 ;
        RECT 68.000 33.750 68.160 33.820 ;
        RECT 70.900 33.750 71.060 33.820 ;
        RECT 73.800 33.750 73.960 33.820 ;
        RECT 76.700 33.750 76.860 33.820 ;
        RECT 79.600 33.750 79.760 33.820 ;
        RECT 82.500 33.750 82.660 33.820 ;
        RECT 85.400 33.750 85.560 33.820 ;
        RECT 88.300 33.750 88.460 33.820 ;
        RECT 91.200 33.750 91.360 33.820 ;
        RECT 1.310 32.470 1.450 32.480 ;
        RECT 4.210 32.470 4.350 32.480 ;
        RECT 7.110 32.470 7.250 32.480 ;
        RECT 10.010 32.470 10.150 32.480 ;
        RECT 12.910 32.470 13.050 32.480 ;
        RECT 15.810 32.470 15.950 32.480 ;
        RECT 18.710 32.470 18.850 32.480 ;
        RECT 21.610 32.470 21.750 32.480 ;
        RECT 24.510 32.470 24.650 32.480 ;
        RECT 27.410 32.470 27.550 32.480 ;
        RECT 30.310 32.470 30.450 32.480 ;
        RECT 33.210 32.470 33.350 32.480 ;
        RECT 36.110 32.470 36.250 32.480 ;
        RECT 39.010 32.470 39.150 32.480 ;
        RECT 41.910 32.470 42.050 32.480 ;
        RECT 44.810 32.470 44.950 32.480 ;
        RECT 47.710 32.470 47.850 32.480 ;
        RECT 50.610 32.470 50.750 32.480 ;
        RECT 53.510 32.470 53.650 32.480 ;
        RECT 56.410 32.470 56.550 32.480 ;
        RECT 59.310 32.470 59.450 32.480 ;
        RECT 62.210 32.470 62.350 32.480 ;
        RECT 65.110 32.470 65.250 32.480 ;
        RECT 68.010 32.470 68.150 32.480 ;
        RECT 70.910 32.470 71.050 32.480 ;
        RECT 73.810 32.470 73.950 32.480 ;
        RECT 76.710 32.470 76.850 32.480 ;
        RECT 79.610 32.470 79.750 32.480 ;
        RECT 82.510 32.470 82.650 32.480 ;
        RECT 85.410 32.470 85.550 32.480 ;
        RECT 88.310 32.470 88.450 32.480 ;
        RECT 91.210 32.470 91.350 32.480 ;
        RECT 1.300 32.400 1.460 32.470 ;
        RECT 4.200 32.400 4.360 32.470 ;
        RECT 7.100 32.400 7.260 32.470 ;
        RECT 10.000 32.400 10.160 32.470 ;
        RECT 12.900 32.400 13.060 32.470 ;
        RECT 15.800 32.400 15.960 32.470 ;
        RECT 18.700 32.400 18.860 32.470 ;
        RECT 21.600 32.400 21.760 32.470 ;
        RECT 24.500 32.400 24.660 32.470 ;
        RECT 27.400 32.400 27.560 32.470 ;
        RECT 30.300 32.400 30.460 32.470 ;
        RECT 33.200 32.400 33.360 32.470 ;
        RECT 36.100 32.400 36.260 32.470 ;
        RECT 39.000 32.400 39.160 32.470 ;
        RECT 41.900 32.400 42.060 32.470 ;
        RECT 44.800 32.400 44.960 32.470 ;
        RECT 47.700 32.400 47.860 32.470 ;
        RECT 50.600 32.400 50.760 32.470 ;
        RECT 53.500 32.400 53.660 32.470 ;
        RECT 56.400 32.400 56.560 32.470 ;
        RECT 59.300 32.400 59.460 32.470 ;
        RECT 62.200 32.400 62.360 32.470 ;
        RECT 65.100 32.400 65.260 32.470 ;
        RECT 68.000 32.400 68.160 32.470 ;
        RECT 70.900 32.400 71.060 32.470 ;
        RECT 73.800 32.400 73.960 32.470 ;
        RECT 76.700 32.400 76.860 32.470 ;
        RECT 79.600 32.400 79.760 32.470 ;
        RECT 82.500 32.400 82.660 32.470 ;
        RECT 85.400 32.400 85.560 32.470 ;
        RECT 88.300 32.400 88.460 32.470 ;
        RECT 91.200 32.400 91.360 32.470 ;
        RECT 1.310 31.120 1.450 31.130 ;
        RECT 4.210 31.120 4.350 31.130 ;
        RECT 7.110 31.120 7.250 31.130 ;
        RECT 10.010 31.120 10.150 31.130 ;
        RECT 12.910 31.120 13.050 31.130 ;
        RECT 15.810 31.120 15.950 31.130 ;
        RECT 18.710 31.120 18.850 31.130 ;
        RECT 21.610 31.120 21.750 31.130 ;
        RECT 24.510 31.120 24.650 31.130 ;
        RECT 27.410 31.120 27.550 31.130 ;
        RECT 30.310 31.120 30.450 31.130 ;
        RECT 33.210 31.120 33.350 31.130 ;
        RECT 36.110 31.120 36.250 31.130 ;
        RECT 39.010 31.120 39.150 31.130 ;
        RECT 41.910 31.120 42.050 31.130 ;
        RECT 44.810 31.120 44.950 31.130 ;
        RECT 47.710 31.120 47.850 31.130 ;
        RECT 50.610 31.120 50.750 31.130 ;
        RECT 53.510 31.120 53.650 31.130 ;
        RECT 56.410 31.120 56.550 31.130 ;
        RECT 59.310 31.120 59.450 31.130 ;
        RECT 62.210 31.120 62.350 31.130 ;
        RECT 65.110 31.120 65.250 31.130 ;
        RECT 68.010 31.120 68.150 31.130 ;
        RECT 70.910 31.120 71.050 31.130 ;
        RECT 73.810 31.120 73.950 31.130 ;
        RECT 76.710 31.120 76.850 31.130 ;
        RECT 79.610 31.120 79.750 31.130 ;
        RECT 82.510 31.120 82.650 31.130 ;
        RECT 85.410 31.120 85.550 31.130 ;
        RECT 88.310 31.120 88.450 31.130 ;
        RECT 91.210 31.120 91.350 31.130 ;
        RECT 1.300 31.050 1.460 31.120 ;
        RECT 4.200 31.050 4.360 31.120 ;
        RECT 7.100 31.050 7.260 31.120 ;
        RECT 10.000 31.050 10.160 31.120 ;
        RECT 12.900 31.050 13.060 31.120 ;
        RECT 15.800 31.050 15.960 31.120 ;
        RECT 18.700 31.050 18.860 31.120 ;
        RECT 21.600 31.050 21.760 31.120 ;
        RECT 24.500 31.050 24.660 31.120 ;
        RECT 27.400 31.050 27.560 31.120 ;
        RECT 30.300 31.050 30.460 31.120 ;
        RECT 33.200 31.050 33.360 31.120 ;
        RECT 36.100 31.050 36.260 31.120 ;
        RECT 39.000 31.050 39.160 31.120 ;
        RECT 41.900 31.050 42.060 31.120 ;
        RECT 44.800 31.050 44.960 31.120 ;
        RECT 47.700 31.050 47.860 31.120 ;
        RECT 50.600 31.050 50.760 31.120 ;
        RECT 53.500 31.050 53.660 31.120 ;
        RECT 56.400 31.050 56.560 31.120 ;
        RECT 59.300 31.050 59.460 31.120 ;
        RECT 62.200 31.050 62.360 31.120 ;
        RECT 65.100 31.050 65.260 31.120 ;
        RECT 68.000 31.050 68.160 31.120 ;
        RECT 70.900 31.050 71.060 31.120 ;
        RECT 73.800 31.050 73.960 31.120 ;
        RECT 76.700 31.050 76.860 31.120 ;
        RECT 79.600 31.050 79.760 31.120 ;
        RECT 82.500 31.050 82.660 31.120 ;
        RECT 85.400 31.050 85.560 31.120 ;
        RECT 88.300 31.050 88.460 31.120 ;
        RECT 91.200 31.050 91.360 31.120 ;
        RECT 1.310 29.770 1.450 29.780 ;
        RECT 4.210 29.770 4.350 29.780 ;
        RECT 7.110 29.770 7.250 29.780 ;
        RECT 10.010 29.770 10.150 29.780 ;
        RECT 12.910 29.770 13.050 29.780 ;
        RECT 15.810 29.770 15.950 29.780 ;
        RECT 18.710 29.770 18.850 29.780 ;
        RECT 21.610 29.770 21.750 29.780 ;
        RECT 24.510 29.770 24.650 29.780 ;
        RECT 27.410 29.770 27.550 29.780 ;
        RECT 30.310 29.770 30.450 29.780 ;
        RECT 33.210 29.770 33.350 29.780 ;
        RECT 36.110 29.770 36.250 29.780 ;
        RECT 39.010 29.770 39.150 29.780 ;
        RECT 41.910 29.770 42.050 29.780 ;
        RECT 44.810 29.770 44.950 29.780 ;
        RECT 47.710 29.770 47.850 29.780 ;
        RECT 50.610 29.770 50.750 29.780 ;
        RECT 53.510 29.770 53.650 29.780 ;
        RECT 56.410 29.770 56.550 29.780 ;
        RECT 59.310 29.770 59.450 29.780 ;
        RECT 62.210 29.770 62.350 29.780 ;
        RECT 65.110 29.770 65.250 29.780 ;
        RECT 68.010 29.770 68.150 29.780 ;
        RECT 70.910 29.770 71.050 29.780 ;
        RECT 73.810 29.770 73.950 29.780 ;
        RECT 76.710 29.770 76.850 29.780 ;
        RECT 79.610 29.770 79.750 29.780 ;
        RECT 82.510 29.770 82.650 29.780 ;
        RECT 85.410 29.770 85.550 29.780 ;
        RECT 88.310 29.770 88.450 29.780 ;
        RECT 91.210 29.770 91.350 29.780 ;
        RECT 1.300 29.700 1.460 29.770 ;
        RECT 4.200 29.700 4.360 29.770 ;
        RECT 7.100 29.700 7.260 29.770 ;
        RECT 10.000 29.700 10.160 29.770 ;
        RECT 12.900 29.700 13.060 29.770 ;
        RECT 15.800 29.700 15.960 29.770 ;
        RECT 18.700 29.700 18.860 29.770 ;
        RECT 21.600 29.700 21.760 29.770 ;
        RECT 24.500 29.700 24.660 29.770 ;
        RECT 27.400 29.700 27.560 29.770 ;
        RECT 30.300 29.700 30.460 29.770 ;
        RECT 33.200 29.700 33.360 29.770 ;
        RECT 36.100 29.700 36.260 29.770 ;
        RECT 39.000 29.700 39.160 29.770 ;
        RECT 41.900 29.700 42.060 29.770 ;
        RECT 44.800 29.700 44.960 29.770 ;
        RECT 47.700 29.700 47.860 29.770 ;
        RECT 50.600 29.700 50.760 29.770 ;
        RECT 53.500 29.700 53.660 29.770 ;
        RECT 56.400 29.700 56.560 29.770 ;
        RECT 59.300 29.700 59.460 29.770 ;
        RECT 62.200 29.700 62.360 29.770 ;
        RECT 65.100 29.700 65.260 29.770 ;
        RECT 68.000 29.700 68.160 29.770 ;
        RECT 70.900 29.700 71.060 29.770 ;
        RECT 73.800 29.700 73.960 29.770 ;
        RECT 76.700 29.700 76.860 29.770 ;
        RECT 79.600 29.700 79.760 29.770 ;
        RECT 82.500 29.700 82.660 29.770 ;
        RECT 85.400 29.700 85.560 29.770 ;
        RECT 88.300 29.700 88.460 29.770 ;
        RECT 91.200 29.700 91.360 29.770 ;
        RECT 1.310 28.420 1.450 28.430 ;
        RECT 4.210 28.420 4.350 28.430 ;
        RECT 7.110 28.420 7.250 28.430 ;
        RECT 10.010 28.420 10.150 28.430 ;
        RECT 12.910 28.420 13.050 28.430 ;
        RECT 15.810 28.420 15.950 28.430 ;
        RECT 18.710 28.420 18.850 28.430 ;
        RECT 21.610 28.420 21.750 28.430 ;
        RECT 24.510 28.420 24.650 28.430 ;
        RECT 27.410 28.420 27.550 28.430 ;
        RECT 30.310 28.420 30.450 28.430 ;
        RECT 33.210 28.420 33.350 28.430 ;
        RECT 36.110 28.420 36.250 28.430 ;
        RECT 39.010 28.420 39.150 28.430 ;
        RECT 41.910 28.420 42.050 28.430 ;
        RECT 44.810 28.420 44.950 28.430 ;
        RECT 47.710 28.420 47.850 28.430 ;
        RECT 50.610 28.420 50.750 28.430 ;
        RECT 53.510 28.420 53.650 28.430 ;
        RECT 56.410 28.420 56.550 28.430 ;
        RECT 59.310 28.420 59.450 28.430 ;
        RECT 62.210 28.420 62.350 28.430 ;
        RECT 65.110 28.420 65.250 28.430 ;
        RECT 68.010 28.420 68.150 28.430 ;
        RECT 70.910 28.420 71.050 28.430 ;
        RECT 73.810 28.420 73.950 28.430 ;
        RECT 76.710 28.420 76.850 28.430 ;
        RECT 79.610 28.420 79.750 28.430 ;
        RECT 82.510 28.420 82.650 28.430 ;
        RECT 85.410 28.420 85.550 28.430 ;
        RECT 88.310 28.420 88.450 28.430 ;
        RECT 91.210 28.420 91.350 28.430 ;
        RECT 1.300 28.350 1.460 28.420 ;
        RECT 4.200 28.350 4.360 28.420 ;
        RECT 7.100 28.350 7.260 28.420 ;
        RECT 10.000 28.350 10.160 28.420 ;
        RECT 12.900 28.350 13.060 28.420 ;
        RECT 15.800 28.350 15.960 28.420 ;
        RECT 18.700 28.350 18.860 28.420 ;
        RECT 21.600 28.350 21.760 28.420 ;
        RECT 24.500 28.350 24.660 28.420 ;
        RECT 27.400 28.350 27.560 28.420 ;
        RECT 30.300 28.350 30.460 28.420 ;
        RECT 33.200 28.350 33.360 28.420 ;
        RECT 36.100 28.350 36.260 28.420 ;
        RECT 39.000 28.350 39.160 28.420 ;
        RECT 41.900 28.350 42.060 28.420 ;
        RECT 44.800 28.350 44.960 28.420 ;
        RECT 47.700 28.350 47.860 28.420 ;
        RECT 50.600 28.350 50.760 28.420 ;
        RECT 53.500 28.350 53.660 28.420 ;
        RECT 56.400 28.350 56.560 28.420 ;
        RECT 59.300 28.350 59.460 28.420 ;
        RECT 62.200 28.350 62.360 28.420 ;
        RECT 65.100 28.350 65.260 28.420 ;
        RECT 68.000 28.350 68.160 28.420 ;
        RECT 70.900 28.350 71.060 28.420 ;
        RECT 73.800 28.350 73.960 28.420 ;
        RECT 76.700 28.350 76.860 28.420 ;
        RECT 79.600 28.350 79.760 28.420 ;
        RECT 82.500 28.350 82.660 28.420 ;
        RECT 85.400 28.350 85.560 28.420 ;
        RECT 88.300 28.350 88.460 28.420 ;
        RECT 91.200 28.350 91.360 28.420 ;
        RECT 1.310 27.070 1.450 27.080 ;
        RECT 4.210 27.070 4.350 27.080 ;
        RECT 7.110 27.070 7.250 27.080 ;
        RECT 10.010 27.070 10.150 27.080 ;
        RECT 12.910 27.070 13.050 27.080 ;
        RECT 15.810 27.070 15.950 27.080 ;
        RECT 18.710 27.070 18.850 27.080 ;
        RECT 21.610 27.070 21.750 27.080 ;
        RECT 24.510 27.070 24.650 27.080 ;
        RECT 27.410 27.070 27.550 27.080 ;
        RECT 30.310 27.070 30.450 27.080 ;
        RECT 33.210 27.070 33.350 27.080 ;
        RECT 36.110 27.070 36.250 27.080 ;
        RECT 39.010 27.070 39.150 27.080 ;
        RECT 41.910 27.070 42.050 27.080 ;
        RECT 44.810 27.070 44.950 27.080 ;
        RECT 47.710 27.070 47.850 27.080 ;
        RECT 50.610 27.070 50.750 27.080 ;
        RECT 53.510 27.070 53.650 27.080 ;
        RECT 56.410 27.070 56.550 27.080 ;
        RECT 59.310 27.070 59.450 27.080 ;
        RECT 62.210 27.070 62.350 27.080 ;
        RECT 65.110 27.070 65.250 27.080 ;
        RECT 68.010 27.070 68.150 27.080 ;
        RECT 70.910 27.070 71.050 27.080 ;
        RECT 73.810 27.070 73.950 27.080 ;
        RECT 76.710 27.070 76.850 27.080 ;
        RECT 79.610 27.070 79.750 27.080 ;
        RECT 82.510 27.070 82.650 27.080 ;
        RECT 85.410 27.070 85.550 27.080 ;
        RECT 88.310 27.070 88.450 27.080 ;
        RECT 91.210 27.070 91.350 27.080 ;
        RECT 1.300 27.000 1.460 27.070 ;
        RECT 4.200 27.000 4.360 27.070 ;
        RECT 7.100 27.000 7.260 27.070 ;
        RECT 10.000 27.000 10.160 27.070 ;
        RECT 12.900 27.000 13.060 27.070 ;
        RECT 15.800 27.000 15.960 27.070 ;
        RECT 18.700 27.000 18.860 27.070 ;
        RECT 21.600 27.000 21.760 27.070 ;
        RECT 24.500 27.000 24.660 27.070 ;
        RECT 27.400 27.000 27.560 27.070 ;
        RECT 30.300 27.000 30.460 27.070 ;
        RECT 33.200 27.000 33.360 27.070 ;
        RECT 36.100 27.000 36.260 27.070 ;
        RECT 39.000 27.000 39.160 27.070 ;
        RECT 41.900 27.000 42.060 27.070 ;
        RECT 44.800 27.000 44.960 27.070 ;
        RECT 47.700 27.000 47.860 27.070 ;
        RECT 50.600 27.000 50.760 27.070 ;
        RECT 53.500 27.000 53.660 27.070 ;
        RECT 56.400 27.000 56.560 27.070 ;
        RECT 59.300 27.000 59.460 27.070 ;
        RECT 62.200 27.000 62.360 27.070 ;
        RECT 65.100 27.000 65.260 27.070 ;
        RECT 68.000 27.000 68.160 27.070 ;
        RECT 70.900 27.000 71.060 27.070 ;
        RECT 73.800 27.000 73.960 27.070 ;
        RECT 76.700 27.000 76.860 27.070 ;
        RECT 79.600 27.000 79.760 27.070 ;
        RECT 82.500 27.000 82.660 27.070 ;
        RECT 85.400 27.000 85.560 27.070 ;
        RECT 88.300 27.000 88.460 27.070 ;
        RECT 91.200 27.000 91.360 27.070 ;
        RECT 1.310 25.720 1.450 25.730 ;
        RECT 4.210 25.720 4.350 25.730 ;
        RECT 7.110 25.720 7.250 25.730 ;
        RECT 10.010 25.720 10.150 25.730 ;
        RECT 12.910 25.720 13.050 25.730 ;
        RECT 15.810 25.720 15.950 25.730 ;
        RECT 18.710 25.720 18.850 25.730 ;
        RECT 21.610 25.720 21.750 25.730 ;
        RECT 24.510 25.720 24.650 25.730 ;
        RECT 27.410 25.720 27.550 25.730 ;
        RECT 30.310 25.720 30.450 25.730 ;
        RECT 33.210 25.720 33.350 25.730 ;
        RECT 36.110 25.720 36.250 25.730 ;
        RECT 39.010 25.720 39.150 25.730 ;
        RECT 41.910 25.720 42.050 25.730 ;
        RECT 44.810 25.720 44.950 25.730 ;
        RECT 47.710 25.720 47.850 25.730 ;
        RECT 50.610 25.720 50.750 25.730 ;
        RECT 53.510 25.720 53.650 25.730 ;
        RECT 56.410 25.720 56.550 25.730 ;
        RECT 59.310 25.720 59.450 25.730 ;
        RECT 62.210 25.720 62.350 25.730 ;
        RECT 65.110 25.720 65.250 25.730 ;
        RECT 68.010 25.720 68.150 25.730 ;
        RECT 70.910 25.720 71.050 25.730 ;
        RECT 73.810 25.720 73.950 25.730 ;
        RECT 76.710 25.720 76.850 25.730 ;
        RECT 79.610 25.720 79.750 25.730 ;
        RECT 82.510 25.720 82.650 25.730 ;
        RECT 85.410 25.720 85.550 25.730 ;
        RECT 88.310 25.720 88.450 25.730 ;
        RECT 91.210 25.720 91.350 25.730 ;
        RECT 1.300 25.650 1.460 25.720 ;
        RECT 4.200 25.650 4.360 25.720 ;
        RECT 7.100 25.650 7.260 25.720 ;
        RECT 10.000 25.650 10.160 25.720 ;
        RECT 12.900 25.650 13.060 25.720 ;
        RECT 15.800 25.650 15.960 25.720 ;
        RECT 18.700 25.650 18.860 25.720 ;
        RECT 21.600 25.650 21.760 25.720 ;
        RECT 24.500 25.650 24.660 25.720 ;
        RECT 27.400 25.650 27.560 25.720 ;
        RECT 30.300 25.650 30.460 25.720 ;
        RECT 33.200 25.650 33.360 25.720 ;
        RECT 36.100 25.650 36.260 25.720 ;
        RECT 39.000 25.650 39.160 25.720 ;
        RECT 41.900 25.650 42.060 25.720 ;
        RECT 44.800 25.650 44.960 25.720 ;
        RECT 47.700 25.650 47.860 25.720 ;
        RECT 50.600 25.650 50.760 25.720 ;
        RECT 53.500 25.650 53.660 25.720 ;
        RECT 56.400 25.650 56.560 25.720 ;
        RECT 59.300 25.650 59.460 25.720 ;
        RECT 62.200 25.650 62.360 25.720 ;
        RECT 65.100 25.650 65.260 25.720 ;
        RECT 68.000 25.650 68.160 25.720 ;
        RECT 70.900 25.650 71.060 25.720 ;
        RECT 73.800 25.650 73.960 25.720 ;
        RECT 76.700 25.650 76.860 25.720 ;
        RECT 79.600 25.650 79.760 25.720 ;
        RECT 82.500 25.650 82.660 25.720 ;
        RECT 85.400 25.650 85.560 25.720 ;
        RECT 88.300 25.650 88.460 25.720 ;
        RECT 91.200 25.650 91.360 25.720 ;
        RECT 1.310 24.370 1.450 24.380 ;
        RECT 4.210 24.370 4.350 24.380 ;
        RECT 7.110 24.370 7.250 24.380 ;
        RECT 10.010 24.370 10.150 24.380 ;
        RECT 12.910 24.370 13.050 24.380 ;
        RECT 15.810 24.370 15.950 24.380 ;
        RECT 18.710 24.370 18.850 24.380 ;
        RECT 21.610 24.370 21.750 24.380 ;
        RECT 24.510 24.370 24.650 24.380 ;
        RECT 27.410 24.370 27.550 24.380 ;
        RECT 30.310 24.370 30.450 24.380 ;
        RECT 33.210 24.370 33.350 24.380 ;
        RECT 36.110 24.370 36.250 24.380 ;
        RECT 39.010 24.370 39.150 24.380 ;
        RECT 41.910 24.370 42.050 24.380 ;
        RECT 44.810 24.370 44.950 24.380 ;
        RECT 47.710 24.370 47.850 24.380 ;
        RECT 50.610 24.370 50.750 24.380 ;
        RECT 53.510 24.370 53.650 24.380 ;
        RECT 56.410 24.370 56.550 24.380 ;
        RECT 59.310 24.370 59.450 24.380 ;
        RECT 62.210 24.370 62.350 24.380 ;
        RECT 65.110 24.370 65.250 24.380 ;
        RECT 68.010 24.370 68.150 24.380 ;
        RECT 70.910 24.370 71.050 24.380 ;
        RECT 73.810 24.370 73.950 24.380 ;
        RECT 76.710 24.370 76.850 24.380 ;
        RECT 79.610 24.370 79.750 24.380 ;
        RECT 82.510 24.370 82.650 24.380 ;
        RECT 85.410 24.370 85.550 24.380 ;
        RECT 88.310 24.370 88.450 24.380 ;
        RECT 91.210 24.370 91.350 24.380 ;
        RECT 1.300 24.300 1.460 24.370 ;
        RECT 4.200 24.300 4.360 24.370 ;
        RECT 7.100 24.300 7.260 24.370 ;
        RECT 10.000 24.300 10.160 24.370 ;
        RECT 12.900 24.300 13.060 24.370 ;
        RECT 15.800 24.300 15.960 24.370 ;
        RECT 18.700 24.300 18.860 24.370 ;
        RECT 21.600 24.300 21.760 24.370 ;
        RECT 24.500 24.300 24.660 24.370 ;
        RECT 27.400 24.300 27.560 24.370 ;
        RECT 30.300 24.300 30.460 24.370 ;
        RECT 33.200 24.300 33.360 24.370 ;
        RECT 36.100 24.300 36.260 24.370 ;
        RECT 39.000 24.300 39.160 24.370 ;
        RECT 41.900 24.300 42.060 24.370 ;
        RECT 44.800 24.300 44.960 24.370 ;
        RECT 47.700 24.300 47.860 24.370 ;
        RECT 50.600 24.300 50.760 24.370 ;
        RECT 53.500 24.300 53.660 24.370 ;
        RECT 56.400 24.300 56.560 24.370 ;
        RECT 59.300 24.300 59.460 24.370 ;
        RECT 62.200 24.300 62.360 24.370 ;
        RECT 65.100 24.300 65.260 24.370 ;
        RECT 68.000 24.300 68.160 24.370 ;
        RECT 70.900 24.300 71.060 24.370 ;
        RECT 73.800 24.300 73.960 24.370 ;
        RECT 76.700 24.300 76.860 24.370 ;
        RECT 79.600 24.300 79.760 24.370 ;
        RECT 82.500 24.300 82.660 24.370 ;
        RECT 85.400 24.300 85.560 24.370 ;
        RECT 88.300 24.300 88.460 24.370 ;
        RECT 91.200 24.300 91.360 24.370 ;
        RECT 1.310 23.020 1.450 23.030 ;
        RECT 4.210 23.020 4.350 23.030 ;
        RECT 7.110 23.020 7.250 23.030 ;
        RECT 10.010 23.020 10.150 23.030 ;
        RECT 12.910 23.020 13.050 23.030 ;
        RECT 15.810 23.020 15.950 23.030 ;
        RECT 18.710 23.020 18.850 23.030 ;
        RECT 21.610 23.020 21.750 23.030 ;
        RECT 24.510 23.020 24.650 23.030 ;
        RECT 27.410 23.020 27.550 23.030 ;
        RECT 30.310 23.020 30.450 23.030 ;
        RECT 33.210 23.020 33.350 23.030 ;
        RECT 36.110 23.020 36.250 23.030 ;
        RECT 39.010 23.020 39.150 23.030 ;
        RECT 41.910 23.020 42.050 23.030 ;
        RECT 44.810 23.020 44.950 23.030 ;
        RECT 47.710 23.020 47.850 23.030 ;
        RECT 50.610 23.020 50.750 23.030 ;
        RECT 53.510 23.020 53.650 23.030 ;
        RECT 56.410 23.020 56.550 23.030 ;
        RECT 59.310 23.020 59.450 23.030 ;
        RECT 62.210 23.020 62.350 23.030 ;
        RECT 65.110 23.020 65.250 23.030 ;
        RECT 68.010 23.020 68.150 23.030 ;
        RECT 70.910 23.020 71.050 23.030 ;
        RECT 73.810 23.020 73.950 23.030 ;
        RECT 76.710 23.020 76.850 23.030 ;
        RECT 79.610 23.020 79.750 23.030 ;
        RECT 82.510 23.020 82.650 23.030 ;
        RECT 85.410 23.020 85.550 23.030 ;
        RECT 88.310 23.020 88.450 23.030 ;
        RECT 91.210 23.020 91.350 23.030 ;
        RECT 1.300 22.950 1.460 23.020 ;
        RECT 4.200 22.950 4.360 23.020 ;
        RECT 7.100 22.950 7.260 23.020 ;
        RECT 10.000 22.950 10.160 23.020 ;
        RECT 12.900 22.950 13.060 23.020 ;
        RECT 15.800 22.950 15.960 23.020 ;
        RECT 18.700 22.950 18.860 23.020 ;
        RECT 21.600 22.950 21.760 23.020 ;
        RECT 24.500 22.950 24.660 23.020 ;
        RECT 27.400 22.950 27.560 23.020 ;
        RECT 30.300 22.950 30.460 23.020 ;
        RECT 33.200 22.950 33.360 23.020 ;
        RECT 36.100 22.950 36.260 23.020 ;
        RECT 39.000 22.950 39.160 23.020 ;
        RECT 41.900 22.950 42.060 23.020 ;
        RECT 44.800 22.950 44.960 23.020 ;
        RECT 47.700 22.950 47.860 23.020 ;
        RECT 50.600 22.950 50.760 23.020 ;
        RECT 53.500 22.950 53.660 23.020 ;
        RECT 56.400 22.950 56.560 23.020 ;
        RECT 59.300 22.950 59.460 23.020 ;
        RECT 62.200 22.950 62.360 23.020 ;
        RECT 65.100 22.950 65.260 23.020 ;
        RECT 68.000 22.950 68.160 23.020 ;
        RECT 70.900 22.950 71.060 23.020 ;
        RECT 73.800 22.950 73.960 23.020 ;
        RECT 76.700 22.950 76.860 23.020 ;
        RECT 79.600 22.950 79.760 23.020 ;
        RECT 82.500 22.950 82.660 23.020 ;
        RECT 85.400 22.950 85.560 23.020 ;
        RECT 88.300 22.950 88.460 23.020 ;
        RECT 91.200 22.950 91.360 23.020 ;
        RECT 1.310 21.670 1.450 21.680 ;
        RECT 4.210 21.670 4.350 21.680 ;
        RECT 7.110 21.670 7.250 21.680 ;
        RECT 10.010 21.670 10.150 21.680 ;
        RECT 12.910 21.670 13.050 21.680 ;
        RECT 15.810 21.670 15.950 21.680 ;
        RECT 18.710 21.670 18.850 21.680 ;
        RECT 21.610 21.670 21.750 21.680 ;
        RECT 24.510 21.670 24.650 21.680 ;
        RECT 27.410 21.670 27.550 21.680 ;
        RECT 30.310 21.670 30.450 21.680 ;
        RECT 33.210 21.670 33.350 21.680 ;
        RECT 36.110 21.670 36.250 21.680 ;
        RECT 39.010 21.670 39.150 21.680 ;
        RECT 41.910 21.670 42.050 21.680 ;
        RECT 44.810 21.670 44.950 21.680 ;
        RECT 47.710 21.670 47.850 21.680 ;
        RECT 50.610 21.670 50.750 21.680 ;
        RECT 53.510 21.670 53.650 21.680 ;
        RECT 56.410 21.670 56.550 21.680 ;
        RECT 59.310 21.670 59.450 21.680 ;
        RECT 62.210 21.670 62.350 21.680 ;
        RECT 65.110 21.670 65.250 21.680 ;
        RECT 68.010 21.670 68.150 21.680 ;
        RECT 70.910 21.670 71.050 21.680 ;
        RECT 73.810 21.670 73.950 21.680 ;
        RECT 76.710 21.670 76.850 21.680 ;
        RECT 79.610 21.670 79.750 21.680 ;
        RECT 82.510 21.670 82.650 21.680 ;
        RECT 85.410 21.670 85.550 21.680 ;
        RECT 88.310 21.670 88.450 21.680 ;
        RECT 91.210 21.670 91.350 21.680 ;
        RECT 1.300 21.600 1.460 21.670 ;
        RECT 4.200 21.600 4.360 21.670 ;
        RECT 7.100 21.600 7.260 21.670 ;
        RECT 10.000 21.600 10.160 21.670 ;
        RECT 12.900 21.600 13.060 21.670 ;
        RECT 15.800 21.600 15.960 21.670 ;
        RECT 18.700 21.600 18.860 21.670 ;
        RECT 21.600 21.600 21.760 21.670 ;
        RECT 24.500 21.600 24.660 21.670 ;
        RECT 27.400 21.600 27.560 21.670 ;
        RECT 30.300 21.600 30.460 21.670 ;
        RECT 33.200 21.600 33.360 21.670 ;
        RECT 36.100 21.600 36.260 21.670 ;
        RECT 39.000 21.600 39.160 21.670 ;
        RECT 41.900 21.600 42.060 21.670 ;
        RECT 44.800 21.600 44.960 21.670 ;
        RECT 47.700 21.600 47.860 21.670 ;
        RECT 50.600 21.600 50.760 21.670 ;
        RECT 53.500 21.600 53.660 21.670 ;
        RECT 56.400 21.600 56.560 21.670 ;
        RECT 59.300 21.600 59.460 21.670 ;
        RECT 62.200 21.600 62.360 21.670 ;
        RECT 65.100 21.600 65.260 21.670 ;
        RECT 68.000 21.600 68.160 21.670 ;
        RECT 70.900 21.600 71.060 21.670 ;
        RECT 73.800 21.600 73.960 21.670 ;
        RECT 76.700 21.600 76.860 21.670 ;
        RECT 79.600 21.600 79.760 21.670 ;
        RECT 82.500 21.600 82.660 21.670 ;
        RECT 85.400 21.600 85.560 21.670 ;
        RECT 88.300 21.600 88.460 21.670 ;
        RECT 91.200 21.600 91.360 21.670 ;
        RECT 1.310 20.320 1.450 20.330 ;
        RECT 4.210 20.320 4.350 20.330 ;
        RECT 7.110 20.320 7.250 20.330 ;
        RECT 10.010 20.320 10.150 20.330 ;
        RECT 12.910 20.320 13.050 20.330 ;
        RECT 15.810 20.320 15.950 20.330 ;
        RECT 18.710 20.320 18.850 20.330 ;
        RECT 21.610 20.320 21.750 20.330 ;
        RECT 24.510 20.320 24.650 20.330 ;
        RECT 27.410 20.320 27.550 20.330 ;
        RECT 30.310 20.320 30.450 20.330 ;
        RECT 33.210 20.320 33.350 20.330 ;
        RECT 36.110 20.320 36.250 20.330 ;
        RECT 39.010 20.320 39.150 20.330 ;
        RECT 41.910 20.320 42.050 20.330 ;
        RECT 44.810 20.320 44.950 20.330 ;
        RECT 47.710 20.320 47.850 20.330 ;
        RECT 50.610 20.320 50.750 20.330 ;
        RECT 53.510 20.320 53.650 20.330 ;
        RECT 56.410 20.320 56.550 20.330 ;
        RECT 59.310 20.320 59.450 20.330 ;
        RECT 62.210 20.320 62.350 20.330 ;
        RECT 65.110 20.320 65.250 20.330 ;
        RECT 68.010 20.320 68.150 20.330 ;
        RECT 70.910 20.320 71.050 20.330 ;
        RECT 73.810 20.320 73.950 20.330 ;
        RECT 76.710 20.320 76.850 20.330 ;
        RECT 79.610 20.320 79.750 20.330 ;
        RECT 82.510 20.320 82.650 20.330 ;
        RECT 85.410 20.320 85.550 20.330 ;
        RECT 88.310 20.320 88.450 20.330 ;
        RECT 91.210 20.320 91.350 20.330 ;
        RECT 1.300 20.250 1.460 20.320 ;
        RECT 4.200 20.250 4.360 20.320 ;
        RECT 7.100 20.250 7.260 20.320 ;
        RECT 10.000 20.250 10.160 20.320 ;
        RECT 12.900 20.250 13.060 20.320 ;
        RECT 15.800 20.250 15.960 20.320 ;
        RECT 18.700 20.250 18.860 20.320 ;
        RECT 21.600 20.250 21.760 20.320 ;
        RECT 24.500 20.250 24.660 20.320 ;
        RECT 27.400 20.250 27.560 20.320 ;
        RECT 30.300 20.250 30.460 20.320 ;
        RECT 33.200 20.250 33.360 20.320 ;
        RECT 36.100 20.250 36.260 20.320 ;
        RECT 39.000 20.250 39.160 20.320 ;
        RECT 41.900 20.250 42.060 20.320 ;
        RECT 44.800 20.250 44.960 20.320 ;
        RECT 47.700 20.250 47.860 20.320 ;
        RECT 50.600 20.250 50.760 20.320 ;
        RECT 53.500 20.250 53.660 20.320 ;
        RECT 56.400 20.250 56.560 20.320 ;
        RECT 59.300 20.250 59.460 20.320 ;
        RECT 62.200 20.250 62.360 20.320 ;
        RECT 65.100 20.250 65.260 20.320 ;
        RECT 68.000 20.250 68.160 20.320 ;
        RECT 70.900 20.250 71.060 20.320 ;
        RECT 73.800 20.250 73.960 20.320 ;
        RECT 76.700 20.250 76.860 20.320 ;
        RECT 79.600 20.250 79.760 20.320 ;
        RECT 82.500 20.250 82.660 20.320 ;
        RECT 85.400 20.250 85.560 20.320 ;
        RECT 88.300 20.250 88.460 20.320 ;
        RECT 91.200 20.250 91.360 20.320 ;
        RECT 1.310 18.970 1.450 18.980 ;
        RECT 4.210 18.970 4.350 18.980 ;
        RECT 7.110 18.970 7.250 18.980 ;
        RECT 10.010 18.970 10.150 18.980 ;
        RECT 12.910 18.970 13.050 18.980 ;
        RECT 15.810 18.970 15.950 18.980 ;
        RECT 18.710 18.970 18.850 18.980 ;
        RECT 21.610 18.970 21.750 18.980 ;
        RECT 24.510 18.970 24.650 18.980 ;
        RECT 27.410 18.970 27.550 18.980 ;
        RECT 30.310 18.970 30.450 18.980 ;
        RECT 33.210 18.970 33.350 18.980 ;
        RECT 36.110 18.970 36.250 18.980 ;
        RECT 39.010 18.970 39.150 18.980 ;
        RECT 41.910 18.970 42.050 18.980 ;
        RECT 44.810 18.970 44.950 18.980 ;
        RECT 47.710 18.970 47.850 18.980 ;
        RECT 50.610 18.970 50.750 18.980 ;
        RECT 53.510 18.970 53.650 18.980 ;
        RECT 56.410 18.970 56.550 18.980 ;
        RECT 59.310 18.970 59.450 18.980 ;
        RECT 62.210 18.970 62.350 18.980 ;
        RECT 65.110 18.970 65.250 18.980 ;
        RECT 68.010 18.970 68.150 18.980 ;
        RECT 70.910 18.970 71.050 18.980 ;
        RECT 73.810 18.970 73.950 18.980 ;
        RECT 76.710 18.970 76.850 18.980 ;
        RECT 79.610 18.970 79.750 18.980 ;
        RECT 82.510 18.970 82.650 18.980 ;
        RECT 85.410 18.970 85.550 18.980 ;
        RECT 88.310 18.970 88.450 18.980 ;
        RECT 91.210 18.970 91.350 18.980 ;
        RECT 1.300 18.900 1.460 18.970 ;
        RECT 4.200 18.900 4.360 18.970 ;
        RECT 7.100 18.900 7.260 18.970 ;
        RECT 10.000 18.900 10.160 18.970 ;
        RECT 12.900 18.900 13.060 18.970 ;
        RECT 15.800 18.900 15.960 18.970 ;
        RECT 18.700 18.900 18.860 18.970 ;
        RECT 21.600 18.900 21.760 18.970 ;
        RECT 24.500 18.900 24.660 18.970 ;
        RECT 27.400 18.900 27.560 18.970 ;
        RECT 30.300 18.900 30.460 18.970 ;
        RECT 33.200 18.900 33.360 18.970 ;
        RECT 36.100 18.900 36.260 18.970 ;
        RECT 39.000 18.900 39.160 18.970 ;
        RECT 41.900 18.900 42.060 18.970 ;
        RECT 44.800 18.900 44.960 18.970 ;
        RECT 47.700 18.900 47.860 18.970 ;
        RECT 50.600 18.900 50.760 18.970 ;
        RECT 53.500 18.900 53.660 18.970 ;
        RECT 56.400 18.900 56.560 18.970 ;
        RECT 59.300 18.900 59.460 18.970 ;
        RECT 62.200 18.900 62.360 18.970 ;
        RECT 65.100 18.900 65.260 18.970 ;
        RECT 68.000 18.900 68.160 18.970 ;
        RECT 70.900 18.900 71.060 18.970 ;
        RECT 73.800 18.900 73.960 18.970 ;
        RECT 76.700 18.900 76.860 18.970 ;
        RECT 79.600 18.900 79.760 18.970 ;
        RECT 82.500 18.900 82.660 18.970 ;
        RECT 85.400 18.900 85.560 18.970 ;
        RECT 88.300 18.900 88.460 18.970 ;
        RECT 91.200 18.900 91.360 18.970 ;
        RECT 1.310 17.620 1.450 17.630 ;
        RECT 4.210 17.620 4.350 17.630 ;
        RECT 7.110 17.620 7.250 17.630 ;
        RECT 10.010 17.620 10.150 17.630 ;
        RECT 12.910 17.620 13.050 17.630 ;
        RECT 15.810 17.620 15.950 17.630 ;
        RECT 18.710 17.620 18.850 17.630 ;
        RECT 21.610 17.620 21.750 17.630 ;
        RECT 24.510 17.620 24.650 17.630 ;
        RECT 27.410 17.620 27.550 17.630 ;
        RECT 30.310 17.620 30.450 17.630 ;
        RECT 33.210 17.620 33.350 17.630 ;
        RECT 36.110 17.620 36.250 17.630 ;
        RECT 39.010 17.620 39.150 17.630 ;
        RECT 41.910 17.620 42.050 17.630 ;
        RECT 44.810 17.620 44.950 17.630 ;
        RECT 47.710 17.620 47.850 17.630 ;
        RECT 50.610 17.620 50.750 17.630 ;
        RECT 53.510 17.620 53.650 17.630 ;
        RECT 56.410 17.620 56.550 17.630 ;
        RECT 59.310 17.620 59.450 17.630 ;
        RECT 62.210 17.620 62.350 17.630 ;
        RECT 65.110 17.620 65.250 17.630 ;
        RECT 68.010 17.620 68.150 17.630 ;
        RECT 70.910 17.620 71.050 17.630 ;
        RECT 73.810 17.620 73.950 17.630 ;
        RECT 76.710 17.620 76.850 17.630 ;
        RECT 79.610 17.620 79.750 17.630 ;
        RECT 82.510 17.620 82.650 17.630 ;
        RECT 85.410 17.620 85.550 17.630 ;
        RECT 88.310 17.620 88.450 17.630 ;
        RECT 91.210 17.620 91.350 17.630 ;
        RECT 1.300 17.550 1.460 17.620 ;
        RECT 4.200 17.550 4.360 17.620 ;
        RECT 7.100 17.550 7.260 17.620 ;
        RECT 10.000 17.550 10.160 17.620 ;
        RECT 12.900 17.550 13.060 17.620 ;
        RECT 15.800 17.550 15.960 17.620 ;
        RECT 18.700 17.550 18.860 17.620 ;
        RECT 21.600 17.550 21.760 17.620 ;
        RECT 24.500 17.550 24.660 17.620 ;
        RECT 27.400 17.550 27.560 17.620 ;
        RECT 30.300 17.550 30.460 17.620 ;
        RECT 33.200 17.550 33.360 17.620 ;
        RECT 36.100 17.550 36.260 17.620 ;
        RECT 39.000 17.550 39.160 17.620 ;
        RECT 41.900 17.550 42.060 17.620 ;
        RECT 44.800 17.550 44.960 17.620 ;
        RECT 47.700 17.550 47.860 17.620 ;
        RECT 50.600 17.550 50.760 17.620 ;
        RECT 53.500 17.550 53.660 17.620 ;
        RECT 56.400 17.550 56.560 17.620 ;
        RECT 59.300 17.550 59.460 17.620 ;
        RECT 62.200 17.550 62.360 17.620 ;
        RECT 65.100 17.550 65.260 17.620 ;
        RECT 68.000 17.550 68.160 17.620 ;
        RECT 70.900 17.550 71.060 17.620 ;
        RECT 73.800 17.550 73.960 17.620 ;
        RECT 76.700 17.550 76.860 17.620 ;
        RECT 79.600 17.550 79.760 17.620 ;
        RECT 82.500 17.550 82.660 17.620 ;
        RECT 85.400 17.550 85.560 17.620 ;
        RECT 88.300 17.550 88.460 17.620 ;
        RECT 91.200 17.550 91.360 17.620 ;
        RECT 1.310 16.270 1.450 16.280 ;
        RECT 4.210 16.270 4.350 16.280 ;
        RECT 7.110 16.270 7.250 16.280 ;
        RECT 10.010 16.270 10.150 16.280 ;
        RECT 12.910 16.270 13.050 16.280 ;
        RECT 15.810 16.270 15.950 16.280 ;
        RECT 18.710 16.270 18.850 16.280 ;
        RECT 21.610 16.270 21.750 16.280 ;
        RECT 24.510 16.270 24.650 16.280 ;
        RECT 27.410 16.270 27.550 16.280 ;
        RECT 30.310 16.270 30.450 16.280 ;
        RECT 33.210 16.270 33.350 16.280 ;
        RECT 36.110 16.270 36.250 16.280 ;
        RECT 39.010 16.270 39.150 16.280 ;
        RECT 41.910 16.270 42.050 16.280 ;
        RECT 44.810 16.270 44.950 16.280 ;
        RECT 47.710 16.270 47.850 16.280 ;
        RECT 50.610 16.270 50.750 16.280 ;
        RECT 53.510 16.270 53.650 16.280 ;
        RECT 56.410 16.270 56.550 16.280 ;
        RECT 59.310 16.270 59.450 16.280 ;
        RECT 62.210 16.270 62.350 16.280 ;
        RECT 65.110 16.270 65.250 16.280 ;
        RECT 68.010 16.270 68.150 16.280 ;
        RECT 70.910 16.270 71.050 16.280 ;
        RECT 73.810 16.270 73.950 16.280 ;
        RECT 76.710 16.270 76.850 16.280 ;
        RECT 79.610 16.270 79.750 16.280 ;
        RECT 82.510 16.270 82.650 16.280 ;
        RECT 85.410 16.270 85.550 16.280 ;
        RECT 88.310 16.270 88.450 16.280 ;
        RECT 91.210 16.270 91.350 16.280 ;
        RECT 1.300 16.200 1.460 16.270 ;
        RECT 4.200 16.200 4.360 16.270 ;
        RECT 7.100 16.200 7.260 16.270 ;
        RECT 10.000 16.200 10.160 16.270 ;
        RECT 12.900 16.200 13.060 16.270 ;
        RECT 15.800 16.200 15.960 16.270 ;
        RECT 18.700 16.200 18.860 16.270 ;
        RECT 21.600 16.200 21.760 16.270 ;
        RECT 24.500 16.200 24.660 16.270 ;
        RECT 27.400 16.200 27.560 16.270 ;
        RECT 30.300 16.200 30.460 16.270 ;
        RECT 33.200 16.200 33.360 16.270 ;
        RECT 36.100 16.200 36.260 16.270 ;
        RECT 39.000 16.200 39.160 16.270 ;
        RECT 41.900 16.200 42.060 16.270 ;
        RECT 44.800 16.200 44.960 16.270 ;
        RECT 47.700 16.200 47.860 16.270 ;
        RECT 50.600 16.200 50.760 16.270 ;
        RECT 53.500 16.200 53.660 16.270 ;
        RECT 56.400 16.200 56.560 16.270 ;
        RECT 59.300 16.200 59.460 16.270 ;
        RECT 62.200 16.200 62.360 16.270 ;
        RECT 65.100 16.200 65.260 16.270 ;
        RECT 68.000 16.200 68.160 16.270 ;
        RECT 70.900 16.200 71.060 16.270 ;
        RECT 73.800 16.200 73.960 16.270 ;
        RECT 76.700 16.200 76.860 16.270 ;
        RECT 79.600 16.200 79.760 16.270 ;
        RECT 82.500 16.200 82.660 16.270 ;
        RECT 85.400 16.200 85.560 16.270 ;
        RECT 88.300 16.200 88.460 16.270 ;
        RECT 91.200 16.200 91.360 16.270 ;
        RECT 1.310 14.920 1.450 14.930 ;
        RECT 4.210 14.920 4.350 14.930 ;
        RECT 7.110 14.920 7.250 14.930 ;
        RECT 10.010 14.920 10.150 14.930 ;
        RECT 12.910 14.920 13.050 14.930 ;
        RECT 15.810 14.920 15.950 14.930 ;
        RECT 18.710 14.920 18.850 14.930 ;
        RECT 21.610 14.920 21.750 14.930 ;
        RECT 24.510 14.920 24.650 14.930 ;
        RECT 27.410 14.920 27.550 14.930 ;
        RECT 30.310 14.920 30.450 14.930 ;
        RECT 33.210 14.920 33.350 14.930 ;
        RECT 36.110 14.920 36.250 14.930 ;
        RECT 39.010 14.920 39.150 14.930 ;
        RECT 41.910 14.920 42.050 14.930 ;
        RECT 44.810 14.920 44.950 14.930 ;
        RECT 47.710 14.920 47.850 14.930 ;
        RECT 50.610 14.920 50.750 14.930 ;
        RECT 53.510 14.920 53.650 14.930 ;
        RECT 56.410 14.920 56.550 14.930 ;
        RECT 59.310 14.920 59.450 14.930 ;
        RECT 62.210 14.920 62.350 14.930 ;
        RECT 65.110 14.920 65.250 14.930 ;
        RECT 68.010 14.920 68.150 14.930 ;
        RECT 70.910 14.920 71.050 14.930 ;
        RECT 73.810 14.920 73.950 14.930 ;
        RECT 76.710 14.920 76.850 14.930 ;
        RECT 79.610 14.920 79.750 14.930 ;
        RECT 82.510 14.920 82.650 14.930 ;
        RECT 85.410 14.920 85.550 14.930 ;
        RECT 88.310 14.920 88.450 14.930 ;
        RECT 91.210 14.920 91.350 14.930 ;
        RECT 1.300 14.850 1.460 14.920 ;
        RECT 4.200 14.850 4.360 14.920 ;
        RECT 7.100 14.850 7.260 14.920 ;
        RECT 10.000 14.850 10.160 14.920 ;
        RECT 12.900 14.850 13.060 14.920 ;
        RECT 15.800 14.850 15.960 14.920 ;
        RECT 18.700 14.850 18.860 14.920 ;
        RECT 21.600 14.850 21.760 14.920 ;
        RECT 24.500 14.850 24.660 14.920 ;
        RECT 27.400 14.850 27.560 14.920 ;
        RECT 30.300 14.850 30.460 14.920 ;
        RECT 33.200 14.850 33.360 14.920 ;
        RECT 36.100 14.850 36.260 14.920 ;
        RECT 39.000 14.850 39.160 14.920 ;
        RECT 41.900 14.850 42.060 14.920 ;
        RECT 44.800 14.850 44.960 14.920 ;
        RECT 47.700 14.850 47.860 14.920 ;
        RECT 50.600 14.850 50.760 14.920 ;
        RECT 53.500 14.850 53.660 14.920 ;
        RECT 56.400 14.850 56.560 14.920 ;
        RECT 59.300 14.850 59.460 14.920 ;
        RECT 62.200 14.850 62.360 14.920 ;
        RECT 65.100 14.850 65.260 14.920 ;
        RECT 68.000 14.850 68.160 14.920 ;
        RECT 70.900 14.850 71.060 14.920 ;
        RECT 73.800 14.850 73.960 14.920 ;
        RECT 76.700 14.850 76.860 14.920 ;
        RECT 79.600 14.850 79.760 14.920 ;
        RECT 82.500 14.850 82.660 14.920 ;
        RECT 85.400 14.850 85.560 14.920 ;
        RECT 88.300 14.850 88.460 14.920 ;
        RECT 91.200 14.850 91.360 14.920 ;
        RECT 1.310 13.570 1.450 13.580 ;
        RECT 4.210 13.570 4.350 13.580 ;
        RECT 7.110 13.570 7.250 13.580 ;
        RECT 10.010 13.570 10.150 13.580 ;
        RECT 12.910 13.570 13.050 13.580 ;
        RECT 15.810 13.570 15.950 13.580 ;
        RECT 18.710 13.570 18.850 13.580 ;
        RECT 21.610 13.570 21.750 13.580 ;
        RECT 24.510 13.570 24.650 13.580 ;
        RECT 27.410 13.570 27.550 13.580 ;
        RECT 30.310 13.570 30.450 13.580 ;
        RECT 33.210 13.570 33.350 13.580 ;
        RECT 36.110 13.570 36.250 13.580 ;
        RECT 39.010 13.570 39.150 13.580 ;
        RECT 41.910 13.570 42.050 13.580 ;
        RECT 44.810 13.570 44.950 13.580 ;
        RECT 47.710 13.570 47.850 13.580 ;
        RECT 50.610 13.570 50.750 13.580 ;
        RECT 53.510 13.570 53.650 13.580 ;
        RECT 56.410 13.570 56.550 13.580 ;
        RECT 59.310 13.570 59.450 13.580 ;
        RECT 62.210 13.570 62.350 13.580 ;
        RECT 65.110 13.570 65.250 13.580 ;
        RECT 68.010 13.570 68.150 13.580 ;
        RECT 70.910 13.570 71.050 13.580 ;
        RECT 73.810 13.570 73.950 13.580 ;
        RECT 76.710 13.570 76.850 13.580 ;
        RECT 79.610 13.570 79.750 13.580 ;
        RECT 82.510 13.570 82.650 13.580 ;
        RECT 85.410 13.570 85.550 13.580 ;
        RECT 88.310 13.570 88.450 13.580 ;
        RECT 91.210 13.570 91.350 13.580 ;
        RECT 1.300 13.500 1.460 13.570 ;
        RECT 4.200 13.500 4.360 13.570 ;
        RECT 7.100 13.500 7.260 13.570 ;
        RECT 10.000 13.500 10.160 13.570 ;
        RECT 12.900 13.500 13.060 13.570 ;
        RECT 15.800 13.500 15.960 13.570 ;
        RECT 18.700 13.500 18.860 13.570 ;
        RECT 21.600 13.500 21.760 13.570 ;
        RECT 24.500 13.500 24.660 13.570 ;
        RECT 27.400 13.500 27.560 13.570 ;
        RECT 30.300 13.500 30.460 13.570 ;
        RECT 33.200 13.500 33.360 13.570 ;
        RECT 36.100 13.500 36.260 13.570 ;
        RECT 39.000 13.500 39.160 13.570 ;
        RECT 41.900 13.500 42.060 13.570 ;
        RECT 44.800 13.500 44.960 13.570 ;
        RECT 47.700 13.500 47.860 13.570 ;
        RECT 50.600 13.500 50.760 13.570 ;
        RECT 53.500 13.500 53.660 13.570 ;
        RECT 56.400 13.500 56.560 13.570 ;
        RECT 59.300 13.500 59.460 13.570 ;
        RECT 62.200 13.500 62.360 13.570 ;
        RECT 65.100 13.500 65.260 13.570 ;
        RECT 68.000 13.500 68.160 13.570 ;
        RECT 70.900 13.500 71.060 13.570 ;
        RECT 73.800 13.500 73.960 13.570 ;
        RECT 76.700 13.500 76.860 13.570 ;
        RECT 79.600 13.500 79.760 13.570 ;
        RECT 82.500 13.500 82.660 13.570 ;
        RECT 85.400 13.500 85.560 13.570 ;
        RECT 88.300 13.500 88.460 13.570 ;
        RECT 91.200 13.500 91.360 13.570 ;
        RECT 1.310 12.220 1.450 12.230 ;
        RECT 4.210 12.220 4.350 12.230 ;
        RECT 7.110 12.220 7.250 12.230 ;
        RECT 10.010 12.220 10.150 12.230 ;
        RECT 12.910 12.220 13.050 12.230 ;
        RECT 15.810 12.220 15.950 12.230 ;
        RECT 18.710 12.220 18.850 12.230 ;
        RECT 21.610 12.220 21.750 12.230 ;
        RECT 24.510 12.220 24.650 12.230 ;
        RECT 27.410 12.220 27.550 12.230 ;
        RECT 30.310 12.220 30.450 12.230 ;
        RECT 33.210 12.220 33.350 12.230 ;
        RECT 36.110 12.220 36.250 12.230 ;
        RECT 39.010 12.220 39.150 12.230 ;
        RECT 41.910 12.220 42.050 12.230 ;
        RECT 44.810 12.220 44.950 12.230 ;
        RECT 47.710 12.220 47.850 12.230 ;
        RECT 50.610 12.220 50.750 12.230 ;
        RECT 53.510 12.220 53.650 12.230 ;
        RECT 56.410 12.220 56.550 12.230 ;
        RECT 59.310 12.220 59.450 12.230 ;
        RECT 62.210 12.220 62.350 12.230 ;
        RECT 65.110 12.220 65.250 12.230 ;
        RECT 68.010 12.220 68.150 12.230 ;
        RECT 70.910 12.220 71.050 12.230 ;
        RECT 73.810 12.220 73.950 12.230 ;
        RECT 76.710 12.220 76.850 12.230 ;
        RECT 79.610 12.220 79.750 12.230 ;
        RECT 82.510 12.220 82.650 12.230 ;
        RECT 85.410 12.220 85.550 12.230 ;
        RECT 88.310 12.220 88.450 12.230 ;
        RECT 91.210 12.220 91.350 12.230 ;
        RECT 1.300 12.150 1.460 12.220 ;
        RECT 4.200 12.150 4.360 12.220 ;
        RECT 7.100 12.150 7.260 12.220 ;
        RECT 10.000 12.150 10.160 12.220 ;
        RECT 12.900 12.150 13.060 12.220 ;
        RECT 15.800 12.150 15.960 12.220 ;
        RECT 18.700 12.150 18.860 12.220 ;
        RECT 21.600 12.150 21.760 12.220 ;
        RECT 24.500 12.150 24.660 12.220 ;
        RECT 27.400 12.150 27.560 12.220 ;
        RECT 30.300 12.150 30.460 12.220 ;
        RECT 33.200 12.150 33.360 12.220 ;
        RECT 36.100 12.150 36.260 12.220 ;
        RECT 39.000 12.150 39.160 12.220 ;
        RECT 41.900 12.150 42.060 12.220 ;
        RECT 44.800 12.150 44.960 12.220 ;
        RECT 47.700 12.150 47.860 12.220 ;
        RECT 50.600 12.150 50.760 12.220 ;
        RECT 53.500 12.150 53.660 12.220 ;
        RECT 56.400 12.150 56.560 12.220 ;
        RECT 59.300 12.150 59.460 12.220 ;
        RECT 62.200 12.150 62.360 12.220 ;
        RECT 65.100 12.150 65.260 12.220 ;
        RECT 68.000 12.150 68.160 12.220 ;
        RECT 70.900 12.150 71.060 12.220 ;
        RECT 73.800 12.150 73.960 12.220 ;
        RECT 76.700 12.150 76.860 12.220 ;
        RECT 79.600 12.150 79.760 12.220 ;
        RECT 82.500 12.150 82.660 12.220 ;
        RECT 85.400 12.150 85.560 12.220 ;
        RECT 88.300 12.150 88.460 12.220 ;
        RECT 91.200 12.150 91.360 12.220 ;
        RECT 1.310 10.870 1.450 10.880 ;
        RECT 4.210 10.870 4.350 10.880 ;
        RECT 7.110 10.870 7.250 10.880 ;
        RECT 10.010 10.870 10.150 10.880 ;
        RECT 12.910 10.870 13.050 10.880 ;
        RECT 15.810 10.870 15.950 10.880 ;
        RECT 18.710 10.870 18.850 10.880 ;
        RECT 21.610 10.870 21.750 10.880 ;
        RECT 24.510 10.870 24.650 10.880 ;
        RECT 27.410 10.870 27.550 10.880 ;
        RECT 30.310 10.870 30.450 10.880 ;
        RECT 33.210 10.870 33.350 10.880 ;
        RECT 36.110 10.870 36.250 10.880 ;
        RECT 39.010 10.870 39.150 10.880 ;
        RECT 41.910 10.870 42.050 10.880 ;
        RECT 44.810 10.870 44.950 10.880 ;
        RECT 47.710 10.870 47.850 10.880 ;
        RECT 50.610 10.870 50.750 10.880 ;
        RECT 53.510 10.870 53.650 10.880 ;
        RECT 56.410 10.870 56.550 10.880 ;
        RECT 59.310 10.870 59.450 10.880 ;
        RECT 62.210 10.870 62.350 10.880 ;
        RECT 65.110 10.870 65.250 10.880 ;
        RECT 68.010 10.870 68.150 10.880 ;
        RECT 70.910 10.870 71.050 10.880 ;
        RECT 73.810 10.870 73.950 10.880 ;
        RECT 76.710 10.870 76.850 10.880 ;
        RECT 79.610 10.870 79.750 10.880 ;
        RECT 82.510 10.870 82.650 10.880 ;
        RECT 85.410 10.870 85.550 10.880 ;
        RECT 88.310 10.870 88.450 10.880 ;
        RECT 91.210 10.870 91.350 10.880 ;
        RECT 1.300 10.800 1.460 10.870 ;
        RECT 4.200 10.800 4.360 10.870 ;
        RECT 7.100 10.800 7.260 10.870 ;
        RECT 10.000 10.800 10.160 10.870 ;
        RECT 12.900 10.800 13.060 10.870 ;
        RECT 15.800 10.800 15.960 10.870 ;
        RECT 18.700 10.800 18.860 10.870 ;
        RECT 21.600 10.800 21.760 10.870 ;
        RECT 24.500 10.800 24.660 10.870 ;
        RECT 27.400 10.800 27.560 10.870 ;
        RECT 30.300 10.800 30.460 10.870 ;
        RECT 33.200 10.800 33.360 10.870 ;
        RECT 36.100 10.800 36.260 10.870 ;
        RECT 39.000 10.800 39.160 10.870 ;
        RECT 41.900 10.800 42.060 10.870 ;
        RECT 44.800 10.800 44.960 10.870 ;
        RECT 47.700 10.800 47.860 10.870 ;
        RECT 50.600 10.800 50.760 10.870 ;
        RECT 53.500 10.800 53.660 10.870 ;
        RECT 56.400 10.800 56.560 10.870 ;
        RECT 59.300 10.800 59.460 10.870 ;
        RECT 62.200 10.800 62.360 10.870 ;
        RECT 65.100 10.800 65.260 10.870 ;
        RECT 68.000 10.800 68.160 10.870 ;
        RECT 70.900 10.800 71.060 10.870 ;
        RECT 73.800 10.800 73.960 10.870 ;
        RECT 76.700 10.800 76.860 10.870 ;
        RECT 79.600 10.800 79.760 10.870 ;
        RECT 82.500 10.800 82.660 10.870 ;
        RECT 85.400 10.800 85.560 10.870 ;
        RECT 88.300 10.800 88.460 10.870 ;
        RECT 91.200 10.800 91.360 10.870 ;
        RECT 1.310 9.520 1.450 9.530 ;
        RECT 4.210 9.520 4.350 9.530 ;
        RECT 7.110 9.520 7.250 9.530 ;
        RECT 10.010 9.520 10.150 9.530 ;
        RECT 12.910 9.520 13.050 9.530 ;
        RECT 15.810 9.520 15.950 9.530 ;
        RECT 18.710 9.520 18.850 9.530 ;
        RECT 21.610 9.520 21.750 9.530 ;
        RECT 24.510 9.520 24.650 9.530 ;
        RECT 27.410 9.520 27.550 9.530 ;
        RECT 30.310 9.520 30.450 9.530 ;
        RECT 33.210 9.520 33.350 9.530 ;
        RECT 36.110 9.520 36.250 9.530 ;
        RECT 39.010 9.520 39.150 9.530 ;
        RECT 41.910 9.520 42.050 9.530 ;
        RECT 44.810 9.520 44.950 9.530 ;
        RECT 47.710 9.520 47.850 9.530 ;
        RECT 50.610 9.520 50.750 9.530 ;
        RECT 53.510 9.520 53.650 9.530 ;
        RECT 56.410 9.520 56.550 9.530 ;
        RECT 59.310 9.520 59.450 9.530 ;
        RECT 62.210 9.520 62.350 9.530 ;
        RECT 65.110 9.520 65.250 9.530 ;
        RECT 68.010 9.520 68.150 9.530 ;
        RECT 70.910 9.520 71.050 9.530 ;
        RECT 73.810 9.520 73.950 9.530 ;
        RECT 76.710 9.520 76.850 9.530 ;
        RECT 79.610 9.520 79.750 9.530 ;
        RECT 82.510 9.520 82.650 9.530 ;
        RECT 85.410 9.520 85.550 9.530 ;
        RECT 88.310 9.520 88.450 9.530 ;
        RECT 91.210 9.520 91.350 9.530 ;
        RECT 1.300 9.450 1.460 9.520 ;
        RECT 4.200 9.450 4.360 9.520 ;
        RECT 7.100 9.450 7.260 9.520 ;
        RECT 10.000 9.450 10.160 9.520 ;
        RECT 12.900 9.450 13.060 9.520 ;
        RECT 15.800 9.450 15.960 9.520 ;
        RECT 18.700 9.450 18.860 9.520 ;
        RECT 21.600 9.450 21.760 9.520 ;
        RECT 24.500 9.450 24.660 9.520 ;
        RECT 27.400 9.450 27.560 9.520 ;
        RECT 30.300 9.450 30.460 9.520 ;
        RECT 33.200 9.450 33.360 9.520 ;
        RECT 36.100 9.450 36.260 9.520 ;
        RECT 39.000 9.450 39.160 9.520 ;
        RECT 41.900 9.450 42.060 9.520 ;
        RECT 44.800 9.450 44.960 9.520 ;
        RECT 47.700 9.450 47.860 9.520 ;
        RECT 50.600 9.450 50.760 9.520 ;
        RECT 53.500 9.450 53.660 9.520 ;
        RECT 56.400 9.450 56.560 9.520 ;
        RECT 59.300 9.450 59.460 9.520 ;
        RECT 62.200 9.450 62.360 9.520 ;
        RECT 65.100 9.450 65.260 9.520 ;
        RECT 68.000 9.450 68.160 9.520 ;
        RECT 70.900 9.450 71.060 9.520 ;
        RECT 73.800 9.450 73.960 9.520 ;
        RECT 76.700 9.450 76.860 9.520 ;
        RECT 79.600 9.450 79.760 9.520 ;
        RECT 82.500 9.450 82.660 9.520 ;
        RECT 85.400 9.450 85.560 9.520 ;
        RECT 88.300 9.450 88.460 9.520 ;
        RECT 91.200 9.450 91.360 9.520 ;
        RECT 1.310 8.170 1.450 8.180 ;
        RECT 4.210 8.170 4.350 8.180 ;
        RECT 7.110 8.170 7.250 8.180 ;
        RECT 10.010 8.170 10.150 8.180 ;
        RECT 12.910 8.170 13.050 8.180 ;
        RECT 15.810 8.170 15.950 8.180 ;
        RECT 18.710 8.170 18.850 8.180 ;
        RECT 21.610 8.170 21.750 8.180 ;
        RECT 24.510 8.170 24.650 8.180 ;
        RECT 27.410 8.170 27.550 8.180 ;
        RECT 30.310 8.170 30.450 8.180 ;
        RECT 33.210 8.170 33.350 8.180 ;
        RECT 36.110 8.170 36.250 8.180 ;
        RECT 39.010 8.170 39.150 8.180 ;
        RECT 41.910 8.170 42.050 8.180 ;
        RECT 44.810 8.170 44.950 8.180 ;
        RECT 47.710 8.170 47.850 8.180 ;
        RECT 50.610 8.170 50.750 8.180 ;
        RECT 53.510 8.170 53.650 8.180 ;
        RECT 56.410 8.170 56.550 8.180 ;
        RECT 59.310 8.170 59.450 8.180 ;
        RECT 62.210 8.170 62.350 8.180 ;
        RECT 65.110 8.170 65.250 8.180 ;
        RECT 68.010 8.170 68.150 8.180 ;
        RECT 70.910 8.170 71.050 8.180 ;
        RECT 73.810 8.170 73.950 8.180 ;
        RECT 76.710 8.170 76.850 8.180 ;
        RECT 79.610 8.170 79.750 8.180 ;
        RECT 82.510 8.170 82.650 8.180 ;
        RECT 85.410 8.170 85.550 8.180 ;
        RECT 88.310 8.170 88.450 8.180 ;
        RECT 91.210 8.170 91.350 8.180 ;
        RECT 1.300 8.100 1.460 8.170 ;
        RECT 4.200 8.100 4.360 8.170 ;
        RECT 7.100 8.100 7.260 8.170 ;
        RECT 10.000 8.100 10.160 8.170 ;
        RECT 12.900 8.100 13.060 8.170 ;
        RECT 15.800 8.100 15.960 8.170 ;
        RECT 18.700 8.100 18.860 8.170 ;
        RECT 21.600 8.100 21.760 8.170 ;
        RECT 24.500 8.100 24.660 8.170 ;
        RECT 27.400 8.100 27.560 8.170 ;
        RECT 30.300 8.100 30.460 8.170 ;
        RECT 33.200 8.100 33.360 8.170 ;
        RECT 36.100 8.100 36.260 8.170 ;
        RECT 39.000 8.100 39.160 8.170 ;
        RECT 41.900 8.100 42.060 8.170 ;
        RECT 44.800 8.100 44.960 8.170 ;
        RECT 47.700 8.100 47.860 8.170 ;
        RECT 50.600 8.100 50.760 8.170 ;
        RECT 53.500 8.100 53.660 8.170 ;
        RECT 56.400 8.100 56.560 8.170 ;
        RECT 59.300 8.100 59.460 8.170 ;
        RECT 62.200 8.100 62.360 8.170 ;
        RECT 65.100 8.100 65.260 8.170 ;
        RECT 68.000 8.100 68.160 8.170 ;
        RECT 70.900 8.100 71.060 8.170 ;
        RECT 73.800 8.100 73.960 8.170 ;
        RECT 76.700 8.100 76.860 8.170 ;
        RECT 79.600 8.100 79.760 8.170 ;
        RECT 82.500 8.100 82.660 8.170 ;
        RECT 85.400 8.100 85.560 8.170 ;
        RECT 88.300 8.100 88.460 8.170 ;
        RECT 91.200 8.100 91.360 8.170 ;
        RECT 1.310 6.820 1.450 6.830 ;
        RECT 4.210 6.820 4.350 6.830 ;
        RECT 7.110 6.820 7.250 6.830 ;
        RECT 10.010 6.820 10.150 6.830 ;
        RECT 12.910 6.820 13.050 6.830 ;
        RECT 15.810 6.820 15.950 6.830 ;
        RECT 18.710 6.820 18.850 6.830 ;
        RECT 21.610 6.820 21.750 6.830 ;
        RECT 24.510 6.820 24.650 6.830 ;
        RECT 27.410 6.820 27.550 6.830 ;
        RECT 30.310 6.820 30.450 6.830 ;
        RECT 33.210 6.820 33.350 6.830 ;
        RECT 36.110 6.820 36.250 6.830 ;
        RECT 39.010 6.820 39.150 6.830 ;
        RECT 41.910 6.820 42.050 6.830 ;
        RECT 44.810 6.820 44.950 6.830 ;
        RECT 47.710 6.820 47.850 6.830 ;
        RECT 50.610 6.820 50.750 6.830 ;
        RECT 53.510 6.820 53.650 6.830 ;
        RECT 56.410 6.820 56.550 6.830 ;
        RECT 59.310 6.820 59.450 6.830 ;
        RECT 62.210 6.820 62.350 6.830 ;
        RECT 65.110 6.820 65.250 6.830 ;
        RECT 68.010 6.820 68.150 6.830 ;
        RECT 70.910 6.820 71.050 6.830 ;
        RECT 73.810 6.820 73.950 6.830 ;
        RECT 76.710 6.820 76.850 6.830 ;
        RECT 79.610 6.820 79.750 6.830 ;
        RECT 82.510 6.820 82.650 6.830 ;
        RECT 85.410 6.820 85.550 6.830 ;
        RECT 88.310 6.820 88.450 6.830 ;
        RECT 91.210 6.820 91.350 6.830 ;
        RECT 1.300 6.750 1.460 6.820 ;
        RECT 4.200 6.750 4.360 6.820 ;
        RECT 7.100 6.750 7.260 6.820 ;
        RECT 10.000 6.750 10.160 6.820 ;
        RECT 12.900 6.750 13.060 6.820 ;
        RECT 15.800 6.750 15.960 6.820 ;
        RECT 18.700 6.750 18.860 6.820 ;
        RECT 21.600 6.750 21.760 6.820 ;
        RECT 24.500 6.750 24.660 6.820 ;
        RECT 27.400 6.750 27.560 6.820 ;
        RECT 30.300 6.750 30.460 6.820 ;
        RECT 33.200 6.750 33.360 6.820 ;
        RECT 36.100 6.750 36.260 6.820 ;
        RECT 39.000 6.750 39.160 6.820 ;
        RECT 41.900 6.750 42.060 6.820 ;
        RECT 44.800 6.750 44.960 6.820 ;
        RECT 47.700 6.750 47.860 6.820 ;
        RECT 50.600 6.750 50.760 6.820 ;
        RECT 53.500 6.750 53.660 6.820 ;
        RECT 56.400 6.750 56.560 6.820 ;
        RECT 59.300 6.750 59.460 6.820 ;
        RECT 62.200 6.750 62.360 6.820 ;
        RECT 65.100 6.750 65.260 6.820 ;
        RECT 68.000 6.750 68.160 6.820 ;
        RECT 70.900 6.750 71.060 6.820 ;
        RECT 73.800 6.750 73.960 6.820 ;
        RECT 76.700 6.750 76.860 6.820 ;
        RECT 79.600 6.750 79.760 6.820 ;
        RECT 82.500 6.750 82.660 6.820 ;
        RECT 85.400 6.750 85.560 6.820 ;
        RECT 88.300 6.750 88.460 6.820 ;
        RECT 91.200 6.750 91.360 6.820 ;
        RECT 1.310 5.470 1.450 5.480 ;
        RECT 4.210 5.470 4.350 5.480 ;
        RECT 7.110 5.470 7.250 5.480 ;
        RECT 10.010 5.470 10.150 5.480 ;
        RECT 12.910 5.470 13.050 5.480 ;
        RECT 15.810 5.470 15.950 5.480 ;
        RECT 18.710 5.470 18.850 5.480 ;
        RECT 21.610 5.470 21.750 5.480 ;
        RECT 24.510 5.470 24.650 5.480 ;
        RECT 27.410 5.470 27.550 5.480 ;
        RECT 30.310 5.470 30.450 5.480 ;
        RECT 33.210 5.470 33.350 5.480 ;
        RECT 36.110 5.470 36.250 5.480 ;
        RECT 39.010 5.470 39.150 5.480 ;
        RECT 41.910 5.470 42.050 5.480 ;
        RECT 44.810 5.470 44.950 5.480 ;
        RECT 47.710 5.470 47.850 5.480 ;
        RECT 50.610 5.470 50.750 5.480 ;
        RECT 53.510 5.470 53.650 5.480 ;
        RECT 56.410 5.470 56.550 5.480 ;
        RECT 59.310 5.470 59.450 5.480 ;
        RECT 62.210 5.470 62.350 5.480 ;
        RECT 65.110 5.470 65.250 5.480 ;
        RECT 68.010 5.470 68.150 5.480 ;
        RECT 70.910 5.470 71.050 5.480 ;
        RECT 73.810 5.470 73.950 5.480 ;
        RECT 76.710 5.470 76.850 5.480 ;
        RECT 79.610 5.470 79.750 5.480 ;
        RECT 82.510 5.470 82.650 5.480 ;
        RECT 85.410 5.470 85.550 5.480 ;
        RECT 88.310 5.470 88.450 5.480 ;
        RECT 91.210 5.470 91.350 5.480 ;
        RECT 1.300 5.400 1.460 5.470 ;
        RECT 4.200 5.400 4.360 5.470 ;
        RECT 7.100 5.400 7.260 5.470 ;
        RECT 10.000 5.400 10.160 5.470 ;
        RECT 12.900 5.400 13.060 5.470 ;
        RECT 15.800 5.400 15.960 5.470 ;
        RECT 18.700 5.400 18.860 5.470 ;
        RECT 21.600 5.400 21.760 5.470 ;
        RECT 24.500 5.400 24.660 5.470 ;
        RECT 27.400 5.400 27.560 5.470 ;
        RECT 30.300 5.400 30.460 5.470 ;
        RECT 33.200 5.400 33.360 5.470 ;
        RECT 36.100 5.400 36.260 5.470 ;
        RECT 39.000 5.400 39.160 5.470 ;
        RECT 41.900 5.400 42.060 5.470 ;
        RECT 44.800 5.400 44.960 5.470 ;
        RECT 47.700 5.400 47.860 5.470 ;
        RECT 50.600 5.400 50.760 5.470 ;
        RECT 53.500 5.400 53.660 5.470 ;
        RECT 56.400 5.400 56.560 5.470 ;
        RECT 59.300 5.400 59.460 5.470 ;
        RECT 62.200 5.400 62.360 5.470 ;
        RECT 65.100 5.400 65.260 5.470 ;
        RECT 68.000 5.400 68.160 5.470 ;
        RECT 70.900 5.400 71.060 5.470 ;
        RECT 73.800 5.400 73.960 5.470 ;
        RECT 76.700 5.400 76.860 5.470 ;
        RECT 79.600 5.400 79.760 5.470 ;
        RECT 82.500 5.400 82.660 5.470 ;
        RECT 85.400 5.400 85.560 5.470 ;
        RECT 88.300 5.400 88.460 5.470 ;
        RECT 91.200 5.400 91.360 5.470 ;
        RECT 1.310 4.120 1.450 4.130 ;
        RECT 4.210 4.120 4.350 4.130 ;
        RECT 7.110 4.120 7.250 4.130 ;
        RECT 10.010 4.120 10.150 4.130 ;
        RECT 12.910 4.120 13.050 4.130 ;
        RECT 15.810 4.120 15.950 4.130 ;
        RECT 18.710 4.120 18.850 4.130 ;
        RECT 21.610 4.120 21.750 4.130 ;
        RECT 24.510 4.120 24.650 4.130 ;
        RECT 27.410 4.120 27.550 4.130 ;
        RECT 30.310 4.120 30.450 4.130 ;
        RECT 33.210 4.120 33.350 4.130 ;
        RECT 36.110 4.120 36.250 4.130 ;
        RECT 39.010 4.120 39.150 4.130 ;
        RECT 41.910 4.120 42.050 4.130 ;
        RECT 44.810 4.120 44.950 4.130 ;
        RECT 47.710 4.120 47.850 4.130 ;
        RECT 50.610 4.120 50.750 4.130 ;
        RECT 53.510 4.120 53.650 4.130 ;
        RECT 56.410 4.120 56.550 4.130 ;
        RECT 59.310 4.120 59.450 4.130 ;
        RECT 62.210 4.120 62.350 4.130 ;
        RECT 65.110 4.120 65.250 4.130 ;
        RECT 68.010 4.120 68.150 4.130 ;
        RECT 70.910 4.120 71.050 4.130 ;
        RECT 73.810 4.120 73.950 4.130 ;
        RECT 76.710 4.120 76.850 4.130 ;
        RECT 79.610 4.120 79.750 4.130 ;
        RECT 82.510 4.120 82.650 4.130 ;
        RECT 85.410 4.120 85.550 4.130 ;
        RECT 88.310 4.120 88.450 4.130 ;
        RECT 91.210 4.120 91.350 4.130 ;
        RECT 1.300 4.050 1.460 4.120 ;
        RECT 4.200 4.050 4.360 4.120 ;
        RECT 7.100 4.050 7.260 4.120 ;
        RECT 10.000 4.050 10.160 4.120 ;
        RECT 12.900 4.050 13.060 4.120 ;
        RECT 15.800 4.050 15.960 4.120 ;
        RECT 18.700 4.050 18.860 4.120 ;
        RECT 21.600 4.050 21.760 4.120 ;
        RECT 24.500 4.050 24.660 4.120 ;
        RECT 27.400 4.050 27.560 4.120 ;
        RECT 30.300 4.050 30.460 4.120 ;
        RECT 33.200 4.050 33.360 4.120 ;
        RECT 36.100 4.050 36.260 4.120 ;
        RECT 39.000 4.050 39.160 4.120 ;
        RECT 41.900 4.050 42.060 4.120 ;
        RECT 44.800 4.050 44.960 4.120 ;
        RECT 47.700 4.050 47.860 4.120 ;
        RECT 50.600 4.050 50.760 4.120 ;
        RECT 53.500 4.050 53.660 4.120 ;
        RECT 56.400 4.050 56.560 4.120 ;
        RECT 59.300 4.050 59.460 4.120 ;
        RECT 62.200 4.050 62.360 4.120 ;
        RECT 65.100 4.050 65.260 4.120 ;
        RECT 68.000 4.050 68.160 4.120 ;
        RECT 70.900 4.050 71.060 4.120 ;
        RECT 73.800 4.050 73.960 4.120 ;
        RECT 76.700 4.050 76.860 4.120 ;
        RECT 79.600 4.050 79.760 4.120 ;
        RECT 82.500 4.050 82.660 4.120 ;
        RECT 85.400 4.050 85.560 4.120 ;
        RECT 88.300 4.050 88.460 4.120 ;
        RECT 91.200 4.050 91.360 4.120 ;
        RECT 1.310 2.770 1.450 2.780 ;
        RECT 4.210 2.770 4.350 2.780 ;
        RECT 7.110 2.770 7.250 2.780 ;
        RECT 10.010 2.770 10.150 2.780 ;
        RECT 12.910 2.770 13.050 2.780 ;
        RECT 15.810 2.770 15.950 2.780 ;
        RECT 18.710 2.770 18.850 2.780 ;
        RECT 21.610 2.770 21.750 2.780 ;
        RECT 24.510 2.770 24.650 2.780 ;
        RECT 27.410 2.770 27.550 2.780 ;
        RECT 30.310 2.770 30.450 2.780 ;
        RECT 33.210 2.770 33.350 2.780 ;
        RECT 36.110 2.770 36.250 2.780 ;
        RECT 39.010 2.770 39.150 2.780 ;
        RECT 41.910 2.770 42.050 2.780 ;
        RECT 44.810 2.770 44.950 2.780 ;
        RECT 47.710 2.770 47.850 2.780 ;
        RECT 50.610 2.770 50.750 2.780 ;
        RECT 53.510 2.770 53.650 2.780 ;
        RECT 56.410 2.770 56.550 2.780 ;
        RECT 59.310 2.770 59.450 2.780 ;
        RECT 62.210 2.770 62.350 2.780 ;
        RECT 65.110 2.770 65.250 2.780 ;
        RECT 68.010 2.770 68.150 2.780 ;
        RECT 70.910 2.770 71.050 2.780 ;
        RECT 73.810 2.770 73.950 2.780 ;
        RECT 76.710 2.770 76.850 2.780 ;
        RECT 79.610 2.770 79.750 2.780 ;
        RECT 82.510 2.770 82.650 2.780 ;
        RECT 85.410 2.770 85.550 2.780 ;
        RECT 88.310 2.770 88.450 2.780 ;
        RECT 91.210 2.770 91.350 2.780 ;
        RECT 1.300 2.700 1.460 2.770 ;
        RECT 4.200 2.700 4.360 2.770 ;
        RECT 7.100 2.700 7.260 2.770 ;
        RECT 10.000 2.700 10.160 2.770 ;
        RECT 12.900 2.700 13.060 2.770 ;
        RECT 15.800 2.700 15.960 2.770 ;
        RECT 18.700 2.700 18.860 2.770 ;
        RECT 21.600 2.700 21.760 2.770 ;
        RECT 24.500 2.700 24.660 2.770 ;
        RECT 27.400 2.700 27.560 2.770 ;
        RECT 30.300 2.700 30.460 2.770 ;
        RECT 33.200 2.700 33.360 2.770 ;
        RECT 36.100 2.700 36.260 2.770 ;
        RECT 39.000 2.700 39.160 2.770 ;
        RECT 41.900 2.700 42.060 2.770 ;
        RECT 44.800 2.700 44.960 2.770 ;
        RECT 47.700 2.700 47.860 2.770 ;
        RECT 50.600 2.700 50.760 2.770 ;
        RECT 53.500 2.700 53.660 2.770 ;
        RECT 56.400 2.700 56.560 2.770 ;
        RECT 59.300 2.700 59.460 2.770 ;
        RECT 62.200 2.700 62.360 2.770 ;
        RECT 65.100 2.700 65.260 2.770 ;
        RECT 68.000 2.700 68.160 2.770 ;
        RECT 70.900 2.700 71.060 2.770 ;
        RECT 73.800 2.700 73.960 2.770 ;
        RECT 76.700 2.700 76.860 2.770 ;
        RECT 79.600 2.700 79.760 2.770 ;
        RECT 82.500 2.700 82.660 2.770 ;
        RECT 85.400 2.700 85.560 2.770 ;
        RECT 88.300 2.700 88.460 2.770 ;
        RECT 91.200 2.700 91.360 2.770 ;
        RECT 1.310 1.420 1.450 1.430 ;
        RECT 4.210 1.420 4.350 1.430 ;
        RECT 7.110 1.420 7.250 1.430 ;
        RECT 10.010 1.420 10.150 1.430 ;
        RECT 12.910 1.420 13.050 1.430 ;
        RECT 15.810 1.420 15.950 1.430 ;
        RECT 18.710 1.420 18.850 1.430 ;
        RECT 21.610 1.420 21.750 1.430 ;
        RECT 24.510 1.425 24.650 1.435 ;
        RECT 27.410 1.425 27.550 1.435 ;
        RECT 30.310 1.425 30.450 1.435 ;
        RECT 33.210 1.425 33.350 1.435 ;
        RECT 36.110 1.425 36.250 1.435 ;
        RECT 39.010 1.425 39.150 1.435 ;
        RECT 41.910 1.425 42.050 1.435 ;
        RECT 44.810 1.425 44.950 1.435 ;
        RECT 47.710 1.425 47.850 1.435 ;
        RECT 50.610 1.425 50.750 1.435 ;
        RECT 53.510 1.425 53.650 1.435 ;
        RECT 56.410 1.425 56.550 1.435 ;
        RECT 59.310 1.425 59.450 1.435 ;
        RECT 62.210 1.425 62.350 1.435 ;
        RECT 65.110 1.425 65.250 1.435 ;
        RECT 68.010 1.425 68.150 1.435 ;
        RECT 70.910 1.425 71.050 1.435 ;
        RECT 73.810 1.425 73.950 1.435 ;
        RECT 76.710 1.425 76.850 1.435 ;
        RECT 79.610 1.425 79.750 1.435 ;
        RECT 82.510 1.425 82.650 1.435 ;
        RECT 85.410 1.425 85.550 1.435 ;
        RECT 88.310 1.425 88.450 1.435 ;
        RECT 91.210 1.425 91.350 1.435 ;
        RECT 1.300 1.350 1.460 1.420 ;
        RECT 4.200 1.350 4.360 1.420 ;
        RECT 7.100 1.350 7.260 1.420 ;
        RECT 10.000 1.350 10.160 1.420 ;
        RECT 12.900 1.350 13.060 1.420 ;
        RECT 15.800 1.350 15.960 1.420 ;
        RECT 18.700 1.350 18.860 1.420 ;
        RECT 21.600 1.350 21.760 1.420 ;
        RECT 24.500 1.355 24.660 1.425 ;
        RECT 27.400 1.355 27.560 1.425 ;
        RECT 30.300 1.355 30.460 1.425 ;
        RECT 33.200 1.355 33.360 1.425 ;
        RECT 36.100 1.355 36.260 1.425 ;
        RECT 39.000 1.355 39.160 1.425 ;
        RECT 41.900 1.355 42.060 1.425 ;
        RECT 44.800 1.355 44.960 1.425 ;
        RECT 47.700 1.355 47.860 1.425 ;
        RECT 50.600 1.355 50.760 1.425 ;
        RECT 53.500 1.355 53.660 1.425 ;
        RECT 56.400 1.355 56.560 1.425 ;
        RECT 59.300 1.355 59.460 1.425 ;
        RECT 62.200 1.355 62.360 1.425 ;
        RECT 65.100 1.355 65.260 1.425 ;
        RECT 68.000 1.355 68.160 1.425 ;
        RECT 70.900 1.355 71.060 1.425 ;
        RECT 73.800 1.355 73.960 1.425 ;
        RECT 76.700 1.355 76.860 1.425 ;
        RECT 79.600 1.355 79.760 1.425 ;
        RECT 82.500 1.355 82.660 1.425 ;
        RECT 85.400 1.355 85.560 1.425 ;
        RECT 88.300 1.355 88.460 1.425 ;
        RECT 91.200 1.355 91.360 1.425 ;
        RECT 1.310 0.070 1.450 0.080 ;
        RECT 4.210 0.070 4.350 0.080 ;
        RECT 7.110 0.070 7.250 0.080 ;
        RECT 10.010 0.070 10.150 0.080 ;
        RECT 12.910 0.070 13.050 0.080 ;
        RECT 15.810 0.070 15.950 0.080 ;
        RECT 18.710 0.070 18.850 0.080 ;
        RECT 21.610 0.070 21.750 0.080 ;
        RECT 24.510 0.075 24.650 0.085 ;
        RECT 27.410 0.075 27.550 0.085 ;
        RECT 30.310 0.075 30.450 0.085 ;
        RECT 33.210 0.075 33.350 0.085 ;
        RECT 36.110 0.075 36.250 0.085 ;
        RECT 39.010 0.075 39.150 0.085 ;
        RECT 41.910 0.075 42.050 0.085 ;
        RECT 44.810 0.075 44.950 0.085 ;
        RECT 47.710 0.075 47.850 0.085 ;
        RECT 50.610 0.075 50.750 0.085 ;
        RECT 53.510 0.075 53.650 0.085 ;
        RECT 56.410 0.075 56.550 0.085 ;
        RECT 59.310 0.075 59.450 0.085 ;
        RECT 62.210 0.075 62.350 0.085 ;
        RECT 65.110 0.075 65.250 0.085 ;
        RECT 68.010 0.075 68.150 0.085 ;
        RECT 70.910 0.075 71.050 0.085 ;
        RECT 73.810 0.075 73.950 0.085 ;
        RECT 76.710 0.075 76.850 0.085 ;
        RECT 79.610 0.075 79.750 0.085 ;
        RECT 82.510 0.075 82.650 0.085 ;
        RECT 85.410 0.075 85.550 0.085 ;
        RECT 88.310 0.075 88.450 0.085 ;
        RECT 91.210 0.075 91.350 0.085 ;
        RECT 1.300 0.000 1.460 0.070 ;
        RECT 4.200 0.000 4.360 0.070 ;
        RECT 7.100 0.000 7.260 0.070 ;
        RECT 10.000 0.000 10.160 0.070 ;
        RECT 12.900 0.000 13.060 0.070 ;
        RECT 15.800 0.000 15.960 0.070 ;
        RECT 18.700 0.000 18.860 0.070 ;
        RECT 21.600 0.000 21.760 0.070 ;
        RECT 24.500 0.005 24.660 0.075 ;
        RECT 27.400 0.005 27.560 0.075 ;
        RECT 30.300 0.005 30.460 0.075 ;
        RECT 33.200 0.005 33.360 0.075 ;
        RECT 36.100 0.005 36.260 0.075 ;
        RECT 39.000 0.005 39.160 0.075 ;
        RECT 41.900 0.005 42.060 0.075 ;
        RECT 44.800 0.005 44.960 0.075 ;
        RECT 47.700 0.005 47.860 0.075 ;
        RECT 50.600 0.005 50.760 0.075 ;
        RECT 53.500 0.005 53.660 0.075 ;
        RECT 56.400 0.005 56.560 0.075 ;
        RECT 59.300 0.005 59.460 0.075 ;
        RECT 62.200 0.005 62.360 0.075 ;
        RECT 65.100 0.005 65.260 0.075 ;
        RECT 68.000 0.005 68.160 0.075 ;
        RECT 70.900 0.005 71.060 0.075 ;
        RECT 73.800 0.005 73.960 0.075 ;
        RECT 76.700 0.005 76.860 0.075 ;
        RECT 79.600 0.005 79.760 0.075 ;
        RECT 82.500 0.005 82.660 0.075 ;
        RECT 85.400 0.005 85.560 0.075 ;
        RECT 88.300 0.005 88.460 0.075 ;
        RECT 91.200 0.005 91.360 0.075 ;
      LAYER met1 ;
        RECT 0.000 41.850 92.660 41.920 ;
        RECT 0.000 40.500 92.660 40.570 ;
        RECT 0.000 39.150 92.660 39.220 ;
        RECT 0.000 37.800 92.660 37.870 ;
        RECT 0.000 36.450 92.660 36.520 ;
        RECT 0.000 35.100 92.660 35.170 ;
        RECT 0.000 33.750 92.660 33.820 ;
        RECT 0.000 32.400 92.660 32.470 ;
        RECT 0.000 31.050 92.660 31.120 ;
        RECT 0.000 29.700 92.660 29.770 ;
        RECT 0.000 28.350 92.660 28.420 ;
        RECT 0.000 27.000 92.660 27.070 ;
        RECT 0.000 25.650 92.660 25.720 ;
        RECT 0.000 24.300 92.660 24.370 ;
        RECT 0.000 22.950 92.660 23.020 ;
        RECT 0.000 21.600 92.660 21.670 ;
        RECT 0.000 20.250 92.660 20.320 ;
        RECT 0.000 18.900 92.660 18.970 ;
        RECT 0.000 17.550 92.660 17.620 ;
        RECT 0.000 16.200 92.660 16.270 ;
        RECT 0.000 14.850 92.660 14.920 ;
        RECT 0.000 13.500 92.660 13.570 ;
        RECT 0.000 12.150 92.660 12.220 ;
        RECT 0.000 10.800 92.660 10.870 ;
        RECT 0.000 9.450 92.660 9.520 ;
        RECT 0.000 8.100 92.660 8.170 ;
        RECT 0.000 6.750 92.660 6.820 ;
        RECT 0.000 5.400 92.660 5.470 ;
        RECT 0.000 4.050 92.660 4.120 ;
        RECT 46.055 2.770 46.650 2.775 ;
        RECT 0.000 2.705 92.660 2.770 ;
        RECT 0.000 2.700 46.260 2.705 ;
        RECT 46.400 2.700 92.660 2.705 ;
        RECT 23.155 1.420 69.460 1.425 ;
        RECT 69.600 1.420 92.660 1.425 ;
        RECT 0.000 1.355 92.660 1.420 ;
        RECT 0.000 1.350 23.155 1.355 ;
        RECT 23.155 0.070 92.660 0.075 ;
        RECT 0.000 0.005 92.660 0.070 ;
        RECT 0.000 0.000 23.155 0.005 ;
    END
  END GND
  OBS
      LAYER li1 ;
        RECT 0.775 42.770 0.850 42.910 ;
        RECT 0.990 42.720 1.065 42.860 ;
        RECT 1.695 42.780 1.755 42.860 ;
        POLYGON 1.695 42.780 1.755 42.780 1.755 42.720 ;
        RECT 1.910 42.770 1.985 42.910 ;
        RECT 3.675 42.770 3.750 42.910 ;
        RECT 3.890 42.720 3.965 42.860 ;
        RECT 4.595 42.780 4.655 42.860 ;
        POLYGON 4.595 42.780 4.655 42.780 4.655 42.720 ;
        RECT 4.810 42.770 4.885 42.910 ;
        RECT 6.575 42.770 6.650 42.910 ;
        RECT 6.790 42.720 6.865 42.860 ;
        RECT 7.495 42.780 7.555 42.860 ;
        POLYGON 7.495 42.780 7.555 42.780 7.555 42.720 ;
        RECT 7.710 42.770 7.785 42.910 ;
        RECT 9.475 42.770 9.550 42.910 ;
        RECT 9.690 42.720 9.765 42.860 ;
        RECT 10.395 42.780 10.455 42.860 ;
        POLYGON 10.395 42.780 10.455 42.780 10.455 42.720 ;
        RECT 10.610 42.770 10.685 42.910 ;
        RECT 12.375 42.770 12.450 42.910 ;
        RECT 12.590 42.720 12.665 42.860 ;
        RECT 13.295 42.780 13.355 42.860 ;
        POLYGON 13.295 42.780 13.355 42.780 13.355 42.720 ;
        RECT 13.510 42.770 13.585 42.910 ;
        RECT 15.275 42.770 15.350 42.910 ;
        RECT 15.490 42.720 15.565 42.860 ;
        RECT 16.195 42.780 16.255 42.860 ;
        POLYGON 16.195 42.780 16.255 42.780 16.255 42.720 ;
        RECT 16.410 42.770 16.485 42.910 ;
        RECT 18.175 42.770 18.250 42.910 ;
        RECT 18.390 42.720 18.465 42.860 ;
        RECT 19.095 42.780 19.155 42.860 ;
        POLYGON 19.095 42.780 19.155 42.780 19.155 42.720 ;
        RECT 19.310 42.770 19.385 42.910 ;
        RECT 21.075 42.770 21.150 42.910 ;
        RECT 21.290 42.720 21.365 42.860 ;
        RECT 21.995 42.780 22.055 42.860 ;
        POLYGON 21.995 42.780 22.055 42.780 22.055 42.720 ;
        RECT 22.210 42.770 22.285 42.910 ;
        RECT 23.975 42.770 24.050 42.910 ;
        RECT 24.190 42.720 24.265 42.860 ;
        RECT 24.895 42.780 24.955 42.860 ;
        POLYGON 24.895 42.780 24.955 42.780 24.955 42.720 ;
        RECT 25.110 42.770 25.185 42.910 ;
        RECT 26.875 42.770 26.950 42.910 ;
        RECT 27.090 42.720 27.165 42.860 ;
        RECT 27.795 42.780 27.855 42.860 ;
        POLYGON 27.795 42.780 27.855 42.780 27.855 42.720 ;
        RECT 28.010 42.770 28.085 42.910 ;
        RECT 29.775 42.770 29.850 42.910 ;
        RECT 29.990 42.720 30.065 42.860 ;
        RECT 30.695 42.780 30.755 42.860 ;
        POLYGON 30.695 42.780 30.755 42.780 30.755 42.720 ;
        RECT 30.910 42.770 30.985 42.910 ;
        RECT 32.675 42.770 32.750 42.910 ;
        RECT 32.890 42.720 32.965 42.860 ;
        RECT 33.595 42.780 33.655 42.860 ;
        POLYGON 33.595 42.780 33.655 42.780 33.655 42.720 ;
        RECT 33.810 42.770 33.885 42.910 ;
        RECT 35.575 42.770 35.650 42.910 ;
        RECT 35.790 42.720 35.865 42.860 ;
        RECT 36.495 42.780 36.555 42.860 ;
        POLYGON 36.495 42.780 36.555 42.780 36.555 42.720 ;
        RECT 36.710 42.770 36.785 42.910 ;
        RECT 38.475 42.770 38.550 42.910 ;
        RECT 38.690 42.720 38.765 42.860 ;
        RECT 39.395 42.780 39.455 42.860 ;
        POLYGON 39.395 42.780 39.455 42.780 39.455 42.720 ;
        RECT 39.610 42.770 39.685 42.910 ;
        RECT 41.375 42.770 41.450 42.910 ;
        RECT 41.590 42.720 41.665 42.860 ;
        RECT 42.295 42.780 42.355 42.860 ;
        POLYGON 42.295 42.780 42.355 42.780 42.355 42.720 ;
        RECT 42.510 42.770 42.585 42.910 ;
        RECT 44.275 42.770 44.350 42.910 ;
        RECT 44.490 42.720 44.565 42.860 ;
        RECT 45.195 42.780 45.255 42.860 ;
        POLYGON 45.195 42.780 45.255 42.780 45.255 42.720 ;
        RECT 45.410 42.770 45.485 42.910 ;
        RECT 47.175 42.770 47.250 42.910 ;
        RECT 47.390 42.720 47.465 42.860 ;
        RECT 48.095 42.780 48.155 42.860 ;
        POLYGON 48.095 42.780 48.155 42.780 48.155 42.720 ;
        RECT 48.310 42.770 48.385 42.910 ;
        RECT 50.075 42.770 50.150 42.910 ;
        RECT 50.290 42.720 50.365 42.860 ;
        RECT 50.995 42.780 51.055 42.860 ;
        POLYGON 50.995 42.780 51.055 42.780 51.055 42.720 ;
        RECT 51.210 42.770 51.285 42.910 ;
        RECT 52.975 42.770 53.050 42.910 ;
        RECT 53.190 42.720 53.265 42.860 ;
        RECT 53.895 42.780 53.955 42.860 ;
        POLYGON 53.895 42.780 53.955 42.780 53.955 42.720 ;
        RECT 54.110 42.770 54.185 42.910 ;
        RECT 55.875 42.770 55.950 42.910 ;
        RECT 56.090 42.720 56.165 42.860 ;
        RECT 56.795 42.780 56.855 42.860 ;
        POLYGON 56.795 42.780 56.855 42.780 56.855 42.720 ;
        RECT 57.010 42.770 57.085 42.910 ;
        RECT 58.775 42.770 58.850 42.910 ;
        RECT 58.990 42.720 59.065 42.860 ;
        RECT 59.695 42.780 59.755 42.860 ;
        POLYGON 59.695 42.780 59.755 42.780 59.755 42.720 ;
        RECT 59.910 42.770 59.985 42.910 ;
        RECT 61.675 42.770 61.750 42.910 ;
        RECT 61.890 42.720 61.965 42.860 ;
        RECT 62.595 42.780 62.655 42.860 ;
        POLYGON 62.595 42.780 62.655 42.780 62.655 42.720 ;
        RECT 62.810 42.770 62.885 42.910 ;
        RECT 64.575 42.770 64.650 42.910 ;
        RECT 64.790 42.720 64.865 42.860 ;
        RECT 65.495 42.780 65.555 42.860 ;
        POLYGON 65.495 42.780 65.555 42.780 65.555 42.720 ;
        RECT 65.710 42.770 65.785 42.910 ;
        RECT 67.475 42.770 67.550 42.910 ;
        RECT 67.690 42.720 67.765 42.860 ;
        RECT 68.395 42.780 68.455 42.860 ;
        POLYGON 68.395 42.780 68.455 42.780 68.455 42.720 ;
        RECT 68.610 42.770 68.685 42.910 ;
        RECT 70.375 42.770 70.450 42.910 ;
        RECT 70.590 42.720 70.665 42.860 ;
        RECT 71.295 42.780 71.355 42.860 ;
        POLYGON 71.295 42.780 71.355 42.780 71.355 42.720 ;
        RECT 71.510 42.770 71.585 42.910 ;
        RECT 73.275 42.770 73.350 42.910 ;
        RECT 73.490 42.720 73.565 42.860 ;
        RECT 74.195 42.780 74.255 42.860 ;
        POLYGON 74.195 42.780 74.255 42.780 74.255 42.720 ;
        RECT 74.410 42.770 74.485 42.910 ;
        RECT 76.175 42.770 76.250 42.910 ;
        RECT 76.390 42.720 76.465 42.860 ;
        RECT 77.095 42.780 77.155 42.860 ;
        POLYGON 77.095 42.780 77.155 42.780 77.155 42.720 ;
        RECT 77.310 42.770 77.385 42.910 ;
        RECT 79.075 42.770 79.150 42.910 ;
        RECT 79.290 42.720 79.365 42.860 ;
        RECT 79.995 42.780 80.055 42.860 ;
        POLYGON 79.995 42.780 80.055 42.780 80.055 42.720 ;
        RECT 80.210 42.770 80.285 42.910 ;
        RECT 81.975 42.770 82.050 42.910 ;
        RECT 82.190 42.720 82.265 42.860 ;
        RECT 82.895 42.780 82.955 42.860 ;
        POLYGON 82.895 42.780 82.955 42.780 82.955 42.720 ;
        RECT 83.110 42.770 83.185 42.910 ;
        RECT 84.875 42.770 84.950 42.910 ;
        RECT 85.090 42.720 85.165 42.860 ;
        RECT 85.795 42.780 85.855 42.860 ;
        POLYGON 85.795 42.780 85.855 42.780 85.855 42.720 ;
        RECT 86.010 42.770 86.085 42.910 ;
        RECT 87.775 42.770 87.850 42.910 ;
        RECT 87.990 42.720 88.065 42.860 ;
        RECT 88.695 42.780 88.755 42.860 ;
        POLYGON 88.695 42.780 88.755 42.780 88.755 42.720 ;
        RECT 88.910 42.770 88.985 42.910 ;
        RECT 90.675 42.770 90.750 42.910 ;
        RECT 90.890 42.720 90.965 42.860 ;
        RECT 91.595 42.780 91.655 42.860 ;
        POLYGON 91.595 42.780 91.655 42.780 91.655 42.720 ;
        RECT 91.810 42.770 91.885 42.910 ;
        RECT 0.720 42.250 0.870 42.420 ;
        RECT 1.110 42.385 1.260 42.555 ;
        RECT 1.500 42.385 1.650 42.555 ;
        RECT 1.890 42.250 2.040 42.420 ;
        RECT 3.620 42.250 3.770 42.420 ;
        RECT 4.010 42.385 4.160 42.555 ;
        RECT 4.400 42.385 4.550 42.555 ;
        RECT 4.790 42.250 4.940 42.420 ;
        RECT 6.520 42.250 6.670 42.420 ;
        RECT 6.910 42.385 7.060 42.555 ;
        RECT 7.300 42.385 7.450 42.555 ;
        RECT 7.690 42.250 7.840 42.420 ;
        RECT 9.420 42.250 9.570 42.420 ;
        RECT 9.810 42.385 9.960 42.555 ;
        RECT 10.200 42.385 10.350 42.555 ;
        RECT 10.590 42.250 10.740 42.420 ;
        RECT 12.320 42.250 12.470 42.420 ;
        RECT 12.710 42.385 12.860 42.555 ;
        RECT 13.100 42.385 13.250 42.555 ;
        RECT 13.490 42.250 13.640 42.420 ;
        RECT 15.220 42.250 15.370 42.420 ;
        RECT 15.610 42.385 15.760 42.555 ;
        RECT 16.000 42.385 16.150 42.555 ;
        RECT 16.390 42.250 16.540 42.420 ;
        RECT 18.120 42.250 18.270 42.420 ;
        RECT 18.510 42.385 18.660 42.555 ;
        RECT 18.900 42.385 19.050 42.555 ;
        RECT 19.290 42.250 19.440 42.420 ;
        RECT 21.020 42.250 21.170 42.420 ;
        RECT 21.410 42.385 21.560 42.555 ;
        RECT 21.800 42.385 21.950 42.555 ;
        RECT 22.190 42.250 22.340 42.420 ;
        RECT 23.920 42.250 24.070 42.420 ;
        RECT 24.310 42.385 24.460 42.555 ;
        RECT 24.700 42.385 24.850 42.555 ;
        RECT 25.090 42.250 25.240 42.420 ;
        RECT 26.820 42.250 26.970 42.420 ;
        RECT 27.210 42.385 27.360 42.555 ;
        RECT 27.600 42.385 27.750 42.555 ;
        RECT 27.990 42.250 28.140 42.420 ;
        RECT 29.720 42.250 29.870 42.420 ;
        RECT 30.110 42.385 30.260 42.555 ;
        RECT 30.500 42.385 30.650 42.555 ;
        RECT 30.890 42.250 31.040 42.420 ;
        RECT 32.620 42.250 32.770 42.420 ;
        RECT 33.010 42.385 33.160 42.555 ;
        RECT 33.400 42.385 33.550 42.555 ;
        RECT 33.790 42.250 33.940 42.420 ;
        RECT 35.520 42.250 35.670 42.420 ;
        RECT 35.910 42.385 36.060 42.555 ;
        RECT 36.300 42.385 36.450 42.555 ;
        RECT 36.690 42.250 36.840 42.420 ;
        RECT 38.420 42.250 38.570 42.420 ;
        RECT 38.810 42.385 38.960 42.555 ;
        RECT 39.200 42.385 39.350 42.555 ;
        RECT 39.590 42.250 39.740 42.420 ;
        RECT 41.320 42.250 41.470 42.420 ;
        RECT 41.710 42.385 41.860 42.555 ;
        RECT 42.100 42.385 42.250 42.555 ;
        RECT 42.490 42.250 42.640 42.420 ;
        RECT 44.220 42.250 44.370 42.420 ;
        RECT 44.610 42.385 44.760 42.555 ;
        RECT 45.000 42.385 45.150 42.555 ;
        RECT 45.390 42.250 45.540 42.420 ;
        RECT 47.120 42.250 47.270 42.420 ;
        RECT 47.510 42.385 47.660 42.555 ;
        RECT 47.900 42.385 48.050 42.555 ;
        RECT 48.290 42.250 48.440 42.420 ;
        RECT 50.020 42.250 50.170 42.420 ;
        RECT 50.410 42.385 50.560 42.555 ;
        RECT 50.800 42.385 50.950 42.555 ;
        RECT 51.190 42.250 51.340 42.420 ;
        RECT 52.920 42.250 53.070 42.420 ;
        RECT 53.310 42.385 53.460 42.555 ;
        RECT 53.700 42.385 53.850 42.555 ;
        RECT 54.090 42.250 54.240 42.420 ;
        RECT 55.820 42.250 55.970 42.420 ;
        RECT 56.210 42.385 56.360 42.555 ;
        RECT 56.600 42.385 56.750 42.555 ;
        RECT 56.990 42.250 57.140 42.420 ;
        RECT 58.720 42.250 58.870 42.420 ;
        RECT 59.110 42.385 59.260 42.555 ;
        RECT 59.500 42.385 59.650 42.555 ;
        RECT 59.890 42.250 60.040 42.420 ;
        RECT 61.620 42.250 61.770 42.420 ;
        RECT 62.010 42.385 62.160 42.555 ;
        RECT 62.400 42.385 62.550 42.555 ;
        RECT 62.790 42.250 62.940 42.420 ;
        RECT 64.520 42.250 64.670 42.420 ;
        RECT 64.910 42.385 65.060 42.555 ;
        RECT 65.300 42.385 65.450 42.555 ;
        RECT 65.690 42.250 65.840 42.420 ;
        RECT 67.420 42.250 67.570 42.420 ;
        RECT 67.810 42.385 67.960 42.555 ;
        RECT 68.200 42.385 68.350 42.555 ;
        RECT 68.590 42.250 68.740 42.420 ;
        RECT 70.320 42.250 70.470 42.420 ;
        RECT 70.710 42.385 70.860 42.555 ;
        RECT 71.100 42.385 71.250 42.555 ;
        RECT 71.490 42.250 71.640 42.420 ;
        RECT 73.220 42.250 73.370 42.420 ;
        RECT 73.610 42.385 73.760 42.555 ;
        RECT 74.000 42.385 74.150 42.555 ;
        RECT 74.390 42.250 74.540 42.420 ;
        RECT 76.120 42.250 76.270 42.420 ;
        RECT 76.510 42.385 76.660 42.555 ;
        RECT 76.900 42.385 77.050 42.555 ;
        RECT 77.290 42.250 77.440 42.420 ;
        RECT 79.020 42.250 79.170 42.420 ;
        RECT 79.410 42.385 79.560 42.555 ;
        RECT 79.800 42.385 79.950 42.555 ;
        RECT 80.190 42.250 80.340 42.420 ;
        RECT 81.920 42.250 82.070 42.420 ;
        RECT 82.310 42.385 82.460 42.555 ;
        RECT 82.700 42.385 82.850 42.555 ;
        RECT 83.090 42.250 83.240 42.420 ;
        RECT 84.820 42.250 84.970 42.420 ;
        RECT 85.210 42.385 85.360 42.555 ;
        RECT 85.600 42.385 85.750 42.555 ;
        RECT 85.990 42.250 86.140 42.420 ;
        RECT 87.720 42.250 87.870 42.420 ;
        RECT 88.110 42.385 88.260 42.555 ;
        RECT 88.500 42.385 88.650 42.555 ;
        RECT 88.890 42.250 89.040 42.420 ;
        RECT 90.620 42.250 90.770 42.420 ;
        RECT 91.010 42.385 91.160 42.555 ;
        RECT 91.400 42.385 91.550 42.555 ;
        RECT 91.790 42.250 91.940 42.420 ;
        RECT 0.985 42.165 1.035 42.200 ;
        POLYGON 1.035 42.200 1.070 42.165 1.035 42.165 ;
        RECT 0.985 42.040 1.070 42.165 ;
        RECT 1.690 42.040 1.775 42.200 ;
        RECT 3.885 42.165 3.935 42.200 ;
        POLYGON 3.935 42.200 3.970 42.165 3.935 42.165 ;
        RECT 3.885 42.040 3.970 42.165 ;
        RECT 4.590 42.040 4.675 42.200 ;
        RECT 6.785 42.165 6.835 42.200 ;
        POLYGON 6.835 42.200 6.870 42.165 6.835 42.165 ;
        RECT 6.785 42.040 6.870 42.165 ;
        RECT 7.490 42.040 7.575 42.200 ;
        RECT 9.685 42.165 9.735 42.200 ;
        POLYGON 9.735 42.200 9.770 42.165 9.735 42.165 ;
        RECT 9.685 42.040 9.770 42.165 ;
        RECT 10.390 42.040 10.475 42.200 ;
        RECT 12.585 42.165 12.635 42.200 ;
        POLYGON 12.635 42.200 12.670 42.165 12.635 42.165 ;
        RECT 12.585 42.040 12.670 42.165 ;
        RECT 13.290 42.040 13.375 42.200 ;
        RECT 15.485 42.165 15.535 42.200 ;
        POLYGON 15.535 42.200 15.570 42.165 15.535 42.165 ;
        RECT 15.485 42.040 15.570 42.165 ;
        RECT 16.190 42.040 16.275 42.200 ;
        RECT 18.385 42.165 18.435 42.200 ;
        POLYGON 18.435 42.200 18.470 42.165 18.435 42.165 ;
        RECT 18.385 42.040 18.470 42.165 ;
        RECT 19.090 42.040 19.175 42.200 ;
        RECT 21.285 42.165 21.335 42.200 ;
        POLYGON 21.335 42.200 21.370 42.165 21.335 42.165 ;
        RECT 21.285 42.040 21.370 42.165 ;
        RECT 21.990 42.040 22.075 42.200 ;
        RECT 24.185 42.165 24.235 42.200 ;
        POLYGON 24.235 42.200 24.270 42.165 24.235 42.165 ;
        RECT 24.185 42.040 24.270 42.165 ;
        RECT 24.890 42.040 24.975 42.200 ;
        RECT 27.085 42.165 27.135 42.200 ;
        POLYGON 27.135 42.200 27.170 42.165 27.135 42.165 ;
        RECT 27.085 42.040 27.170 42.165 ;
        RECT 27.790 42.040 27.875 42.200 ;
        RECT 29.985 42.165 30.035 42.200 ;
        POLYGON 30.035 42.200 30.070 42.165 30.035 42.165 ;
        RECT 29.985 42.040 30.070 42.165 ;
        RECT 30.690 42.040 30.775 42.200 ;
        RECT 32.885 42.165 32.935 42.200 ;
        POLYGON 32.935 42.200 32.970 42.165 32.935 42.165 ;
        RECT 32.885 42.040 32.970 42.165 ;
        RECT 33.590 42.040 33.675 42.200 ;
        RECT 35.785 42.165 35.835 42.200 ;
        POLYGON 35.835 42.200 35.870 42.165 35.835 42.165 ;
        RECT 35.785 42.040 35.870 42.165 ;
        RECT 36.490 42.040 36.575 42.200 ;
        RECT 38.685 42.165 38.735 42.200 ;
        POLYGON 38.735 42.200 38.770 42.165 38.735 42.165 ;
        RECT 38.685 42.040 38.770 42.165 ;
        RECT 39.390 42.040 39.475 42.200 ;
        RECT 41.585 42.165 41.635 42.200 ;
        POLYGON 41.635 42.200 41.670 42.165 41.635 42.165 ;
        RECT 41.585 42.040 41.670 42.165 ;
        RECT 42.290 42.040 42.375 42.200 ;
        RECT 44.485 42.165 44.535 42.200 ;
        POLYGON 44.535 42.200 44.570 42.165 44.535 42.165 ;
        RECT 44.485 42.040 44.570 42.165 ;
        RECT 45.190 42.040 45.275 42.200 ;
        RECT 47.385 42.165 47.435 42.200 ;
        POLYGON 47.435 42.200 47.470 42.165 47.435 42.165 ;
        RECT 47.385 42.040 47.470 42.165 ;
        RECT 48.090 42.040 48.175 42.200 ;
        RECT 50.285 42.165 50.335 42.200 ;
        POLYGON 50.335 42.200 50.370 42.165 50.335 42.165 ;
        RECT 50.285 42.040 50.370 42.165 ;
        RECT 50.990 42.040 51.075 42.200 ;
        RECT 53.185 42.165 53.235 42.200 ;
        POLYGON 53.235 42.200 53.270 42.165 53.235 42.165 ;
        RECT 53.185 42.040 53.270 42.165 ;
        RECT 53.890 42.040 53.975 42.200 ;
        RECT 56.085 42.165 56.135 42.200 ;
        POLYGON 56.135 42.200 56.170 42.165 56.135 42.165 ;
        RECT 56.085 42.040 56.170 42.165 ;
        RECT 56.790 42.040 56.875 42.200 ;
        RECT 58.985 42.165 59.035 42.200 ;
        POLYGON 59.035 42.200 59.070 42.165 59.035 42.165 ;
        RECT 58.985 42.040 59.070 42.165 ;
        RECT 59.690 42.040 59.775 42.200 ;
        RECT 61.885 42.165 61.935 42.200 ;
        POLYGON 61.935 42.200 61.970 42.165 61.935 42.165 ;
        RECT 61.885 42.040 61.970 42.165 ;
        RECT 62.590 42.040 62.675 42.200 ;
        RECT 64.785 42.165 64.835 42.200 ;
        POLYGON 64.835 42.200 64.870 42.165 64.835 42.165 ;
        RECT 64.785 42.040 64.870 42.165 ;
        RECT 65.490 42.040 65.575 42.200 ;
        RECT 67.685 42.165 67.735 42.200 ;
        POLYGON 67.735 42.200 67.770 42.165 67.735 42.165 ;
        RECT 67.685 42.040 67.770 42.165 ;
        RECT 68.390 42.040 68.475 42.200 ;
        RECT 70.585 42.165 70.635 42.200 ;
        POLYGON 70.635 42.200 70.670 42.165 70.635 42.165 ;
        RECT 70.585 42.040 70.670 42.165 ;
        RECT 71.290 42.040 71.375 42.200 ;
        RECT 73.485 42.165 73.535 42.200 ;
        POLYGON 73.535 42.200 73.570 42.165 73.535 42.165 ;
        RECT 73.485 42.040 73.570 42.165 ;
        RECT 74.190 42.040 74.275 42.200 ;
        RECT 76.385 42.165 76.435 42.200 ;
        POLYGON 76.435 42.200 76.470 42.165 76.435 42.165 ;
        RECT 76.385 42.040 76.470 42.165 ;
        RECT 77.090 42.040 77.175 42.200 ;
        RECT 79.285 42.165 79.335 42.200 ;
        POLYGON 79.335 42.200 79.370 42.165 79.335 42.165 ;
        RECT 79.285 42.040 79.370 42.165 ;
        RECT 79.990 42.040 80.075 42.200 ;
        RECT 82.185 42.165 82.235 42.200 ;
        POLYGON 82.235 42.200 82.270 42.165 82.235 42.165 ;
        RECT 82.185 42.040 82.270 42.165 ;
        RECT 82.890 42.040 82.975 42.200 ;
        RECT 85.085 42.165 85.135 42.200 ;
        POLYGON 85.135 42.200 85.170 42.165 85.135 42.165 ;
        RECT 85.085 42.040 85.170 42.165 ;
        RECT 85.790 42.040 85.875 42.200 ;
        RECT 87.985 42.165 88.035 42.200 ;
        POLYGON 88.035 42.200 88.070 42.165 88.035 42.165 ;
        RECT 87.985 42.040 88.070 42.165 ;
        RECT 88.690 42.040 88.775 42.200 ;
        RECT 90.885 42.165 90.935 42.200 ;
        POLYGON 90.935 42.200 90.970 42.165 90.935 42.165 ;
        RECT 90.885 42.040 90.970 42.165 ;
        RECT 91.590 42.040 91.675 42.200 ;
        RECT 0.775 41.420 0.850 41.560 ;
        RECT 0.990 41.370 1.065 41.510 ;
        RECT 1.695 41.430 1.755 41.510 ;
        POLYGON 1.695 41.430 1.755 41.430 1.755 41.370 ;
        RECT 1.910 41.420 1.985 41.560 ;
        RECT 3.675 41.420 3.750 41.560 ;
        RECT 3.890 41.370 3.965 41.510 ;
        RECT 4.595 41.430 4.655 41.510 ;
        POLYGON 4.595 41.430 4.655 41.430 4.655 41.370 ;
        RECT 4.810 41.420 4.885 41.560 ;
        RECT 6.575 41.420 6.650 41.560 ;
        RECT 6.790 41.370 6.865 41.510 ;
        RECT 7.495 41.430 7.555 41.510 ;
        POLYGON 7.495 41.430 7.555 41.430 7.555 41.370 ;
        RECT 7.710 41.420 7.785 41.560 ;
        RECT 9.475 41.420 9.550 41.560 ;
        RECT 9.690 41.370 9.765 41.510 ;
        RECT 10.395 41.430 10.455 41.510 ;
        POLYGON 10.395 41.430 10.455 41.430 10.455 41.370 ;
        RECT 10.610 41.420 10.685 41.560 ;
        RECT 12.375 41.420 12.450 41.560 ;
        RECT 12.590 41.370 12.665 41.510 ;
        RECT 13.295 41.430 13.355 41.510 ;
        POLYGON 13.295 41.430 13.355 41.430 13.355 41.370 ;
        RECT 13.510 41.420 13.585 41.560 ;
        RECT 15.275 41.420 15.350 41.560 ;
        RECT 15.490 41.370 15.565 41.510 ;
        RECT 16.195 41.430 16.255 41.510 ;
        POLYGON 16.195 41.430 16.255 41.430 16.255 41.370 ;
        RECT 16.410 41.420 16.485 41.560 ;
        RECT 18.175 41.420 18.250 41.560 ;
        RECT 18.390 41.370 18.465 41.510 ;
        RECT 19.095 41.430 19.155 41.510 ;
        POLYGON 19.095 41.430 19.155 41.430 19.155 41.370 ;
        RECT 19.310 41.420 19.385 41.560 ;
        RECT 21.075 41.420 21.150 41.560 ;
        RECT 21.290 41.370 21.365 41.510 ;
        RECT 21.995 41.430 22.055 41.510 ;
        POLYGON 21.995 41.430 22.055 41.430 22.055 41.370 ;
        RECT 22.210 41.420 22.285 41.560 ;
        RECT 23.975 41.420 24.050 41.560 ;
        RECT 24.190 41.370 24.265 41.510 ;
        RECT 24.895 41.430 24.955 41.510 ;
        POLYGON 24.895 41.430 24.955 41.430 24.955 41.370 ;
        RECT 25.110 41.420 25.185 41.560 ;
        RECT 26.875 41.420 26.950 41.560 ;
        RECT 27.090 41.370 27.165 41.510 ;
        RECT 27.795 41.430 27.855 41.510 ;
        POLYGON 27.795 41.430 27.855 41.430 27.855 41.370 ;
        RECT 28.010 41.420 28.085 41.560 ;
        RECT 29.775 41.420 29.850 41.560 ;
        RECT 29.990 41.370 30.065 41.510 ;
        RECT 30.695 41.430 30.755 41.510 ;
        POLYGON 30.695 41.430 30.755 41.430 30.755 41.370 ;
        RECT 30.910 41.420 30.985 41.560 ;
        RECT 32.675 41.420 32.750 41.560 ;
        RECT 32.890 41.370 32.965 41.510 ;
        RECT 33.595 41.430 33.655 41.510 ;
        POLYGON 33.595 41.430 33.655 41.430 33.655 41.370 ;
        RECT 33.810 41.420 33.885 41.560 ;
        RECT 35.575 41.420 35.650 41.560 ;
        RECT 35.790 41.370 35.865 41.510 ;
        RECT 36.495 41.430 36.555 41.510 ;
        POLYGON 36.495 41.430 36.555 41.430 36.555 41.370 ;
        RECT 36.710 41.420 36.785 41.560 ;
        RECT 38.475 41.420 38.550 41.560 ;
        RECT 38.690 41.370 38.765 41.510 ;
        RECT 39.395 41.430 39.455 41.510 ;
        POLYGON 39.395 41.430 39.455 41.430 39.455 41.370 ;
        RECT 39.610 41.420 39.685 41.560 ;
        RECT 41.375 41.420 41.450 41.560 ;
        RECT 41.590 41.370 41.665 41.510 ;
        RECT 42.295 41.430 42.355 41.510 ;
        POLYGON 42.295 41.430 42.355 41.430 42.355 41.370 ;
        RECT 42.510 41.420 42.585 41.560 ;
        RECT 44.275 41.420 44.350 41.560 ;
        RECT 44.490 41.370 44.565 41.510 ;
        RECT 45.195 41.430 45.255 41.510 ;
        POLYGON 45.195 41.430 45.255 41.430 45.255 41.370 ;
        RECT 45.410 41.420 45.485 41.560 ;
        RECT 47.175 41.420 47.250 41.560 ;
        RECT 47.390 41.370 47.465 41.510 ;
        RECT 48.095 41.430 48.155 41.510 ;
        POLYGON 48.095 41.430 48.155 41.430 48.155 41.370 ;
        RECT 48.310 41.420 48.385 41.560 ;
        RECT 50.075 41.420 50.150 41.560 ;
        RECT 50.290 41.370 50.365 41.510 ;
        RECT 50.995 41.430 51.055 41.510 ;
        POLYGON 50.995 41.430 51.055 41.430 51.055 41.370 ;
        RECT 51.210 41.420 51.285 41.560 ;
        RECT 52.975 41.420 53.050 41.560 ;
        RECT 53.190 41.370 53.265 41.510 ;
        RECT 53.895 41.430 53.955 41.510 ;
        POLYGON 53.895 41.430 53.955 41.430 53.955 41.370 ;
        RECT 54.110 41.420 54.185 41.560 ;
        RECT 55.875 41.420 55.950 41.560 ;
        RECT 56.090 41.370 56.165 41.510 ;
        RECT 56.795 41.430 56.855 41.510 ;
        POLYGON 56.795 41.430 56.855 41.430 56.855 41.370 ;
        RECT 57.010 41.420 57.085 41.560 ;
        RECT 58.775 41.420 58.850 41.560 ;
        RECT 58.990 41.370 59.065 41.510 ;
        RECT 59.695 41.430 59.755 41.510 ;
        POLYGON 59.695 41.430 59.755 41.430 59.755 41.370 ;
        RECT 59.910 41.420 59.985 41.560 ;
        RECT 61.675 41.420 61.750 41.560 ;
        RECT 61.890 41.370 61.965 41.510 ;
        RECT 62.595 41.430 62.655 41.510 ;
        POLYGON 62.595 41.430 62.655 41.430 62.655 41.370 ;
        RECT 62.810 41.420 62.885 41.560 ;
        RECT 64.575 41.420 64.650 41.560 ;
        RECT 64.790 41.370 64.865 41.510 ;
        RECT 65.495 41.430 65.555 41.510 ;
        POLYGON 65.495 41.430 65.555 41.430 65.555 41.370 ;
        RECT 65.710 41.420 65.785 41.560 ;
        RECT 67.475 41.420 67.550 41.560 ;
        RECT 67.690 41.370 67.765 41.510 ;
        RECT 68.395 41.430 68.455 41.510 ;
        POLYGON 68.395 41.430 68.455 41.430 68.455 41.370 ;
        RECT 68.610 41.420 68.685 41.560 ;
        RECT 70.375 41.420 70.450 41.560 ;
        RECT 70.590 41.370 70.665 41.510 ;
        RECT 71.295 41.430 71.355 41.510 ;
        POLYGON 71.295 41.430 71.355 41.430 71.355 41.370 ;
        RECT 71.510 41.420 71.585 41.560 ;
        RECT 73.275 41.420 73.350 41.560 ;
        RECT 73.490 41.370 73.565 41.510 ;
        RECT 74.195 41.430 74.255 41.510 ;
        POLYGON 74.195 41.430 74.255 41.430 74.255 41.370 ;
        RECT 74.410 41.420 74.485 41.560 ;
        RECT 76.175 41.420 76.250 41.560 ;
        RECT 76.390 41.370 76.465 41.510 ;
        RECT 77.095 41.430 77.155 41.510 ;
        POLYGON 77.095 41.430 77.155 41.430 77.155 41.370 ;
        RECT 77.310 41.420 77.385 41.560 ;
        RECT 79.075 41.420 79.150 41.560 ;
        RECT 79.290 41.370 79.365 41.510 ;
        RECT 79.995 41.430 80.055 41.510 ;
        POLYGON 79.995 41.430 80.055 41.430 80.055 41.370 ;
        RECT 80.210 41.420 80.285 41.560 ;
        RECT 81.975 41.420 82.050 41.560 ;
        RECT 82.190 41.370 82.265 41.510 ;
        RECT 82.895 41.430 82.955 41.510 ;
        POLYGON 82.895 41.430 82.955 41.430 82.955 41.370 ;
        RECT 83.110 41.420 83.185 41.560 ;
        RECT 84.875 41.420 84.950 41.560 ;
        RECT 85.090 41.370 85.165 41.510 ;
        RECT 85.795 41.430 85.855 41.510 ;
        POLYGON 85.795 41.430 85.855 41.430 85.855 41.370 ;
        RECT 86.010 41.420 86.085 41.560 ;
        RECT 87.775 41.420 87.850 41.560 ;
        RECT 87.990 41.370 88.065 41.510 ;
        RECT 88.695 41.430 88.755 41.510 ;
        POLYGON 88.695 41.430 88.755 41.430 88.755 41.370 ;
        RECT 88.910 41.420 88.985 41.560 ;
        RECT 90.675 41.420 90.750 41.560 ;
        RECT 90.890 41.370 90.965 41.510 ;
        RECT 91.595 41.430 91.655 41.510 ;
        POLYGON 91.595 41.430 91.655 41.430 91.655 41.370 ;
        RECT 91.810 41.420 91.885 41.560 ;
        RECT 0.720 40.900 0.870 41.070 ;
        RECT 1.110 41.035 1.260 41.205 ;
        RECT 1.500 41.035 1.650 41.205 ;
        RECT 1.890 40.900 2.040 41.070 ;
        RECT 3.620 40.900 3.770 41.070 ;
        RECT 4.010 41.035 4.160 41.205 ;
        RECT 4.400 41.035 4.550 41.205 ;
        RECT 4.790 40.900 4.940 41.070 ;
        RECT 6.520 40.900 6.670 41.070 ;
        RECT 6.910 41.035 7.060 41.205 ;
        RECT 7.300 41.035 7.450 41.205 ;
        RECT 7.690 40.900 7.840 41.070 ;
        RECT 9.420 40.900 9.570 41.070 ;
        RECT 9.810 41.035 9.960 41.205 ;
        RECT 10.200 41.035 10.350 41.205 ;
        RECT 10.590 40.900 10.740 41.070 ;
        RECT 12.320 40.900 12.470 41.070 ;
        RECT 12.710 41.035 12.860 41.205 ;
        RECT 13.100 41.035 13.250 41.205 ;
        RECT 13.490 40.900 13.640 41.070 ;
        RECT 15.220 40.900 15.370 41.070 ;
        RECT 15.610 41.035 15.760 41.205 ;
        RECT 16.000 41.035 16.150 41.205 ;
        RECT 16.390 40.900 16.540 41.070 ;
        RECT 18.120 40.900 18.270 41.070 ;
        RECT 18.510 41.035 18.660 41.205 ;
        RECT 18.900 41.035 19.050 41.205 ;
        RECT 19.290 40.900 19.440 41.070 ;
        RECT 21.020 40.900 21.170 41.070 ;
        RECT 21.410 41.035 21.560 41.205 ;
        RECT 21.800 41.035 21.950 41.205 ;
        RECT 22.190 40.900 22.340 41.070 ;
        RECT 23.920 40.900 24.070 41.070 ;
        RECT 24.310 41.035 24.460 41.205 ;
        RECT 24.700 41.035 24.850 41.205 ;
        RECT 25.090 40.900 25.240 41.070 ;
        RECT 26.820 40.900 26.970 41.070 ;
        RECT 27.210 41.035 27.360 41.205 ;
        RECT 27.600 41.035 27.750 41.205 ;
        RECT 27.990 40.900 28.140 41.070 ;
        RECT 29.720 40.900 29.870 41.070 ;
        RECT 30.110 41.035 30.260 41.205 ;
        RECT 30.500 41.035 30.650 41.205 ;
        RECT 30.890 40.900 31.040 41.070 ;
        RECT 32.620 40.900 32.770 41.070 ;
        RECT 33.010 41.035 33.160 41.205 ;
        RECT 33.400 41.035 33.550 41.205 ;
        RECT 33.790 40.900 33.940 41.070 ;
        RECT 35.520 40.900 35.670 41.070 ;
        RECT 35.910 41.035 36.060 41.205 ;
        RECT 36.300 41.035 36.450 41.205 ;
        RECT 36.690 40.900 36.840 41.070 ;
        RECT 38.420 40.900 38.570 41.070 ;
        RECT 38.810 41.035 38.960 41.205 ;
        RECT 39.200 41.035 39.350 41.205 ;
        RECT 39.590 40.900 39.740 41.070 ;
        RECT 41.320 40.900 41.470 41.070 ;
        RECT 41.710 41.035 41.860 41.205 ;
        RECT 42.100 41.035 42.250 41.205 ;
        RECT 42.490 40.900 42.640 41.070 ;
        RECT 44.220 40.900 44.370 41.070 ;
        RECT 44.610 41.035 44.760 41.205 ;
        RECT 45.000 41.035 45.150 41.205 ;
        RECT 45.390 40.900 45.540 41.070 ;
        RECT 47.120 40.900 47.270 41.070 ;
        RECT 47.510 41.035 47.660 41.205 ;
        RECT 47.900 41.035 48.050 41.205 ;
        RECT 48.290 40.900 48.440 41.070 ;
        RECT 50.020 40.900 50.170 41.070 ;
        RECT 50.410 41.035 50.560 41.205 ;
        RECT 50.800 41.035 50.950 41.205 ;
        RECT 51.190 40.900 51.340 41.070 ;
        RECT 52.920 40.900 53.070 41.070 ;
        RECT 53.310 41.035 53.460 41.205 ;
        RECT 53.700 41.035 53.850 41.205 ;
        RECT 54.090 40.900 54.240 41.070 ;
        RECT 55.820 40.900 55.970 41.070 ;
        RECT 56.210 41.035 56.360 41.205 ;
        RECT 56.600 41.035 56.750 41.205 ;
        RECT 56.990 40.900 57.140 41.070 ;
        RECT 58.720 40.900 58.870 41.070 ;
        RECT 59.110 41.035 59.260 41.205 ;
        RECT 59.500 41.035 59.650 41.205 ;
        RECT 59.890 40.900 60.040 41.070 ;
        RECT 61.620 40.900 61.770 41.070 ;
        RECT 62.010 41.035 62.160 41.205 ;
        RECT 62.400 41.035 62.550 41.205 ;
        RECT 62.790 40.900 62.940 41.070 ;
        RECT 64.520 40.900 64.670 41.070 ;
        RECT 64.910 41.035 65.060 41.205 ;
        RECT 65.300 41.035 65.450 41.205 ;
        RECT 65.690 40.900 65.840 41.070 ;
        RECT 67.420 40.900 67.570 41.070 ;
        RECT 67.810 41.035 67.960 41.205 ;
        RECT 68.200 41.035 68.350 41.205 ;
        RECT 68.590 40.900 68.740 41.070 ;
        RECT 70.320 40.900 70.470 41.070 ;
        RECT 70.710 41.035 70.860 41.205 ;
        RECT 71.100 41.035 71.250 41.205 ;
        RECT 71.490 40.900 71.640 41.070 ;
        RECT 73.220 40.900 73.370 41.070 ;
        RECT 73.610 41.035 73.760 41.205 ;
        RECT 74.000 41.035 74.150 41.205 ;
        RECT 74.390 40.900 74.540 41.070 ;
        RECT 76.120 40.900 76.270 41.070 ;
        RECT 76.510 41.035 76.660 41.205 ;
        RECT 76.900 41.035 77.050 41.205 ;
        RECT 77.290 40.900 77.440 41.070 ;
        RECT 79.020 40.900 79.170 41.070 ;
        RECT 79.410 41.035 79.560 41.205 ;
        RECT 79.800 41.035 79.950 41.205 ;
        RECT 80.190 40.900 80.340 41.070 ;
        RECT 81.920 40.900 82.070 41.070 ;
        RECT 82.310 41.035 82.460 41.205 ;
        RECT 82.700 41.035 82.850 41.205 ;
        RECT 83.090 40.900 83.240 41.070 ;
        RECT 84.820 40.900 84.970 41.070 ;
        RECT 85.210 41.035 85.360 41.205 ;
        RECT 85.600 41.035 85.750 41.205 ;
        RECT 85.990 40.900 86.140 41.070 ;
        RECT 87.720 40.900 87.870 41.070 ;
        RECT 88.110 41.035 88.260 41.205 ;
        RECT 88.500 41.035 88.650 41.205 ;
        RECT 88.890 40.900 89.040 41.070 ;
        RECT 90.620 40.900 90.770 41.070 ;
        RECT 91.010 41.035 91.160 41.205 ;
        RECT 91.400 41.035 91.550 41.205 ;
        RECT 91.790 40.900 91.940 41.070 ;
        RECT 0.985 40.815 1.035 40.850 ;
        POLYGON 1.035 40.850 1.070 40.815 1.035 40.815 ;
        RECT 0.985 40.690 1.070 40.815 ;
        RECT 1.690 40.690 1.775 40.850 ;
        RECT 3.885 40.815 3.935 40.850 ;
        POLYGON 3.935 40.850 3.970 40.815 3.935 40.815 ;
        RECT 3.885 40.690 3.970 40.815 ;
        RECT 4.590 40.690 4.675 40.850 ;
        RECT 6.785 40.815 6.835 40.850 ;
        POLYGON 6.835 40.850 6.870 40.815 6.835 40.815 ;
        RECT 6.785 40.690 6.870 40.815 ;
        RECT 7.490 40.690 7.575 40.850 ;
        RECT 9.685 40.815 9.735 40.850 ;
        POLYGON 9.735 40.850 9.770 40.815 9.735 40.815 ;
        RECT 9.685 40.690 9.770 40.815 ;
        RECT 10.390 40.690 10.475 40.850 ;
        RECT 12.585 40.815 12.635 40.850 ;
        POLYGON 12.635 40.850 12.670 40.815 12.635 40.815 ;
        RECT 12.585 40.690 12.670 40.815 ;
        RECT 13.290 40.690 13.375 40.850 ;
        RECT 15.485 40.815 15.535 40.850 ;
        POLYGON 15.535 40.850 15.570 40.815 15.535 40.815 ;
        RECT 15.485 40.690 15.570 40.815 ;
        RECT 16.190 40.690 16.275 40.850 ;
        RECT 18.385 40.815 18.435 40.850 ;
        POLYGON 18.435 40.850 18.470 40.815 18.435 40.815 ;
        RECT 18.385 40.690 18.470 40.815 ;
        RECT 19.090 40.690 19.175 40.850 ;
        RECT 21.285 40.815 21.335 40.850 ;
        POLYGON 21.335 40.850 21.370 40.815 21.335 40.815 ;
        RECT 21.285 40.690 21.370 40.815 ;
        RECT 21.990 40.690 22.075 40.850 ;
        RECT 24.185 40.815 24.235 40.850 ;
        POLYGON 24.235 40.850 24.270 40.815 24.235 40.815 ;
        RECT 24.185 40.690 24.270 40.815 ;
        RECT 24.890 40.690 24.975 40.850 ;
        RECT 27.085 40.815 27.135 40.850 ;
        POLYGON 27.135 40.850 27.170 40.815 27.135 40.815 ;
        RECT 27.085 40.690 27.170 40.815 ;
        RECT 27.790 40.690 27.875 40.850 ;
        RECT 29.985 40.815 30.035 40.850 ;
        POLYGON 30.035 40.850 30.070 40.815 30.035 40.815 ;
        RECT 29.985 40.690 30.070 40.815 ;
        RECT 30.690 40.690 30.775 40.850 ;
        RECT 32.885 40.815 32.935 40.850 ;
        POLYGON 32.935 40.850 32.970 40.815 32.935 40.815 ;
        RECT 32.885 40.690 32.970 40.815 ;
        RECT 33.590 40.690 33.675 40.850 ;
        RECT 35.785 40.815 35.835 40.850 ;
        POLYGON 35.835 40.850 35.870 40.815 35.835 40.815 ;
        RECT 35.785 40.690 35.870 40.815 ;
        RECT 36.490 40.690 36.575 40.850 ;
        RECT 38.685 40.815 38.735 40.850 ;
        POLYGON 38.735 40.850 38.770 40.815 38.735 40.815 ;
        RECT 38.685 40.690 38.770 40.815 ;
        RECT 39.390 40.690 39.475 40.850 ;
        RECT 41.585 40.815 41.635 40.850 ;
        POLYGON 41.635 40.850 41.670 40.815 41.635 40.815 ;
        RECT 41.585 40.690 41.670 40.815 ;
        RECT 42.290 40.690 42.375 40.850 ;
        RECT 44.485 40.815 44.535 40.850 ;
        POLYGON 44.535 40.850 44.570 40.815 44.535 40.815 ;
        RECT 44.485 40.690 44.570 40.815 ;
        RECT 45.190 40.690 45.275 40.850 ;
        RECT 47.385 40.815 47.435 40.850 ;
        POLYGON 47.435 40.850 47.470 40.815 47.435 40.815 ;
        RECT 47.385 40.690 47.470 40.815 ;
        RECT 48.090 40.690 48.175 40.850 ;
        RECT 50.285 40.815 50.335 40.850 ;
        POLYGON 50.335 40.850 50.370 40.815 50.335 40.815 ;
        RECT 50.285 40.690 50.370 40.815 ;
        RECT 50.990 40.690 51.075 40.850 ;
        RECT 53.185 40.815 53.235 40.850 ;
        POLYGON 53.235 40.850 53.270 40.815 53.235 40.815 ;
        RECT 53.185 40.690 53.270 40.815 ;
        RECT 53.890 40.690 53.975 40.850 ;
        RECT 56.085 40.815 56.135 40.850 ;
        POLYGON 56.135 40.850 56.170 40.815 56.135 40.815 ;
        RECT 56.085 40.690 56.170 40.815 ;
        RECT 56.790 40.690 56.875 40.850 ;
        RECT 58.985 40.815 59.035 40.850 ;
        POLYGON 59.035 40.850 59.070 40.815 59.035 40.815 ;
        RECT 58.985 40.690 59.070 40.815 ;
        RECT 59.690 40.690 59.775 40.850 ;
        RECT 61.885 40.815 61.935 40.850 ;
        POLYGON 61.935 40.850 61.970 40.815 61.935 40.815 ;
        RECT 61.885 40.690 61.970 40.815 ;
        RECT 62.590 40.690 62.675 40.850 ;
        RECT 64.785 40.815 64.835 40.850 ;
        POLYGON 64.835 40.850 64.870 40.815 64.835 40.815 ;
        RECT 64.785 40.690 64.870 40.815 ;
        RECT 65.490 40.690 65.575 40.850 ;
        RECT 67.685 40.815 67.735 40.850 ;
        POLYGON 67.735 40.850 67.770 40.815 67.735 40.815 ;
        RECT 67.685 40.690 67.770 40.815 ;
        RECT 68.390 40.690 68.475 40.850 ;
        RECT 70.585 40.815 70.635 40.850 ;
        POLYGON 70.635 40.850 70.670 40.815 70.635 40.815 ;
        RECT 70.585 40.690 70.670 40.815 ;
        RECT 71.290 40.690 71.375 40.850 ;
        RECT 73.485 40.815 73.535 40.850 ;
        POLYGON 73.535 40.850 73.570 40.815 73.535 40.815 ;
        RECT 73.485 40.690 73.570 40.815 ;
        RECT 74.190 40.690 74.275 40.850 ;
        RECT 76.385 40.815 76.435 40.850 ;
        POLYGON 76.435 40.850 76.470 40.815 76.435 40.815 ;
        RECT 76.385 40.690 76.470 40.815 ;
        RECT 77.090 40.690 77.175 40.850 ;
        RECT 79.285 40.815 79.335 40.850 ;
        POLYGON 79.335 40.850 79.370 40.815 79.335 40.815 ;
        RECT 79.285 40.690 79.370 40.815 ;
        RECT 79.990 40.690 80.075 40.850 ;
        RECT 82.185 40.815 82.235 40.850 ;
        POLYGON 82.235 40.850 82.270 40.815 82.235 40.815 ;
        RECT 82.185 40.690 82.270 40.815 ;
        RECT 82.890 40.690 82.975 40.850 ;
        RECT 85.085 40.815 85.135 40.850 ;
        POLYGON 85.135 40.850 85.170 40.815 85.135 40.815 ;
        RECT 85.085 40.690 85.170 40.815 ;
        RECT 85.790 40.690 85.875 40.850 ;
        RECT 87.985 40.815 88.035 40.850 ;
        POLYGON 88.035 40.850 88.070 40.815 88.035 40.815 ;
        RECT 87.985 40.690 88.070 40.815 ;
        RECT 88.690 40.690 88.775 40.850 ;
        RECT 90.885 40.815 90.935 40.850 ;
        POLYGON 90.935 40.850 90.970 40.815 90.935 40.815 ;
        RECT 90.885 40.690 90.970 40.815 ;
        RECT 91.590 40.690 91.675 40.850 ;
        RECT 0.775 40.070 0.850 40.210 ;
        RECT 0.990 40.020 1.065 40.160 ;
        RECT 1.695 40.080 1.755 40.160 ;
        POLYGON 1.695 40.080 1.755 40.080 1.755 40.020 ;
        RECT 1.910 40.070 1.985 40.210 ;
        RECT 3.675 40.070 3.750 40.210 ;
        RECT 3.890 40.020 3.965 40.160 ;
        RECT 4.595 40.080 4.655 40.160 ;
        POLYGON 4.595 40.080 4.655 40.080 4.655 40.020 ;
        RECT 4.810 40.070 4.885 40.210 ;
        RECT 6.575 40.070 6.650 40.210 ;
        RECT 6.790 40.020 6.865 40.160 ;
        RECT 7.495 40.080 7.555 40.160 ;
        POLYGON 7.495 40.080 7.555 40.080 7.555 40.020 ;
        RECT 7.710 40.070 7.785 40.210 ;
        RECT 9.475 40.070 9.550 40.210 ;
        RECT 9.690 40.020 9.765 40.160 ;
        RECT 10.395 40.080 10.455 40.160 ;
        POLYGON 10.395 40.080 10.455 40.080 10.455 40.020 ;
        RECT 10.610 40.070 10.685 40.210 ;
        RECT 12.375 40.070 12.450 40.210 ;
        RECT 12.590 40.020 12.665 40.160 ;
        RECT 13.295 40.080 13.355 40.160 ;
        POLYGON 13.295 40.080 13.355 40.080 13.355 40.020 ;
        RECT 13.510 40.070 13.585 40.210 ;
        RECT 15.275 40.070 15.350 40.210 ;
        RECT 15.490 40.020 15.565 40.160 ;
        RECT 16.195 40.080 16.255 40.160 ;
        POLYGON 16.195 40.080 16.255 40.080 16.255 40.020 ;
        RECT 16.410 40.070 16.485 40.210 ;
        RECT 18.175 40.070 18.250 40.210 ;
        RECT 18.390 40.020 18.465 40.160 ;
        RECT 19.095 40.080 19.155 40.160 ;
        POLYGON 19.095 40.080 19.155 40.080 19.155 40.020 ;
        RECT 19.310 40.070 19.385 40.210 ;
        RECT 21.075 40.070 21.150 40.210 ;
        RECT 21.290 40.020 21.365 40.160 ;
        RECT 21.995 40.080 22.055 40.160 ;
        POLYGON 21.995 40.080 22.055 40.080 22.055 40.020 ;
        RECT 22.210 40.070 22.285 40.210 ;
        RECT 23.975 40.070 24.050 40.210 ;
        RECT 24.190 40.020 24.265 40.160 ;
        RECT 24.895 40.080 24.955 40.160 ;
        POLYGON 24.895 40.080 24.955 40.080 24.955 40.020 ;
        RECT 25.110 40.070 25.185 40.210 ;
        RECT 26.875 40.070 26.950 40.210 ;
        RECT 27.090 40.020 27.165 40.160 ;
        RECT 27.795 40.080 27.855 40.160 ;
        POLYGON 27.795 40.080 27.855 40.080 27.855 40.020 ;
        RECT 28.010 40.070 28.085 40.210 ;
        RECT 29.775 40.070 29.850 40.210 ;
        RECT 29.990 40.020 30.065 40.160 ;
        RECT 30.695 40.080 30.755 40.160 ;
        POLYGON 30.695 40.080 30.755 40.080 30.755 40.020 ;
        RECT 30.910 40.070 30.985 40.210 ;
        RECT 32.675 40.070 32.750 40.210 ;
        RECT 32.890 40.020 32.965 40.160 ;
        RECT 33.595 40.080 33.655 40.160 ;
        POLYGON 33.595 40.080 33.655 40.080 33.655 40.020 ;
        RECT 33.810 40.070 33.885 40.210 ;
        RECT 35.575 40.070 35.650 40.210 ;
        RECT 35.790 40.020 35.865 40.160 ;
        RECT 36.495 40.080 36.555 40.160 ;
        POLYGON 36.495 40.080 36.555 40.080 36.555 40.020 ;
        RECT 36.710 40.070 36.785 40.210 ;
        RECT 38.475 40.070 38.550 40.210 ;
        RECT 38.690 40.020 38.765 40.160 ;
        RECT 39.395 40.080 39.455 40.160 ;
        POLYGON 39.395 40.080 39.455 40.080 39.455 40.020 ;
        RECT 39.610 40.070 39.685 40.210 ;
        RECT 41.375 40.070 41.450 40.210 ;
        RECT 41.590 40.020 41.665 40.160 ;
        RECT 42.295 40.080 42.355 40.160 ;
        POLYGON 42.295 40.080 42.355 40.080 42.355 40.020 ;
        RECT 42.510 40.070 42.585 40.210 ;
        RECT 44.275 40.070 44.350 40.210 ;
        RECT 44.490 40.020 44.565 40.160 ;
        RECT 45.195 40.080 45.255 40.160 ;
        POLYGON 45.195 40.080 45.255 40.080 45.255 40.020 ;
        RECT 45.410 40.070 45.485 40.210 ;
        RECT 47.175 40.070 47.250 40.210 ;
        RECT 47.390 40.020 47.465 40.160 ;
        RECT 48.095 40.080 48.155 40.160 ;
        POLYGON 48.095 40.080 48.155 40.080 48.155 40.020 ;
        RECT 48.310 40.070 48.385 40.210 ;
        RECT 50.075 40.070 50.150 40.210 ;
        RECT 50.290 40.020 50.365 40.160 ;
        RECT 50.995 40.080 51.055 40.160 ;
        POLYGON 50.995 40.080 51.055 40.080 51.055 40.020 ;
        RECT 51.210 40.070 51.285 40.210 ;
        RECT 52.975 40.070 53.050 40.210 ;
        RECT 53.190 40.020 53.265 40.160 ;
        RECT 53.895 40.080 53.955 40.160 ;
        POLYGON 53.895 40.080 53.955 40.080 53.955 40.020 ;
        RECT 54.110 40.070 54.185 40.210 ;
        RECT 55.875 40.070 55.950 40.210 ;
        RECT 56.090 40.020 56.165 40.160 ;
        RECT 56.795 40.080 56.855 40.160 ;
        POLYGON 56.795 40.080 56.855 40.080 56.855 40.020 ;
        RECT 57.010 40.070 57.085 40.210 ;
        RECT 58.775 40.070 58.850 40.210 ;
        RECT 58.990 40.020 59.065 40.160 ;
        RECT 59.695 40.080 59.755 40.160 ;
        POLYGON 59.695 40.080 59.755 40.080 59.755 40.020 ;
        RECT 59.910 40.070 59.985 40.210 ;
        RECT 61.675 40.070 61.750 40.210 ;
        RECT 61.890 40.020 61.965 40.160 ;
        RECT 62.595 40.080 62.655 40.160 ;
        POLYGON 62.595 40.080 62.655 40.080 62.655 40.020 ;
        RECT 62.810 40.070 62.885 40.210 ;
        RECT 64.575 40.070 64.650 40.210 ;
        RECT 64.790 40.020 64.865 40.160 ;
        RECT 65.495 40.080 65.555 40.160 ;
        POLYGON 65.495 40.080 65.555 40.080 65.555 40.020 ;
        RECT 65.710 40.070 65.785 40.210 ;
        RECT 67.475 40.070 67.550 40.210 ;
        RECT 67.690 40.020 67.765 40.160 ;
        RECT 68.395 40.080 68.455 40.160 ;
        POLYGON 68.395 40.080 68.455 40.080 68.455 40.020 ;
        RECT 68.610 40.070 68.685 40.210 ;
        RECT 70.375 40.070 70.450 40.210 ;
        RECT 70.590 40.020 70.665 40.160 ;
        RECT 71.295 40.080 71.355 40.160 ;
        POLYGON 71.295 40.080 71.355 40.080 71.355 40.020 ;
        RECT 71.510 40.070 71.585 40.210 ;
        RECT 73.275 40.070 73.350 40.210 ;
        RECT 73.490 40.020 73.565 40.160 ;
        RECT 74.195 40.080 74.255 40.160 ;
        POLYGON 74.195 40.080 74.255 40.080 74.255 40.020 ;
        RECT 74.410 40.070 74.485 40.210 ;
        RECT 76.175 40.070 76.250 40.210 ;
        RECT 76.390 40.020 76.465 40.160 ;
        RECT 77.095 40.080 77.155 40.160 ;
        POLYGON 77.095 40.080 77.155 40.080 77.155 40.020 ;
        RECT 77.310 40.070 77.385 40.210 ;
        RECT 79.075 40.070 79.150 40.210 ;
        RECT 79.290 40.020 79.365 40.160 ;
        RECT 79.995 40.080 80.055 40.160 ;
        POLYGON 79.995 40.080 80.055 40.080 80.055 40.020 ;
        RECT 80.210 40.070 80.285 40.210 ;
        RECT 81.975 40.070 82.050 40.210 ;
        RECT 82.190 40.020 82.265 40.160 ;
        RECT 82.895 40.080 82.955 40.160 ;
        POLYGON 82.895 40.080 82.955 40.080 82.955 40.020 ;
        RECT 83.110 40.070 83.185 40.210 ;
        RECT 84.875 40.070 84.950 40.210 ;
        RECT 85.090 40.020 85.165 40.160 ;
        RECT 85.795 40.080 85.855 40.160 ;
        POLYGON 85.795 40.080 85.855 40.080 85.855 40.020 ;
        RECT 86.010 40.070 86.085 40.210 ;
        RECT 87.775 40.070 87.850 40.210 ;
        RECT 87.990 40.020 88.065 40.160 ;
        RECT 88.695 40.080 88.755 40.160 ;
        POLYGON 88.695 40.080 88.755 40.080 88.755 40.020 ;
        RECT 88.910 40.070 88.985 40.210 ;
        RECT 90.675 40.070 90.750 40.210 ;
        RECT 90.890 40.020 90.965 40.160 ;
        RECT 91.595 40.080 91.655 40.160 ;
        POLYGON 91.595 40.080 91.655 40.080 91.655 40.020 ;
        RECT 91.810 40.070 91.885 40.210 ;
        RECT 0.720 39.550 0.870 39.720 ;
        RECT 1.110 39.685 1.260 39.855 ;
        RECT 1.500 39.685 1.650 39.855 ;
        RECT 1.890 39.550 2.040 39.720 ;
        RECT 3.620 39.550 3.770 39.720 ;
        RECT 4.010 39.685 4.160 39.855 ;
        RECT 4.400 39.685 4.550 39.855 ;
        RECT 4.790 39.550 4.940 39.720 ;
        RECT 6.520 39.550 6.670 39.720 ;
        RECT 6.910 39.685 7.060 39.855 ;
        RECT 7.300 39.685 7.450 39.855 ;
        RECT 7.690 39.550 7.840 39.720 ;
        RECT 9.420 39.550 9.570 39.720 ;
        RECT 9.810 39.685 9.960 39.855 ;
        RECT 10.200 39.685 10.350 39.855 ;
        RECT 10.590 39.550 10.740 39.720 ;
        RECT 12.320 39.550 12.470 39.720 ;
        RECT 12.710 39.685 12.860 39.855 ;
        RECT 13.100 39.685 13.250 39.855 ;
        RECT 13.490 39.550 13.640 39.720 ;
        RECT 15.220 39.550 15.370 39.720 ;
        RECT 15.610 39.685 15.760 39.855 ;
        RECT 16.000 39.685 16.150 39.855 ;
        RECT 16.390 39.550 16.540 39.720 ;
        RECT 18.120 39.550 18.270 39.720 ;
        RECT 18.510 39.685 18.660 39.855 ;
        RECT 18.900 39.685 19.050 39.855 ;
        RECT 19.290 39.550 19.440 39.720 ;
        RECT 21.020 39.550 21.170 39.720 ;
        RECT 21.410 39.685 21.560 39.855 ;
        RECT 21.800 39.685 21.950 39.855 ;
        RECT 22.190 39.550 22.340 39.720 ;
        RECT 23.920 39.550 24.070 39.720 ;
        RECT 24.310 39.685 24.460 39.855 ;
        RECT 24.700 39.685 24.850 39.855 ;
        RECT 25.090 39.550 25.240 39.720 ;
        RECT 26.820 39.550 26.970 39.720 ;
        RECT 27.210 39.685 27.360 39.855 ;
        RECT 27.600 39.685 27.750 39.855 ;
        RECT 27.990 39.550 28.140 39.720 ;
        RECT 29.720 39.550 29.870 39.720 ;
        RECT 30.110 39.685 30.260 39.855 ;
        RECT 30.500 39.685 30.650 39.855 ;
        RECT 30.890 39.550 31.040 39.720 ;
        RECT 32.620 39.550 32.770 39.720 ;
        RECT 33.010 39.685 33.160 39.855 ;
        RECT 33.400 39.685 33.550 39.855 ;
        RECT 33.790 39.550 33.940 39.720 ;
        RECT 35.520 39.550 35.670 39.720 ;
        RECT 35.910 39.685 36.060 39.855 ;
        RECT 36.300 39.685 36.450 39.855 ;
        RECT 36.690 39.550 36.840 39.720 ;
        RECT 38.420 39.550 38.570 39.720 ;
        RECT 38.810 39.685 38.960 39.855 ;
        RECT 39.200 39.685 39.350 39.855 ;
        RECT 39.590 39.550 39.740 39.720 ;
        RECT 41.320 39.550 41.470 39.720 ;
        RECT 41.710 39.685 41.860 39.855 ;
        RECT 42.100 39.685 42.250 39.855 ;
        RECT 42.490 39.550 42.640 39.720 ;
        RECT 44.220 39.550 44.370 39.720 ;
        RECT 44.610 39.685 44.760 39.855 ;
        RECT 45.000 39.685 45.150 39.855 ;
        RECT 45.390 39.550 45.540 39.720 ;
        RECT 47.120 39.550 47.270 39.720 ;
        RECT 47.510 39.685 47.660 39.855 ;
        RECT 47.900 39.685 48.050 39.855 ;
        RECT 48.290 39.550 48.440 39.720 ;
        RECT 50.020 39.550 50.170 39.720 ;
        RECT 50.410 39.685 50.560 39.855 ;
        RECT 50.800 39.685 50.950 39.855 ;
        RECT 51.190 39.550 51.340 39.720 ;
        RECT 52.920 39.550 53.070 39.720 ;
        RECT 53.310 39.685 53.460 39.855 ;
        RECT 53.700 39.685 53.850 39.855 ;
        RECT 54.090 39.550 54.240 39.720 ;
        RECT 55.820 39.550 55.970 39.720 ;
        RECT 56.210 39.685 56.360 39.855 ;
        RECT 56.600 39.685 56.750 39.855 ;
        RECT 56.990 39.550 57.140 39.720 ;
        RECT 58.720 39.550 58.870 39.720 ;
        RECT 59.110 39.685 59.260 39.855 ;
        RECT 59.500 39.685 59.650 39.855 ;
        RECT 59.890 39.550 60.040 39.720 ;
        RECT 61.620 39.550 61.770 39.720 ;
        RECT 62.010 39.685 62.160 39.855 ;
        RECT 62.400 39.685 62.550 39.855 ;
        RECT 62.790 39.550 62.940 39.720 ;
        RECT 64.520 39.550 64.670 39.720 ;
        RECT 64.910 39.685 65.060 39.855 ;
        RECT 65.300 39.685 65.450 39.855 ;
        RECT 65.690 39.550 65.840 39.720 ;
        RECT 67.420 39.550 67.570 39.720 ;
        RECT 67.810 39.685 67.960 39.855 ;
        RECT 68.200 39.685 68.350 39.855 ;
        RECT 68.590 39.550 68.740 39.720 ;
        RECT 70.320 39.550 70.470 39.720 ;
        RECT 70.710 39.685 70.860 39.855 ;
        RECT 71.100 39.685 71.250 39.855 ;
        RECT 71.490 39.550 71.640 39.720 ;
        RECT 73.220 39.550 73.370 39.720 ;
        RECT 73.610 39.685 73.760 39.855 ;
        RECT 74.000 39.685 74.150 39.855 ;
        RECT 74.390 39.550 74.540 39.720 ;
        RECT 76.120 39.550 76.270 39.720 ;
        RECT 76.510 39.685 76.660 39.855 ;
        RECT 76.900 39.685 77.050 39.855 ;
        RECT 77.290 39.550 77.440 39.720 ;
        RECT 79.020 39.550 79.170 39.720 ;
        RECT 79.410 39.685 79.560 39.855 ;
        RECT 79.800 39.685 79.950 39.855 ;
        RECT 80.190 39.550 80.340 39.720 ;
        RECT 81.920 39.550 82.070 39.720 ;
        RECT 82.310 39.685 82.460 39.855 ;
        RECT 82.700 39.685 82.850 39.855 ;
        RECT 83.090 39.550 83.240 39.720 ;
        RECT 84.820 39.550 84.970 39.720 ;
        RECT 85.210 39.685 85.360 39.855 ;
        RECT 85.600 39.685 85.750 39.855 ;
        RECT 85.990 39.550 86.140 39.720 ;
        RECT 87.720 39.550 87.870 39.720 ;
        RECT 88.110 39.685 88.260 39.855 ;
        RECT 88.500 39.685 88.650 39.855 ;
        RECT 88.890 39.550 89.040 39.720 ;
        RECT 90.620 39.550 90.770 39.720 ;
        RECT 91.010 39.685 91.160 39.855 ;
        RECT 91.400 39.685 91.550 39.855 ;
        RECT 91.790 39.550 91.940 39.720 ;
        RECT 0.985 39.465 1.035 39.500 ;
        POLYGON 1.035 39.500 1.070 39.465 1.035 39.465 ;
        RECT 0.985 39.340 1.070 39.465 ;
        RECT 1.690 39.340 1.775 39.500 ;
        RECT 3.885 39.465 3.935 39.500 ;
        POLYGON 3.935 39.500 3.970 39.465 3.935 39.465 ;
        RECT 3.885 39.340 3.970 39.465 ;
        RECT 4.590 39.340 4.675 39.500 ;
        RECT 6.785 39.465 6.835 39.500 ;
        POLYGON 6.835 39.500 6.870 39.465 6.835 39.465 ;
        RECT 6.785 39.340 6.870 39.465 ;
        RECT 7.490 39.340 7.575 39.500 ;
        RECT 9.685 39.465 9.735 39.500 ;
        POLYGON 9.735 39.500 9.770 39.465 9.735 39.465 ;
        RECT 9.685 39.340 9.770 39.465 ;
        RECT 10.390 39.340 10.475 39.500 ;
        RECT 12.585 39.465 12.635 39.500 ;
        POLYGON 12.635 39.500 12.670 39.465 12.635 39.465 ;
        RECT 12.585 39.340 12.670 39.465 ;
        RECT 13.290 39.340 13.375 39.500 ;
        RECT 15.485 39.465 15.535 39.500 ;
        POLYGON 15.535 39.500 15.570 39.465 15.535 39.465 ;
        RECT 15.485 39.340 15.570 39.465 ;
        RECT 16.190 39.340 16.275 39.500 ;
        RECT 18.385 39.465 18.435 39.500 ;
        POLYGON 18.435 39.500 18.470 39.465 18.435 39.465 ;
        RECT 18.385 39.340 18.470 39.465 ;
        RECT 19.090 39.340 19.175 39.500 ;
        RECT 21.285 39.465 21.335 39.500 ;
        POLYGON 21.335 39.500 21.370 39.465 21.335 39.465 ;
        RECT 21.285 39.340 21.370 39.465 ;
        RECT 21.990 39.340 22.075 39.500 ;
        RECT 24.185 39.465 24.235 39.500 ;
        POLYGON 24.235 39.500 24.270 39.465 24.235 39.465 ;
        RECT 24.185 39.340 24.270 39.465 ;
        RECT 24.890 39.340 24.975 39.500 ;
        RECT 27.085 39.465 27.135 39.500 ;
        POLYGON 27.135 39.500 27.170 39.465 27.135 39.465 ;
        RECT 27.085 39.340 27.170 39.465 ;
        RECT 27.790 39.340 27.875 39.500 ;
        RECT 29.985 39.465 30.035 39.500 ;
        POLYGON 30.035 39.500 30.070 39.465 30.035 39.465 ;
        RECT 29.985 39.340 30.070 39.465 ;
        RECT 30.690 39.340 30.775 39.500 ;
        RECT 32.885 39.465 32.935 39.500 ;
        POLYGON 32.935 39.500 32.970 39.465 32.935 39.465 ;
        RECT 32.885 39.340 32.970 39.465 ;
        RECT 33.590 39.340 33.675 39.500 ;
        RECT 35.785 39.465 35.835 39.500 ;
        POLYGON 35.835 39.500 35.870 39.465 35.835 39.465 ;
        RECT 35.785 39.340 35.870 39.465 ;
        RECT 36.490 39.340 36.575 39.500 ;
        RECT 38.685 39.465 38.735 39.500 ;
        POLYGON 38.735 39.500 38.770 39.465 38.735 39.465 ;
        RECT 38.685 39.340 38.770 39.465 ;
        RECT 39.390 39.340 39.475 39.500 ;
        RECT 41.585 39.465 41.635 39.500 ;
        POLYGON 41.635 39.500 41.670 39.465 41.635 39.465 ;
        RECT 41.585 39.340 41.670 39.465 ;
        RECT 42.290 39.340 42.375 39.500 ;
        RECT 44.485 39.465 44.535 39.500 ;
        POLYGON 44.535 39.500 44.570 39.465 44.535 39.465 ;
        RECT 44.485 39.340 44.570 39.465 ;
        RECT 45.190 39.340 45.275 39.500 ;
        RECT 47.385 39.465 47.435 39.500 ;
        POLYGON 47.435 39.500 47.470 39.465 47.435 39.465 ;
        RECT 47.385 39.340 47.470 39.465 ;
        RECT 48.090 39.340 48.175 39.500 ;
        RECT 50.285 39.465 50.335 39.500 ;
        POLYGON 50.335 39.500 50.370 39.465 50.335 39.465 ;
        RECT 50.285 39.340 50.370 39.465 ;
        RECT 50.990 39.340 51.075 39.500 ;
        RECT 53.185 39.465 53.235 39.500 ;
        POLYGON 53.235 39.500 53.270 39.465 53.235 39.465 ;
        RECT 53.185 39.340 53.270 39.465 ;
        RECT 53.890 39.340 53.975 39.500 ;
        RECT 56.085 39.465 56.135 39.500 ;
        POLYGON 56.135 39.500 56.170 39.465 56.135 39.465 ;
        RECT 56.085 39.340 56.170 39.465 ;
        RECT 56.790 39.340 56.875 39.500 ;
        RECT 58.985 39.465 59.035 39.500 ;
        POLYGON 59.035 39.500 59.070 39.465 59.035 39.465 ;
        RECT 58.985 39.340 59.070 39.465 ;
        RECT 59.690 39.340 59.775 39.500 ;
        RECT 61.885 39.465 61.935 39.500 ;
        POLYGON 61.935 39.500 61.970 39.465 61.935 39.465 ;
        RECT 61.885 39.340 61.970 39.465 ;
        RECT 62.590 39.340 62.675 39.500 ;
        RECT 64.785 39.465 64.835 39.500 ;
        POLYGON 64.835 39.500 64.870 39.465 64.835 39.465 ;
        RECT 64.785 39.340 64.870 39.465 ;
        RECT 65.490 39.340 65.575 39.500 ;
        RECT 67.685 39.465 67.735 39.500 ;
        POLYGON 67.735 39.500 67.770 39.465 67.735 39.465 ;
        RECT 67.685 39.340 67.770 39.465 ;
        RECT 68.390 39.340 68.475 39.500 ;
        RECT 70.585 39.465 70.635 39.500 ;
        POLYGON 70.635 39.500 70.670 39.465 70.635 39.465 ;
        RECT 70.585 39.340 70.670 39.465 ;
        RECT 71.290 39.340 71.375 39.500 ;
        RECT 73.485 39.465 73.535 39.500 ;
        POLYGON 73.535 39.500 73.570 39.465 73.535 39.465 ;
        RECT 73.485 39.340 73.570 39.465 ;
        RECT 74.190 39.340 74.275 39.500 ;
        RECT 76.385 39.465 76.435 39.500 ;
        POLYGON 76.435 39.500 76.470 39.465 76.435 39.465 ;
        RECT 76.385 39.340 76.470 39.465 ;
        RECT 77.090 39.340 77.175 39.500 ;
        RECT 79.285 39.465 79.335 39.500 ;
        POLYGON 79.335 39.500 79.370 39.465 79.335 39.465 ;
        RECT 79.285 39.340 79.370 39.465 ;
        RECT 79.990 39.340 80.075 39.500 ;
        RECT 82.185 39.465 82.235 39.500 ;
        POLYGON 82.235 39.500 82.270 39.465 82.235 39.465 ;
        RECT 82.185 39.340 82.270 39.465 ;
        RECT 82.890 39.340 82.975 39.500 ;
        RECT 85.085 39.465 85.135 39.500 ;
        POLYGON 85.135 39.500 85.170 39.465 85.135 39.465 ;
        RECT 85.085 39.340 85.170 39.465 ;
        RECT 85.790 39.340 85.875 39.500 ;
        RECT 87.985 39.465 88.035 39.500 ;
        POLYGON 88.035 39.500 88.070 39.465 88.035 39.465 ;
        RECT 87.985 39.340 88.070 39.465 ;
        RECT 88.690 39.340 88.775 39.500 ;
        RECT 90.885 39.465 90.935 39.500 ;
        POLYGON 90.935 39.500 90.970 39.465 90.935 39.465 ;
        RECT 90.885 39.340 90.970 39.465 ;
        RECT 91.590 39.340 91.675 39.500 ;
        RECT 0.775 38.720 0.850 38.860 ;
        RECT 0.990 38.670 1.065 38.810 ;
        RECT 1.695 38.730 1.755 38.810 ;
        POLYGON 1.695 38.730 1.755 38.730 1.755 38.670 ;
        RECT 1.910 38.720 1.985 38.860 ;
        RECT 3.675 38.720 3.750 38.860 ;
        RECT 3.890 38.670 3.965 38.810 ;
        RECT 4.595 38.730 4.655 38.810 ;
        POLYGON 4.595 38.730 4.655 38.730 4.655 38.670 ;
        RECT 4.810 38.720 4.885 38.860 ;
        RECT 6.575 38.720 6.650 38.860 ;
        RECT 6.790 38.670 6.865 38.810 ;
        RECT 7.495 38.730 7.555 38.810 ;
        POLYGON 7.495 38.730 7.555 38.730 7.555 38.670 ;
        RECT 7.710 38.720 7.785 38.860 ;
        RECT 9.475 38.720 9.550 38.860 ;
        RECT 9.690 38.670 9.765 38.810 ;
        RECT 10.395 38.730 10.455 38.810 ;
        POLYGON 10.395 38.730 10.455 38.730 10.455 38.670 ;
        RECT 10.610 38.720 10.685 38.860 ;
        RECT 12.375 38.720 12.450 38.860 ;
        RECT 12.590 38.670 12.665 38.810 ;
        RECT 13.295 38.730 13.355 38.810 ;
        POLYGON 13.295 38.730 13.355 38.730 13.355 38.670 ;
        RECT 13.510 38.720 13.585 38.860 ;
        RECT 15.275 38.720 15.350 38.860 ;
        RECT 15.490 38.670 15.565 38.810 ;
        RECT 16.195 38.730 16.255 38.810 ;
        POLYGON 16.195 38.730 16.255 38.730 16.255 38.670 ;
        RECT 16.410 38.720 16.485 38.860 ;
        RECT 18.175 38.720 18.250 38.860 ;
        RECT 18.390 38.670 18.465 38.810 ;
        RECT 19.095 38.730 19.155 38.810 ;
        POLYGON 19.095 38.730 19.155 38.730 19.155 38.670 ;
        RECT 19.310 38.720 19.385 38.860 ;
        RECT 21.075 38.720 21.150 38.860 ;
        RECT 21.290 38.670 21.365 38.810 ;
        RECT 21.995 38.730 22.055 38.810 ;
        POLYGON 21.995 38.730 22.055 38.730 22.055 38.670 ;
        RECT 22.210 38.720 22.285 38.860 ;
        RECT 23.975 38.720 24.050 38.860 ;
        RECT 24.190 38.670 24.265 38.810 ;
        RECT 24.895 38.730 24.955 38.810 ;
        POLYGON 24.895 38.730 24.955 38.730 24.955 38.670 ;
        RECT 25.110 38.720 25.185 38.860 ;
        RECT 26.875 38.720 26.950 38.860 ;
        RECT 27.090 38.670 27.165 38.810 ;
        RECT 27.795 38.730 27.855 38.810 ;
        POLYGON 27.795 38.730 27.855 38.730 27.855 38.670 ;
        RECT 28.010 38.720 28.085 38.860 ;
        RECT 29.775 38.720 29.850 38.860 ;
        RECT 29.990 38.670 30.065 38.810 ;
        RECT 30.695 38.730 30.755 38.810 ;
        POLYGON 30.695 38.730 30.755 38.730 30.755 38.670 ;
        RECT 30.910 38.720 30.985 38.860 ;
        RECT 32.675 38.720 32.750 38.860 ;
        RECT 32.890 38.670 32.965 38.810 ;
        RECT 33.595 38.730 33.655 38.810 ;
        POLYGON 33.595 38.730 33.655 38.730 33.655 38.670 ;
        RECT 33.810 38.720 33.885 38.860 ;
        RECT 35.575 38.720 35.650 38.860 ;
        RECT 35.790 38.670 35.865 38.810 ;
        RECT 36.495 38.730 36.555 38.810 ;
        POLYGON 36.495 38.730 36.555 38.730 36.555 38.670 ;
        RECT 36.710 38.720 36.785 38.860 ;
        RECT 38.475 38.720 38.550 38.860 ;
        RECT 38.690 38.670 38.765 38.810 ;
        RECT 39.395 38.730 39.455 38.810 ;
        POLYGON 39.395 38.730 39.455 38.730 39.455 38.670 ;
        RECT 39.610 38.720 39.685 38.860 ;
        RECT 41.375 38.720 41.450 38.860 ;
        RECT 41.590 38.670 41.665 38.810 ;
        RECT 42.295 38.730 42.355 38.810 ;
        POLYGON 42.295 38.730 42.355 38.730 42.355 38.670 ;
        RECT 42.510 38.720 42.585 38.860 ;
        RECT 44.275 38.720 44.350 38.860 ;
        RECT 44.490 38.670 44.565 38.810 ;
        RECT 45.195 38.730 45.255 38.810 ;
        POLYGON 45.195 38.730 45.255 38.730 45.255 38.670 ;
        RECT 45.410 38.720 45.485 38.860 ;
        RECT 47.175 38.720 47.250 38.860 ;
        RECT 47.390 38.670 47.465 38.810 ;
        RECT 48.095 38.730 48.155 38.810 ;
        POLYGON 48.095 38.730 48.155 38.730 48.155 38.670 ;
        RECT 48.310 38.720 48.385 38.860 ;
        RECT 50.075 38.720 50.150 38.860 ;
        RECT 50.290 38.670 50.365 38.810 ;
        RECT 50.995 38.730 51.055 38.810 ;
        POLYGON 50.995 38.730 51.055 38.730 51.055 38.670 ;
        RECT 51.210 38.720 51.285 38.860 ;
        RECT 52.975 38.720 53.050 38.860 ;
        RECT 53.190 38.670 53.265 38.810 ;
        RECT 53.895 38.730 53.955 38.810 ;
        POLYGON 53.895 38.730 53.955 38.730 53.955 38.670 ;
        RECT 54.110 38.720 54.185 38.860 ;
        RECT 55.875 38.720 55.950 38.860 ;
        RECT 56.090 38.670 56.165 38.810 ;
        RECT 56.795 38.730 56.855 38.810 ;
        POLYGON 56.795 38.730 56.855 38.730 56.855 38.670 ;
        RECT 57.010 38.720 57.085 38.860 ;
        RECT 58.775 38.720 58.850 38.860 ;
        RECT 58.990 38.670 59.065 38.810 ;
        RECT 59.695 38.730 59.755 38.810 ;
        POLYGON 59.695 38.730 59.755 38.730 59.755 38.670 ;
        RECT 59.910 38.720 59.985 38.860 ;
        RECT 61.675 38.720 61.750 38.860 ;
        RECT 61.890 38.670 61.965 38.810 ;
        RECT 62.595 38.730 62.655 38.810 ;
        POLYGON 62.595 38.730 62.655 38.730 62.655 38.670 ;
        RECT 62.810 38.720 62.885 38.860 ;
        RECT 64.575 38.720 64.650 38.860 ;
        RECT 64.790 38.670 64.865 38.810 ;
        RECT 65.495 38.730 65.555 38.810 ;
        POLYGON 65.495 38.730 65.555 38.730 65.555 38.670 ;
        RECT 65.710 38.720 65.785 38.860 ;
        RECT 67.475 38.720 67.550 38.860 ;
        RECT 67.690 38.670 67.765 38.810 ;
        RECT 68.395 38.730 68.455 38.810 ;
        POLYGON 68.395 38.730 68.455 38.730 68.455 38.670 ;
        RECT 68.610 38.720 68.685 38.860 ;
        RECT 70.375 38.720 70.450 38.860 ;
        RECT 70.590 38.670 70.665 38.810 ;
        RECT 71.295 38.730 71.355 38.810 ;
        POLYGON 71.295 38.730 71.355 38.730 71.355 38.670 ;
        RECT 71.510 38.720 71.585 38.860 ;
        RECT 73.275 38.720 73.350 38.860 ;
        RECT 73.490 38.670 73.565 38.810 ;
        RECT 74.195 38.730 74.255 38.810 ;
        POLYGON 74.195 38.730 74.255 38.730 74.255 38.670 ;
        RECT 74.410 38.720 74.485 38.860 ;
        RECT 76.175 38.720 76.250 38.860 ;
        RECT 76.390 38.670 76.465 38.810 ;
        RECT 77.095 38.730 77.155 38.810 ;
        POLYGON 77.095 38.730 77.155 38.730 77.155 38.670 ;
        RECT 77.310 38.720 77.385 38.860 ;
        RECT 79.075 38.720 79.150 38.860 ;
        RECT 79.290 38.670 79.365 38.810 ;
        RECT 79.995 38.730 80.055 38.810 ;
        POLYGON 79.995 38.730 80.055 38.730 80.055 38.670 ;
        RECT 80.210 38.720 80.285 38.860 ;
        RECT 81.975 38.720 82.050 38.860 ;
        RECT 82.190 38.670 82.265 38.810 ;
        RECT 82.895 38.730 82.955 38.810 ;
        POLYGON 82.895 38.730 82.955 38.730 82.955 38.670 ;
        RECT 83.110 38.720 83.185 38.860 ;
        RECT 84.875 38.720 84.950 38.860 ;
        RECT 85.090 38.670 85.165 38.810 ;
        RECT 85.795 38.730 85.855 38.810 ;
        POLYGON 85.795 38.730 85.855 38.730 85.855 38.670 ;
        RECT 86.010 38.720 86.085 38.860 ;
        RECT 87.775 38.720 87.850 38.860 ;
        RECT 87.990 38.670 88.065 38.810 ;
        RECT 88.695 38.730 88.755 38.810 ;
        POLYGON 88.695 38.730 88.755 38.730 88.755 38.670 ;
        RECT 88.910 38.720 88.985 38.860 ;
        RECT 90.675 38.720 90.750 38.860 ;
        RECT 90.890 38.670 90.965 38.810 ;
        RECT 91.595 38.730 91.655 38.810 ;
        POLYGON 91.595 38.730 91.655 38.730 91.655 38.670 ;
        RECT 91.810 38.720 91.885 38.860 ;
        RECT 0.720 38.200 0.870 38.370 ;
        RECT 1.110 38.335 1.260 38.505 ;
        RECT 1.500 38.335 1.650 38.505 ;
        RECT 1.890 38.200 2.040 38.370 ;
        RECT 3.620 38.200 3.770 38.370 ;
        RECT 4.010 38.335 4.160 38.505 ;
        RECT 4.400 38.335 4.550 38.505 ;
        RECT 4.790 38.200 4.940 38.370 ;
        RECT 6.520 38.200 6.670 38.370 ;
        RECT 6.910 38.335 7.060 38.505 ;
        RECT 7.300 38.335 7.450 38.505 ;
        RECT 7.690 38.200 7.840 38.370 ;
        RECT 9.420 38.200 9.570 38.370 ;
        RECT 9.810 38.335 9.960 38.505 ;
        RECT 10.200 38.335 10.350 38.505 ;
        RECT 10.590 38.200 10.740 38.370 ;
        RECT 12.320 38.200 12.470 38.370 ;
        RECT 12.710 38.335 12.860 38.505 ;
        RECT 13.100 38.335 13.250 38.505 ;
        RECT 13.490 38.200 13.640 38.370 ;
        RECT 15.220 38.200 15.370 38.370 ;
        RECT 15.610 38.335 15.760 38.505 ;
        RECT 16.000 38.335 16.150 38.505 ;
        RECT 16.390 38.200 16.540 38.370 ;
        RECT 18.120 38.200 18.270 38.370 ;
        RECT 18.510 38.335 18.660 38.505 ;
        RECT 18.900 38.335 19.050 38.505 ;
        RECT 19.290 38.200 19.440 38.370 ;
        RECT 21.020 38.200 21.170 38.370 ;
        RECT 21.410 38.335 21.560 38.505 ;
        RECT 21.800 38.335 21.950 38.505 ;
        RECT 22.190 38.200 22.340 38.370 ;
        RECT 23.415 38.310 23.565 38.480 ;
        RECT 23.920 38.200 24.070 38.370 ;
        RECT 24.310 38.335 24.460 38.505 ;
        RECT 24.700 38.335 24.850 38.505 ;
        RECT 25.090 38.200 25.240 38.370 ;
        RECT 25.595 38.310 25.745 38.480 ;
        RECT 26.315 38.310 26.465 38.480 ;
        RECT 26.820 38.200 26.970 38.370 ;
        RECT 27.210 38.335 27.360 38.505 ;
        RECT 27.600 38.335 27.750 38.505 ;
        RECT 27.990 38.200 28.140 38.370 ;
        RECT 28.495 38.310 28.645 38.480 ;
        RECT 29.215 38.310 29.365 38.480 ;
        RECT 29.720 38.200 29.870 38.370 ;
        RECT 30.110 38.335 30.260 38.505 ;
        RECT 30.500 38.335 30.650 38.505 ;
        RECT 30.890 38.200 31.040 38.370 ;
        RECT 31.395 38.310 31.545 38.480 ;
        RECT 32.115 38.310 32.265 38.480 ;
        RECT 32.620 38.200 32.770 38.370 ;
        RECT 33.010 38.335 33.160 38.505 ;
        RECT 33.400 38.335 33.550 38.505 ;
        RECT 33.790 38.200 33.940 38.370 ;
        RECT 34.295 38.310 34.445 38.480 ;
        RECT 35.015 38.310 35.165 38.480 ;
        RECT 35.520 38.200 35.670 38.370 ;
        RECT 35.910 38.335 36.060 38.505 ;
        RECT 36.300 38.335 36.450 38.505 ;
        RECT 36.690 38.200 36.840 38.370 ;
        RECT 37.195 38.310 37.345 38.480 ;
        RECT 37.915 38.310 38.065 38.480 ;
        RECT 38.420 38.200 38.570 38.370 ;
        RECT 38.810 38.335 38.960 38.505 ;
        RECT 39.200 38.335 39.350 38.505 ;
        RECT 39.590 38.200 39.740 38.370 ;
        RECT 40.095 38.310 40.245 38.480 ;
        RECT 40.815 38.310 40.965 38.480 ;
        RECT 41.320 38.200 41.470 38.370 ;
        RECT 41.710 38.335 41.860 38.505 ;
        RECT 42.100 38.335 42.250 38.505 ;
        RECT 42.490 38.200 42.640 38.370 ;
        RECT 42.995 38.310 43.145 38.480 ;
        RECT 43.715 38.310 43.865 38.480 ;
        RECT 44.220 38.200 44.370 38.370 ;
        RECT 44.610 38.335 44.760 38.505 ;
        RECT 45.000 38.335 45.150 38.505 ;
        RECT 45.390 38.200 45.540 38.370 ;
        RECT 45.895 38.310 46.045 38.480 ;
        RECT 46.615 38.310 46.765 38.480 ;
        RECT 47.120 38.200 47.270 38.370 ;
        RECT 47.510 38.335 47.660 38.505 ;
        RECT 47.900 38.335 48.050 38.505 ;
        RECT 48.290 38.200 48.440 38.370 ;
        RECT 48.795 38.310 48.945 38.480 ;
        RECT 49.515 38.310 49.665 38.480 ;
        RECT 50.020 38.200 50.170 38.370 ;
        RECT 50.410 38.335 50.560 38.505 ;
        RECT 50.800 38.335 50.950 38.505 ;
        RECT 51.190 38.200 51.340 38.370 ;
        RECT 51.695 38.310 51.845 38.480 ;
        RECT 52.415 38.310 52.565 38.480 ;
        RECT 52.920 38.200 53.070 38.370 ;
        RECT 53.310 38.335 53.460 38.505 ;
        RECT 53.700 38.335 53.850 38.505 ;
        RECT 54.090 38.200 54.240 38.370 ;
        RECT 54.595 38.310 54.745 38.480 ;
        RECT 55.315 38.310 55.465 38.480 ;
        RECT 55.820 38.200 55.970 38.370 ;
        RECT 56.210 38.335 56.360 38.505 ;
        RECT 56.600 38.335 56.750 38.505 ;
        RECT 56.990 38.200 57.140 38.370 ;
        RECT 57.495 38.310 57.645 38.480 ;
        RECT 58.215 38.310 58.365 38.480 ;
        RECT 58.720 38.200 58.870 38.370 ;
        RECT 59.110 38.335 59.260 38.505 ;
        RECT 59.500 38.335 59.650 38.505 ;
        RECT 59.890 38.200 60.040 38.370 ;
        RECT 60.395 38.310 60.545 38.480 ;
        RECT 61.115 38.310 61.265 38.480 ;
        RECT 61.620 38.200 61.770 38.370 ;
        RECT 62.010 38.335 62.160 38.505 ;
        RECT 62.400 38.335 62.550 38.505 ;
        RECT 62.790 38.200 62.940 38.370 ;
        RECT 63.295 38.310 63.445 38.480 ;
        RECT 64.015 38.310 64.165 38.480 ;
        RECT 64.520 38.200 64.670 38.370 ;
        RECT 64.910 38.335 65.060 38.505 ;
        RECT 65.300 38.335 65.450 38.505 ;
        RECT 65.690 38.200 65.840 38.370 ;
        RECT 66.195 38.310 66.345 38.480 ;
        RECT 66.915 38.310 67.065 38.480 ;
        RECT 67.420 38.200 67.570 38.370 ;
        RECT 67.810 38.335 67.960 38.505 ;
        RECT 68.200 38.335 68.350 38.505 ;
        RECT 68.590 38.200 68.740 38.370 ;
        RECT 69.095 38.310 69.245 38.480 ;
        RECT 69.815 38.310 69.965 38.480 ;
        RECT 70.320 38.200 70.470 38.370 ;
        RECT 70.710 38.335 70.860 38.505 ;
        RECT 71.100 38.335 71.250 38.505 ;
        RECT 71.490 38.200 71.640 38.370 ;
        RECT 71.995 38.310 72.145 38.480 ;
        RECT 72.715 38.310 72.865 38.480 ;
        RECT 73.220 38.200 73.370 38.370 ;
        RECT 73.610 38.335 73.760 38.505 ;
        RECT 74.000 38.335 74.150 38.505 ;
        RECT 74.390 38.200 74.540 38.370 ;
        RECT 74.895 38.310 75.045 38.480 ;
        RECT 75.615 38.310 75.765 38.480 ;
        RECT 76.120 38.200 76.270 38.370 ;
        RECT 76.510 38.335 76.660 38.505 ;
        RECT 76.900 38.335 77.050 38.505 ;
        RECT 77.290 38.200 77.440 38.370 ;
        RECT 77.795 38.310 77.945 38.480 ;
        RECT 78.515 38.310 78.665 38.480 ;
        RECT 79.020 38.200 79.170 38.370 ;
        RECT 79.410 38.335 79.560 38.505 ;
        RECT 79.800 38.335 79.950 38.505 ;
        RECT 80.190 38.200 80.340 38.370 ;
        RECT 80.695 38.310 80.845 38.480 ;
        RECT 81.415 38.310 81.565 38.480 ;
        RECT 81.920 38.200 82.070 38.370 ;
        RECT 82.310 38.335 82.460 38.505 ;
        RECT 82.700 38.335 82.850 38.505 ;
        RECT 83.090 38.200 83.240 38.370 ;
        RECT 83.595 38.310 83.745 38.480 ;
        RECT 84.315 38.310 84.465 38.480 ;
        RECT 84.820 38.200 84.970 38.370 ;
        RECT 85.210 38.335 85.360 38.505 ;
        RECT 85.600 38.335 85.750 38.505 ;
        RECT 85.990 38.200 86.140 38.370 ;
        RECT 86.495 38.310 86.645 38.480 ;
        RECT 87.215 38.310 87.365 38.480 ;
        RECT 87.720 38.200 87.870 38.370 ;
        RECT 88.110 38.335 88.260 38.505 ;
        RECT 88.500 38.335 88.650 38.505 ;
        RECT 88.890 38.200 89.040 38.370 ;
        RECT 89.395 38.310 89.545 38.480 ;
        RECT 90.115 38.310 90.265 38.480 ;
        RECT 90.620 38.200 90.770 38.370 ;
        RECT 91.010 38.335 91.160 38.505 ;
        RECT 91.400 38.335 91.550 38.505 ;
        RECT 91.790 38.200 91.940 38.370 ;
        RECT 92.295 38.310 92.445 38.480 ;
        RECT 0.985 38.115 1.035 38.150 ;
        POLYGON 1.035 38.150 1.070 38.115 1.035 38.115 ;
        RECT 0.985 37.990 1.070 38.115 ;
        RECT 1.690 37.990 1.775 38.150 ;
        RECT 3.885 38.115 3.935 38.150 ;
        POLYGON 3.935 38.150 3.970 38.115 3.935 38.115 ;
        RECT 3.885 37.990 3.970 38.115 ;
        RECT 4.590 37.990 4.675 38.150 ;
        RECT 6.785 38.115 6.835 38.150 ;
        POLYGON 6.835 38.150 6.870 38.115 6.835 38.115 ;
        RECT 6.785 37.990 6.870 38.115 ;
        RECT 7.490 37.990 7.575 38.150 ;
        RECT 9.685 38.115 9.735 38.150 ;
        POLYGON 9.735 38.150 9.770 38.115 9.735 38.115 ;
        RECT 9.685 37.990 9.770 38.115 ;
        RECT 10.390 37.990 10.475 38.150 ;
        RECT 12.585 38.115 12.635 38.150 ;
        POLYGON 12.635 38.150 12.670 38.115 12.635 38.115 ;
        RECT 12.585 37.990 12.670 38.115 ;
        RECT 13.290 37.990 13.375 38.150 ;
        RECT 15.485 38.115 15.535 38.150 ;
        POLYGON 15.535 38.150 15.570 38.115 15.535 38.115 ;
        RECT 15.485 37.990 15.570 38.115 ;
        RECT 16.190 37.990 16.275 38.150 ;
        RECT 18.385 38.115 18.435 38.150 ;
        POLYGON 18.435 38.150 18.470 38.115 18.435 38.115 ;
        RECT 18.385 37.990 18.470 38.115 ;
        RECT 19.090 37.990 19.175 38.150 ;
        RECT 21.285 38.115 21.335 38.150 ;
        POLYGON 21.335 38.150 21.370 38.115 21.335 38.115 ;
        RECT 21.285 37.990 21.370 38.115 ;
        RECT 21.990 37.990 22.075 38.150 ;
        RECT 24.185 38.115 24.235 38.150 ;
        POLYGON 24.235 38.150 24.270 38.115 24.235 38.115 ;
        RECT 24.185 37.990 24.270 38.115 ;
        RECT 24.890 37.990 24.975 38.150 ;
        RECT 27.085 38.115 27.135 38.150 ;
        POLYGON 27.135 38.150 27.170 38.115 27.135 38.115 ;
        RECT 27.085 37.990 27.170 38.115 ;
        RECT 27.790 37.990 27.875 38.150 ;
        RECT 29.985 38.115 30.035 38.150 ;
        POLYGON 30.035 38.150 30.070 38.115 30.035 38.115 ;
        RECT 29.985 37.990 30.070 38.115 ;
        RECT 30.690 37.990 30.775 38.150 ;
        RECT 32.885 38.115 32.935 38.150 ;
        POLYGON 32.935 38.150 32.970 38.115 32.935 38.115 ;
        RECT 32.885 37.990 32.970 38.115 ;
        RECT 33.590 37.990 33.675 38.150 ;
        RECT 35.785 38.115 35.835 38.150 ;
        POLYGON 35.835 38.150 35.870 38.115 35.835 38.115 ;
        RECT 35.785 37.990 35.870 38.115 ;
        RECT 36.490 37.990 36.575 38.150 ;
        RECT 38.685 38.115 38.735 38.150 ;
        POLYGON 38.735 38.150 38.770 38.115 38.735 38.115 ;
        RECT 38.685 37.990 38.770 38.115 ;
        RECT 39.390 37.990 39.475 38.150 ;
        RECT 41.585 38.115 41.635 38.150 ;
        POLYGON 41.635 38.150 41.670 38.115 41.635 38.115 ;
        RECT 41.585 37.990 41.670 38.115 ;
        RECT 42.290 37.990 42.375 38.150 ;
        RECT 44.485 38.115 44.535 38.150 ;
        POLYGON 44.535 38.150 44.570 38.115 44.535 38.115 ;
        RECT 44.485 37.990 44.570 38.115 ;
        RECT 45.190 37.990 45.275 38.150 ;
        RECT 47.385 38.115 47.435 38.150 ;
        POLYGON 47.435 38.150 47.470 38.115 47.435 38.115 ;
        RECT 47.385 37.990 47.470 38.115 ;
        RECT 48.090 37.990 48.175 38.150 ;
        RECT 50.285 38.115 50.335 38.150 ;
        POLYGON 50.335 38.150 50.370 38.115 50.335 38.115 ;
        RECT 50.285 37.990 50.370 38.115 ;
        RECT 50.990 37.990 51.075 38.150 ;
        RECT 53.185 38.115 53.235 38.150 ;
        POLYGON 53.235 38.150 53.270 38.115 53.235 38.115 ;
        RECT 53.185 37.990 53.270 38.115 ;
        RECT 53.890 37.990 53.975 38.150 ;
        RECT 56.085 38.115 56.135 38.150 ;
        POLYGON 56.135 38.150 56.170 38.115 56.135 38.115 ;
        RECT 56.085 37.990 56.170 38.115 ;
        RECT 56.790 37.990 56.875 38.150 ;
        RECT 58.985 38.115 59.035 38.150 ;
        POLYGON 59.035 38.150 59.070 38.115 59.035 38.115 ;
        RECT 58.985 37.990 59.070 38.115 ;
        RECT 59.690 37.990 59.775 38.150 ;
        RECT 61.885 38.115 61.935 38.150 ;
        POLYGON 61.935 38.150 61.970 38.115 61.935 38.115 ;
        RECT 61.885 37.990 61.970 38.115 ;
        RECT 62.590 37.990 62.675 38.150 ;
        RECT 64.785 38.115 64.835 38.150 ;
        POLYGON 64.835 38.150 64.870 38.115 64.835 38.115 ;
        RECT 64.785 37.990 64.870 38.115 ;
        RECT 65.490 37.990 65.575 38.150 ;
        RECT 67.685 38.115 67.735 38.150 ;
        POLYGON 67.735 38.150 67.770 38.115 67.735 38.115 ;
        RECT 67.685 37.990 67.770 38.115 ;
        RECT 68.390 37.990 68.475 38.150 ;
        RECT 70.585 38.115 70.635 38.150 ;
        POLYGON 70.635 38.150 70.670 38.115 70.635 38.115 ;
        RECT 70.585 37.990 70.670 38.115 ;
        RECT 71.290 37.990 71.375 38.150 ;
        RECT 73.485 38.115 73.535 38.150 ;
        POLYGON 73.535 38.150 73.570 38.115 73.535 38.115 ;
        RECT 73.485 37.990 73.570 38.115 ;
        RECT 74.190 37.990 74.275 38.150 ;
        RECT 76.385 38.115 76.435 38.150 ;
        POLYGON 76.435 38.150 76.470 38.115 76.435 38.115 ;
        RECT 76.385 37.990 76.470 38.115 ;
        RECT 77.090 37.990 77.175 38.150 ;
        RECT 79.285 38.115 79.335 38.150 ;
        POLYGON 79.335 38.150 79.370 38.115 79.335 38.115 ;
        RECT 79.285 37.990 79.370 38.115 ;
        RECT 79.990 37.990 80.075 38.150 ;
        RECT 82.185 38.115 82.235 38.150 ;
        POLYGON 82.235 38.150 82.270 38.115 82.235 38.115 ;
        RECT 82.185 37.990 82.270 38.115 ;
        RECT 82.890 37.990 82.975 38.150 ;
        RECT 85.085 38.115 85.135 38.150 ;
        POLYGON 85.135 38.150 85.170 38.115 85.135 38.115 ;
        RECT 85.085 37.990 85.170 38.115 ;
        RECT 85.790 37.990 85.875 38.150 ;
        RECT 87.985 38.115 88.035 38.150 ;
        POLYGON 88.035 38.150 88.070 38.115 88.035 38.115 ;
        RECT 87.985 37.990 88.070 38.115 ;
        RECT 88.690 37.990 88.775 38.150 ;
        RECT 90.885 38.115 90.935 38.150 ;
        POLYGON 90.935 38.150 90.970 38.115 90.935 38.115 ;
        RECT 90.885 37.990 90.970 38.115 ;
        RECT 91.590 37.990 91.675 38.150 ;
        RECT 0.775 37.370 0.850 37.510 ;
        RECT 0.990 37.320 1.065 37.460 ;
        RECT 1.695 37.380 1.755 37.460 ;
        POLYGON 1.695 37.380 1.755 37.380 1.755 37.320 ;
        RECT 1.910 37.370 1.985 37.510 ;
        RECT 3.675 37.370 3.750 37.510 ;
        RECT 3.890 37.320 3.965 37.460 ;
        RECT 4.595 37.380 4.655 37.460 ;
        POLYGON 4.595 37.380 4.655 37.380 4.655 37.320 ;
        RECT 4.810 37.370 4.885 37.510 ;
        RECT 6.575 37.370 6.650 37.510 ;
        RECT 6.790 37.320 6.865 37.460 ;
        RECT 7.495 37.380 7.555 37.460 ;
        POLYGON 7.495 37.380 7.555 37.380 7.555 37.320 ;
        RECT 7.710 37.370 7.785 37.510 ;
        RECT 9.475 37.370 9.550 37.510 ;
        RECT 9.690 37.320 9.765 37.460 ;
        RECT 10.395 37.380 10.455 37.460 ;
        POLYGON 10.395 37.380 10.455 37.380 10.455 37.320 ;
        RECT 10.610 37.370 10.685 37.510 ;
        RECT 12.375 37.370 12.450 37.510 ;
        RECT 12.590 37.320 12.665 37.460 ;
        RECT 13.295 37.380 13.355 37.460 ;
        POLYGON 13.295 37.380 13.355 37.380 13.355 37.320 ;
        RECT 13.510 37.370 13.585 37.510 ;
        RECT 15.275 37.370 15.350 37.510 ;
        RECT 15.490 37.320 15.565 37.460 ;
        RECT 16.195 37.380 16.255 37.460 ;
        POLYGON 16.195 37.380 16.255 37.380 16.255 37.320 ;
        RECT 16.410 37.370 16.485 37.510 ;
        RECT 18.175 37.370 18.250 37.510 ;
        RECT 18.390 37.320 18.465 37.460 ;
        RECT 19.095 37.380 19.155 37.460 ;
        POLYGON 19.095 37.380 19.155 37.380 19.155 37.320 ;
        RECT 19.310 37.370 19.385 37.510 ;
        RECT 21.075 37.370 21.150 37.510 ;
        RECT 21.290 37.320 21.365 37.460 ;
        RECT 21.995 37.380 22.055 37.460 ;
        POLYGON 21.995 37.380 22.055 37.380 22.055 37.320 ;
        RECT 22.210 37.370 22.285 37.510 ;
        RECT 23.975 37.370 24.050 37.510 ;
        RECT 24.190 37.320 24.265 37.460 ;
        RECT 24.895 37.380 24.955 37.460 ;
        POLYGON 24.895 37.380 24.955 37.380 24.955 37.320 ;
        RECT 25.110 37.370 25.185 37.510 ;
        RECT 26.875 37.370 26.950 37.510 ;
        RECT 27.090 37.320 27.165 37.460 ;
        RECT 27.795 37.380 27.855 37.460 ;
        POLYGON 27.795 37.380 27.855 37.380 27.855 37.320 ;
        RECT 28.010 37.370 28.085 37.510 ;
        RECT 29.775 37.370 29.850 37.510 ;
        RECT 29.990 37.320 30.065 37.460 ;
        RECT 30.695 37.380 30.755 37.460 ;
        POLYGON 30.695 37.380 30.755 37.380 30.755 37.320 ;
        RECT 30.910 37.370 30.985 37.510 ;
        RECT 32.675 37.370 32.750 37.510 ;
        RECT 32.890 37.320 32.965 37.460 ;
        RECT 33.595 37.380 33.655 37.460 ;
        POLYGON 33.595 37.380 33.655 37.380 33.655 37.320 ;
        RECT 33.810 37.370 33.885 37.510 ;
        RECT 35.575 37.370 35.650 37.510 ;
        RECT 35.790 37.320 35.865 37.460 ;
        RECT 36.495 37.380 36.555 37.460 ;
        POLYGON 36.495 37.380 36.555 37.380 36.555 37.320 ;
        RECT 36.710 37.370 36.785 37.510 ;
        RECT 38.475 37.370 38.550 37.510 ;
        RECT 38.690 37.320 38.765 37.460 ;
        RECT 39.395 37.380 39.455 37.460 ;
        POLYGON 39.395 37.380 39.455 37.380 39.455 37.320 ;
        RECT 39.610 37.370 39.685 37.510 ;
        RECT 41.375 37.370 41.450 37.510 ;
        RECT 41.590 37.320 41.665 37.460 ;
        RECT 42.295 37.380 42.355 37.460 ;
        POLYGON 42.295 37.380 42.355 37.380 42.355 37.320 ;
        RECT 42.510 37.370 42.585 37.510 ;
        RECT 44.275 37.370 44.350 37.510 ;
        RECT 44.490 37.320 44.565 37.460 ;
        RECT 45.195 37.380 45.255 37.460 ;
        POLYGON 45.195 37.380 45.255 37.380 45.255 37.320 ;
        RECT 45.410 37.370 45.485 37.510 ;
        RECT 47.175 37.370 47.250 37.510 ;
        RECT 47.390 37.320 47.465 37.460 ;
        RECT 48.095 37.380 48.155 37.460 ;
        POLYGON 48.095 37.380 48.155 37.380 48.155 37.320 ;
        RECT 48.310 37.370 48.385 37.510 ;
        RECT 50.075 37.370 50.150 37.510 ;
        RECT 50.290 37.320 50.365 37.460 ;
        RECT 50.995 37.380 51.055 37.460 ;
        POLYGON 50.995 37.380 51.055 37.380 51.055 37.320 ;
        RECT 51.210 37.370 51.285 37.510 ;
        RECT 52.975 37.370 53.050 37.510 ;
        RECT 53.190 37.320 53.265 37.460 ;
        RECT 53.895 37.380 53.955 37.460 ;
        POLYGON 53.895 37.380 53.955 37.380 53.955 37.320 ;
        RECT 54.110 37.370 54.185 37.510 ;
        RECT 55.875 37.370 55.950 37.510 ;
        RECT 56.090 37.320 56.165 37.460 ;
        RECT 56.795 37.380 56.855 37.460 ;
        POLYGON 56.795 37.380 56.855 37.380 56.855 37.320 ;
        RECT 57.010 37.370 57.085 37.510 ;
        RECT 58.775 37.370 58.850 37.510 ;
        RECT 58.990 37.320 59.065 37.460 ;
        RECT 59.695 37.380 59.755 37.460 ;
        POLYGON 59.695 37.380 59.755 37.380 59.755 37.320 ;
        RECT 59.910 37.370 59.985 37.510 ;
        RECT 61.675 37.370 61.750 37.510 ;
        RECT 61.890 37.320 61.965 37.460 ;
        RECT 62.595 37.380 62.655 37.460 ;
        POLYGON 62.595 37.380 62.655 37.380 62.655 37.320 ;
        RECT 62.810 37.370 62.885 37.510 ;
        RECT 64.575 37.370 64.650 37.510 ;
        RECT 64.790 37.320 64.865 37.460 ;
        RECT 65.495 37.380 65.555 37.460 ;
        POLYGON 65.495 37.380 65.555 37.380 65.555 37.320 ;
        RECT 65.710 37.370 65.785 37.510 ;
        RECT 67.475 37.370 67.550 37.510 ;
        RECT 67.690 37.320 67.765 37.460 ;
        RECT 68.395 37.380 68.455 37.460 ;
        POLYGON 68.395 37.380 68.455 37.380 68.455 37.320 ;
        RECT 68.610 37.370 68.685 37.510 ;
        RECT 70.375 37.370 70.450 37.510 ;
        RECT 70.590 37.320 70.665 37.460 ;
        RECT 71.295 37.380 71.355 37.460 ;
        POLYGON 71.295 37.380 71.355 37.380 71.355 37.320 ;
        RECT 71.510 37.370 71.585 37.510 ;
        RECT 73.275 37.370 73.350 37.510 ;
        RECT 73.490 37.320 73.565 37.460 ;
        RECT 74.195 37.380 74.255 37.460 ;
        POLYGON 74.195 37.380 74.255 37.380 74.255 37.320 ;
        RECT 74.410 37.370 74.485 37.510 ;
        RECT 76.175 37.370 76.250 37.510 ;
        RECT 76.390 37.320 76.465 37.460 ;
        RECT 77.095 37.380 77.155 37.460 ;
        POLYGON 77.095 37.380 77.155 37.380 77.155 37.320 ;
        RECT 77.310 37.370 77.385 37.510 ;
        RECT 79.075 37.370 79.150 37.510 ;
        RECT 79.290 37.320 79.365 37.460 ;
        RECT 79.995 37.380 80.055 37.460 ;
        POLYGON 79.995 37.380 80.055 37.380 80.055 37.320 ;
        RECT 80.210 37.370 80.285 37.510 ;
        RECT 81.975 37.370 82.050 37.510 ;
        RECT 82.190 37.320 82.265 37.460 ;
        RECT 82.895 37.380 82.955 37.460 ;
        POLYGON 82.895 37.380 82.955 37.380 82.955 37.320 ;
        RECT 83.110 37.370 83.185 37.510 ;
        RECT 84.875 37.370 84.950 37.510 ;
        RECT 85.090 37.320 85.165 37.460 ;
        RECT 85.795 37.380 85.855 37.460 ;
        POLYGON 85.795 37.380 85.855 37.380 85.855 37.320 ;
        RECT 86.010 37.370 86.085 37.510 ;
        RECT 87.775 37.370 87.850 37.510 ;
        RECT 87.990 37.320 88.065 37.460 ;
        RECT 88.695 37.380 88.755 37.460 ;
        POLYGON 88.695 37.380 88.755 37.380 88.755 37.320 ;
        RECT 88.910 37.370 88.985 37.510 ;
        RECT 90.675 37.370 90.750 37.510 ;
        RECT 90.890 37.320 90.965 37.460 ;
        RECT 91.595 37.380 91.655 37.460 ;
        POLYGON 91.595 37.380 91.655 37.380 91.655 37.320 ;
        RECT 91.810 37.370 91.885 37.510 ;
        RECT 0.720 36.850 0.870 37.020 ;
        RECT 1.110 36.985 1.260 37.155 ;
        RECT 1.500 36.985 1.650 37.155 ;
        RECT 1.890 36.850 2.040 37.020 ;
        RECT 3.620 36.850 3.770 37.020 ;
        RECT 4.010 36.985 4.160 37.155 ;
        RECT 4.400 36.985 4.550 37.155 ;
        RECT 4.790 36.850 4.940 37.020 ;
        RECT 6.520 36.850 6.670 37.020 ;
        RECT 6.910 36.985 7.060 37.155 ;
        RECT 7.300 36.985 7.450 37.155 ;
        RECT 7.690 36.850 7.840 37.020 ;
        RECT 9.420 36.850 9.570 37.020 ;
        RECT 9.810 36.985 9.960 37.155 ;
        RECT 10.200 36.985 10.350 37.155 ;
        RECT 10.590 36.850 10.740 37.020 ;
        RECT 12.320 36.850 12.470 37.020 ;
        RECT 12.710 36.985 12.860 37.155 ;
        RECT 13.100 36.985 13.250 37.155 ;
        RECT 13.490 36.850 13.640 37.020 ;
        RECT 15.220 36.850 15.370 37.020 ;
        RECT 15.610 36.985 15.760 37.155 ;
        RECT 16.000 36.985 16.150 37.155 ;
        RECT 16.390 36.850 16.540 37.020 ;
        RECT 18.120 36.850 18.270 37.020 ;
        RECT 18.510 36.985 18.660 37.155 ;
        RECT 18.900 36.985 19.050 37.155 ;
        RECT 19.290 36.850 19.440 37.020 ;
        RECT 21.020 36.850 21.170 37.020 ;
        RECT 21.410 36.985 21.560 37.155 ;
        RECT 21.800 36.985 21.950 37.155 ;
        RECT 22.190 36.850 22.340 37.020 ;
        RECT 23.920 36.850 24.070 37.020 ;
        RECT 24.310 36.985 24.460 37.155 ;
        RECT 24.700 36.985 24.850 37.155 ;
        RECT 25.090 36.850 25.240 37.020 ;
        RECT 26.820 36.850 26.970 37.020 ;
        RECT 27.210 36.985 27.360 37.155 ;
        RECT 27.600 36.985 27.750 37.155 ;
        RECT 27.990 36.850 28.140 37.020 ;
        RECT 29.720 36.850 29.870 37.020 ;
        RECT 30.110 36.985 30.260 37.155 ;
        RECT 30.500 36.985 30.650 37.155 ;
        RECT 30.890 36.850 31.040 37.020 ;
        RECT 32.620 36.850 32.770 37.020 ;
        RECT 33.010 36.985 33.160 37.155 ;
        RECT 33.400 36.985 33.550 37.155 ;
        RECT 33.790 36.850 33.940 37.020 ;
        RECT 35.520 36.850 35.670 37.020 ;
        RECT 35.910 36.985 36.060 37.155 ;
        RECT 36.300 36.985 36.450 37.155 ;
        RECT 36.690 36.850 36.840 37.020 ;
        RECT 38.420 36.850 38.570 37.020 ;
        RECT 38.810 36.985 38.960 37.155 ;
        RECT 39.200 36.985 39.350 37.155 ;
        RECT 39.590 36.850 39.740 37.020 ;
        RECT 41.320 36.850 41.470 37.020 ;
        RECT 41.710 36.985 41.860 37.155 ;
        RECT 42.100 36.985 42.250 37.155 ;
        RECT 42.490 36.850 42.640 37.020 ;
        RECT 44.220 36.850 44.370 37.020 ;
        RECT 44.610 36.985 44.760 37.155 ;
        RECT 45.000 36.985 45.150 37.155 ;
        RECT 45.390 36.850 45.540 37.020 ;
        RECT 47.120 36.850 47.270 37.020 ;
        RECT 47.510 36.985 47.660 37.155 ;
        RECT 47.900 36.985 48.050 37.155 ;
        RECT 48.290 36.850 48.440 37.020 ;
        RECT 50.020 36.850 50.170 37.020 ;
        RECT 50.410 36.985 50.560 37.155 ;
        RECT 50.800 36.985 50.950 37.155 ;
        RECT 51.190 36.850 51.340 37.020 ;
        RECT 52.920 36.850 53.070 37.020 ;
        RECT 53.310 36.985 53.460 37.155 ;
        RECT 53.700 36.985 53.850 37.155 ;
        RECT 54.090 36.850 54.240 37.020 ;
        RECT 55.820 36.850 55.970 37.020 ;
        RECT 56.210 36.985 56.360 37.155 ;
        RECT 56.600 36.985 56.750 37.155 ;
        RECT 56.990 36.850 57.140 37.020 ;
        RECT 58.720 36.850 58.870 37.020 ;
        RECT 59.110 36.985 59.260 37.155 ;
        RECT 59.500 36.985 59.650 37.155 ;
        RECT 59.890 36.850 60.040 37.020 ;
        RECT 61.620 36.850 61.770 37.020 ;
        RECT 62.010 36.985 62.160 37.155 ;
        RECT 62.400 36.985 62.550 37.155 ;
        RECT 62.790 36.850 62.940 37.020 ;
        RECT 64.520 36.850 64.670 37.020 ;
        RECT 64.910 36.985 65.060 37.155 ;
        RECT 65.300 36.985 65.450 37.155 ;
        RECT 65.690 36.850 65.840 37.020 ;
        RECT 67.420 36.850 67.570 37.020 ;
        RECT 67.810 36.985 67.960 37.155 ;
        RECT 68.200 36.985 68.350 37.155 ;
        RECT 68.590 36.850 68.740 37.020 ;
        RECT 70.320 36.850 70.470 37.020 ;
        RECT 70.710 36.985 70.860 37.155 ;
        RECT 71.100 36.985 71.250 37.155 ;
        RECT 71.490 36.850 71.640 37.020 ;
        RECT 73.220 36.850 73.370 37.020 ;
        RECT 73.610 36.985 73.760 37.155 ;
        RECT 74.000 36.985 74.150 37.155 ;
        RECT 74.390 36.850 74.540 37.020 ;
        RECT 76.120 36.850 76.270 37.020 ;
        RECT 76.510 36.985 76.660 37.155 ;
        RECT 76.900 36.985 77.050 37.155 ;
        RECT 77.290 36.850 77.440 37.020 ;
        RECT 79.020 36.850 79.170 37.020 ;
        RECT 79.410 36.985 79.560 37.155 ;
        RECT 79.800 36.985 79.950 37.155 ;
        RECT 80.190 36.850 80.340 37.020 ;
        RECT 81.920 36.850 82.070 37.020 ;
        RECT 82.310 36.985 82.460 37.155 ;
        RECT 82.700 36.985 82.850 37.155 ;
        RECT 83.090 36.850 83.240 37.020 ;
        RECT 84.820 36.850 84.970 37.020 ;
        RECT 85.210 36.985 85.360 37.155 ;
        RECT 85.600 36.985 85.750 37.155 ;
        RECT 85.990 36.850 86.140 37.020 ;
        RECT 87.720 36.850 87.870 37.020 ;
        RECT 88.110 36.985 88.260 37.155 ;
        RECT 88.500 36.985 88.650 37.155 ;
        RECT 88.890 36.850 89.040 37.020 ;
        RECT 90.620 36.850 90.770 37.020 ;
        RECT 91.010 36.985 91.160 37.155 ;
        RECT 91.400 36.985 91.550 37.155 ;
        RECT 91.790 36.850 91.940 37.020 ;
        RECT 0.985 36.765 1.035 36.800 ;
        POLYGON 1.035 36.800 1.070 36.765 1.035 36.765 ;
        RECT 0.985 36.640 1.070 36.765 ;
        RECT 1.690 36.640 1.775 36.800 ;
        RECT 3.885 36.765 3.935 36.800 ;
        POLYGON 3.935 36.800 3.970 36.765 3.935 36.765 ;
        RECT 3.885 36.640 3.970 36.765 ;
        RECT 4.590 36.640 4.675 36.800 ;
        RECT 6.785 36.765 6.835 36.800 ;
        POLYGON 6.835 36.800 6.870 36.765 6.835 36.765 ;
        RECT 6.785 36.640 6.870 36.765 ;
        RECT 7.490 36.640 7.575 36.800 ;
        RECT 9.685 36.765 9.735 36.800 ;
        POLYGON 9.735 36.800 9.770 36.765 9.735 36.765 ;
        RECT 9.685 36.640 9.770 36.765 ;
        RECT 10.390 36.640 10.475 36.800 ;
        RECT 12.585 36.765 12.635 36.800 ;
        POLYGON 12.635 36.800 12.670 36.765 12.635 36.765 ;
        RECT 12.585 36.640 12.670 36.765 ;
        RECT 13.290 36.640 13.375 36.800 ;
        RECT 15.485 36.765 15.535 36.800 ;
        POLYGON 15.535 36.800 15.570 36.765 15.535 36.765 ;
        RECT 15.485 36.640 15.570 36.765 ;
        RECT 16.190 36.640 16.275 36.800 ;
        RECT 18.385 36.765 18.435 36.800 ;
        POLYGON 18.435 36.800 18.470 36.765 18.435 36.765 ;
        RECT 18.385 36.640 18.470 36.765 ;
        RECT 19.090 36.640 19.175 36.800 ;
        RECT 21.285 36.765 21.335 36.800 ;
        POLYGON 21.335 36.800 21.370 36.765 21.335 36.765 ;
        RECT 21.285 36.640 21.370 36.765 ;
        RECT 21.990 36.640 22.075 36.800 ;
        RECT 24.185 36.765 24.235 36.800 ;
        POLYGON 24.235 36.800 24.270 36.765 24.235 36.765 ;
        RECT 24.185 36.640 24.270 36.765 ;
        RECT 24.890 36.640 24.975 36.800 ;
        RECT 27.085 36.765 27.135 36.800 ;
        POLYGON 27.135 36.800 27.170 36.765 27.135 36.765 ;
        RECT 27.085 36.640 27.170 36.765 ;
        RECT 27.790 36.640 27.875 36.800 ;
        RECT 29.985 36.765 30.035 36.800 ;
        POLYGON 30.035 36.800 30.070 36.765 30.035 36.765 ;
        RECT 29.985 36.640 30.070 36.765 ;
        RECT 30.690 36.640 30.775 36.800 ;
        RECT 32.885 36.765 32.935 36.800 ;
        POLYGON 32.935 36.800 32.970 36.765 32.935 36.765 ;
        RECT 32.885 36.640 32.970 36.765 ;
        RECT 33.590 36.640 33.675 36.800 ;
        RECT 35.785 36.765 35.835 36.800 ;
        POLYGON 35.835 36.800 35.870 36.765 35.835 36.765 ;
        RECT 35.785 36.640 35.870 36.765 ;
        RECT 36.490 36.640 36.575 36.800 ;
        RECT 38.685 36.765 38.735 36.800 ;
        POLYGON 38.735 36.800 38.770 36.765 38.735 36.765 ;
        RECT 38.685 36.640 38.770 36.765 ;
        RECT 39.390 36.640 39.475 36.800 ;
        RECT 41.585 36.765 41.635 36.800 ;
        POLYGON 41.635 36.800 41.670 36.765 41.635 36.765 ;
        RECT 41.585 36.640 41.670 36.765 ;
        RECT 42.290 36.640 42.375 36.800 ;
        RECT 44.485 36.765 44.535 36.800 ;
        POLYGON 44.535 36.800 44.570 36.765 44.535 36.765 ;
        RECT 44.485 36.640 44.570 36.765 ;
        RECT 45.190 36.640 45.275 36.800 ;
        RECT 47.385 36.765 47.435 36.800 ;
        POLYGON 47.435 36.800 47.470 36.765 47.435 36.765 ;
        RECT 47.385 36.640 47.470 36.765 ;
        RECT 48.090 36.640 48.175 36.800 ;
        RECT 50.285 36.765 50.335 36.800 ;
        POLYGON 50.335 36.800 50.370 36.765 50.335 36.765 ;
        RECT 50.285 36.640 50.370 36.765 ;
        RECT 50.990 36.640 51.075 36.800 ;
        RECT 53.185 36.765 53.235 36.800 ;
        POLYGON 53.235 36.800 53.270 36.765 53.235 36.765 ;
        RECT 53.185 36.640 53.270 36.765 ;
        RECT 53.890 36.640 53.975 36.800 ;
        RECT 56.085 36.765 56.135 36.800 ;
        POLYGON 56.135 36.800 56.170 36.765 56.135 36.765 ;
        RECT 56.085 36.640 56.170 36.765 ;
        RECT 56.790 36.640 56.875 36.800 ;
        RECT 58.985 36.765 59.035 36.800 ;
        POLYGON 59.035 36.800 59.070 36.765 59.035 36.765 ;
        RECT 58.985 36.640 59.070 36.765 ;
        RECT 59.690 36.640 59.775 36.800 ;
        RECT 61.885 36.765 61.935 36.800 ;
        POLYGON 61.935 36.800 61.970 36.765 61.935 36.765 ;
        RECT 61.885 36.640 61.970 36.765 ;
        RECT 62.590 36.640 62.675 36.800 ;
        RECT 64.785 36.765 64.835 36.800 ;
        POLYGON 64.835 36.800 64.870 36.765 64.835 36.765 ;
        RECT 64.785 36.640 64.870 36.765 ;
        RECT 65.490 36.640 65.575 36.800 ;
        RECT 67.685 36.765 67.735 36.800 ;
        POLYGON 67.735 36.800 67.770 36.765 67.735 36.765 ;
        RECT 67.685 36.640 67.770 36.765 ;
        RECT 68.390 36.640 68.475 36.800 ;
        RECT 70.585 36.765 70.635 36.800 ;
        POLYGON 70.635 36.800 70.670 36.765 70.635 36.765 ;
        RECT 70.585 36.640 70.670 36.765 ;
        RECT 71.290 36.640 71.375 36.800 ;
        RECT 73.485 36.765 73.535 36.800 ;
        POLYGON 73.535 36.800 73.570 36.765 73.535 36.765 ;
        RECT 73.485 36.640 73.570 36.765 ;
        RECT 74.190 36.640 74.275 36.800 ;
        RECT 76.385 36.765 76.435 36.800 ;
        POLYGON 76.435 36.800 76.470 36.765 76.435 36.765 ;
        RECT 76.385 36.640 76.470 36.765 ;
        RECT 77.090 36.640 77.175 36.800 ;
        RECT 79.285 36.765 79.335 36.800 ;
        POLYGON 79.335 36.800 79.370 36.765 79.335 36.765 ;
        RECT 79.285 36.640 79.370 36.765 ;
        RECT 79.990 36.640 80.075 36.800 ;
        RECT 82.185 36.765 82.235 36.800 ;
        POLYGON 82.235 36.800 82.270 36.765 82.235 36.765 ;
        RECT 82.185 36.640 82.270 36.765 ;
        RECT 82.890 36.640 82.975 36.800 ;
        RECT 85.085 36.765 85.135 36.800 ;
        POLYGON 85.135 36.800 85.170 36.765 85.135 36.765 ;
        RECT 85.085 36.640 85.170 36.765 ;
        RECT 85.790 36.640 85.875 36.800 ;
        RECT 87.985 36.765 88.035 36.800 ;
        POLYGON 88.035 36.800 88.070 36.765 88.035 36.765 ;
        RECT 87.985 36.640 88.070 36.765 ;
        RECT 88.690 36.640 88.775 36.800 ;
        RECT 90.885 36.765 90.935 36.800 ;
        POLYGON 90.935 36.800 90.970 36.765 90.935 36.765 ;
        RECT 90.885 36.640 90.970 36.765 ;
        RECT 91.590 36.640 91.675 36.800 ;
        RECT 0.775 36.020 0.850 36.160 ;
        RECT 0.990 35.970 1.065 36.110 ;
        RECT 1.695 36.030 1.755 36.110 ;
        POLYGON 1.695 36.030 1.755 36.030 1.755 35.970 ;
        RECT 1.910 36.020 1.985 36.160 ;
        RECT 3.675 36.020 3.750 36.160 ;
        RECT 3.890 35.970 3.965 36.110 ;
        RECT 4.595 36.030 4.655 36.110 ;
        POLYGON 4.595 36.030 4.655 36.030 4.655 35.970 ;
        RECT 4.810 36.020 4.885 36.160 ;
        RECT 6.575 36.020 6.650 36.160 ;
        RECT 6.790 35.970 6.865 36.110 ;
        RECT 7.495 36.030 7.555 36.110 ;
        POLYGON 7.495 36.030 7.555 36.030 7.555 35.970 ;
        RECT 7.710 36.020 7.785 36.160 ;
        RECT 9.475 36.020 9.550 36.160 ;
        RECT 9.690 35.970 9.765 36.110 ;
        RECT 10.395 36.030 10.455 36.110 ;
        POLYGON 10.395 36.030 10.455 36.030 10.455 35.970 ;
        RECT 10.610 36.020 10.685 36.160 ;
        RECT 12.375 36.020 12.450 36.160 ;
        RECT 12.590 35.970 12.665 36.110 ;
        RECT 13.295 36.030 13.355 36.110 ;
        POLYGON 13.295 36.030 13.355 36.030 13.355 35.970 ;
        RECT 13.510 36.020 13.585 36.160 ;
        RECT 15.275 36.020 15.350 36.160 ;
        RECT 15.490 35.970 15.565 36.110 ;
        RECT 16.195 36.030 16.255 36.110 ;
        POLYGON 16.195 36.030 16.255 36.030 16.255 35.970 ;
        RECT 16.410 36.020 16.485 36.160 ;
        RECT 18.175 36.020 18.250 36.160 ;
        RECT 18.390 35.970 18.465 36.110 ;
        RECT 19.095 36.030 19.155 36.110 ;
        POLYGON 19.095 36.030 19.155 36.030 19.155 35.970 ;
        RECT 19.310 36.020 19.385 36.160 ;
        RECT 21.075 36.020 21.150 36.160 ;
        RECT 21.290 35.970 21.365 36.110 ;
        RECT 21.995 36.030 22.055 36.110 ;
        POLYGON 21.995 36.030 22.055 36.030 22.055 35.970 ;
        RECT 22.210 36.020 22.285 36.160 ;
        RECT 23.975 36.020 24.050 36.160 ;
        RECT 24.190 35.970 24.265 36.110 ;
        RECT 24.895 36.030 24.955 36.110 ;
        POLYGON 24.895 36.030 24.955 36.030 24.955 35.970 ;
        RECT 25.110 36.020 25.185 36.160 ;
        RECT 26.875 36.020 26.950 36.160 ;
        RECT 27.090 35.970 27.165 36.110 ;
        RECT 27.795 36.030 27.855 36.110 ;
        POLYGON 27.795 36.030 27.855 36.030 27.855 35.970 ;
        RECT 28.010 36.020 28.085 36.160 ;
        RECT 29.775 36.020 29.850 36.160 ;
        RECT 29.990 35.970 30.065 36.110 ;
        RECT 30.695 36.030 30.755 36.110 ;
        POLYGON 30.695 36.030 30.755 36.030 30.755 35.970 ;
        RECT 30.910 36.020 30.985 36.160 ;
        RECT 32.675 36.020 32.750 36.160 ;
        RECT 32.890 35.970 32.965 36.110 ;
        RECT 33.595 36.030 33.655 36.110 ;
        POLYGON 33.595 36.030 33.655 36.030 33.655 35.970 ;
        RECT 33.810 36.020 33.885 36.160 ;
        RECT 35.575 36.020 35.650 36.160 ;
        RECT 35.790 35.970 35.865 36.110 ;
        RECT 36.495 36.030 36.555 36.110 ;
        POLYGON 36.495 36.030 36.555 36.030 36.555 35.970 ;
        RECT 36.710 36.020 36.785 36.160 ;
        RECT 38.475 36.020 38.550 36.160 ;
        RECT 38.690 35.970 38.765 36.110 ;
        RECT 39.395 36.030 39.455 36.110 ;
        POLYGON 39.395 36.030 39.455 36.030 39.455 35.970 ;
        RECT 39.610 36.020 39.685 36.160 ;
        RECT 41.375 36.020 41.450 36.160 ;
        RECT 41.590 35.970 41.665 36.110 ;
        RECT 42.295 36.030 42.355 36.110 ;
        POLYGON 42.295 36.030 42.355 36.030 42.355 35.970 ;
        RECT 42.510 36.020 42.585 36.160 ;
        RECT 44.275 36.020 44.350 36.160 ;
        RECT 44.490 35.970 44.565 36.110 ;
        RECT 45.195 36.030 45.255 36.110 ;
        POLYGON 45.195 36.030 45.255 36.030 45.255 35.970 ;
        RECT 45.410 36.020 45.485 36.160 ;
        RECT 47.175 36.020 47.250 36.160 ;
        RECT 47.390 35.970 47.465 36.110 ;
        RECT 48.095 36.030 48.155 36.110 ;
        POLYGON 48.095 36.030 48.155 36.030 48.155 35.970 ;
        RECT 48.310 36.020 48.385 36.160 ;
        RECT 50.075 36.020 50.150 36.160 ;
        RECT 50.290 35.970 50.365 36.110 ;
        RECT 50.995 36.030 51.055 36.110 ;
        POLYGON 50.995 36.030 51.055 36.030 51.055 35.970 ;
        RECT 51.210 36.020 51.285 36.160 ;
        RECT 52.975 36.020 53.050 36.160 ;
        RECT 53.190 35.970 53.265 36.110 ;
        RECT 53.895 36.030 53.955 36.110 ;
        POLYGON 53.895 36.030 53.955 36.030 53.955 35.970 ;
        RECT 54.110 36.020 54.185 36.160 ;
        RECT 55.875 36.020 55.950 36.160 ;
        RECT 56.090 35.970 56.165 36.110 ;
        RECT 56.795 36.030 56.855 36.110 ;
        POLYGON 56.795 36.030 56.855 36.030 56.855 35.970 ;
        RECT 57.010 36.020 57.085 36.160 ;
        RECT 58.775 36.020 58.850 36.160 ;
        RECT 58.990 35.970 59.065 36.110 ;
        RECT 59.695 36.030 59.755 36.110 ;
        POLYGON 59.695 36.030 59.755 36.030 59.755 35.970 ;
        RECT 59.910 36.020 59.985 36.160 ;
        RECT 61.675 36.020 61.750 36.160 ;
        RECT 61.890 35.970 61.965 36.110 ;
        RECT 62.595 36.030 62.655 36.110 ;
        POLYGON 62.595 36.030 62.655 36.030 62.655 35.970 ;
        RECT 62.810 36.020 62.885 36.160 ;
        RECT 64.575 36.020 64.650 36.160 ;
        RECT 64.790 35.970 64.865 36.110 ;
        RECT 65.495 36.030 65.555 36.110 ;
        POLYGON 65.495 36.030 65.555 36.030 65.555 35.970 ;
        RECT 65.710 36.020 65.785 36.160 ;
        RECT 67.475 36.020 67.550 36.160 ;
        RECT 67.690 35.970 67.765 36.110 ;
        RECT 68.395 36.030 68.455 36.110 ;
        POLYGON 68.395 36.030 68.455 36.030 68.455 35.970 ;
        RECT 68.610 36.020 68.685 36.160 ;
        RECT 70.375 36.020 70.450 36.160 ;
        RECT 70.590 35.970 70.665 36.110 ;
        RECT 71.295 36.030 71.355 36.110 ;
        POLYGON 71.295 36.030 71.355 36.030 71.355 35.970 ;
        RECT 71.510 36.020 71.585 36.160 ;
        RECT 73.275 36.020 73.350 36.160 ;
        RECT 73.490 35.970 73.565 36.110 ;
        RECT 74.195 36.030 74.255 36.110 ;
        POLYGON 74.195 36.030 74.255 36.030 74.255 35.970 ;
        RECT 74.410 36.020 74.485 36.160 ;
        RECT 76.175 36.020 76.250 36.160 ;
        RECT 76.390 35.970 76.465 36.110 ;
        RECT 77.095 36.030 77.155 36.110 ;
        POLYGON 77.095 36.030 77.155 36.030 77.155 35.970 ;
        RECT 77.310 36.020 77.385 36.160 ;
        RECT 79.075 36.020 79.150 36.160 ;
        RECT 79.290 35.970 79.365 36.110 ;
        RECT 79.995 36.030 80.055 36.110 ;
        POLYGON 79.995 36.030 80.055 36.030 80.055 35.970 ;
        RECT 80.210 36.020 80.285 36.160 ;
        RECT 81.975 36.020 82.050 36.160 ;
        RECT 82.190 35.970 82.265 36.110 ;
        RECT 82.895 36.030 82.955 36.110 ;
        POLYGON 82.895 36.030 82.955 36.030 82.955 35.970 ;
        RECT 83.110 36.020 83.185 36.160 ;
        RECT 84.875 36.020 84.950 36.160 ;
        RECT 85.090 35.970 85.165 36.110 ;
        RECT 85.795 36.030 85.855 36.110 ;
        POLYGON 85.795 36.030 85.855 36.030 85.855 35.970 ;
        RECT 86.010 36.020 86.085 36.160 ;
        RECT 87.775 36.020 87.850 36.160 ;
        RECT 87.990 35.970 88.065 36.110 ;
        RECT 88.695 36.030 88.755 36.110 ;
        POLYGON 88.695 36.030 88.755 36.030 88.755 35.970 ;
        RECT 88.910 36.020 88.985 36.160 ;
        RECT 90.675 36.020 90.750 36.160 ;
        RECT 90.890 35.970 90.965 36.110 ;
        RECT 91.595 36.030 91.655 36.110 ;
        POLYGON 91.595 36.030 91.655 36.030 91.655 35.970 ;
        RECT 91.810 36.020 91.885 36.160 ;
        RECT 0.720 35.500 0.870 35.670 ;
        RECT 1.110 35.635 1.260 35.805 ;
        RECT 1.500 35.635 1.650 35.805 ;
        RECT 1.890 35.500 2.040 35.670 ;
        RECT 3.620 35.500 3.770 35.670 ;
        RECT 4.010 35.635 4.160 35.805 ;
        RECT 4.400 35.635 4.550 35.805 ;
        RECT 4.790 35.500 4.940 35.670 ;
        RECT 6.520 35.500 6.670 35.670 ;
        RECT 6.910 35.635 7.060 35.805 ;
        RECT 7.300 35.635 7.450 35.805 ;
        RECT 7.690 35.500 7.840 35.670 ;
        RECT 9.420 35.500 9.570 35.670 ;
        RECT 9.810 35.635 9.960 35.805 ;
        RECT 10.200 35.635 10.350 35.805 ;
        RECT 10.590 35.500 10.740 35.670 ;
        RECT 12.320 35.500 12.470 35.670 ;
        RECT 12.710 35.635 12.860 35.805 ;
        RECT 13.100 35.635 13.250 35.805 ;
        RECT 13.490 35.500 13.640 35.670 ;
        RECT 15.220 35.500 15.370 35.670 ;
        RECT 15.610 35.635 15.760 35.805 ;
        RECT 16.000 35.635 16.150 35.805 ;
        RECT 16.390 35.500 16.540 35.670 ;
        RECT 18.120 35.500 18.270 35.670 ;
        RECT 18.510 35.635 18.660 35.805 ;
        RECT 18.900 35.635 19.050 35.805 ;
        RECT 19.290 35.500 19.440 35.670 ;
        RECT 21.020 35.500 21.170 35.670 ;
        RECT 21.410 35.635 21.560 35.805 ;
        RECT 21.800 35.635 21.950 35.805 ;
        RECT 22.190 35.500 22.340 35.670 ;
        RECT 23.920 35.500 24.070 35.670 ;
        RECT 24.310 35.635 24.460 35.805 ;
        RECT 24.700 35.635 24.850 35.805 ;
        RECT 25.090 35.500 25.240 35.670 ;
        RECT 26.820 35.500 26.970 35.670 ;
        RECT 27.210 35.635 27.360 35.805 ;
        RECT 27.600 35.635 27.750 35.805 ;
        RECT 27.990 35.500 28.140 35.670 ;
        RECT 29.720 35.500 29.870 35.670 ;
        RECT 30.110 35.635 30.260 35.805 ;
        RECT 30.500 35.635 30.650 35.805 ;
        RECT 30.890 35.500 31.040 35.670 ;
        RECT 32.620 35.500 32.770 35.670 ;
        RECT 33.010 35.635 33.160 35.805 ;
        RECT 33.400 35.635 33.550 35.805 ;
        RECT 33.790 35.500 33.940 35.670 ;
        RECT 35.520 35.500 35.670 35.670 ;
        RECT 35.910 35.635 36.060 35.805 ;
        RECT 36.300 35.635 36.450 35.805 ;
        RECT 36.690 35.500 36.840 35.670 ;
        RECT 38.420 35.500 38.570 35.670 ;
        RECT 38.810 35.635 38.960 35.805 ;
        RECT 39.200 35.635 39.350 35.805 ;
        RECT 39.590 35.500 39.740 35.670 ;
        RECT 41.320 35.500 41.470 35.670 ;
        RECT 41.710 35.635 41.860 35.805 ;
        RECT 42.100 35.635 42.250 35.805 ;
        RECT 42.490 35.500 42.640 35.670 ;
        RECT 44.220 35.500 44.370 35.670 ;
        RECT 44.610 35.635 44.760 35.805 ;
        RECT 45.000 35.635 45.150 35.805 ;
        RECT 45.390 35.500 45.540 35.670 ;
        RECT 47.120 35.500 47.270 35.670 ;
        RECT 47.510 35.635 47.660 35.805 ;
        RECT 47.900 35.635 48.050 35.805 ;
        RECT 48.290 35.500 48.440 35.670 ;
        RECT 50.020 35.500 50.170 35.670 ;
        RECT 50.410 35.635 50.560 35.805 ;
        RECT 50.800 35.635 50.950 35.805 ;
        RECT 51.190 35.500 51.340 35.670 ;
        RECT 52.920 35.500 53.070 35.670 ;
        RECT 53.310 35.635 53.460 35.805 ;
        RECT 53.700 35.635 53.850 35.805 ;
        RECT 54.090 35.500 54.240 35.670 ;
        RECT 55.820 35.500 55.970 35.670 ;
        RECT 56.210 35.635 56.360 35.805 ;
        RECT 56.600 35.635 56.750 35.805 ;
        RECT 56.990 35.500 57.140 35.670 ;
        RECT 58.720 35.500 58.870 35.670 ;
        RECT 59.110 35.635 59.260 35.805 ;
        RECT 59.500 35.635 59.650 35.805 ;
        RECT 59.890 35.500 60.040 35.670 ;
        RECT 61.620 35.500 61.770 35.670 ;
        RECT 62.010 35.635 62.160 35.805 ;
        RECT 62.400 35.635 62.550 35.805 ;
        RECT 62.790 35.500 62.940 35.670 ;
        RECT 64.520 35.500 64.670 35.670 ;
        RECT 64.910 35.635 65.060 35.805 ;
        RECT 65.300 35.635 65.450 35.805 ;
        RECT 65.690 35.500 65.840 35.670 ;
        RECT 67.420 35.500 67.570 35.670 ;
        RECT 67.810 35.635 67.960 35.805 ;
        RECT 68.200 35.635 68.350 35.805 ;
        RECT 68.590 35.500 68.740 35.670 ;
        RECT 70.320 35.500 70.470 35.670 ;
        RECT 70.710 35.635 70.860 35.805 ;
        RECT 71.100 35.635 71.250 35.805 ;
        RECT 71.490 35.500 71.640 35.670 ;
        RECT 73.220 35.500 73.370 35.670 ;
        RECT 73.610 35.635 73.760 35.805 ;
        RECT 74.000 35.635 74.150 35.805 ;
        RECT 74.390 35.500 74.540 35.670 ;
        RECT 76.120 35.500 76.270 35.670 ;
        RECT 76.510 35.635 76.660 35.805 ;
        RECT 76.900 35.635 77.050 35.805 ;
        RECT 77.290 35.500 77.440 35.670 ;
        RECT 79.020 35.500 79.170 35.670 ;
        RECT 79.410 35.635 79.560 35.805 ;
        RECT 79.800 35.635 79.950 35.805 ;
        RECT 80.190 35.500 80.340 35.670 ;
        RECT 81.920 35.500 82.070 35.670 ;
        RECT 82.310 35.635 82.460 35.805 ;
        RECT 82.700 35.635 82.850 35.805 ;
        RECT 83.090 35.500 83.240 35.670 ;
        RECT 84.820 35.500 84.970 35.670 ;
        RECT 85.210 35.635 85.360 35.805 ;
        RECT 85.600 35.635 85.750 35.805 ;
        RECT 85.990 35.500 86.140 35.670 ;
        RECT 87.720 35.500 87.870 35.670 ;
        RECT 88.110 35.635 88.260 35.805 ;
        RECT 88.500 35.635 88.650 35.805 ;
        RECT 88.890 35.500 89.040 35.670 ;
        RECT 90.620 35.500 90.770 35.670 ;
        RECT 91.010 35.635 91.160 35.805 ;
        RECT 91.400 35.635 91.550 35.805 ;
        RECT 91.790 35.500 91.940 35.670 ;
        RECT 0.985 35.415 1.035 35.450 ;
        POLYGON 1.035 35.450 1.070 35.415 1.035 35.415 ;
        RECT 0.985 35.290 1.070 35.415 ;
        RECT 1.690 35.290 1.775 35.450 ;
        RECT 3.885 35.415 3.935 35.450 ;
        POLYGON 3.935 35.450 3.970 35.415 3.935 35.415 ;
        RECT 3.885 35.290 3.970 35.415 ;
        RECT 4.590 35.290 4.675 35.450 ;
        RECT 6.785 35.415 6.835 35.450 ;
        POLYGON 6.835 35.450 6.870 35.415 6.835 35.415 ;
        RECT 6.785 35.290 6.870 35.415 ;
        RECT 7.490 35.290 7.575 35.450 ;
        RECT 9.685 35.415 9.735 35.450 ;
        POLYGON 9.735 35.450 9.770 35.415 9.735 35.415 ;
        RECT 9.685 35.290 9.770 35.415 ;
        RECT 10.390 35.290 10.475 35.450 ;
        RECT 12.585 35.415 12.635 35.450 ;
        POLYGON 12.635 35.450 12.670 35.415 12.635 35.415 ;
        RECT 12.585 35.290 12.670 35.415 ;
        RECT 13.290 35.290 13.375 35.450 ;
        RECT 15.485 35.415 15.535 35.450 ;
        POLYGON 15.535 35.450 15.570 35.415 15.535 35.415 ;
        RECT 15.485 35.290 15.570 35.415 ;
        RECT 16.190 35.290 16.275 35.450 ;
        RECT 18.385 35.415 18.435 35.450 ;
        POLYGON 18.435 35.450 18.470 35.415 18.435 35.415 ;
        RECT 18.385 35.290 18.470 35.415 ;
        RECT 19.090 35.290 19.175 35.450 ;
        RECT 21.285 35.415 21.335 35.450 ;
        POLYGON 21.335 35.450 21.370 35.415 21.335 35.415 ;
        RECT 21.285 35.290 21.370 35.415 ;
        RECT 21.990 35.290 22.075 35.450 ;
        RECT 24.185 35.415 24.235 35.450 ;
        POLYGON 24.235 35.450 24.270 35.415 24.235 35.415 ;
        RECT 24.185 35.290 24.270 35.415 ;
        RECT 24.890 35.290 24.975 35.450 ;
        RECT 27.085 35.415 27.135 35.450 ;
        POLYGON 27.135 35.450 27.170 35.415 27.135 35.415 ;
        RECT 27.085 35.290 27.170 35.415 ;
        RECT 27.790 35.290 27.875 35.450 ;
        RECT 29.985 35.415 30.035 35.450 ;
        POLYGON 30.035 35.450 30.070 35.415 30.035 35.415 ;
        RECT 29.985 35.290 30.070 35.415 ;
        RECT 30.690 35.290 30.775 35.450 ;
        RECT 32.885 35.415 32.935 35.450 ;
        POLYGON 32.935 35.450 32.970 35.415 32.935 35.415 ;
        RECT 32.885 35.290 32.970 35.415 ;
        RECT 33.590 35.290 33.675 35.450 ;
        RECT 35.785 35.415 35.835 35.450 ;
        POLYGON 35.835 35.450 35.870 35.415 35.835 35.415 ;
        RECT 35.785 35.290 35.870 35.415 ;
        RECT 36.490 35.290 36.575 35.450 ;
        RECT 38.685 35.415 38.735 35.450 ;
        POLYGON 38.735 35.450 38.770 35.415 38.735 35.415 ;
        RECT 38.685 35.290 38.770 35.415 ;
        RECT 39.390 35.290 39.475 35.450 ;
        RECT 41.585 35.415 41.635 35.450 ;
        POLYGON 41.635 35.450 41.670 35.415 41.635 35.415 ;
        RECT 41.585 35.290 41.670 35.415 ;
        RECT 42.290 35.290 42.375 35.450 ;
        RECT 44.485 35.415 44.535 35.450 ;
        POLYGON 44.535 35.450 44.570 35.415 44.535 35.415 ;
        RECT 44.485 35.290 44.570 35.415 ;
        RECT 45.190 35.290 45.275 35.450 ;
        RECT 47.385 35.415 47.435 35.450 ;
        POLYGON 47.435 35.450 47.470 35.415 47.435 35.415 ;
        RECT 47.385 35.290 47.470 35.415 ;
        RECT 48.090 35.290 48.175 35.450 ;
        RECT 50.285 35.415 50.335 35.450 ;
        POLYGON 50.335 35.450 50.370 35.415 50.335 35.415 ;
        RECT 50.285 35.290 50.370 35.415 ;
        RECT 50.990 35.290 51.075 35.450 ;
        RECT 53.185 35.415 53.235 35.450 ;
        POLYGON 53.235 35.450 53.270 35.415 53.235 35.415 ;
        RECT 53.185 35.290 53.270 35.415 ;
        RECT 53.890 35.290 53.975 35.450 ;
        RECT 56.085 35.415 56.135 35.450 ;
        POLYGON 56.135 35.450 56.170 35.415 56.135 35.415 ;
        RECT 56.085 35.290 56.170 35.415 ;
        RECT 56.790 35.290 56.875 35.450 ;
        RECT 58.985 35.415 59.035 35.450 ;
        POLYGON 59.035 35.450 59.070 35.415 59.035 35.415 ;
        RECT 58.985 35.290 59.070 35.415 ;
        RECT 59.690 35.290 59.775 35.450 ;
        RECT 61.885 35.415 61.935 35.450 ;
        POLYGON 61.935 35.450 61.970 35.415 61.935 35.415 ;
        RECT 61.885 35.290 61.970 35.415 ;
        RECT 62.590 35.290 62.675 35.450 ;
        RECT 64.785 35.415 64.835 35.450 ;
        POLYGON 64.835 35.450 64.870 35.415 64.835 35.415 ;
        RECT 64.785 35.290 64.870 35.415 ;
        RECT 65.490 35.290 65.575 35.450 ;
        RECT 67.685 35.415 67.735 35.450 ;
        POLYGON 67.735 35.450 67.770 35.415 67.735 35.415 ;
        RECT 67.685 35.290 67.770 35.415 ;
        RECT 68.390 35.290 68.475 35.450 ;
        RECT 70.585 35.415 70.635 35.450 ;
        POLYGON 70.635 35.450 70.670 35.415 70.635 35.415 ;
        RECT 70.585 35.290 70.670 35.415 ;
        RECT 71.290 35.290 71.375 35.450 ;
        RECT 73.485 35.415 73.535 35.450 ;
        POLYGON 73.535 35.450 73.570 35.415 73.535 35.415 ;
        RECT 73.485 35.290 73.570 35.415 ;
        RECT 74.190 35.290 74.275 35.450 ;
        RECT 76.385 35.415 76.435 35.450 ;
        POLYGON 76.435 35.450 76.470 35.415 76.435 35.415 ;
        RECT 76.385 35.290 76.470 35.415 ;
        RECT 77.090 35.290 77.175 35.450 ;
        RECT 79.285 35.415 79.335 35.450 ;
        POLYGON 79.335 35.450 79.370 35.415 79.335 35.415 ;
        RECT 79.285 35.290 79.370 35.415 ;
        RECT 79.990 35.290 80.075 35.450 ;
        RECT 82.185 35.415 82.235 35.450 ;
        POLYGON 82.235 35.450 82.270 35.415 82.235 35.415 ;
        RECT 82.185 35.290 82.270 35.415 ;
        RECT 82.890 35.290 82.975 35.450 ;
        RECT 85.085 35.415 85.135 35.450 ;
        POLYGON 85.135 35.450 85.170 35.415 85.135 35.415 ;
        RECT 85.085 35.290 85.170 35.415 ;
        RECT 85.790 35.290 85.875 35.450 ;
        RECT 87.985 35.415 88.035 35.450 ;
        POLYGON 88.035 35.450 88.070 35.415 88.035 35.415 ;
        RECT 87.985 35.290 88.070 35.415 ;
        RECT 88.690 35.290 88.775 35.450 ;
        RECT 90.885 35.415 90.935 35.450 ;
        POLYGON 90.935 35.450 90.970 35.415 90.935 35.415 ;
        RECT 90.885 35.290 90.970 35.415 ;
        RECT 91.590 35.290 91.675 35.450 ;
        RECT 0.775 34.670 0.850 34.810 ;
        RECT 0.990 34.620 1.065 34.760 ;
        RECT 1.695 34.680 1.755 34.760 ;
        POLYGON 1.695 34.680 1.755 34.680 1.755 34.620 ;
        RECT 1.910 34.670 1.985 34.810 ;
        RECT 3.675 34.670 3.750 34.810 ;
        RECT 3.890 34.620 3.965 34.760 ;
        RECT 4.595 34.680 4.655 34.760 ;
        POLYGON 4.595 34.680 4.655 34.680 4.655 34.620 ;
        RECT 4.810 34.670 4.885 34.810 ;
        RECT 6.575 34.670 6.650 34.810 ;
        RECT 6.790 34.620 6.865 34.760 ;
        RECT 7.495 34.680 7.555 34.760 ;
        POLYGON 7.495 34.680 7.555 34.680 7.555 34.620 ;
        RECT 7.710 34.670 7.785 34.810 ;
        RECT 9.475 34.670 9.550 34.810 ;
        RECT 9.690 34.620 9.765 34.760 ;
        RECT 10.395 34.680 10.455 34.760 ;
        POLYGON 10.395 34.680 10.455 34.680 10.455 34.620 ;
        RECT 10.610 34.670 10.685 34.810 ;
        RECT 12.375 34.670 12.450 34.810 ;
        RECT 12.590 34.620 12.665 34.760 ;
        RECT 13.295 34.680 13.355 34.760 ;
        POLYGON 13.295 34.680 13.355 34.680 13.355 34.620 ;
        RECT 13.510 34.670 13.585 34.810 ;
        RECT 15.275 34.670 15.350 34.810 ;
        RECT 15.490 34.620 15.565 34.760 ;
        RECT 16.195 34.680 16.255 34.760 ;
        POLYGON 16.195 34.680 16.255 34.680 16.255 34.620 ;
        RECT 16.410 34.670 16.485 34.810 ;
        RECT 18.175 34.670 18.250 34.810 ;
        RECT 18.390 34.620 18.465 34.760 ;
        RECT 19.095 34.680 19.155 34.760 ;
        POLYGON 19.095 34.680 19.155 34.680 19.155 34.620 ;
        RECT 19.310 34.670 19.385 34.810 ;
        RECT 21.075 34.670 21.150 34.810 ;
        RECT 21.290 34.620 21.365 34.760 ;
        RECT 21.995 34.680 22.055 34.760 ;
        POLYGON 21.995 34.680 22.055 34.680 22.055 34.620 ;
        RECT 22.210 34.670 22.285 34.810 ;
        RECT 23.975 34.670 24.050 34.810 ;
        RECT 24.190 34.620 24.265 34.760 ;
        RECT 24.895 34.680 24.955 34.760 ;
        POLYGON 24.895 34.680 24.955 34.680 24.955 34.620 ;
        RECT 25.110 34.670 25.185 34.810 ;
        RECT 26.875 34.670 26.950 34.810 ;
        RECT 27.090 34.620 27.165 34.760 ;
        RECT 27.795 34.680 27.855 34.760 ;
        POLYGON 27.795 34.680 27.855 34.680 27.855 34.620 ;
        RECT 28.010 34.670 28.085 34.810 ;
        RECT 29.775 34.670 29.850 34.810 ;
        RECT 29.990 34.620 30.065 34.760 ;
        RECT 30.695 34.680 30.755 34.760 ;
        POLYGON 30.695 34.680 30.755 34.680 30.755 34.620 ;
        RECT 30.910 34.670 30.985 34.810 ;
        RECT 32.675 34.670 32.750 34.810 ;
        RECT 32.890 34.620 32.965 34.760 ;
        RECT 33.595 34.680 33.655 34.760 ;
        POLYGON 33.595 34.680 33.655 34.680 33.655 34.620 ;
        RECT 33.810 34.670 33.885 34.810 ;
        RECT 35.575 34.670 35.650 34.810 ;
        RECT 35.790 34.620 35.865 34.760 ;
        RECT 36.495 34.680 36.555 34.760 ;
        POLYGON 36.495 34.680 36.555 34.680 36.555 34.620 ;
        RECT 36.710 34.670 36.785 34.810 ;
        RECT 38.475 34.670 38.550 34.810 ;
        RECT 38.690 34.620 38.765 34.760 ;
        RECT 39.395 34.680 39.455 34.760 ;
        POLYGON 39.395 34.680 39.455 34.680 39.455 34.620 ;
        RECT 39.610 34.670 39.685 34.810 ;
        RECT 41.375 34.670 41.450 34.810 ;
        RECT 41.590 34.620 41.665 34.760 ;
        RECT 42.295 34.680 42.355 34.760 ;
        POLYGON 42.295 34.680 42.355 34.680 42.355 34.620 ;
        RECT 42.510 34.670 42.585 34.810 ;
        RECT 44.275 34.670 44.350 34.810 ;
        RECT 44.490 34.620 44.565 34.760 ;
        RECT 45.195 34.680 45.255 34.760 ;
        POLYGON 45.195 34.680 45.255 34.680 45.255 34.620 ;
        RECT 45.410 34.670 45.485 34.810 ;
        RECT 47.175 34.670 47.250 34.810 ;
        RECT 47.390 34.620 47.465 34.760 ;
        RECT 48.095 34.680 48.155 34.760 ;
        POLYGON 48.095 34.680 48.155 34.680 48.155 34.620 ;
        RECT 48.310 34.670 48.385 34.810 ;
        RECT 50.075 34.670 50.150 34.810 ;
        RECT 50.290 34.620 50.365 34.760 ;
        RECT 50.995 34.680 51.055 34.760 ;
        POLYGON 50.995 34.680 51.055 34.680 51.055 34.620 ;
        RECT 51.210 34.670 51.285 34.810 ;
        RECT 52.975 34.670 53.050 34.810 ;
        RECT 53.190 34.620 53.265 34.760 ;
        RECT 53.895 34.680 53.955 34.760 ;
        POLYGON 53.895 34.680 53.955 34.680 53.955 34.620 ;
        RECT 54.110 34.670 54.185 34.810 ;
        RECT 55.875 34.670 55.950 34.810 ;
        RECT 56.090 34.620 56.165 34.760 ;
        RECT 56.795 34.680 56.855 34.760 ;
        POLYGON 56.795 34.680 56.855 34.680 56.855 34.620 ;
        RECT 57.010 34.670 57.085 34.810 ;
        RECT 58.775 34.670 58.850 34.810 ;
        RECT 58.990 34.620 59.065 34.760 ;
        RECT 59.695 34.680 59.755 34.760 ;
        POLYGON 59.695 34.680 59.755 34.680 59.755 34.620 ;
        RECT 59.910 34.670 59.985 34.810 ;
        RECT 61.675 34.670 61.750 34.810 ;
        RECT 61.890 34.620 61.965 34.760 ;
        RECT 62.595 34.680 62.655 34.760 ;
        POLYGON 62.595 34.680 62.655 34.680 62.655 34.620 ;
        RECT 62.810 34.670 62.885 34.810 ;
        RECT 64.575 34.670 64.650 34.810 ;
        RECT 64.790 34.620 64.865 34.760 ;
        RECT 65.495 34.680 65.555 34.760 ;
        POLYGON 65.495 34.680 65.555 34.680 65.555 34.620 ;
        RECT 65.710 34.670 65.785 34.810 ;
        RECT 67.475 34.670 67.550 34.810 ;
        RECT 67.690 34.620 67.765 34.760 ;
        RECT 68.395 34.680 68.455 34.760 ;
        POLYGON 68.395 34.680 68.455 34.680 68.455 34.620 ;
        RECT 68.610 34.670 68.685 34.810 ;
        RECT 70.375 34.670 70.450 34.810 ;
        RECT 70.590 34.620 70.665 34.760 ;
        RECT 71.295 34.680 71.355 34.760 ;
        POLYGON 71.295 34.680 71.355 34.680 71.355 34.620 ;
        RECT 71.510 34.670 71.585 34.810 ;
        RECT 73.275 34.670 73.350 34.810 ;
        RECT 73.490 34.620 73.565 34.760 ;
        RECT 74.195 34.680 74.255 34.760 ;
        POLYGON 74.195 34.680 74.255 34.680 74.255 34.620 ;
        RECT 74.410 34.670 74.485 34.810 ;
        RECT 76.175 34.670 76.250 34.810 ;
        RECT 76.390 34.620 76.465 34.760 ;
        RECT 77.095 34.680 77.155 34.760 ;
        POLYGON 77.095 34.680 77.155 34.680 77.155 34.620 ;
        RECT 77.310 34.670 77.385 34.810 ;
        RECT 79.075 34.670 79.150 34.810 ;
        RECT 79.290 34.620 79.365 34.760 ;
        RECT 79.995 34.680 80.055 34.760 ;
        POLYGON 79.995 34.680 80.055 34.680 80.055 34.620 ;
        RECT 80.210 34.670 80.285 34.810 ;
        RECT 81.975 34.670 82.050 34.810 ;
        RECT 82.190 34.620 82.265 34.760 ;
        RECT 82.895 34.680 82.955 34.760 ;
        POLYGON 82.895 34.680 82.955 34.680 82.955 34.620 ;
        RECT 83.110 34.670 83.185 34.810 ;
        RECT 84.875 34.670 84.950 34.810 ;
        RECT 85.090 34.620 85.165 34.760 ;
        RECT 85.795 34.680 85.855 34.760 ;
        POLYGON 85.795 34.680 85.855 34.680 85.855 34.620 ;
        RECT 86.010 34.670 86.085 34.810 ;
        RECT 87.775 34.670 87.850 34.810 ;
        RECT 87.990 34.620 88.065 34.760 ;
        RECT 88.695 34.680 88.755 34.760 ;
        POLYGON 88.695 34.680 88.755 34.680 88.755 34.620 ;
        RECT 88.910 34.670 88.985 34.810 ;
        RECT 90.675 34.670 90.750 34.810 ;
        RECT 90.890 34.620 90.965 34.760 ;
        RECT 91.595 34.680 91.655 34.760 ;
        POLYGON 91.595 34.680 91.655 34.680 91.655 34.620 ;
        RECT 91.810 34.670 91.885 34.810 ;
        RECT 0.720 34.150 0.870 34.320 ;
        RECT 1.110 34.285 1.260 34.455 ;
        RECT 1.500 34.285 1.650 34.455 ;
        RECT 1.890 34.150 2.040 34.320 ;
        RECT 3.620 34.150 3.770 34.320 ;
        RECT 4.010 34.285 4.160 34.455 ;
        RECT 4.400 34.285 4.550 34.455 ;
        RECT 4.790 34.150 4.940 34.320 ;
        RECT 6.520 34.150 6.670 34.320 ;
        RECT 6.910 34.285 7.060 34.455 ;
        RECT 7.300 34.285 7.450 34.455 ;
        RECT 7.690 34.150 7.840 34.320 ;
        RECT 9.420 34.150 9.570 34.320 ;
        RECT 9.810 34.285 9.960 34.455 ;
        RECT 10.200 34.285 10.350 34.455 ;
        RECT 10.590 34.150 10.740 34.320 ;
        RECT 12.320 34.150 12.470 34.320 ;
        RECT 12.710 34.285 12.860 34.455 ;
        RECT 13.100 34.285 13.250 34.455 ;
        RECT 13.490 34.150 13.640 34.320 ;
        RECT 15.220 34.150 15.370 34.320 ;
        RECT 15.610 34.285 15.760 34.455 ;
        RECT 16.000 34.285 16.150 34.455 ;
        RECT 16.390 34.150 16.540 34.320 ;
        RECT 18.120 34.150 18.270 34.320 ;
        RECT 18.510 34.285 18.660 34.455 ;
        RECT 18.900 34.285 19.050 34.455 ;
        RECT 19.290 34.150 19.440 34.320 ;
        RECT 21.020 34.150 21.170 34.320 ;
        RECT 21.410 34.285 21.560 34.455 ;
        RECT 21.800 34.285 21.950 34.455 ;
        RECT 22.190 34.150 22.340 34.320 ;
        RECT 23.920 34.150 24.070 34.320 ;
        RECT 24.310 34.285 24.460 34.455 ;
        RECT 24.700 34.285 24.850 34.455 ;
        RECT 25.090 34.150 25.240 34.320 ;
        RECT 26.820 34.150 26.970 34.320 ;
        RECT 27.210 34.285 27.360 34.455 ;
        RECT 27.600 34.285 27.750 34.455 ;
        RECT 27.990 34.150 28.140 34.320 ;
        RECT 29.720 34.150 29.870 34.320 ;
        RECT 30.110 34.285 30.260 34.455 ;
        RECT 30.500 34.285 30.650 34.455 ;
        RECT 30.890 34.150 31.040 34.320 ;
        RECT 32.620 34.150 32.770 34.320 ;
        RECT 33.010 34.285 33.160 34.455 ;
        RECT 33.400 34.285 33.550 34.455 ;
        RECT 33.790 34.150 33.940 34.320 ;
        RECT 35.520 34.150 35.670 34.320 ;
        RECT 35.910 34.285 36.060 34.455 ;
        RECT 36.300 34.285 36.450 34.455 ;
        RECT 36.690 34.150 36.840 34.320 ;
        RECT 38.420 34.150 38.570 34.320 ;
        RECT 38.810 34.285 38.960 34.455 ;
        RECT 39.200 34.285 39.350 34.455 ;
        RECT 39.590 34.150 39.740 34.320 ;
        RECT 41.320 34.150 41.470 34.320 ;
        RECT 41.710 34.285 41.860 34.455 ;
        RECT 42.100 34.285 42.250 34.455 ;
        RECT 42.490 34.150 42.640 34.320 ;
        RECT 44.220 34.150 44.370 34.320 ;
        RECT 44.610 34.285 44.760 34.455 ;
        RECT 45.000 34.285 45.150 34.455 ;
        RECT 45.390 34.150 45.540 34.320 ;
        RECT 47.120 34.150 47.270 34.320 ;
        RECT 47.510 34.285 47.660 34.455 ;
        RECT 47.900 34.285 48.050 34.455 ;
        RECT 48.290 34.150 48.440 34.320 ;
        RECT 50.020 34.150 50.170 34.320 ;
        RECT 50.410 34.285 50.560 34.455 ;
        RECT 50.800 34.285 50.950 34.455 ;
        RECT 51.190 34.150 51.340 34.320 ;
        RECT 52.920 34.150 53.070 34.320 ;
        RECT 53.310 34.285 53.460 34.455 ;
        RECT 53.700 34.285 53.850 34.455 ;
        RECT 54.090 34.150 54.240 34.320 ;
        RECT 55.820 34.150 55.970 34.320 ;
        RECT 56.210 34.285 56.360 34.455 ;
        RECT 56.600 34.285 56.750 34.455 ;
        RECT 56.990 34.150 57.140 34.320 ;
        RECT 58.720 34.150 58.870 34.320 ;
        RECT 59.110 34.285 59.260 34.455 ;
        RECT 59.500 34.285 59.650 34.455 ;
        RECT 59.890 34.150 60.040 34.320 ;
        RECT 61.620 34.150 61.770 34.320 ;
        RECT 62.010 34.285 62.160 34.455 ;
        RECT 62.400 34.285 62.550 34.455 ;
        RECT 62.790 34.150 62.940 34.320 ;
        RECT 64.520 34.150 64.670 34.320 ;
        RECT 64.910 34.285 65.060 34.455 ;
        RECT 65.300 34.285 65.450 34.455 ;
        RECT 65.690 34.150 65.840 34.320 ;
        RECT 67.420 34.150 67.570 34.320 ;
        RECT 67.810 34.285 67.960 34.455 ;
        RECT 68.200 34.285 68.350 34.455 ;
        RECT 68.590 34.150 68.740 34.320 ;
        RECT 70.320 34.150 70.470 34.320 ;
        RECT 70.710 34.285 70.860 34.455 ;
        RECT 71.100 34.285 71.250 34.455 ;
        RECT 71.490 34.150 71.640 34.320 ;
        RECT 73.220 34.150 73.370 34.320 ;
        RECT 73.610 34.285 73.760 34.455 ;
        RECT 74.000 34.285 74.150 34.455 ;
        RECT 74.390 34.150 74.540 34.320 ;
        RECT 76.120 34.150 76.270 34.320 ;
        RECT 76.510 34.285 76.660 34.455 ;
        RECT 76.900 34.285 77.050 34.455 ;
        RECT 77.290 34.150 77.440 34.320 ;
        RECT 79.020 34.150 79.170 34.320 ;
        RECT 79.410 34.285 79.560 34.455 ;
        RECT 79.800 34.285 79.950 34.455 ;
        RECT 80.190 34.150 80.340 34.320 ;
        RECT 81.920 34.150 82.070 34.320 ;
        RECT 82.310 34.285 82.460 34.455 ;
        RECT 82.700 34.285 82.850 34.455 ;
        RECT 83.090 34.150 83.240 34.320 ;
        RECT 84.820 34.150 84.970 34.320 ;
        RECT 85.210 34.285 85.360 34.455 ;
        RECT 85.600 34.285 85.750 34.455 ;
        RECT 85.990 34.150 86.140 34.320 ;
        RECT 87.720 34.150 87.870 34.320 ;
        RECT 88.110 34.285 88.260 34.455 ;
        RECT 88.500 34.285 88.650 34.455 ;
        RECT 88.890 34.150 89.040 34.320 ;
        RECT 90.620 34.150 90.770 34.320 ;
        RECT 91.010 34.285 91.160 34.455 ;
        RECT 91.400 34.285 91.550 34.455 ;
        RECT 91.790 34.150 91.940 34.320 ;
        RECT 0.985 34.065 1.035 34.100 ;
        POLYGON 1.035 34.100 1.070 34.065 1.035 34.065 ;
        RECT 0.985 33.940 1.070 34.065 ;
        RECT 1.690 33.940 1.775 34.100 ;
        RECT 3.885 34.065 3.935 34.100 ;
        POLYGON 3.935 34.100 3.970 34.065 3.935 34.065 ;
        RECT 3.885 33.940 3.970 34.065 ;
        RECT 4.590 33.940 4.675 34.100 ;
        RECT 6.785 34.065 6.835 34.100 ;
        POLYGON 6.835 34.100 6.870 34.065 6.835 34.065 ;
        RECT 6.785 33.940 6.870 34.065 ;
        RECT 7.490 33.940 7.575 34.100 ;
        RECT 9.685 34.065 9.735 34.100 ;
        POLYGON 9.735 34.100 9.770 34.065 9.735 34.065 ;
        RECT 9.685 33.940 9.770 34.065 ;
        RECT 10.390 33.940 10.475 34.100 ;
        RECT 12.585 34.065 12.635 34.100 ;
        POLYGON 12.635 34.100 12.670 34.065 12.635 34.065 ;
        RECT 12.585 33.940 12.670 34.065 ;
        RECT 13.290 33.940 13.375 34.100 ;
        RECT 15.485 34.065 15.535 34.100 ;
        POLYGON 15.535 34.100 15.570 34.065 15.535 34.065 ;
        RECT 15.485 33.940 15.570 34.065 ;
        RECT 16.190 33.940 16.275 34.100 ;
        RECT 18.385 34.065 18.435 34.100 ;
        POLYGON 18.435 34.100 18.470 34.065 18.435 34.065 ;
        RECT 18.385 33.940 18.470 34.065 ;
        RECT 19.090 33.940 19.175 34.100 ;
        RECT 21.285 34.065 21.335 34.100 ;
        POLYGON 21.335 34.100 21.370 34.065 21.335 34.065 ;
        RECT 21.285 33.940 21.370 34.065 ;
        RECT 21.990 33.940 22.075 34.100 ;
        RECT 24.185 34.065 24.235 34.100 ;
        POLYGON 24.235 34.100 24.270 34.065 24.235 34.065 ;
        RECT 24.185 33.940 24.270 34.065 ;
        RECT 24.890 33.940 24.975 34.100 ;
        RECT 27.085 34.065 27.135 34.100 ;
        POLYGON 27.135 34.100 27.170 34.065 27.135 34.065 ;
        RECT 27.085 33.940 27.170 34.065 ;
        RECT 27.790 33.940 27.875 34.100 ;
        RECT 29.985 34.065 30.035 34.100 ;
        POLYGON 30.035 34.100 30.070 34.065 30.035 34.065 ;
        RECT 29.985 33.940 30.070 34.065 ;
        RECT 30.690 33.940 30.775 34.100 ;
        RECT 32.885 34.065 32.935 34.100 ;
        POLYGON 32.935 34.100 32.970 34.065 32.935 34.065 ;
        RECT 32.885 33.940 32.970 34.065 ;
        RECT 33.590 33.940 33.675 34.100 ;
        RECT 35.785 34.065 35.835 34.100 ;
        POLYGON 35.835 34.100 35.870 34.065 35.835 34.065 ;
        RECT 35.785 33.940 35.870 34.065 ;
        RECT 36.490 33.940 36.575 34.100 ;
        RECT 38.685 34.065 38.735 34.100 ;
        POLYGON 38.735 34.100 38.770 34.065 38.735 34.065 ;
        RECT 38.685 33.940 38.770 34.065 ;
        RECT 39.390 33.940 39.475 34.100 ;
        RECT 41.585 34.065 41.635 34.100 ;
        POLYGON 41.635 34.100 41.670 34.065 41.635 34.065 ;
        RECT 41.585 33.940 41.670 34.065 ;
        RECT 42.290 33.940 42.375 34.100 ;
        RECT 44.485 34.065 44.535 34.100 ;
        POLYGON 44.535 34.100 44.570 34.065 44.535 34.065 ;
        RECT 44.485 33.940 44.570 34.065 ;
        RECT 45.190 33.940 45.275 34.100 ;
        RECT 47.385 34.065 47.435 34.100 ;
        POLYGON 47.435 34.100 47.470 34.065 47.435 34.065 ;
        RECT 47.385 33.940 47.470 34.065 ;
        RECT 48.090 33.940 48.175 34.100 ;
        RECT 50.285 34.065 50.335 34.100 ;
        POLYGON 50.335 34.100 50.370 34.065 50.335 34.065 ;
        RECT 50.285 33.940 50.370 34.065 ;
        RECT 50.990 33.940 51.075 34.100 ;
        RECT 53.185 34.065 53.235 34.100 ;
        POLYGON 53.235 34.100 53.270 34.065 53.235 34.065 ;
        RECT 53.185 33.940 53.270 34.065 ;
        RECT 53.890 33.940 53.975 34.100 ;
        RECT 56.085 34.065 56.135 34.100 ;
        POLYGON 56.135 34.100 56.170 34.065 56.135 34.065 ;
        RECT 56.085 33.940 56.170 34.065 ;
        RECT 56.790 33.940 56.875 34.100 ;
        RECT 58.985 34.065 59.035 34.100 ;
        POLYGON 59.035 34.100 59.070 34.065 59.035 34.065 ;
        RECT 58.985 33.940 59.070 34.065 ;
        RECT 59.690 33.940 59.775 34.100 ;
        RECT 61.885 34.065 61.935 34.100 ;
        POLYGON 61.935 34.100 61.970 34.065 61.935 34.065 ;
        RECT 61.885 33.940 61.970 34.065 ;
        RECT 62.590 33.940 62.675 34.100 ;
        RECT 64.785 34.065 64.835 34.100 ;
        POLYGON 64.835 34.100 64.870 34.065 64.835 34.065 ;
        RECT 64.785 33.940 64.870 34.065 ;
        RECT 65.490 33.940 65.575 34.100 ;
        RECT 67.685 34.065 67.735 34.100 ;
        POLYGON 67.735 34.100 67.770 34.065 67.735 34.065 ;
        RECT 67.685 33.940 67.770 34.065 ;
        RECT 68.390 33.940 68.475 34.100 ;
        RECT 70.585 34.065 70.635 34.100 ;
        POLYGON 70.635 34.100 70.670 34.065 70.635 34.065 ;
        RECT 70.585 33.940 70.670 34.065 ;
        RECT 71.290 33.940 71.375 34.100 ;
        RECT 73.485 34.065 73.535 34.100 ;
        POLYGON 73.535 34.100 73.570 34.065 73.535 34.065 ;
        RECT 73.485 33.940 73.570 34.065 ;
        RECT 74.190 33.940 74.275 34.100 ;
        RECT 76.385 34.065 76.435 34.100 ;
        POLYGON 76.435 34.100 76.470 34.065 76.435 34.065 ;
        RECT 76.385 33.940 76.470 34.065 ;
        RECT 77.090 33.940 77.175 34.100 ;
        RECT 79.285 34.065 79.335 34.100 ;
        POLYGON 79.335 34.100 79.370 34.065 79.335 34.065 ;
        RECT 79.285 33.940 79.370 34.065 ;
        RECT 79.990 33.940 80.075 34.100 ;
        RECT 82.185 34.065 82.235 34.100 ;
        POLYGON 82.235 34.100 82.270 34.065 82.235 34.065 ;
        RECT 82.185 33.940 82.270 34.065 ;
        RECT 82.890 33.940 82.975 34.100 ;
        RECT 85.085 34.065 85.135 34.100 ;
        POLYGON 85.135 34.100 85.170 34.065 85.135 34.065 ;
        RECT 85.085 33.940 85.170 34.065 ;
        RECT 85.790 33.940 85.875 34.100 ;
        RECT 87.985 34.065 88.035 34.100 ;
        POLYGON 88.035 34.100 88.070 34.065 88.035 34.065 ;
        RECT 87.985 33.940 88.070 34.065 ;
        RECT 88.690 33.940 88.775 34.100 ;
        RECT 90.885 34.065 90.935 34.100 ;
        POLYGON 90.935 34.100 90.970 34.065 90.935 34.065 ;
        RECT 90.885 33.940 90.970 34.065 ;
        RECT 91.590 33.940 91.675 34.100 ;
        RECT 0.775 33.320 0.850 33.460 ;
        RECT 0.990 33.270 1.065 33.410 ;
        RECT 1.695 33.330 1.755 33.410 ;
        POLYGON 1.695 33.330 1.755 33.330 1.755 33.270 ;
        RECT 1.910 33.320 1.985 33.460 ;
        RECT 3.675 33.320 3.750 33.460 ;
        RECT 3.890 33.270 3.965 33.410 ;
        RECT 4.595 33.330 4.655 33.410 ;
        POLYGON 4.595 33.330 4.655 33.330 4.655 33.270 ;
        RECT 4.810 33.320 4.885 33.460 ;
        RECT 6.575 33.320 6.650 33.460 ;
        RECT 6.790 33.270 6.865 33.410 ;
        RECT 7.495 33.330 7.555 33.410 ;
        POLYGON 7.495 33.330 7.555 33.330 7.555 33.270 ;
        RECT 7.710 33.320 7.785 33.460 ;
        RECT 9.475 33.320 9.550 33.460 ;
        RECT 9.690 33.270 9.765 33.410 ;
        RECT 10.395 33.330 10.455 33.410 ;
        POLYGON 10.395 33.330 10.455 33.330 10.455 33.270 ;
        RECT 10.610 33.320 10.685 33.460 ;
        RECT 12.375 33.320 12.450 33.460 ;
        RECT 12.590 33.270 12.665 33.410 ;
        RECT 13.295 33.330 13.355 33.410 ;
        POLYGON 13.295 33.330 13.355 33.330 13.355 33.270 ;
        RECT 13.510 33.320 13.585 33.460 ;
        RECT 15.275 33.320 15.350 33.460 ;
        RECT 15.490 33.270 15.565 33.410 ;
        RECT 16.195 33.330 16.255 33.410 ;
        POLYGON 16.195 33.330 16.255 33.330 16.255 33.270 ;
        RECT 16.410 33.320 16.485 33.460 ;
        RECT 18.175 33.320 18.250 33.460 ;
        RECT 18.390 33.270 18.465 33.410 ;
        RECT 19.095 33.330 19.155 33.410 ;
        POLYGON 19.095 33.330 19.155 33.330 19.155 33.270 ;
        RECT 19.310 33.320 19.385 33.460 ;
        RECT 21.075 33.320 21.150 33.460 ;
        RECT 21.290 33.270 21.365 33.410 ;
        RECT 21.995 33.330 22.055 33.410 ;
        POLYGON 21.995 33.330 22.055 33.330 22.055 33.270 ;
        RECT 22.210 33.320 22.285 33.460 ;
        RECT 23.975 33.320 24.050 33.460 ;
        RECT 24.190 33.270 24.265 33.410 ;
        RECT 24.895 33.330 24.955 33.410 ;
        POLYGON 24.895 33.330 24.955 33.330 24.955 33.270 ;
        RECT 25.110 33.320 25.185 33.460 ;
        RECT 26.875 33.320 26.950 33.460 ;
        RECT 27.090 33.270 27.165 33.410 ;
        RECT 27.795 33.330 27.855 33.410 ;
        POLYGON 27.795 33.330 27.855 33.330 27.855 33.270 ;
        RECT 28.010 33.320 28.085 33.460 ;
        RECT 29.775 33.320 29.850 33.460 ;
        RECT 29.990 33.270 30.065 33.410 ;
        RECT 30.695 33.330 30.755 33.410 ;
        POLYGON 30.695 33.330 30.755 33.330 30.755 33.270 ;
        RECT 30.910 33.320 30.985 33.460 ;
        RECT 32.675 33.320 32.750 33.460 ;
        RECT 32.890 33.270 32.965 33.410 ;
        RECT 33.595 33.330 33.655 33.410 ;
        POLYGON 33.595 33.330 33.655 33.330 33.655 33.270 ;
        RECT 33.810 33.320 33.885 33.460 ;
        RECT 35.575 33.320 35.650 33.460 ;
        RECT 35.790 33.270 35.865 33.410 ;
        RECT 36.495 33.330 36.555 33.410 ;
        POLYGON 36.495 33.330 36.555 33.330 36.555 33.270 ;
        RECT 36.710 33.320 36.785 33.460 ;
        RECT 38.475 33.320 38.550 33.460 ;
        RECT 38.690 33.270 38.765 33.410 ;
        RECT 39.395 33.330 39.455 33.410 ;
        POLYGON 39.395 33.330 39.455 33.330 39.455 33.270 ;
        RECT 39.610 33.320 39.685 33.460 ;
        RECT 41.375 33.320 41.450 33.460 ;
        RECT 41.590 33.270 41.665 33.410 ;
        RECT 42.295 33.330 42.355 33.410 ;
        POLYGON 42.295 33.330 42.355 33.330 42.355 33.270 ;
        RECT 42.510 33.320 42.585 33.460 ;
        RECT 44.275 33.320 44.350 33.460 ;
        RECT 44.490 33.270 44.565 33.410 ;
        RECT 45.195 33.330 45.255 33.410 ;
        POLYGON 45.195 33.330 45.255 33.330 45.255 33.270 ;
        RECT 45.410 33.320 45.485 33.460 ;
        RECT 47.175 33.320 47.250 33.460 ;
        RECT 47.390 33.270 47.465 33.410 ;
        RECT 48.095 33.330 48.155 33.410 ;
        POLYGON 48.095 33.330 48.155 33.330 48.155 33.270 ;
        RECT 48.310 33.320 48.385 33.460 ;
        RECT 50.075 33.320 50.150 33.460 ;
        RECT 50.290 33.270 50.365 33.410 ;
        RECT 50.995 33.330 51.055 33.410 ;
        POLYGON 50.995 33.330 51.055 33.330 51.055 33.270 ;
        RECT 51.210 33.320 51.285 33.460 ;
        RECT 52.975 33.320 53.050 33.460 ;
        RECT 53.190 33.270 53.265 33.410 ;
        RECT 53.895 33.330 53.955 33.410 ;
        POLYGON 53.895 33.330 53.955 33.330 53.955 33.270 ;
        RECT 54.110 33.320 54.185 33.460 ;
        RECT 55.875 33.320 55.950 33.460 ;
        RECT 56.090 33.270 56.165 33.410 ;
        RECT 56.795 33.330 56.855 33.410 ;
        POLYGON 56.795 33.330 56.855 33.330 56.855 33.270 ;
        RECT 57.010 33.320 57.085 33.460 ;
        RECT 58.775 33.320 58.850 33.460 ;
        RECT 58.990 33.270 59.065 33.410 ;
        RECT 59.695 33.330 59.755 33.410 ;
        POLYGON 59.695 33.330 59.755 33.330 59.755 33.270 ;
        RECT 59.910 33.320 59.985 33.460 ;
        RECT 61.675 33.320 61.750 33.460 ;
        RECT 61.890 33.270 61.965 33.410 ;
        RECT 62.595 33.330 62.655 33.410 ;
        POLYGON 62.595 33.330 62.655 33.330 62.655 33.270 ;
        RECT 62.810 33.320 62.885 33.460 ;
        RECT 64.575 33.320 64.650 33.460 ;
        RECT 64.790 33.270 64.865 33.410 ;
        RECT 65.495 33.330 65.555 33.410 ;
        POLYGON 65.495 33.330 65.555 33.330 65.555 33.270 ;
        RECT 65.710 33.320 65.785 33.460 ;
        RECT 67.475 33.320 67.550 33.460 ;
        RECT 67.690 33.270 67.765 33.410 ;
        RECT 68.395 33.330 68.455 33.410 ;
        POLYGON 68.395 33.330 68.455 33.330 68.455 33.270 ;
        RECT 68.610 33.320 68.685 33.460 ;
        RECT 70.375 33.320 70.450 33.460 ;
        RECT 70.590 33.270 70.665 33.410 ;
        RECT 71.295 33.330 71.355 33.410 ;
        POLYGON 71.295 33.330 71.355 33.330 71.355 33.270 ;
        RECT 71.510 33.320 71.585 33.460 ;
        RECT 73.275 33.320 73.350 33.460 ;
        RECT 73.490 33.270 73.565 33.410 ;
        RECT 74.195 33.330 74.255 33.410 ;
        POLYGON 74.195 33.330 74.255 33.330 74.255 33.270 ;
        RECT 74.410 33.320 74.485 33.460 ;
        RECT 76.175 33.320 76.250 33.460 ;
        RECT 76.390 33.270 76.465 33.410 ;
        RECT 77.095 33.330 77.155 33.410 ;
        POLYGON 77.095 33.330 77.155 33.330 77.155 33.270 ;
        RECT 77.310 33.320 77.385 33.460 ;
        RECT 79.075 33.320 79.150 33.460 ;
        RECT 79.290 33.270 79.365 33.410 ;
        RECT 79.995 33.330 80.055 33.410 ;
        POLYGON 79.995 33.330 80.055 33.330 80.055 33.270 ;
        RECT 80.210 33.320 80.285 33.460 ;
        RECT 81.975 33.320 82.050 33.460 ;
        RECT 82.190 33.270 82.265 33.410 ;
        RECT 82.895 33.330 82.955 33.410 ;
        POLYGON 82.895 33.330 82.955 33.330 82.955 33.270 ;
        RECT 83.110 33.320 83.185 33.460 ;
        RECT 84.875 33.320 84.950 33.460 ;
        RECT 85.090 33.270 85.165 33.410 ;
        RECT 85.795 33.330 85.855 33.410 ;
        POLYGON 85.795 33.330 85.855 33.330 85.855 33.270 ;
        RECT 86.010 33.320 86.085 33.460 ;
        RECT 87.775 33.320 87.850 33.460 ;
        RECT 87.990 33.270 88.065 33.410 ;
        RECT 88.695 33.330 88.755 33.410 ;
        POLYGON 88.695 33.330 88.755 33.330 88.755 33.270 ;
        RECT 88.910 33.320 88.985 33.460 ;
        RECT 90.675 33.320 90.750 33.460 ;
        RECT 90.890 33.270 90.965 33.410 ;
        RECT 91.595 33.330 91.655 33.410 ;
        POLYGON 91.595 33.330 91.655 33.330 91.655 33.270 ;
        RECT 91.810 33.320 91.885 33.460 ;
        RECT 0.720 32.800 0.870 32.970 ;
        RECT 1.110 32.935 1.260 33.105 ;
        RECT 1.500 32.935 1.650 33.105 ;
        RECT 1.890 32.800 2.040 32.970 ;
        RECT 3.620 32.800 3.770 32.970 ;
        RECT 4.010 32.935 4.160 33.105 ;
        RECT 4.400 32.935 4.550 33.105 ;
        RECT 4.790 32.800 4.940 32.970 ;
        RECT 6.520 32.800 6.670 32.970 ;
        RECT 6.910 32.935 7.060 33.105 ;
        RECT 7.300 32.935 7.450 33.105 ;
        RECT 7.690 32.800 7.840 32.970 ;
        RECT 9.420 32.800 9.570 32.970 ;
        RECT 9.810 32.935 9.960 33.105 ;
        RECT 10.200 32.935 10.350 33.105 ;
        RECT 10.590 32.800 10.740 32.970 ;
        RECT 12.320 32.800 12.470 32.970 ;
        RECT 12.710 32.935 12.860 33.105 ;
        RECT 13.100 32.935 13.250 33.105 ;
        RECT 13.490 32.800 13.640 32.970 ;
        RECT 15.220 32.800 15.370 32.970 ;
        RECT 15.610 32.935 15.760 33.105 ;
        RECT 16.000 32.935 16.150 33.105 ;
        RECT 16.390 32.800 16.540 32.970 ;
        RECT 18.120 32.800 18.270 32.970 ;
        RECT 18.510 32.935 18.660 33.105 ;
        RECT 18.900 32.935 19.050 33.105 ;
        RECT 19.290 32.800 19.440 32.970 ;
        RECT 21.020 32.800 21.170 32.970 ;
        RECT 21.410 32.935 21.560 33.105 ;
        RECT 21.800 32.935 21.950 33.105 ;
        RECT 22.190 32.800 22.340 32.970 ;
        RECT 23.920 32.800 24.070 32.970 ;
        RECT 24.310 32.935 24.460 33.105 ;
        RECT 24.700 32.935 24.850 33.105 ;
        RECT 25.090 32.800 25.240 32.970 ;
        RECT 26.820 32.800 26.970 32.970 ;
        RECT 27.210 32.935 27.360 33.105 ;
        RECT 27.600 32.935 27.750 33.105 ;
        RECT 27.990 32.800 28.140 32.970 ;
        RECT 29.720 32.800 29.870 32.970 ;
        RECT 30.110 32.935 30.260 33.105 ;
        RECT 30.500 32.935 30.650 33.105 ;
        RECT 30.890 32.800 31.040 32.970 ;
        RECT 32.620 32.800 32.770 32.970 ;
        RECT 33.010 32.935 33.160 33.105 ;
        RECT 33.400 32.935 33.550 33.105 ;
        RECT 33.790 32.800 33.940 32.970 ;
        RECT 35.520 32.800 35.670 32.970 ;
        RECT 35.910 32.935 36.060 33.105 ;
        RECT 36.300 32.935 36.450 33.105 ;
        RECT 36.690 32.800 36.840 32.970 ;
        RECT 38.420 32.800 38.570 32.970 ;
        RECT 38.810 32.935 38.960 33.105 ;
        RECT 39.200 32.935 39.350 33.105 ;
        RECT 39.590 32.800 39.740 32.970 ;
        RECT 41.320 32.800 41.470 32.970 ;
        RECT 41.710 32.935 41.860 33.105 ;
        RECT 42.100 32.935 42.250 33.105 ;
        RECT 42.490 32.800 42.640 32.970 ;
        RECT 44.220 32.800 44.370 32.970 ;
        RECT 44.610 32.935 44.760 33.105 ;
        RECT 45.000 32.935 45.150 33.105 ;
        RECT 45.390 32.800 45.540 32.970 ;
        RECT 47.120 32.800 47.270 32.970 ;
        RECT 47.510 32.935 47.660 33.105 ;
        RECT 47.900 32.935 48.050 33.105 ;
        RECT 48.290 32.800 48.440 32.970 ;
        RECT 50.020 32.800 50.170 32.970 ;
        RECT 50.410 32.935 50.560 33.105 ;
        RECT 50.800 32.935 50.950 33.105 ;
        RECT 51.190 32.800 51.340 32.970 ;
        RECT 52.920 32.800 53.070 32.970 ;
        RECT 53.310 32.935 53.460 33.105 ;
        RECT 53.700 32.935 53.850 33.105 ;
        RECT 54.090 32.800 54.240 32.970 ;
        RECT 55.820 32.800 55.970 32.970 ;
        RECT 56.210 32.935 56.360 33.105 ;
        RECT 56.600 32.935 56.750 33.105 ;
        RECT 56.990 32.800 57.140 32.970 ;
        RECT 58.720 32.800 58.870 32.970 ;
        RECT 59.110 32.935 59.260 33.105 ;
        RECT 59.500 32.935 59.650 33.105 ;
        RECT 59.890 32.800 60.040 32.970 ;
        RECT 61.620 32.800 61.770 32.970 ;
        RECT 62.010 32.935 62.160 33.105 ;
        RECT 62.400 32.935 62.550 33.105 ;
        RECT 62.790 32.800 62.940 32.970 ;
        RECT 64.520 32.800 64.670 32.970 ;
        RECT 64.910 32.935 65.060 33.105 ;
        RECT 65.300 32.935 65.450 33.105 ;
        RECT 65.690 32.800 65.840 32.970 ;
        RECT 67.420 32.800 67.570 32.970 ;
        RECT 67.810 32.935 67.960 33.105 ;
        RECT 68.200 32.935 68.350 33.105 ;
        RECT 68.590 32.800 68.740 32.970 ;
        RECT 70.320 32.800 70.470 32.970 ;
        RECT 70.710 32.935 70.860 33.105 ;
        RECT 71.100 32.935 71.250 33.105 ;
        RECT 71.490 32.800 71.640 32.970 ;
        RECT 73.220 32.800 73.370 32.970 ;
        RECT 73.610 32.935 73.760 33.105 ;
        RECT 74.000 32.935 74.150 33.105 ;
        RECT 74.390 32.800 74.540 32.970 ;
        RECT 76.120 32.800 76.270 32.970 ;
        RECT 76.510 32.935 76.660 33.105 ;
        RECT 76.900 32.935 77.050 33.105 ;
        RECT 77.290 32.800 77.440 32.970 ;
        RECT 79.020 32.800 79.170 32.970 ;
        RECT 79.410 32.935 79.560 33.105 ;
        RECT 79.800 32.935 79.950 33.105 ;
        RECT 80.190 32.800 80.340 32.970 ;
        RECT 81.920 32.800 82.070 32.970 ;
        RECT 82.310 32.935 82.460 33.105 ;
        RECT 82.700 32.935 82.850 33.105 ;
        RECT 83.090 32.800 83.240 32.970 ;
        RECT 84.820 32.800 84.970 32.970 ;
        RECT 85.210 32.935 85.360 33.105 ;
        RECT 85.600 32.935 85.750 33.105 ;
        RECT 85.990 32.800 86.140 32.970 ;
        RECT 87.720 32.800 87.870 32.970 ;
        RECT 88.110 32.935 88.260 33.105 ;
        RECT 88.500 32.935 88.650 33.105 ;
        RECT 88.890 32.800 89.040 32.970 ;
        RECT 90.620 32.800 90.770 32.970 ;
        RECT 91.010 32.935 91.160 33.105 ;
        RECT 91.400 32.935 91.550 33.105 ;
        RECT 91.790 32.800 91.940 32.970 ;
        RECT 0.985 32.715 1.035 32.750 ;
        POLYGON 1.035 32.750 1.070 32.715 1.035 32.715 ;
        RECT 0.985 32.590 1.070 32.715 ;
        RECT 1.690 32.590 1.775 32.750 ;
        RECT 3.885 32.715 3.935 32.750 ;
        POLYGON 3.935 32.750 3.970 32.715 3.935 32.715 ;
        RECT 3.885 32.590 3.970 32.715 ;
        RECT 4.590 32.590 4.675 32.750 ;
        RECT 6.785 32.715 6.835 32.750 ;
        POLYGON 6.835 32.750 6.870 32.715 6.835 32.715 ;
        RECT 6.785 32.590 6.870 32.715 ;
        RECT 7.490 32.590 7.575 32.750 ;
        RECT 9.685 32.715 9.735 32.750 ;
        POLYGON 9.735 32.750 9.770 32.715 9.735 32.715 ;
        RECT 9.685 32.590 9.770 32.715 ;
        RECT 10.390 32.590 10.475 32.750 ;
        RECT 12.585 32.715 12.635 32.750 ;
        POLYGON 12.635 32.750 12.670 32.715 12.635 32.715 ;
        RECT 12.585 32.590 12.670 32.715 ;
        RECT 13.290 32.590 13.375 32.750 ;
        RECT 15.485 32.715 15.535 32.750 ;
        POLYGON 15.535 32.750 15.570 32.715 15.535 32.715 ;
        RECT 15.485 32.590 15.570 32.715 ;
        RECT 16.190 32.590 16.275 32.750 ;
        RECT 18.385 32.715 18.435 32.750 ;
        POLYGON 18.435 32.750 18.470 32.715 18.435 32.715 ;
        RECT 18.385 32.590 18.470 32.715 ;
        RECT 19.090 32.590 19.175 32.750 ;
        RECT 21.285 32.715 21.335 32.750 ;
        POLYGON 21.335 32.750 21.370 32.715 21.335 32.715 ;
        RECT 21.285 32.590 21.370 32.715 ;
        RECT 21.990 32.590 22.075 32.750 ;
        RECT 24.185 32.715 24.235 32.750 ;
        POLYGON 24.235 32.750 24.270 32.715 24.235 32.715 ;
        RECT 24.185 32.590 24.270 32.715 ;
        RECT 24.890 32.590 24.975 32.750 ;
        RECT 27.085 32.715 27.135 32.750 ;
        POLYGON 27.135 32.750 27.170 32.715 27.135 32.715 ;
        RECT 27.085 32.590 27.170 32.715 ;
        RECT 27.790 32.590 27.875 32.750 ;
        RECT 29.985 32.715 30.035 32.750 ;
        POLYGON 30.035 32.750 30.070 32.715 30.035 32.715 ;
        RECT 29.985 32.590 30.070 32.715 ;
        RECT 30.690 32.590 30.775 32.750 ;
        RECT 32.885 32.715 32.935 32.750 ;
        POLYGON 32.935 32.750 32.970 32.715 32.935 32.715 ;
        RECT 32.885 32.590 32.970 32.715 ;
        RECT 33.590 32.590 33.675 32.750 ;
        RECT 35.785 32.715 35.835 32.750 ;
        POLYGON 35.835 32.750 35.870 32.715 35.835 32.715 ;
        RECT 35.785 32.590 35.870 32.715 ;
        RECT 36.490 32.590 36.575 32.750 ;
        RECT 38.685 32.715 38.735 32.750 ;
        POLYGON 38.735 32.750 38.770 32.715 38.735 32.715 ;
        RECT 38.685 32.590 38.770 32.715 ;
        RECT 39.390 32.590 39.475 32.750 ;
        RECT 41.585 32.715 41.635 32.750 ;
        POLYGON 41.635 32.750 41.670 32.715 41.635 32.715 ;
        RECT 41.585 32.590 41.670 32.715 ;
        RECT 42.290 32.590 42.375 32.750 ;
        RECT 44.485 32.715 44.535 32.750 ;
        POLYGON 44.535 32.750 44.570 32.715 44.535 32.715 ;
        RECT 44.485 32.590 44.570 32.715 ;
        RECT 45.190 32.590 45.275 32.750 ;
        RECT 47.385 32.715 47.435 32.750 ;
        POLYGON 47.435 32.750 47.470 32.715 47.435 32.715 ;
        RECT 47.385 32.590 47.470 32.715 ;
        RECT 48.090 32.590 48.175 32.750 ;
        RECT 50.285 32.715 50.335 32.750 ;
        POLYGON 50.335 32.750 50.370 32.715 50.335 32.715 ;
        RECT 50.285 32.590 50.370 32.715 ;
        RECT 50.990 32.590 51.075 32.750 ;
        RECT 53.185 32.715 53.235 32.750 ;
        POLYGON 53.235 32.750 53.270 32.715 53.235 32.715 ;
        RECT 53.185 32.590 53.270 32.715 ;
        RECT 53.890 32.590 53.975 32.750 ;
        RECT 56.085 32.715 56.135 32.750 ;
        POLYGON 56.135 32.750 56.170 32.715 56.135 32.715 ;
        RECT 56.085 32.590 56.170 32.715 ;
        RECT 56.790 32.590 56.875 32.750 ;
        RECT 58.985 32.715 59.035 32.750 ;
        POLYGON 59.035 32.750 59.070 32.715 59.035 32.715 ;
        RECT 58.985 32.590 59.070 32.715 ;
        RECT 59.690 32.590 59.775 32.750 ;
        RECT 61.885 32.715 61.935 32.750 ;
        POLYGON 61.935 32.750 61.970 32.715 61.935 32.715 ;
        RECT 61.885 32.590 61.970 32.715 ;
        RECT 62.590 32.590 62.675 32.750 ;
        RECT 64.785 32.715 64.835 32.750 ;
        POLYGON 64.835 32.750 64.870 32.715 64.835 32.715 ;
        RECT 64.785 32.590 64.870 32.715 ;
        RECT 65.490 32.590 65.575 32.750 ;
        RECT 67.685 32.715 67.735 32.750 ;
        POLYGON 67.735 32.750 67.770 32.715 67.735 32.715 ;
        RECT 67.685 32.590 67.770 32.715 ;
        RECT 68.390 32.590 68.475 32.750 ;
        RECT 70.585 32.715 70.635 32.750 ;
        POLYGON 70.635 32.750 70.670 32.715 70.635 32.715 ;
        RECT 70.585 32.590 70.670 32.715 ;
        RECT 71.290 32.590 71.375 32.750 ;
        RECT 73.485 32.715 73.535 32.750 ;
        POLYGON 73.535 32.750 73.570 32.715 73.535 32.715 ;
        RECT 73.485 32.590 73.570 32.715 ;
        RECT 74.190 32.590 74.275 32.750 ;
        RECT 76.385 32.715 76.435 32.750 ;
        POLYGON 76.435 32.750 76.470 32.715 76.435 32.715 ;
        RECT 76.385 32.590 76.470 32.715 ;
        RECT 77.090 32.590 77.175 32.750 ;
        RECT 79.285 32.715 79.335 32.750 ;
        POLYGON 79.335 32.750 79.370 32.715 79.335 32.715 ;
        RECT 79.285 32.590 79.370 32.715 ;
        RECT 79.990 32.590 80.075 32.750 ;
        RECT 82.185 32.715 82.235 32.750 ;
        POLYGON 82.235 32.750 82.270 32.715 82.235 32.715 ;
        RECT 82.185 32.590 82.270 32.715 ;
        RECT 82.890 32.590 82.975 32.750 ;
        RECT 85.085 32.715 85.135 32.750 ;
        POLYGON 85.135 32.750 85.170 32.715 85.135 32.715 ;
        RECT 85.085 32.590 85.170 32.715 ;
        RECT 85.790 32.590 85.875 32.750 ;
        RECT 87.985 32.715 88.035 32.750 ;
        POLYGON 88.035 32.750 88.070 32.715 88.035 32.715 ;
        RECT 87.985 32.590 88.070 32.715 ;
        RECT 88.690 32.590 88.775 32.750 ;
        RECT 90.885 32.715 90.935 32.750 ;
        POLYGON 90.935 32.750 90.970 32.715 90.935 32.715 ;
        RECT 90.885 32.590 90.970 32.715 ;
        RECT 91.590 32.590 91.675 32.750 ;
        RECT 0.775 31.970 0.850 32.110 ;
        RECT 0.990 31.920 1.065 32.060 ;
        RECT 1.695 31.980 1.755 32.060 ;
        POLYGON 1.695 31.980 1.755 31.980 1.755 31.920 ;
        RECT 1.910 31.970 1.985 32.110 ;
        RECT 3.675 31.970 3.750 32.110 ;
        RECT 3.890 31.920 3.965 32.060 ;
        RECT 4.595 31.980 4.655 32.060 ;
        POLYGON 4.595 31.980 4.655 31.980 4.655 31.920 ;
        RECT 4.810 31.970 4.885 32.110 ;
        RECT 6.575 31.970 6.650 32.110 ;
        RECT 6.790 31.920 6.865 32.060 ;
        RECT 7.495 31.980 7.555 32.060 ;
        POLYGON 7.495 31.980 7.555 31.980 7.555 31.920 ;
        RECT 7.710 31.970 7.785 32.110 ;
        RECT 9.475 31.970 9.550 32.110 ;
        RECT 9.690 31.920 9.765 32.060 ;
        RECT 10.395 31.980 10.455 32.060 ;
        POLYGON 10.395 31.980 10.455 31.980 10.455 31.920 ;
        RECT 10.610 31.970 10.685 32.110 ;
        RECT 12.375 31.970 12.450 32.110 ;
        RECT 12.590 31.920 12.665 32.060 ;
        RECT 13.295 31.980 13.355 32.060 ;
        POLYGON 13.295 31.980 13.355 31.980 13.355 31.920 ;
        RECT 13.510 31.970 13.585 32.110 ;
        RECT 15.275 31.970 15.350 32.110 ;
        RECT 15.490 31.920 15.565 32.060 ;
        RECT 16.195 31.980 16.255 32.060 ;
        POLYGON 16.195 31.980 16.255 31.980 16.255 31.920 ;
        RECT 16.410 31.970 16.485 32.110 ;
        RECT 18.175 31.970 18.250 32.110 ;
        RECT 18.390 31.920 18.465 32.060 ;
        RECT 19.095 31.980 19.155 32.060 ;
        POLYGON 19.095 31.980 19.155 31.980 19.155 31.920 ;
        RECT 19.310 31.970 19.385 32.110 ;
        RECT 21.075 31.970 21.150 32.110 ;
        RECT 21.290 31.920 21.365 32.060 ;
        RECT 21.995 31.980 22.055 32.060 ;
        POLYGON 21.995 31.980 22.055 31.980 22.055 31.920 ;
        RECT 22.210 31.970 22.285 32.110 ;
        RECT 23.975 31.970 24.050 32.110 ;
        RECT 24.190 31.920 24.265 32.060 ;
        RECT 24.895 31.980 24.955 32.060 ;
        POLYGON 24.895 31.980 24.955 31.980 24.955 31.920 ;
        RECT 25.110 31.970 25.185 32.110 ;
        RECT 26.875 31.970 26.950 32.110 ;
        RECT 27.090 31.920 27.165 32.060 ;
        RECT 27.795 31.980 27.855 32.060 ;
        POLYGON 27.795 31.980 27.855 31.980 27.855 31.920 ;
        RECT 28.010 31.970 28.085 32.110 ;
        RECT 29.775 31.970 29.850 32.110 ;
        RECT 29.990 31.920 30.065 32.060 ;
        RECT 30.695 31.980 30.755 32.060 ;
        POLYGON 30.695 31.980 30.755 31.980 30.755 31.920 ;
        RECT 30.910 31.970 30.985 32.110 ;
        RECT 32.675 31.970 32.750 32.110 ;
        RECT 32.890 31.920 32.965 32.060 ;
        RECT 33.595 31.980 33.655 32.060 ;
        POLYGON 33.595 31.980 33.655 31.980 33.655 31.920 ;
        RECT 33.810 31.970 33.885 32.110 ;
        RECT 35.575 31.970 35.650 32.110 ;
        RECT 35.790 31.920 35.865 32.060 ;
        RECT 36.495 31.980 36.555 32.060 ;
        POLYGON 36.495 31.980 36.555 31.980 36.555 31.920 ;
        RECT 36.710 31.970 36.785 32.110 ;
        RECT 38.475 31.970 38.550 32.110 ;
        RECT 38.690 31.920 38.765 32.060 ;
        RECT 39.395 31.980 39.455 32.060 ;
        POLYGON 39.395 31.980 39.455 31.980 39.455 31.920 ;
        RECT 39.610 31.970 39.685 32.110 ;
        RECT 41.375 31.970 41.450 32.110 ;
        RECT 41.590 31.920 41.665 32.060 ;
        RECT 42.295 31.980 42.355 32.060 ;
        POLYGON 42.295 31.980 42.355 31.980 42.355 31.920 ;
        RECT 42.510 31.970 42.585 32.110 ;
        RECT 44.275 31.970 44.350 32.110 ;
        RECT 44.490 31.920 44.565 32.060 ;
        RECT 45.195 31.980 45.255 32.060 ;
        POLYGON 45.195 31.980 45.255 31.980 45.255 31.920 ;
        RECT 45.410 31.970 45.485 32.110 ;
        RECT 47.175 31.970 47.250 32.110 ;
        RECT 47.390 31.920 47.465 32.060 ;
        RECT 48.095 31.980 48.155 32.060 ;
        POLYGON 48.095 31.980 48.155 31.980 48.155 31.920 ;
        RECT 48.310 31.970 48.385 32.110 ;
        RECT 50.075 31.970 50.150 32.110 ;
        RECT 50.290 31.920 50.365 32.060 ;
        RECT 50.995 31.980 51.055 32.060 ;
        POLYGON 50.995 31.980 51.055 31.980 51.055 31.920 ;
        RECT 51.210 31.970 51.285 32.110 ;
        RECT 52.975 31.970 53.050 32.110 ;
        RECT 53.190 31.920 53.265 32.060 ;
        RECT 53.895 31.980 53.955 32.060 ;
        POLYGON 53.895 31.980 53.955 31.980 53.955 31.920 ;
        RECT 54.110 31.970 54.185 32.110 ;
        RECT 55.875 31.970 55.950 32.110 ;
        RECT 56.090 31.920 56.165 32.060 ;
        RECT 56.795 31.980 56.855 32.060 ;
        POLYGON 56.795 31.980 56.855 31.980 56.855 31.920 ;
        RECT 57.010 31.970 57.085 32.110 ;
        RECT 58.775 31.970 58.850 32.110 ;
        RECT 58.990 31.920 59.065 32.060 ;
        RECT 59.695 31.980 59.755 32.060 ;
        POLYGON 59.695 31.980 59.755 31.980 59.755 31.920 ;
        RECT 59.910 31.970 59.985 32.110 ;
        RECT 61.675 31.970 61.750 32.110 ;
        RECT 61.890 31.920 61.965 32.060 ;
        RECT 62.595 31.980 62.655 32.060 ;
        POLYGON 62.595 31.980 62.655 31.980 62.655 31.920 ;
        RECT 62.810 31.970 62.885 32.110 ;
        RECT 64.575 31.970 64.650 32.110 ;
        RECT 64.790 31.920 64.865 32.060 ;
        RECT 65.495 31.980 65.555 32.060 ;
        POLYGON 65.495 31.980 65.555 31.980 65.555 31.920 ;
        RECT 65.710 31.970 65.785 32.110 ;
        RECT 67.475 31.970 67.550 32.110 ;
        RECT 67.690 31.920 67.765 32.060 ;
        RECT 68.395 31.980 68.455 32.060 ;
        POLYGON 68.395 31.980 68.455 31.980 68.455 31.920 ;
        RECT 68.610 31.970 68.685 32.110 ;
        RECT 70.375 31.970 70.450 32.110 ;
        RECT 70.590 31.920 70.665 32.060 ;
        RECT 71.295 31.980 71.355 32.060 ;
        POLYGON 71.295 31.980 71.355 31.980 71.355 31.920 ;
        RECT 71.510 31.970 71.585 32.110 ;
        RECT 73.275 31.970 73.350 32.110 ;
        RECT 73.490 31.920 73.565 32.060 ;
        RECT 74.195 31.980 74.255 32.060 ;
        POLYGON 74.195 31.980 74.255 31.980 74.255 31.920 ;
        RECT 74.410 31.970 74.485 32.110 ;
        RECT 76.175 31.970 76.250 32.110 ;
        RECT 76.390 31.920 76.465 32.060 ;
        RECT 77.095 31.980 77.155 32.060 ;
        POLYGON 77.095 31.980 77.155 31.980 77.155 31.920 ;
        RECT 77.310 31.970 77.385 32.110 ;
        RECT 79.075 31.970 79.150 32.110 ;
        RECT 79.290 31.920 79.365 32.060 ;
        RECT 79.995 31.980 80.055 32.060 ;
        POLYGON 79.995 31.980 80.055 31.980 80.055 31.920 ;
        RECT 80.210 31.970 80.285 32.110 ;
        RECT 81.975 31.970 82.050 32.110 ;
        RECT 82.190 31.920 82.265 32.060 ;
        RECT 82.895 31.980 82.955 32.060 ;
        POLYGON 82.895 31.980 82.955 31.980 82.955 31.920 ;
        RECT 83.110 31.970 83.185 32.110 ;
        RECT 84.875 31.970 84.950 32.110 ;
        RECT 85.090 31.920 85.165 32.060 ;
        RECT 85.795 31.980 85.855 32.060 ;
        POLYGON 85.795 31.980 85.855 31.980 85.855 31.920 ;
        RECT 86.010 31.970 86.085 32.110 ;
        RECT 87.775 31.970 87.850 32.110 ;
        RECT 87.990 31.920 88.065 32.060 ;
        RECT 88.695 31.980 88.755 32.060 ;
        POLYGON 88.695 31.980 88.755 31.980 88.755 31.920 ;
        RECT 88.910 31.970 88.985 32.110 ;
        RECT 90.675 31.970 90.750 32.110 ;
        RECT 90.890 31.920 90.965 32.060 ;
        RECT 91.595 31.980 91.655 32.060 ;
        POLYGON 91.595 31.980 91.655 31.980 91.655 31.920 ;
        RECT 91.810 31.970 91.885 32.110 ;
        RECT 0.720 31.450 0.870 31.620 ;
        RECT 1.110 31.585 1.260 31.755 ;
        RECT 1.500 31.585 1.650 31.755 ;
        RECT 1.890 31.450 2.040 31.620 ;
        RECT 3.620 31.450 3.770 31.620 ;
        RECT 4.010 31.585 4.160 31.755 ;
        RECT 4.400 31.585 4.550 31.755 ;
        RECT 4.790 31.450 4.940 31.620 ;
        RECT 6.520 31.450 6.670 31.620 ;
        RECT 6.910 31.585 7.060 31.755 ;
        RECT 7.300 31.585 7.450 31.755 ;
        RECT 7.690 31.450 7.840 31.620 ;
        RECT 9.420 31.450 9.570 31.620 ;
        RECT 9.810 31.585 9.960 31.755 ;
        RECT 10.200 31.585 10.350 31.755 ;
        RECT 10.590 31.450 10.740 31.620 ;
        RECT 12.320 31.450 12.470 31.620 ;
        RECT 12.710 31.585 12.860 31.755 ;
        RECT 13.100 31.585 13.250 31.755 ;
        RECT 13.490 31.450 13.640 31.620 ;
        RECT 15.220 31.450 15.370 31.620 ;
        RECT 15.610 31.585 15.760 31.755 ;
        RECT 16.000 31.585 16.150 31.755 ;
        RECT 16.390 31.450 16.540 31.620 ;
        RECT 18.120 31.450 18.270 31.620 ;
        RECT 18.510 31.585 18.660 31.755 ;
        RECT 18.900 31.585 19.050 31.755 ;
        RECT 19.290 31.450 19.440 31.620 ;
        RECT 21.020 31.450 21.170 31.620 ;
        RECT 21.410 31.585 21.560 31.755 ;
        RECT 21.800 31.585 21.950 31.755 ;
        RECT 22.190 31.450 22.340 31.620 ;
        RECT 23.920 31.450 24.070 31.620 ;
        RECT 24.310 31.585 24.460 31.755 ;
        RECT 24.700 31.585 24.850 31.755 ;
        RECT 25.090 31.450 25.240 31.620 ;
        RECT 26.820 31.450 26.970 31.620 ;
        RECT 27.210 31.585 27.360 31.755 ;
        RECT 27.600 31.585 27.750 31.755 ;
        RECT 27.990 31.450 28.140 31.620 ;
        RECT 29.720 31.450 29.870 31.620 ;
        RECT 30.110 31.585 30.260 31.755 ;
        RECT 30.500 31.585 30.650 31.755 ;
        RECT 30.890 31.450 31.040 31.620 ;
        RECT 32.620 31.450 32.770 31.620 ;
        RECT 33.010 31.585 33.160 31.755 ;
        RECT 33.400 31.585 33.550 31.755 ;
        RECT 33.790 31.450 33.940 31.620 ;
        RECT 35.520 31.450 35.670 31.620 ;
        RECT 35.910 31.585 36.060 31.755 ;
        RECT 36.300 31.585 36.450 31.755 ;
        RECT 36.690 31.450 36.840 31.620 ;
        RECT 38.420 31.450 38.570 31.620 ;
        RECT 38.810 31.585 38.960 31.755 ;
        RECT 39.200 31.585 39.350 31.755 ;
        RECT 39.590 31.450 39.740 31.620 ;
        RECT 41.320 31.450 41.470 31.620 ;
        RECT 41.710 31.585 41.860 31.755 ;
        RECT 42.100 31.585 42.250 31.755 ;
        RECT 42.490 31.450 42.640 31.620 ;
        RECT 44.220 31.450 44.370 31.620 ;
        RECT 44.610 31.585 44.760 31.755 ;
        RECT 45.000 31.585 45.150 31.755 ;
        RECT 45.390 31.450 45.540 31.620 ;
        RECT 47.120 31.450 47.270 31.620 ;
        RECT 47.510 31.585 47.660 31.755 ;
        RECT 47.900 31.585 48.050 31.755 ;
        RECT 48.290 31.450 48.440 31.620 ;
        RECT 50.020 31.450 50.170 31.620 ;
        RECT 50.410 31.585 50.560 31.755 ;
        RECT 50.800 31.585 50.950 31.755 ;
        RECT 51.190 31.450 51.340 31.620 ;
        RECT 52.920 31.450 53.070 31.620 ;
        RECT 53.310 31.585 53.460 31.755 ;
        RECT 53.700 31.585 53.850 31.755 ;
        RECT 54.090 31.450 54.240 31.620 ;
        RECT 55.820 31.450 55.970 31.620 ;
        RECT 56.210 31.585 56.360 31.755 ;
        RECT 56.600 31.585 56.750 31.755 ;
        RECT 56.990 31.450 57.140 31.620 ;
        RECT 58.720 31.450 58.870 31.620 ;
        RECT 59.110 31.585 59.260 31.755 ;
        RECT 59.500 31.585 59.650 31.755 ;
        RECT 59.890 31.450 60.040 31.620 ;
        RECT 61.620 31.450 61.770 31.620 ;
        RECT 62.010 31.585 62.160 31.755 ;
        RECT 62.400 31.585 62.550 31.755 ;
        RECT 62.790 31.450 62.940 31.620 ;
        RECT 64.520 31.450 64.670 31.620 ;
        RECT 64.910 31.585 65.060 31.755 ;
        RECT 65.300 31.585 65.450 31.755 ;
        RECT 65.690 31.450 65.840 31.620 ;
        RECT 67.420 31.450 67.570 31.620 ;
        RECT 67.810 31.585 67.960 31.755 ;
        RECT 68.200 31.585 68.350 31.755 ;
        RECT 68.590 31.450 68.740 31.620 ;
        RECT 70.320 31.450 70.470 31.620 ;
        RECT 70.710 31.585 70.860 31.755 ;
        RECT 71.100 31.585 71.250 31.755 ;
        RECT 71.490 31.450 71.640 31.620 ;
        RECT 73.220 31.450 73.370 31.620 ;
        RECT 73.610 31.585 73.760 31.755 ;
        RECT 74.000 31.585 74.150 31.755 ;
        RECT 74.390 31.450 74.540 31.620 ;
        RECT 76.120 31.450 76.270 31.620 ;
        RECT 76.510 31.585 76.660 31.755 ;
        RECT 76.900 31.585 77.050 31.755 ;
        RECT 77.290 31.450 77.440 31.620 ;
        RECT 79.020 31.450 79.170 31.620 ;
        RECT 79.410 31.585 79.560 31.755 ;
        RECT 79.800 31.585 79.950 31.755 ;
        RECT 80.190 31.450 80.340 31.620 ;
        RECT 81.920 31.450 82.070 31.620 ;
        RECT 82.310 31.585 82.460 31.755 ;
        RECT 82.700 31.585 82.850 31.755 ;
        RECT 83.090 31.450 83.240 31.620 ;
        RECT 84.820 31.450 84.970 31.620 ;
        RECT 85.210 31.585 85.360 31.755 ;
        RECT 85.600 31.585 85.750 31.755 ;
        RECT 85.990 31.450 86.140 31.620 ;
        RECT 87.720 31.450 87.870 31.620 ;
        RECT 88.110 31.585 88.260 31.755 ;
        RECT 88.500 31.585 88.650 31.755 ;
        RECT 88.890 31.450 89.040 31.620 ;
        RECT 90.620 31.450 90.770 31.620 ;
        RECT 91.010 31.585 91.160 31.755 ;
        RECT 91.400 31.585 91.550 31.755 ;
        RECT 91.790 31.450 91.940 31.620 ;
        RECT 0.985 31.365 1.035 31.400 ;
        POLYGON 1.035 31.400 1.070 31.365 1.035 31.365 ;
        RECT 0.985 31.240 1.070 31.365 ;
        RECT 1.690 31.240 1.775 31.400 ;
        RECT 3.885 31.365 3.935 31.400 ;
        POLYGON 3.935 31.400 3.970 31.365 3.935 31.365 ;
        RECT 3.885 31.240 3.970 31.365 ;
        RECT 4.590 31.240 4.675 31.400 ;
        RECT 6.785 31.365 6.835 31.400 ;
        POLYGON 6.835 31.400 6.870 31.365 6.835 31.365 ;
        RECT 6.785 31.240 6.870 31.365 ;
        RECT 7.490 31.240 7.575 31.400 ;
        RECT 9.685 31.365 9.735 31.400 ;
        POLYGON 9.735 31.400 9.770 31.365 9.735 31.365 ;
        RECT 9.685 31.240 9.770 31.365 ;
        RECT 10.390 31.240 10.475 31.400 ;
        RECT 12.585 31.365 12.635 31.400 ;
        POLYGON 12.635 31.400 12.670 31.365 12.635 31.365 ;
        RECT 12.585 31.240 12.670 31.365 ;
        RECT 13.290 31.240 13.375 31.400 ;
        RECT 15.485 31.365 15.535 31.400 ;
        POLYGON 15.535 31.400 15.570 31.365 15.535 31.365 ;
        RECT 15.485 31.240 15.570 31.365 ;
        RECT 16.190 31.240 16.275 31.400 ;
        RECT 18.385 31.365 18.435 31.400 ;
        POLYGON 18.435 31.400 18.470 31.365 18.435 31.365 ;
        RECT 18.385 31.240 18.470 31.365 ;
        RECT 19.090 31.240 19.175 31.400 ;
        RECT 21.285 31.365 21.335 31.400 ;
        POLYGON 21.335 31.400 21.370 31.365 21.335 31.365 ;
        RECT 21.285 31.240 21.370 31.365 ;
        RECT 21.990 31.240 22.075 31.400 ;
        RECT 24.185 31.365 24.235 31.400 ;
        POLYGON 24.235 31.400 24.270 31.365 24.235 31.365 ;
        RECT 24.185 31.240 24.270 31.365 ;
        RECT 24.890 31.240 24.975 31.400 ;
        RECT 27.085 31.365 27.135 31.400 ;
        POLYGON 27.135 31.400 27.170 31.365 27.135 31.365 ;
        RECT 27.085 31.240 27.170 31.365 ;
        RECT 27.790 31.240 27.875 31.400 ;
        RECT 29.985 31.365 30.035 31.400 ;
        POLYGON 30.035 31.400 30.070 31.365 30.035 31.365 ;
        RECT 29.985 31.240 30.070 31.365 ;
        RECT 30.690 31.240 30.775 31.400 ;
        RECT 32.885 31.365 32.935 31.400 ;
        POLYGON 32.935 31.400 32.970 31.365 32.935 31.365 ;
        RECT 32.885 31.240 32.970 31.365 ;
        RECT 33.590 31.240 33.675 31.400 ;
        RECT 35.785 31.365 35.835 31.400 ;
        POLYGON 35.835 31.400 35.870 31.365 35.835 31.365 ;
        RECT 35.785 31.240 35.870 31.365 ;
        RECT 36.490 31.240 36.575 31.400 ;
        RECT 38.685 31.365 38.735 31.400 ;
        POLYGON 38.735 31.400 38.770 31.365 38.735 31.365 ;
        RECT 38.685 31.240 38.770 31.365 ;
        RECT 39.390 31.240 39.475 31.400 ;
        RECT 41.585 31.365 41.635 31.400 ;
        POLYGON 41.635 31.400 41.670 31.365 41.635 31.365 ;
        RECT 41.585 31.240 41.670 31.365 ;
        RECT 42.290 31.240 42.375 31.400 ;
        RECT 44.485 31.365 44.535 31.400 ;
        POLYGON 44.535 31.400 44.570 31.365 44.535 31.365 ;
        RECT 44.485 31.240 44.570 31.365 ;
        RECT 45.190 31.240 45.275 31.400 ;
        RECT 47.385 31.365 47.435 31.400 ;
        POLYGON 47.435 31.400 47.470 31.365 47.435 31.365 ;
        RECT 47.385 31.240 47.470 31.365 ;
        RECT 48.090 31.240 48.175 31.400 ;
        RECT 50.285 31.365 50.335 31.400 ;
        POLYGON 50.335 31.400 50.370 31.365 50.335 31.365 ;
        RECT 50.285 31.240 50.370 31.365 ;
        RECT 50.990 31.240 51.075 31.400 ;
        RECT 53.185 31.365 53.235 31.400 ;
        POLYGON 53.235 31.400 53.270 31.365 53.235 31.365 ;
        RECT 53.185 31.240 53.270 31.365 ;
        RECT 53.890 31.240 53.975 31.400 ;
        RECT 56.085 31.365 56.135 31.400 ;
        POLYGON 56.135 31.400 56.170 31.365 56.135 31.365 ;
        RECT 56.085 31.240 56.170 31.365 ;
        RECT 56.790 31.240 56.875 31.400 ;
        RECT 58.985 31.365 59.035 31.400 ;
        POLYGON 59.035 31.400 59.070 31.365 59.035 31.365 ;
        RECT 58.985 31.240 59.070 31.365 ;
        RECT 59.690 31.240 59.775 31.400 ;
        RECT 61.885 31.365 61.935 31.400 ;
        POLYGON 61.935 31.400 61.970 31.365 61.935 31.365 ;
        RECT 61.885 31.240 61.970 31.365 ;
        RECT 62.590 31.240 62.675 31.400 ;
        RECT 64.785 31.365 64.835 31.400 ;
        POLYGON 64.835 31.400 64.870 31.365 64.835 31.365 ;
        RECT 64.785 31.240 64.870 31.365 ;
        RECT 65.490 31.240 65.575 31.400 ;
        RECT 67.685 31.365 67.735 31.400 ;
        POLYGON 67.735 31.400 67.770 31.365 67.735 31.365 ;
        RECT 67.685 31.240 67.770 31.365 ;
        RECT 68.390 31.240 68.475 31.400 ;
        RECT 70.585 31.365 70.635 31.400 ;
        POLYGON 70.635 31.400 70.670 31.365 70.635 31.365 ;
        RECT 70.585 31.240 70.670 31.365 ;
        RECT 71.290 31.240 71.375 31.400 ;
        RECT 73.485 31.365 73.535 31.400 ;
        POLYGON 73.535 31.400 73.570 31.365 73.535 31.365 ;
        RECT 73.485 31.240 73.570 31.365 ;
        RECT 74.190 31.240 74.275 31.400 ;
        RECT 76.385 31.365 76.435 31.400 ;
        POLYGON 76.435 31.400 76.470 31.365 76.435 31.365 ;
        RECT 76.385 31.240 76.470 31.365 ;
        RECT 77.090 31.240 77.175 31.400 ;
        RECT 79.285 31.365 79.335 31.400 ;
        POLYGON 79.335 31.400 79.370 31.365 79.335 31.365 ;
        RECT 79.285 31.240 79.370 31.365 ;
        RECT 79.990 31.240 80.075 31.400 ;
        RECT 82.185 31.365 82.235 31.400 ;
        POLYGON 82.235 31.400 82.270 31.365 82.235 31.365 ;
        RECT 82.185 31.240 82.270 31.365 ;
        RECT 82.890 31.240 82.975 31.400 ;
        RECT 85.085 31.365 85.135 31.400 ;
        POLYGON 85.135 31.400 85.170 31.365 85.135 31.365 ;
        RECT 85.085 31.240 85.170 31.365 ;
        RECT 85.790 31.240 85.875 31.400 ;
        RECT 87.985 31.365 88.035 31.400 ;
        POLYGON 88.035 31.400 88.070 31.365 88.035 31.365 ;
        RECT 87.985 31.240 88.070 31.365 ;
        RECT 88.690 31.240 88.775 31.400 ;
        RECT 90.885 31.365 90.935 31.400 ;
        POLYGON 90.935 31.400 90.970 31.365 90.935 31.365 ;
        RECT 90.885 31.240 90.970 31.365 ;
        RECT 91.590 31.240 91.675 31.400 ;
        RECT 0.775 30.620 0.850 30.760 ;
        RECT 0.990 30.570 1.065 30.710 ;
        RECT 1.695 30.630 1.755 30.710 ;
        POLYGON 1.695 30.630 1.755 30.630 1.755 30.570 ;
        RECT 1.910 30.620 1.985 30.760 ;
        RECT 3.675 30.620 3.750 30.760 ;
        RECT 3.890 30.570 3.965 30.710 ;
        RECT 4.595 30.630 4.655 30.710 ;
        POLYGON 4.595 30.630 4.655 30.630 4.655 30.570 ;
        RECT 4.810 30.620 4.885 30.760 ;
        RECT 6.575 30.620 6.650 30.760 ;
        RECT 6.790 30.570 6.865 30.710 ;
        RECT 7.495 30.630 7.555 30.710 ;
        POLYGON 7.495 30.630 7.555 30.630 7.555 30.570 ;
        RECT 7.710 30.620 7.785 30.760 ;
        RECT 9.475 30.620 9.550 30.760 ;
        RECT 9.690 30.570 9.765 30.710 ;
        RECT 10.395 30.630 10.455 30.710 ;
        POLYGON 10.395 30.630 10.455 30.630 10.455 30.570 ;
        RECT 10.610 30.620 10.685 30.760 ;
        RECT 12.375 30.620 12.450 30.760 ;
        RECT 12.590 30.570 12.665 30.710 ;
        RECT 13.295 30.630 13.355 30.710 ;
        POLYGON 13.295 30.630 13.355 30.630 13.355 30.570 ;
        RECT 13.510 30.620 13.585 30.760 ;
        RECT 15.275 30.620 15.350 30.760 ;
        RECT 15.490 30.570 15.565 30.710 ;
        RECT 16.195 30.630 16.255 30.710 ;
        POLYGON 16.195 30.630 16.255 30.630 16.255 30.570 ;
        RECT 16.410 30.620 16.485 30.760 ;
        RECT 18.175 30.620 18.250 30.760 ;
        RECT 18.390 30.570 18.465 30.710 ;
        RECT 19.095 30.630 19.155 30.710 ;
        POLYGON 19.095 30.630 19.155 30.630 19.155 30.570 ;
        RECT 19.310 30.620 19.385 30.760 ;
        RECT 21.075 30.620 21.150 30.760 ;
        RECT 21.290 30.570 21.365 30.710 ;
        RECT 21.995 30.630 22.055 30.710 ;
        POLYGON 21.995 30.630 22.055 30.630 22.055 30.570 ;
        RECT 22.210 30.620 22.285 30.760 ;
        RECT 23.975 30.620 24.050 30.760 ;
        RECT 24.190 30.570 24.265 30.710 ;
        RECT 24.895 30.630 24.955 30.710 ;
        POLYGON 24.895 30.630 24.955 30.630 24.955 30.570 ;
        RECT 25.110 30.620 25.185 30.760 ;
        RECT 26.875 30.620 26.950 30.760 ;
        RECT 27.090 30.570 27.165 30.710 ;
        RECT 27.795 30.630 27.855 30.710 ;
        POLYGON 27.795 30.630 27.855 30.630 27.855 30.570 ;
        RECT 28.010 30.620 28.085 30.760 ;
        RECT 29.775 30.620 29.850 30.760 ;
        RECT 29.990 30.570 30.065 30.710 ;
        RECT 30.695 30.630 30.755 30.710 ;
        POLYGON 30.695 30.630 30.755 30.630 30.755 30.570 ;
        RECT 30.910 30.620 30.985 30.760 ;
        RECT 32.675 30.620 32.750 30.760 ;
        RECT 32.890 30.570 32.965 30.710 ;
        RECT 33.595 30.630 33.655 30.710 ;
        POLYGON 33.595 30.630 33.655 30.630 33.655 30.570 ;
        RECT 33.810 30.620 33.885 30.760 ;
        RECT 35.575 30.620 35.650 30.760 ;
        RECT 35.790 30.570 35.865 30.710 ;
        RECT 36.495 30.630 36.555 30.710 ;
        POLYGON 36.495 30.630 36.555 30.630 36.555 30.570 ;
        RECT 36.710 30.620 36.785 30.760 ;
        RECT 38.475 30.620 38.550 30.760 ;
        RECT 38.690 30.570 38.765 30.710 ;
        RECT 39.395 30.630 39.455 30.710 ;
        POLYGON 39.395 30.630 39.455 30.630 39.455 30.570 ;
        RECT 39.610 30.620 39.685 30.760 ;
        RECT 41.375 30.620 41.450 30.760 ;
        RECT 41.590 30.570 41.665 30.710 ;
        RECT 42.295 30.630 42.355 30.710 ;
        POLYGON 42.295 30.630 42.355 30.630 42.355 30.570 ;
        RECT 42.510 30.620 42.585 30.760 ;
        RECT 44.275 30.620 44.350 30.760 ;
        RECT 44.490 30.570 44.565 30.710 ;
        RECT 45.195 30.630 45.255 30.710 ;
        POLYGON 45.195 30.630 45.255 30.630 45.255 30.570 ;
        RECT 45.410 30.620 45.485 30.760 ;
        RECT 47.175 30.620 47.250 30.760 ;
        RECT 47.390 30.570 47.465 30.710 ;
        RECT 48.095 30.630 48.155 30.710 ;
        POLYGON 48.095 30.630 48.155 30.630 48.155 30.570 ;
        RECT 48.310 30.620 48.385 30.760 ;
        RECT 50.075 30.620 50.150 30.760 ;
        RECT 50.290 30.570 50.365 30.710 ;
        RECT 50.995 30.630 51.055 30.710 ;
        POLYGON 50.995 30.630 51.055 30.630 51.055 30.570 ;
        RECT 51.210 30.620 51.285 30.760 ;
        RECT 52.975 30.620 53.050 30.760 ;
        RECT 53.190 30.570 53.265 30.710 ;
        RECT 53.895 30.630 53.955 30.710 ;
        POLYGON 53.895 30.630 53.955 30.630 53.955 30.570 ;
        RECT 54.110 30.620 54.185 30.760 ;
        RECT 55.875 30.620 55.950 30.760 ;
        RECT 56.090 30.570 56.165 30.710 ;
        RECT 56.795 30.630 56.855 30.710 ;
        POLYGON 56.795 30.630 56.855 30.630 56.855 30.570 ;
        RECT 57.010 30.620 57.085 30.760 ;
        RECT 58.775 30.620 58.850 30.760 ;
        RECT 58.990 30.570 59.065 30.710 ;
        RECT 59.695 30.630 59.755 30.710 ;
        POLYGON 59.695 30.630 59.755 30.630 59.755 30.570 ;
        RECT 59.910 30.620 59.985 30.760 ;
        RECT 61.675 30.620 61.750 30.760 ;
        RECT 61.890 30.570 61.965 30.710 ;
        RECT 62.595 30.630 62.655 30.710 ;
        POLYGON 62.595 30.630 62.655 30.630 62.655 30.570 ;
        RECT 62.810 30.620 62.885 30.760 ;
        RECT 64.575 30.620 64.650 30.760 ;
        RECT 64.790 30.570 64.865 30.710 ;
        RECT 65.495 30.630 65.555 30.710 ;
        POLYGON 65.495 30.630 65.555 30.630 65.555 30.570 ;
        RECT 65.710 30.620 65.785 30.760 ;
        RECT 67.475 30.620 67.550 30.760 ;
        RECT 67.690 30.570 67.765 30.710 ;
        RECT 68.395 30.630 68.455 30.710 ;
        POLYGON 68.395 30.630 68.455 30.630 68.455 30.570 ;
        RECT 68.610 30.620 68.685 30.760 ;
        RECT 70.375 30.620 70.450 30.760 ;
        RECT 70.590 30.570 70.665 30.710 ;
        RECT 71.295 30.630 71.355 30.710 ;
        POLYGON 71.295 30.630 71.355 30.630 71.355 30.570 ;
        RECT 71.510 30.620 71.585 30.760 ;
        RECT 73.275 30.620 73.350 30.760 ;
        RECT 73.490 30.570 73.565 30.710 ;
        RECT 74.195 30.630 74.255 30.710 ;
        POLYGON 74.195 30.630 74.255 30.630 74.255 30.570 ;
        RECT 74.410 30.620 74.485 30.760 ;
        RECT 76.175 30.620 76.250 30.760 ;
        RECT 76.390 30.570 76.465 30.710 ;
        RECT 77.095 30.630 77.155 30.710 ;
        POLYGON 77.095 30.630 77.155 30.630 77.155 30.570 ;
        RECT 77.310 30.620 77.385 30.760 ;
        RECT 79.075 30.620 79.150 30.760 ;
        RECT 79.290 30.570 79.365 30.710 ;
        RECT 79.995 30.630 80.055 30.710 ;
        POLYGON 79.995 30.630 80.055 30.630 80.055 30.570 ;
        RECT 80.210 30.620 80.285 30.760 ;
        RECT 81.975 30.620 82.050 30.760 ;
        RECT 82.190 30.570 82.265 30.710 ;
        RECT 82.895 30.630 82.955 30.710 ;
        POLYGON 82.895 30.630 82.955 30.630 82.955 30.570 ;
        RECT 83.110 30.620 83.185 30.760 ;
        RECT 84.875 30.620 84.950 30.760 ;
        RECT 85.090 30.570 85.165 30.710 ;
        RECT 85.795 30.630 85.855 30.710 ;
        POLYGON 85.795 30.630 85.855 30.630 85.855 30.570 ;
        RECT 86.010 30.620 86.085 30.760 ;
        RECT 87.775 30.620 87.850 30.760 ;
        RECT 87.990 30.570 88.065 30.710 ;
        RECT 88.695 30.630 88.755 30.710 ;
        POLYGON 88.695 30.630 88.755 30.630 88.755 30.570 ;
        RECT 88.910 30.620 88.985 30.760 ;
        RECT 90.675 30.620 90.750 30.760 ;
        RECT 90.890 30.570 90.965 30.710 ;
        RECT 91.595 30.630 91.655 30.710 ;
        POLYGON 91.595 30.630 91.655 30.630 91.655 30.570 ;
        RECT 91.810 30.620 91.885 30.760 ;
        RECT 0.720 30.100 0.870 30.270 ;
        RECT 1.110 30.235 1.260 30.405 ;
        RECT 1.500 30.235 1.650 30.405 ;
        RECT 1.890 30.100 2.040 30.270 ;
        RECT 3.620 30.100 3.770 30.270 ;
        RECT 4.010 30.235 4.160 30.405 ;
        RECT 4.400 30.235 4.550 30.405 ;
        RECT 4.790 30.100 4.940 30.270 ;
        RECT 6.520 30.100 6.670 30.270 ;
        RECT 6.910 30.235 7.060 30.405 ;
        RECT 7.300 30.235 7.450 30.405 ;
        RECT 7.690 30.100 7.840 30.270 ;
        RECT 9.420 30.100 9.570 30.270 ;
        RECT 9.810 30.235 9.960 30.405 ;
        RECT 10.200 30.235 10.350 30.405 ;
        RECT 10.590 30.100 10.740 30.270 ;
        RECT 12.320 30.100 12.470 30.270 ;
        RECT 12.710 30.235 12.860 30.405 ;
        RECT 13.100 30.235 13.250 30.405 ;
        RECT 13.490 30.100 13.640 30.270 ;
        RECT 15.220 30.100 15.370 30.270 ;
        RECT 15.610 30.235 15.760 30.405 ;
        RECT 16.000 30.235 16.150 30.405 ;
        RECT 16.390 30.100 16.540 30.270 ;
        RECT 18.120 30.100 18.270 30.270 ;
        RECT 18.510 30.235 18.660 30.405 ;
        RECT 18.900 30.235 19.050 30.405 ;
        RECT 19.290 30.100 19.440 30.270 ;
        RECT 21.020 30.100 21.170 30.270 ;
        RECT 21.410 30.235 21.560 30.405 ;
        RECT 21.800 30.235 21.950 30.405 ;
        RECT 22.190 30.100 22.340 30.270 ;
        RECT 23.920 30.100 24.070 30.270 ;
        RECT 24.310 30.235 24.460 30.405 ;
        RECT 24.700 30.235 24.850 30.405 ;
        RECT 25.090 30.100 25.240 30.270 ;
        RECT 26.820 30.100 26.970 30.270 ;
        RECT 27.210 30.235 27.360 30.405 ;
        RECT 27.600 30.235 27.750 30.405 ;
        RECT 27.990 30.100 28.140 30.270 ;
        RECT 29.720 30.100 29.870 30.270 ;
        RECT 30.110 30.235 30.260 30.405 ;
        RECT 30.500 30.235 30.650 30.405 ;
        RECT 30.890 30.100 31.040 30.270 ;
        RECT 32.620 30.100 32.770 30.270 ;
        RECT 33.010 30.235 33.160 30.405 ;
        RECT 33.400 30.235 33.550 30.405 ;
        RECT 33.790 30.100 33.940 30.270 ;
        RECT 35.520 30.100 35.670 30.270 ;
        RECT 35.910 30.235 36.060 30.405 ;
        RECT 36.300 30.235 36.450 30.405 ;
        RECT 36.690 30.100 36.840 30.270 ;
        RECT 38.420 30.100 38.570 30.270 ;
        RECT 38.810 30.235 38.960 30.405 ;
        RECT 39.200 30.235 39.350 30.405 ;
        RECT 39.590 30.100 39.740 30.270 ;
        RECT 41.320 30.100 41.470 30.270 ;
        RECT 41.710 30.235 41.860 30.405 ;
        RECT 42.100 30.235 42.250 30.405 ;
        RECT 42.490 30.100 42.640 30.270 ;
        RECT 44.220 30.100 44.370 30.270 ;
        RECT 44.610 30.235 44.760 30.405 ;
        RECT 45.000 30.235 45.150 30.405 ;
        RECT 45.390 30.100 45.540 30.270 ;
        RECT 47.120 30.100 47.270 30.270 ;
        RECT 47.510 30.235 47.660 30.405 ;
        RECT 47.900 30.235 48.050 30.405 ;
        RECT 48.290 30.100 48.440 30.270 ;
        RECT 50.020 30.100 50.170 30.270 ;
        RECT 50.410 30.235 50.560 30.405 ;
        RECT 50.800 30.235 50.950 30.405 ;
        RECT 51.190 30.100 51.340 30.270 ;
        RECT 52.920 30.100 53.070 30.270 ;
        RECT 53.310 30.235 53.460 30.405 ;
        RECT 53.700 30.235 53.850 30.405 ;
        RECT 54.090 30.100 54.240 30.270 ;
        RECT 55.820 30.100 55.970 30.270 ;
        RECT 56.210 30.235 56.360 30.405 ;
        RECT 56.600 30.235 56.750 30.405 ;
        RECT 56.990 30.100 57.140 30.270 ;
        RECT 58.720 30.100 58.870 30.270 ;
        RECT 59.110 30.235 59.260 30.405 ;
        RECT 59.500 30.235 59.650 30.405 ;
        RECT 59.890 30.100 60.040 30.270 ;
        RECT 61.620 30.100 61.770 30.270 ;
        RECT 62.010 30.235 62.160 30.405 ;
        RECT 62.400 30.235 62.550 30.405 ;
        RECT 62.790 30.100 62.940 30.270 ;
        RECT 64.520 30.100 64.670 30.270 ;
        RECT 64.910 30.235 65.060 30.405 ;
        RECT 65.300 30.235 65.450 30.405 ;
        RECT 65.690 30.100 65.840 30.270 ;
        RECT 67.420 30.100 67.570 30.270 ;
        RECT 67.810 30.235 67.960 30.405 ;
        RECT 68.200 30.235 68.350 30.405 ;
        RECT 68.590 30.100 68.740 30.270 ;
        RECT 70.320 30.100 70.470 30.270 ;
        RECT 70.710 30.235 70.860 30.405 ;
        RECT 71.100 30.235 71.250 30.405 ;
        RECT 71.490 30.100 71.640 30.270 ;
        RECT 73.220 30.100 73.370 30.270 ;
        RECT 73.610 30.235 73.760 30.405 ;
        RECT 74.000 30.235 74.150 30.405 ;
        RECT 74.390 30.100 74.540 30.270 ;
        RECT 76.120 30.100 76.270 30.270 ;
        RECT 76.510 30.235 76.660 30.405 ;
        RECT 76.900 30.235 77.050 30.405 ;
        RECT 77.290 30.100 77.440 30.270 ;
        RECT 79.020 30.100 79.170 30.270 ;
        RECT 79.410 30.235 79.560 30.405 ;
        RECT 79.800 30.235 79.950 30.405 ;
        RECT 80.190 30.100 80.340 30.270 ;
        RECT 81.920 30.100 82.070 30.270 ;
        RECT 82.310 30.235 82.460 30.405 ;
        RECT 82.700 30.235 82.850 30.405 ;
        RECT 83.090 30.100 83.240 30.270 ;
        RECT 84.820 30.100 84.970 30.270 ;
        RECT 85.210 30.235 85.360 30.405 ;
        RECT 85.600 30.235 85.750 30.405 ;
        RECT 85.990 30.100 86.140 30.270 ;
        RECT 87.720 30.100 87.870 30.270 ;
        RECT 88.110 30.235 88.260 30.405 ;
        RECT 88.500 30.235 88.650 30.405 ;
        RECT 88.890 30.100 89.040 30.270 ;
        RECT 90.620 30.100 90.770 30.270 ;
        RECT 91.010 30.235 91.160 30.405 ;
        RECT 91.400 30.235 91.550 30.405 ;
        RECT 91.790 30.100 91.940 30.270 ;
        RECT 0.985 30.015 1.035 30.050 ;
        POLYGON 1.035 30.050 1.070 30.015 1.035 30.015 ;
        RECT 0.985 29.890 1.070 30.015 ;
        RECT 1.690 29.890 1.775 30.050 ;
        RECT 3.885 30.015 3.935 30.050 ;
        POLYGON 3.935 30.050 3.970 30.015 3.935 30.015 ;
        RECT 3.885 29.890 3.970 30.015 ;
        RECT 4.590 29.890 4.675 30.050 ;
        RECT 6.785 30.015 6.835 30.050 ;
        POLYGON 6.835 30.050 6.870 30.015 6.835 30.015 ;
        RECT 6.785 29.890 6.870 30.015 ;
        RECT 7.490 29.890 7.575 30.050 ;
        RECT 9.685 30.015 9.735 30.050 ;
        POLYGON 9.735 30.050 9.770 30.015 9.735 30.015 ;
        RECT 9.685 29.890 9.770 30.015 ;
        RECT 10.390 29.890 10.475 30.050 ;
        RECT 12.585 30.015 12.635 30.050 ;
        POLYGON 12.635 30.050 12.670 30.015 12.635 30.015 ;
        RECT 12.585 29.890 12.670 30.015 ;
        RECT 13.290 29.890 13.375 30.050 ;
        RECT 15.485 30.015 15.535 30.050 ;
        POLYGON 15.535 30.050 15.570 30.015 15.535 30.015 ;
        RECT 15.485 29.890 15.570 30.015 ;
        RECT 16.190 29.890 16.275 30.050 ;
        RECT 18.385 30.015 18.435 30.050 ;
        POLYGON 18.435 30.050 18.470 30.015 18.435 30.015 ;
        RECT 18.385 29.890 18.470 30.015 ;
        RECT 19.090 29.890 19.175 30.050 ;
        RECT 21.285 30.015 21.335 30.050 ;
        POLYGON 21.335 30.050 21.370 30.015 21.335 30.015 ;
        RECT 21.285 29.890 21.370 30.015 ;
        RECT 21.990 29.890 22.075 30.050 ;
        RECT 24.185 30.015 24.235 30.050 ;
        POLYGON 24.235 30.050 24.270 30.015 24.235 30.015 ;
        RECT 24.185 29.890 24.270 30.015 ;
        RECT 24.890 29.890 24.975 30.050 ;
        RECT 27.085 30.015 27.135 30.050 ;
        POLYGON 27.135 30.050 27.170 30.015 27.135 30.015 ;
        RECT 27.085 29.890 27.170 30.015 ;
        RECT 27.790 29.890 27.875 30.050 ;
        RECT 29.985 30.015 30.035 30.050 ;
        POLYGON 30.035 30.050 30.070 30.015 30.035 30.015 ;
        RECT 29.985 29.890 30.070 30.015 ;
        RECT 30.690 29.890 30.775 30.050 ;
        RECT 32.885 30.015 32.935 30.050 ;
        POLYGON 32.935 30.050 32.970 30.015 32.935 30.015 ;
        RECT 32.885 29.890 32.970 30.015 ;
        RECT 33.590 29.890 33.675 30.050 ;
        RECT 35.785 30.015 35.835 30.050 ;
        POLYGON 35.835 30.050 35.870 30.015 35.835 30.015 ;
        RECT 35.785 29.890 35.870 30.015 ;
        RECT 36.490 29.890 36.575 30.050 ;
        RECT 38.685 30.015 38.735 30.050 ;
        POLYGON 38.735 30.050 38.770 30.015 38.735 30.015 ;
        RECT 38.685 29.890 38.770 30.015 ;
        RECT 39.390 29.890 39.475 30.050 ;
        RECT 41.585 30.015 41.635 30.050 ;
        POLYGON 41.635 30.050 41.670 30.015 41.635 30.015 ;
        RECT 41.585 29.890 41.670 30.015 ;
        RECT 42.290 29.890 42.375 30.050 ;
        RECT 44.485 30.015 44.535 30.050 ;
        POLYGON 44.535 30.050 44.570 30.015 44.535 30.015 ;
        RECT 44.485 29.890 44.570 30.015 ;
        RECT 45.190 29.890 45.275 30.050 ;
        RECT 47.385 30.015 47.435 30.050 ;
        POLYGON 47.435 30.050 47.470 30.015 47.435 30.015 ;
        RECT 47.385 29.890 47.470 30.015 ;
        RECT 48.090 29.890 48.175 30.050 ;
        RECT 50.285 30.015 50.335 30.050 ;
        POLYGON 50.335 30.050 50.370 30.015 50.335 30.015 ;
        RECT 50.285 29.890 50.370 30.015 ;
        RECT 50.990 29.890 51.075 30.050 ;
        RECT 53.185 30.015 53.235 30.050 ;
        POLYGON 53.235 30.050 53.270 30.015 53.235 30.015 ;
        RECT 53.185 29.890 53.270 30.015 ;
        RECT 53.890 29.890 53.975 30.050 ;
        RECT 56.085 30.015 56.135 30.050 ;
        POLYGON 56.135 30.050 56.170 30.015 56.135 30.015 ;
        RECT 56.085 29.890 56.170 30.015 ;
        RECT 56.790 29.890 56.875 30.050 ;
        RECT 58.985 30.015 59.035 30.050 ;
        POLYGON 59.035 30.050 59.070 30.015 59.035 30.015 ;
        RECT 58.985 29.890 59.070 30.015 ;
        RECT 59.690 29.890 59.775 30.050 ;
        RECT 61.885 30.015 61.935 30.050 ;
        POLYGON 61.935 30.050 61.970 30.015 61.935 30.015 ;
        RECT 61.885 29.890 61.970 30.015 ;
        RECT 62.590 29.890 62.675 30.050 ;
        RECT 64.785 30.015 64.835 30.050 ;
        POLYGON 64.835 30.050 64.870 30.015 64.835 30.015 ;
        RECT 64.785 29.890 64.870 30.015 ;
        RECT 65.490 29.890 65.575 30.050 ;
        RECT 67.685 30.015 67.735 30.050 ;
        POLYGON 67.735 30.050 67.770 30.015 67.735 30.015 ;
        RECT 67.685 29.890 67.770 30.015 ;
        RECT 68.390 29.890 68.475 30.050 ;
        RECT 70.585 30.015 70.635 30.050 ;
        POLYGON 70.635 30.050 70.670 30.015 70.635 30.015 ;
        RECT 70.585 29.890 70.670 30.015 ;
        RECT 71.290 29.890 71.375 30.050 ;
        RECT 73.485 30.015 73.535 30.050 ;
        POLYGON 73.535 30.050 73.570 30.015 73.535 30.015 ;
        RECT 73.485 29.890 73.570 30.015 ;
        RECT 74.190 29.890 74.275 30.050 ;
        RECT 76.385 30.015 76.435 30.050 ;
        POLYGON 76.435 30.050 76.470 30.015 76.435 30.015 ;
        RECT 76.385 29.890 76.470 30.015 ;
        RECT 77.090 29.890 77.175 30.050 ;
        RECT 79.285 30.015 79.335 30.050 ;
        POLYGON 79.335 30.050 79.370 30.015 79.335 30.015 ;
        RECT 79.285 29.890 79.370 30.015 ;
        RECT 79.990 29.890 80.075 30.050 ;
        RECT 82.185 30.015 82.235 30.050 ;
        POLYGON 82.235 30.050 82.270 30.015 82.235 30.015 ;
        RECT 82.185 29.890 82.270 30.015 ;
        RECT 82.890 29.890 82.975 30.050 ;
        RECT 85.085 30.015 85.135 30.050 ;
        POLYGON 85.135 30.050 85.170 30.015 85.135 30.015 ;
        RECT 85.085 29.890 85.170 30.015 ;
        RECT 85.790 29.890 85.875 30.050 ;
        RECT 87.985 30.015 88.035 30.050 ;
        POLYGON 88.035 30.050 88.070 30.015 88.035 30.015 ;
        RECT 87.985 29.890 88.070 30.015 ;
        RECT 88.690 29.890 88.775 30.050 ;
        RECT 90.885 30.015 90.935 30.050 ;
        POLYGON 90.935 30.050 90.970 30.015 90.935 30.015 ;
        RECT 90.885 29.890 90.970 30.015 ;
        RECT 91.590 29.890 91.675 30.050 ;
        RECT 0.775 29.270 0.850 29.410 ;
        RECT 0.990 29.220 1.065 29.360 ;
        RECT 1.695 29.280 1.755 29.360 ;
        POLYGON 1.695 29.280 1.755 29.280 1.755 29.220 ;
        RECT 1.910 29.270 1.985 29.410 ;
        RECT 3.675 29.270 3.750 29.410 ;
        RECT 3.890 29.220 3.965 29.360 ;
        RECT 4.595 29.280 4.655 29.360 ;
        POLYGON 4.595 29.280 4.655 29.280 4.655 29.220 ;
        RECT 4.810 29.270 4.885 29.410 ;
        RECT 6.575 29.270 6.650 29.410 ;
        RECT 6.790 29.220 6.865 29.360 ;
        RECT 7.495 29.280 7.555 29.360 ;
        POLYGON 7.495 29.280 7.555 29.280 7.555 29.220 ;
        RECT 7.710 29.270 7.785 29.410 ;
        RECT 9.475 29.270 9.550 29.410 ;
        RECT 9.690 29.220 9.765 29.360 ;
        RECT 10.395 29.280 10.455 29.360 ;
        POLYGON 10.395 29.280 10.455 29.280 10.455 29.220 ;
        RECT 10.610 29.270 10.685 29.410 ;
        RECT 12.375 29.270 12.450 29.410 ;
        RECT 12.590 29.220 12.665 29.360 ;
        RECT 13.295 29.280 13.355 29.360 ;
        POLYGON 13.295 29.280 13.355 29.280 13.355 29.220 ;
        RECT 13.510 29.270 13.585 29.410 ;
        RECT 15.275 29.270 15.350 29.410 ;
        RECT 15.490 29.220 15.565 29.360 ;
        RECT 16.195 29.280 16.255 29.360 ;
        POLYGON 16.195 29.280 16.255 29.280 16.255 29.220 ;
        RECT 16.410 29.270 16.485 29.410 ;
        RECT 18.175 29.270 18.250 29.410 ;
        RECT 18.390 29.220 18.465 29.360 ;
        RECT 19.095 29.280 19.155 29.360 ;
        POLYGON 19.095 29.280 19.155 29.280 19.155 29.220 ;
        RECT 19.310 29.270 19.385 29.410 ;
        RECT 21.075 29.270 21.150 29.410 ;
        RECT 21.290 29.220 21.365 29.360 ;
        RECT 21.995 29.280 22.055 29.360 ;
        POLYGON 21.995 29.280 22.055 29.280 22.055 29.220 ;
        RECT 22.210 29.270 22.285 29.410 ;
        RECT 23.975 29.270 24.050 29.410 ;
        RECT 24.190 29.220 24.265 29.360 ;
        RECT 24.895 29.280 24.955 29.360 ;
        POLYGON 24.895 29.280 24.955 29.280 24.955 29.220 ;
        RECT 25.110 29.270 25.185 29.410 ;
        RECT 26.875 29.270 26.950 29.410 ;
        RECT 27.090 29.220 27.165 29.360 ;
        RECT 27.795 29.280 27.855 29.360 ;
        POLYGON 27.795 29.280 27.855 29.280 27.855 29.220 ;
        RECT 28.010 29.270 28.085 29.410 ;
        RECT 29.775 29.270 29.850 29.410 ;
        RECT 29.990 29.220 30.065 29.360 ;
        RECT 30.695 29.280 30.755 29.360 ;
        POLYGON 30.695 29.280 30.755 29.280 30.755 29.220 ;
        RECT 30.910 29.270 30.985 29.410 ;
        RECT 32.675 29.270 32.750 29.410 ;
        RECT 32.890 29.220 32.965 29.360 ;
        RECT 33.595 29.280 33.655 29.360 ;
        POLYGON 33.595 29.280 33.655 29.280 33.655 29.220 ;
        RECT 33.810 29.270 33.885 29.410 ;
        RECT 35.575 29.270 35.650 29.410 ;
        RECT 35.790 29.220 35.865 29.360 ;
        RECT 36.495 29.280 36.555 29.360 ;
        POLYGON 36.495 29.280 36.555 29.280 36.555 29.220 ;
        RECT 36.710 29.270 36.785 29.410 ;
        RECT 38.475 29.270 38.550 29.410 ;
        RECT 38.690 29.220 38.765 29.360 ;
        RECT 39.395 29.280 39.455 29.360 ;
        POLYGON 39.395 29.280 39.455 29.280 39.455 29.220 ;
        RECT 39.610 29.270 39.685 29.410 ;
        RECT 41.375 29.270 41.450 29.410 ;
        RECT 41.590 29.220 41.665 29.360 ;
        RECT 42.295 29.280 42.355 29.360 ;
        POLYGON 42.295 29.280 42.355 29.280 42.355 29.220 ;
        RECT 42.510 29.270 42.585 29.410 ;
        RECT 44.275 29.270 44.350 29.410 ;
        RECT 44.490 29.220 44.565 29.360 ;
        RECT 45.195 29.280 45.255 29.360 ;
        POLYGON 45.195 29.280 45.255 29.280 45.255 29.220 ;
        RECT 45.410 29.270 45.485 29.410 ;
        RECT 47.175 29.270 47.250 29.410 ;
        RECT 47.390 29.220 47.465 29.360 ;
        RECT 48.095 29.280 48.155 29.360 ;
        POLYGON 48.095 29.280 48.155 29.280 48.155 29.220 ;
        RECT 48.310 29.270 48.385 29.410 ;
        RECT 50.075 29.270 50.150 29.410 ;
        RECT 50.290 29.220 50.365 29.360 ;
        RECT 50.995 29.280 51.055 29.360 ;
        POLYGON 50.995 29.280 51.055 29.280 51.055 29.220 ;
        RECT 51.210 29.270 51.285 29.410 ;
        RECT 52.975 29.270 53.050 29.410 ;
        RECT 53.190 29.220 53.265 29.360 ;
        RECT 53.895 29.280 53.955 29.360 ;
        POLYGON 53.895 29.280 53.955 29.280 53.955 29.220 ;
        RECT 54.110 29.270 54.185 29.410 ;
        RECT 55.875 29.270 55.950 29.410 ;
        RECT 56.090 29.220 56.165 29.360 ;
        RECT 56.795 29.280 56.855 29.360 ;
        POLYGON 56.795 29.280 56.855 29.280 56.855 29.220 ;
        RECT 57.010 29.270 57.085 29.410 ;
        RECT 58.775 29.270 58.850 29.410 ;
        RECT 58.990 29.220 59.065 29.360 ;
        RECT 59.695 29.280 59.755 29.360 ;
        POLYGON 59.695 29.280 59.755 29.280 59.755 29.220 ;
        RECT 59.910 29.270 59.985 29.410 ;
        RECT 61.675 29.270 61.750 29.410 ;
        RECT 61.890 29.220 61.965 29.360 ;
        RECT 62.595 29.280 62.655 29.360 ;
        POLYGON 62.595 29.280 62.655 29.280 62.655 29.220 ;
        RECT 62.810 29.270 62.885 29.410 ;
        RECT 64.575 29.270 64.650 29.410 ;
        RECT 64.790 29.220 64.865 29.360 ;
        RECT 65.495 29.280 65.555 29.360 ;
        POLYGON 65.495 29.280 65.555 29.280 65.555 29.220 ;
        RECT 65.710 29.270 65.785 29.410 ;
        RECT 67.475 29.270 67.550 29.410 ;
        RECT 67.690 29.220 67.765 29.360 ;
        RECT 68.395 29.280 68.455 29.360 ;
        POLYGON 68.395 29.280 68.455 29.280 68.455 29.220 ;
        RECT 68.610 29.270 68.685 29.410 ;
        RECT 70.375 29.270 70.450 29.410 ;
        RECT 70.590 29.220 70.665 29.360 ;
        RECT 71.295 29.280 71.355 29.360 ;
        POLYGON 71.295 29.280 71.355 29.280 71.355 29.220 ;
        RECT 71.510 29.270 71.585 29.410 ;
        RECT 73.275 29.270 73.350 29.410 ;
        RECT 73.490 29.220 73.565 29.360 ;
        RECT 74.195 29.280 74.255 29.360 ;
        POLYGON 74.195 29.280 74.255 29.280 74.255 29.220 ;
        RECT 74.410 29.270 74.485 29.410 ;
        RECT 76.175 29.270 76.250 29.410 ;
        RECT 76.390 29.220 76.465 29.360 ;
        RECT 77.095 29.280 77.155 29.360 ;
        POLYGON 77.095 29.280 77.155 29.280 77.155 29.220 ;
        RECT 77.310 29.270 77.385 29.410 ;
        RECT 79.075 29.270 79.150 29.410 ;
        RECT 79.290 29.220 79.365 29.360 ;
        RECT 79.995 29.280 80.055 29.360 ;
        POLYGON 79.995 29.280 80.055 29.280 80.055 29.220 ;
        RECT 80.210 29.270 80.285 29.410 ;
        RECT 81.975 29.270 82.050 29.410 ;
        RECT 82.190 29.220 82.265 29.360 ;
        RECT 82.895 29.280 82.955 29.360 ;
        POLYGON 82.895 29.280 82.955 29.280 82.955 29.220 ;
        RECT 83.110 29.270 83.185 29.410 ;
        RECT 84.875 29.270 84.950 29.410 ;
        RECT 85.090 29.220 85.165 29.360 ;
        RECT 85.795 29.280 85.855 29.360 ;
        POLYGON 85.795 29.280 85.855 29.280 85.855 29.220 ;
        RECT 86.010 29.270 86.085 29.410 ;
        RECT 87.775 29.270 87.850 29.410 ;
        RECT 87.990 29.220 88.065 29.360 ;
        RECT 88.695 29.280 88.755 29.360 ;
        POLYGON 88.695 29.280 88.755 29.280 88.755 29.220 ;
        RECT 88.910 29.270 88.985 29.410 ;
        RECT 90.675 29.270 90.750 29.410 ;
        RECT 90.890 29.220 90.965 29.360 ;
        RECT 91.595 29.280 91.655 29.360 ;
        POLYGON 91.595 29.280 91.655 29.280 91.655 29.220 ;
        RECT 91.810 29.270 91.885 29.410 ;
        RECT 0.720 28.750 0.870 28.920 ;
        RECT 1.110 28.885 1.260 29.055 ;
        RECT 1.500 28.885 1.650 29.055 ;
        RECT 1.890 28.750 2.040 28.920 ;
        RECT 3.620 28.750 3.770 28.920 ;
        RECT 4.010 28.885 4.160 29.055 ;
        RECT 4.400 28.885 4.550 29.055 ;
        RECT 4.790 28.750 4.940 28.920 ;
        RECT 6.520 28.750 6.670 28.920 ;
        RECT 6.910 28.885 7.060 29.055 ;
        RECT 7.300 28.885 7.450 29.055 ;
        RECT 7.690 28.750 7.840 28.920 ;
        RECT 9.420 28.750 9.570 28.920 ;
        RECT 9.810 28.885 9.960 29.055 ;
        RECT 10.200 28.885 10.350 29.055 ;
        RECT 10.590 28.750 10.740 28.920 ;
        RECT 12.320 28.750 12.470 28.920 ;
        RECT 12.710 28.885 12.860 29.055 ;
        RECT 13.100 28.885 13.250 29.055 ;
        RECT 13.490 28.750 13.640 28.920 ;
        RECT 15.220 28.750 15.370 28.920 ;
        RECT 15.610 28.885 15.760 29.055 ;
        RECT 16.000 28.885 16.150 29.055 ;
        RECT 16.390 28.750 16.540 28.920 ;
        RECT 18.120 28.750 18.270 28.920 ;
        RECT 18.510 28.885 18.660 29.055 ;
        RECT 18.900 28.885 19.050 29.055 ;
        RECT 19.290 28.750 19.440 28.920 ;
        RECT 21.020 28.750 21.170 28.920 ;
        RECT 21.410 28.885 21.560 29.055 ;
        RECT 21.800 28.885 21.950 29.055 ;
        RECT 22.190 28.750 22.340 28.920 ;
        RECT 23.920 28.750 24.070 28.920 ;
        RECT 24.310 28.885 24.460 29.055 ;
        RECT 24.700 28.885 24.850 29.055 ;
        RECT 25.090 28.750 25.240 28.920 ;
        RECT 26.820 28.750 26.970 28.920 ;
        RECT 27.210 28.885 27.360 29.055 ;
        RECT 27.600 28.885 27.750 29.055 ;
        RECT 27.990 28.750 28.140 28.920 ;
        RECT 29.720 28.750 29.870 28.920 ;
        RECT 30.110 28.885 30.260 29.055 ;
        RECT 30.500 28.885 30.650 29.055 ;
        RECT 30.890 28.750 31.040 28.920 ;
        RECT 32.620 28.750 32.770 28.920 ;
        RECT 33.010 28.885 33.160 29.055 ;
        RECT 33.400 28.885 33.550 29.055 ;
        RECT 33.790 28.750 33.940 28.920 ;
        RECT 35.520 28.750 35.670 28.920 ;
        RECT 35.910 28.885 36.060 29.055 ;
        RECT 36.300 28.885 36.450 29.055 ;
        RECT 36.690 28.750 36.840 28.920 ;
        RECT 38.420 28.750 38.570 28.920 ;
        RECT 38.810 28.885 38.960 29.055 ;
        RECT 39.200 28.885 39.350 29.055 ;
        RECT 39.590 28.750 39.740 28.920 ;
        RECT 41.320 28.750 41.470 28.920 ;
        RECT 41.710 28.885 41.860 29.055 ;
        RECT 42.100 28.885 42.250 29.055 ;
        RECT 42.490 28.750 42.640 28.920 ;
        RECT 44.220 28.750 44.370 28.920 ;
        RECT 44.610 28.885 44.760 29.055 ;
        RECT 45.000 28.885 45.150 29.055 ;
        RECT 45.390 28.750 45.540 28.920 ;
        RECT 47.120 28.750 47.270 28.920 ;
        RECT 47.510 28.885 47.660 29.055 ;
        RECT 47.900 28.885 48.050 29.055 ;
        RECT 48.290 28.750 48.440 28.920 ;
        RECT 50.020 28.750 50.170 28.920 ;
        RECT 50.410 28.885 50.560 29.055 ;
        RECT 50.800 28.885 50.950 29.055 ;
        RECT 51.190 28.750 51.340 28.920 ;
        RECT 52.920 28.750 53.070 28.920 ;
        RECT 53.310 28.885 53.460 29.055 ;
        RECT 53.700 28.885 53.850 29.055 ;
        RECT 54.090 28.750 54.240 28.920 ;
        RECT 55.820 28.750 55.970 28.920 ;
        RECT 56.210 28.885 56.360 29.055 ;
        RECT 56.600 28.885 56.750 29.055 ;
        RECT 56.990 28.750 57.140 28.920 ;
        RECT 58.720 28.750 58.870 28.920 ;
        RECT 59.110 28.885 59.260 29.055 ;
        RECT 59.500 28.885 59.650 29.055 ;
        RECT 59.890 28.750 60.040 28.920 ;
        RECT 61.620 28.750 61.770 28.920 ;
        RECT 62.010 28.885 62.160 29.055 ;
        RECT 62.400 28.885 62.550 29.055 ;
        RECT 62.790 28.750 62.940 28.920 ;
        RECT 64.520 28.750 64.670 28.920 ;
        RECT 64.910 28.885 65.060 29.055 ;
        RECT 65.300 28.885 65.450 29.055 ;
        RECT 65.690 28.750 65.840 28.920 ;
        RECT 67.420 28.750 67.570 28.920 ;
        RECT 67.810 28.885 67.960 29.055 ;
        RECT 68.200 28.885 68.350 29.055 ;
        RECT 68.590 28.750 68.740 28.920 ;
        RECT 70.320 28.750 70.470 28.920 ;
        RECT 70.710 28.885 70.860 29.055 ;
        RECT 71.100 28.885 71.250 29.055 ;
        RECT 71.490 28.750 71.640 28.920 ;
        RECT 73.220 28.750 73.370 28.920 ;
        RECT 73.610 28.885 73.760 29.055 ;
        RECT 74.000 28.885 74.150 29.055 ;
        RECT 74.390 28.750 74.540 28.920 ;
        RECT 76.120 28.750 76.270 28.920 ;
        RECT 76.510 28.885 76.660 29.055 ;
        RECT 76.900 28.885 77.050 29.055 ;
        RECT 77.290 28.750 77.440 28.920 ;
        RECT 79.020 28.750 79.170 28.920 ;
        RECT 79.410 28.885 79.560 29.055 ;
        RECT 79.800 28.885 79.950 29.055 ;
        RECT 80.190 28.750 80.340 28.920 ;
        RECT 81.920 28.750 82.070 28.920 ;
        RECT 82.310 28.885 82.460 29.055 ;
        RECT 82.700 28.885 82.850 29.055 ;
        RECT 83.090 28.750 83.240 28.920 ;
        RECT 84.820 28.750 84.970 28.920 ;
        RECT 85.210 28.885 85.360 29.055 ;
        RECT 85.600 28.885 85.750 29.055 ;
        RECT 85.990 28.750 86.140 28.920 ;
        RECT 87.720 28.750 87.870 28.920 ;
        RECT 88.110 28.885 88.260 29.055 ;
        RECT 88.500 28.885 88.650 29.055 ;
        RECT 88.890 28.750 89.040 28.920 ;
        RECT 90.620 28.750 90.770 28.920 ;
        RECT 91.010 28.885 91.160 29.055 ;
        RECT 91.400 28.885 91.550 29.055 ;
        RECT 91.790 28.750 91.940 28.920 ;
        RECT 0.985 28.665 1.035 28.700 ;
        POLYGON 1.035 28.700 1.070 28.665 1.035 28.665 ;
        RECT 0.985 28.540 1.070 28.665 ;
        RECT 1.690 28.540 1.775 28.700 ;
        RECT 3.885 28.665 3.935 28.700 ;
        POLYGON 3.935 28.700 3.970 28.665 3.935 28.665 ;
        RECT 3.885 28.540 3.970 28.665 ;
        RECT 4.590 28.540 4.675 28.700 ;
        RECT 6.785 28.665 6.835 28.700 ;
        POLYGON 6.835 28.700 6.870 28.665 6.835 28.665 ;
        RECT 6.785 28.540 6.870 28.665 ;
        RECT 7.490 28.540 7.575 28.700 ;
        RECT 9.685 28.665 9.735 28.700 ;
        POLYGON 9.735 28.700 9.770 28.665 9.735 28.665 ;
        RECT 9.685 28.540 9.770 28.665 ;
        RECT 10.390 28.540 10.475 28.700 ;
        RECT 12.585 28.665 12.635 28.700 ;
        POLYGON 12.635 28.700 12.670 28.665 12.635 28.665 ;
        RECT 12.585 28.540 12.670 28.665 ;
        RECT 13.290 28.540 13.375 28.700 ;
        RECT 15.485 28.665 15.535 28.700 ;
        POLYGON 15.535 28.700 15.570 28.665 15.535 28.665 ;
        RECT 15.485 28.540 15.570 28.665 ;
        RECT 16.190 28.540 16.275 28.700 ;
        RECT 18.385 28.665 18.435 28.700 ;
        POLYGON 18.435 28.700 18.470 28.665 18.435 28.665 ;
        RECT 18.385 28.540 18.470 28.665 ;
        RECT 19.090 28.540 19.175 28.700 ;
        RECT 21.285 28.665 21.335 28.700 ;
        POLYGON 21.335 28.700 21.370 28.665 21.335 28.665 ;
        RECT 21.285 28.540 21.370 28.665 ;
        RECT 21.990 28.540 22.075 28.700 ;
        RECT 24.185 28.665 24.235 28.700 ;
        POLYGON 24.235 28.700 24.270 28.665 24.235 28.665 ;
        RECT 24.185 28.540 24.270 28.665 ;
        RECT 24.890 28.540 24.975 28.700 ;
        RECT 27.085 28.665 27.135 28.700 ;
        POLYGON 27.135 28.700 27.170 28.665 27.135 28.665 ;
        RECT 27.085 28.540 27.170 28.665 ;
        RECT 27.790 28.540 27.875 28.700 ;
        RECT 29.985 28.665 30.035 28.700 ;
        POLYGON 30.035 28.700 30.070 28.665 30.035 28.665 ;
        RECT 29.985 28.540 30.070 28.665 ;
        RECT 30.690 28.540 30.775 28.700 ;
        RECT 32.885 28.665 32.935 28.700 ;
        POLYGON 32.935 28.700 32.970 28.665 32.935 28.665 ;
        RECT 32.885 28.540 32.970 28.665 ;
        RECT 33.590 28.540 33.675 28.700 ;
        RECT 35.785 28.665 35.835 28.700 ;
        POLYGON 35.835 28.700 35.870 28.665 35.835 28.665 ;
        RECT 35.785 28.540 35.870 28.665 ;
        RECT 36.490 28.540 36.575 28.700 ;
        RECT 38.685 28.665 38.735 28.700 ;
        POLYGON 38.735 28.700 38.770 28.665 38.735 28.665 ;
        RECT 38.685 28.540 38.770 28.665 ;
        RECT 39.390 28.540 39.475 28.700 ;
        RECT 41.585 28.665 41.635 28.700 ;
        POLYGON 41.635 28.700 41.670 28.665 41.635 28.665 ;
        RECT 41.585 28.540 41.670 28.665 ;
        RECT 42.290 28.540 42.375 28.700 ;
        RECT 44.485 28.665 44.535 28.700 ;
        POLYGON 44.535 28.700 44.570 28.665 44.535 28.665 ;
        RECT 44.485 28.540 44.570 28.665 ;
        RECT 45.190 28.540 45.275 28.700 ;
        RECT 47.385 28.665 47.435 28.700 ;
        POLYGON 47.435 28.700 47.470 28.665 47.435 28.665 ;
        RECT 47.385 28.540 47.470 28.665 ;
        RECT 48.090 28.540 48.175 28.700 ;
        RECT 50.285 28.665 50.335 28.700 ;
        POLYGON 50.335 28.700 50.370 28.665 50.335 28.665 ;
        RECT 50.285 28.540 50.370 28.665 ;
        RECT 50.990 28.540 51.075 28.700 ;
        RECT 53.185 28.665 53.235 28.700 ;
        POLYGON 53.235 28.700 53.270 28.665 53.235 28.665 ;
        RECT 53.185 28.540 53.270 28.665 ;
        RECT 53.890 28.540 53.975 28.700 ;
        RECT 56.085 28.665 56.135 28.700 ;
        POLYGON 56.135 28.700 56.170 28.665 56.135 28.665 ;
        RECT 56.085 28.540 56.170 28.665 ;
        RECT 56.790 28.540 56.875 28.700 ;
        RECT 58.985 28.665 59.035 28.700 ;
        POLYGON 59.035 28.700 59.070 28.665 59.035 28.665 ;
        RECT 58.985 28.540 59.070 28.665 ;
        RECT 59.690 28.540 59.775 28.700 ;
        RECT 61.885 28.665 61.935 28.700 ;
        POLYGON 61.935 28.700 61.970 28.665 61.935 28.665 ;
        RECT 61.885 28.540 61.970 28.665 ;
        RECT 62.590 28.540 62.675 28.700 ;
        RECT 64.785 28.665 64.835 28.700 ;
        POLYGON 64.835 28.700 64.870 28.665 64.835 28.665 ;
        RECT 64.785 28.540 64.870 28.665 ;
        RECT 65.490 28.540 65.575 28.700 ;
        RECT 67.685 28.665 67.735 28.700 ;
        POLYGON 67.735 28.700 67.770 28.665 67.735 28.665 ;
        RECT 67.685 28.540 67.770 28.665 ;
        RECT 68.390 28.540 68.475 28.700 ;
        RECT 70.585 28.665 70.635 28.700 ;
        POLYGON 70.635 28.700 70.670 28.665 70.635 28.665 ;
        RECT 70.585 28.540 70.670 28.665 ;
        RECT 71.290 28.540 71.375 28.700 ;
        RECT 73.485 28.665 73.535 28.700 ;
        POLYGON 73.535 28.700 73.570 28.665 73.535 28.665 ;
        RECT 73.485 28.540 73.570 28.665 ;
        RECT 74.190 28.540 74.275 28.700 ;
        RECT 76.385 28.665 76.435 28.700 ;
        POLYGON 76.435 28.700 76.470 28.665 76.435 28.665 ;
        RECT 76.385 28.540 76.470 28.665 ;
        RECT 77.090 28.540 77.175 28.700 ;
        RECT 79.285 28.665 79.335 28.700 ;
        POLYGON 79.335 28.700 79.370 28.665 79.335 28.665 ;
        RECT 79.285 28.540 79.370 28.665 ;
        RECT 79.990 28.540 80.075 28.700 ;
        RECT 82.185 28.665 82.235 28.700 ;
        POLYGON 82.235 28.700 82.270 28.665 82.235 28.665 ;
        RECT 82.185 28.540 82.270 28.665 ;
        RECT 82.890 28.540 82.975 28.700 ;
        RECT 85.085 28.665 85.135 28.700 ;
        POLYGON 85.135 28.700 85.170 28.665 85.135 28.665 ;
        RECT 85.085 28.540 85.170 28.665 ;
        RECT 85.790 28.540 85.875 28.700 ;
        RECT 87.985 28.665 88.035 28.700 ;
        POLYGON 88.035 28.700 88.070 28.665 88.035 28.665 ;
        RECT 87.985 28.540 88.070 28.665 ;
        RECT 88.690 28.540 88.775 28.700 ;
        RECT 90.885 28.665 90.935 28.700 ;
        POLYGON 90.935 28.700 90.970 28.665 90.935 28.665 ;
        RECT 90.885 28.540 90.970 28.665 ;
        RECT 91.590 28.540 91.675 28.700 ;
        RECT 0.775 27.920 0.850 28.060 ;
        RECT 0.990 27.870 1.065 28.010 ;
        RECT 1.695 27.930 1.755 28.010 ;
        POLYGON 1.695 27.930 1.755 27.930 1.755 27.870 ;
        RECT 1.910 27.920 1.985 28.060 ;
        RECT 3.675 27.920 3.750 28.060 ;
        RECT 3.890 27.870 3.965 28.010 ;
        RECT 4.595 27.930 4.655 28.010 ;
        POLYGON 4.595 27.930 4.655 27.930 4.655 27.870 ;
        RECT 4.810 27.920 4.885 28.060 ;
        RECT 6.575 27.920 6.650 28.060 ;
        RECT 6.790 27.870 6.865 28.010 ;
        RECT 7.495 27.930 7.555 28.010 ;
        POLYGON 7.495 27.930 7.555 27.930 7.555 27.870 ;
        RECT 7.710 27.920 7.785 28.060 ;
        RECT 9.475 27.920 9.550 28.060 ;
        RECT 9.690 27.870 9.765 28.010 ;
        RECT 10.395 27.930 10.455 28.010 ;
        POLYGON 10.395 27.930 10.455 27.930 10.455 27.870 ;
        RECT 10.610 27.920 10.685 28.060 ;
        RECT 12.375 27.920 12.450 28.060 ;
        RECT 12.590 27.870 12.665 28.010 ;
        RECT 13.295 27.930 13.355 28.010 ;
        POLYGON 13.295 27.930 13.355 27.930 13.355 27.870 ;
        RECT 13.510 27.920 13.585 28.060 ;
        RECT 15.275 27.920 15.350 28.060 ;
        RECT 15.490 27.870 15.565 28.010 ;
        RECT 16.195 27.930 16.255 28.010 ;
        POLYGON 16.195 27.930 16.255 27.930 16.255 27.870 ;
        RECT 16.410 27.920 16.485 28.060 ;
        RECT 18.175 27.920 18.250 28.060 ;
        RECT 18.390 27.870 18.465 28.010 ;
        RECT 19.095 27.930 19.155 28.010 ;
        POLYGON 19.095 27.930 19.155 27.930 19.155 27.870 ;
        RECT 19.310 27.920 19.385 28.060 ;
        RECT 21.075 27.920 21.150 28.060 ;
        RECT 21.290 27.870 21.365 28.010 ;
        RECT 21.995 27.930 22.055 28.010 ;
        POLYGON 21.995 27.930 22.055 27.930 22.055 27.870 ;
        RECT 22.210 27.920 22.285 28.060 ;
        RECT 23.975 27.920 24.050 28.060 ;
        RECT 24.190 27.870 24.265 28.010 ;
        RECT 24.895 27.930 24.955 28.010 ;
        POLYGON 24.895 27.930 24.955 27.930 24.955 27.870 ;
        RECT 25.110 27.920 25.185 28.060 ;
        RECT 26.875 27.920 26.950 28.060 ;
        RECT 27.090 27.870 27.165 28.010 ;
        RECT 27.795 27.930 27.855 28.010 ;
        POLYGON 27.795 27.930 27.855 27.930 27.855 27.870 ;
        RECT 28.010 27.920 28.085 28.060 ;
        RECT 29.775 27.920 29.850 28.060 ;
        RECT 29.990 27.870 30.065 28.010 ;
        RECT 30.695 27.930 30.755 28.010 ;
        POLYGON 30.695 27.930 30.755 27.930 30.755 27.870 ;
        RECT 30.910 27.920 30.985 28.060 ;
        RECT 32.675 27.920 32.750 28.060 ;
        RECT 32.890 27.870 32.965 28.010 ;
        RECT 33.595 27.930 33.655 28.010 ;
        POLYGON 33.595 27.930 33.655 27.930 33.655 27.870 ;
        RECT 33.810 27.920 33.885 28.060 ;
        RECT 35.575 27.920 35.650 28.060 ;
        RECT 35.790 27.870 35.865 28.010 ;
        RECT 36.495 27.930 36.555 28.010 ;
        POLYGON 36.495 27.930 36.555 27.930 36.555 27.870 ;
        RECT 36.710 27.920 36.785 28.060 ;
        RECT 38.475 27.920 38.550 28.060 ;
        RECT 38.690 27.870 38.765 28.010 ;
        RECT 39.395 27.930 39.455 28.010 ;
        POLYGON 39.395 27.930 39.455 27.930 39.455 27.870 ;
        RECT 39.610 27.920 39.685 28.060 ;
        RECT 41.375 27.920 41.450 28.060 ;
        RECT 41.590 27.870 41.665 28.010 ;
        RECT 42.295 27.930 42.355 28.010 ;
        POLYGON 42.295 27.930 42.355 27.930 42.355 27.870 ;
        RECT 42.510 27.920 42.585 28.060 ;
        RECT 44.275 27.920 44.350 28.060 ;
        RECT 44.490 27.870 44.565 28.010 ;
        RECT 45.195 27.930 45.255 28.010 ;
        POLYGON 45.195 27.930 45.255 27.930 45.255 27.870 ;
        RECT 45.410 27.920 45.485 28.060 ;
        RECT 47.175 27.920 47.250 28.060 ;
        RECT 47.390 27.870 47.465 28.010 ;
        RECT 48.095 27.930 48.155 28.010 ;
        POLYGON 48.095 27.930 48.155 27.930 48.155 27.870 ;
        RECT 48.310 27.920 48.385 28.060 ;
        RECT 50.075 27.920 50.150 28.060 ;
        RECT 50.290 27.870 50.365 28.010 ;
        RECT 50.995 27.930 51.055 28.010 ;
        POLYGON 50.995 27.930 51.055 27.930 51.055 27.870 ;
        RECT 51.210 27.920 51.285 28.060 ;
        RECT 52.975 27.920 53.050 28.060 ;
        RECT 53.190 27.870 53.265 28.010 ;
        RECT 53.895 27.930 53.955 28.010 ;
        POLYGON 53.895 27.930 53.955 27.930 53.955 27.870 ;
        RECT 54.110 27.920 54.185 28.060 ;
        RECT 55.875 27.920 55.950 28.060 ;
        RECT 56.090 27.870 56.165 28.010 ;
        RECT 56.795 27.930 56.855 28.010 ;
        POLYGON 56.795 27.930 56.855 27.930 56.855 27.870 ;
        RECT 57.010 27.920 57.085 28.060 ;
        RECT 58.775 27.920 58.850 28.060 ;
        RECT 58.990 27.870 59.065 28.010 ;
        RECT 59.695 27.930 59.755 28.010 ;
        POLYGON 59.695 27.930 59.755 27.930 59.755 27.870 ;
        RECT 59.910 27.920 59.985 28.060 ;
        RECT 61.675 27.920 61.750 28.060 ;
        RECT 61.890 27.870 61.965 28.010 ;
        RECT 62.595 27.930 62.655 28.010 ;
        POLYGON 62.595 27.930 62.655 27.930 62.655 27.870 ;
        RECT 62.810 27.920 62.885 28.060 ;
        RECT 64.575 27.920 64.650 28.060 ;
        RECT 64.790 27.870 64.865 28.010 ;
        RECT 65.495 27.930 65.555 28.010 ;
        POLYGON 65.495 27.930 65.555 27.930 65.555 27.870 ;
        RECT 65.710 27.920 65.785 28.060 ;
        RECT 67.475 27.920 67.550 28.060 ;
        RECT 67.690 27.870 67.765 28.010 ;
        RECT 68.395 27.930 68.455 28.010 ;
        POLYGON 68.395 27.930 68.455 27.930 68.455 27.870 ;
        RECT 68.610 27.920 68.685 28.060 ;
        RECT 70.375 27.920 70.450 28.060 ;
        RECT 70.590 27.870 70.665 28.010 ;
        RECT 71.295 27.930 71.355 28.010 ;
        POLYGON 71.295 27.930 71.355 27.930 71.355 27.870 ;
        RECT 71.510 27.920 71.585 28.060 ;
        RECT 73.275 27.920 73.350 28.060 ;
        RECT 73.490 27.870 73.565 28.010 ;
        RECT 74.195 27.930 74.255 28.010 ;
        POLYGON 74.195 27.930 74.255 27.930 74.255 27.870 ;
        RECT 74.410 27.920 74.485 28.060 ;
        RECT 76.175 27.920 76.250 28.060 ;
        RECT 76.390 27.870 76.465 28.010 ;
        RECT 77.095 27.930 77.155 28.010 ;
        POLYGON 77.095 27.930 77.155 27.930 77.155 27.870 ;
        RECT 77.310 27.920 77.385 28.060 ;
        RECT 79.075 27.920 79.150 28.060 ;
        RECT 79.290 27.870 79.365 28.010 ;
        RECT 79.995 27.930 80.055 28.010 ;
        POLYGON 79.995 27.930 80.055 27.930 80.055 27.870 ;
        RECT 80.210 27.920 80.285 28.060 ;
        RECT 81.975 27.920 82.050 28.060 ;
        RECT 82.190 27.870 82.265 28.010 ;
        RECT 82.895 27.930 82.955 28.010 ;
        POLYGON 82.895 27.930 82.955 27.930 82.955 27.870 ;
        RECT 83.110 27.920 83.185 28.060 ;
        RECT 84.875 27.920 84.950 28.060 ;
        RECT 85.090 27.870 85.165 28.010 ;
        RECT 85.795 27.930 85.855 28.010 ;
        POLYGON 85.795 27.930 85.855 27.930 85.855 27.870 ;
        RECT 86.010 27.920 86.085 28.060 ;
        RECT 87.775 27.920 87.850 28.060 ;
        RECT 87.990 27.870 88.065 28.010 ;
        RECT 88.695 27.930 88.755 28.010 ;
        POLYGON 88.695 27.930 88.755 27.930 88.755 27.870 ;
        RECT 88.910 27.920 88.985 28.060 ;
        RECT 90.675 27.920 90.750 28.060 ;
        RECT 90.890 27.870 90.965 28.010 ;
        RECT 91.595 27.930 91.655 28.010 ;
        POLYGON 91.595 27.930 91.655 27.930 91.655 27.870 ;
        RECT 91.810 27.920 91.885 28.060 ;
        RECT 0.720 27.400 0.870 27.570 ;
        RECT 1.110 27.535 1.260 27.705 ;
        RECT 1.500 27.535 1.650 27.705 ;
        RECT 1.890 27.400 2.040 27.570 ;
        RECT 3.620 27.400 3.770 27.570 ;
        RECT 4.010 27.535 4.160 27.705 ;
        RECT 4.400 27.535 4.550 27.705 ;
        RECT 4.790 27.400 4.940 27.570 ;
        RECT 6.520 27.400 6.670 27.570 ;
        RECT 6.910 27.535 7.060 27.705 ;
        RECT 7.300 27.535 7.450 27.705 ;
        RECT 7.690 27.400 7.840 27.570 ;
        RECT 9.420 27.400 9.570 27.570 ;
        RECT 9.810 27.535 9.960 27.705 ;
        RECT 10.200 27.535 10.350 27.705 ;
        RECT 10.590 27.400 10.740 27.570 ;
        RECT 12.320 27.400 12.470 27.570 ;
        RECT 12.710 27.535 12.860 27.705 ;
        RECT 13.100 27.535 13.250 27.705 ;
        RECT 13.490 27.400 13.640 27.570 ;
        RECT 15.220 27.400 15.370 27.570 ;
        RECT 15.610 27.535 15.760 27.705 ;
        RECT 16.000 27.535 16.150 27.705 ;
        RECT 16.390 27.400 16.540 27.570 ;
        RECT 18.120 27.400 18.270 27.570 ;
        RECT 18.510 27.535 18.660 27.705 ;
        RECT 18.900 27.535 19.050 27.705 ;
        RECT 19.290 27.400 19.440 27.570 ;
        RECT 21.020 27.400 21.170 27.570 ;
        RECT 21.410 27.535 21.560 27.705 ;
        RECT 21.800 27.535 21.950 27.705 ;
        RECT 22.190 27.400 22.340 27.570 ;
        RECT 23.920 27.400 24.070 27.570 ;
        RECT 24.310 27.535 24.460 27.705 ;
        RECT 24.700 27.535 24.850 27.705 ;
        RECT 25.090 27.400 25.240 27.570 ;
        RECT 26.820 27.400 26.970 27.570 ;
        RECT 27.210 27.535 27.360 27.705 ;
        RECT 27.600 27.535 27.750 27.705 ;
        RECT 27.990 27.400 28.140 27.570 ;
        RECT 29.720 27.400 29.870 27.570 ;
        RECT 30.110 27.535 30.260 27.705 ;
        RECT 30.500 27.535 30.650 27.705 ;
        RECT 30.890 27.400 31.040 27.570 ;
        RECT 32.620 27.400 32.770 27.570 ;
        RECT 33.010 27.535 33.160 27.705 ;
        RECT 33.400 27.535 33.550 27.705 ;
        RECT 33.790 27.400 33.940 27.570 ;
        RECT 35.520 27.400 35.670 27.570 ;
        RECT 35.910 27.535 36.060 27.705 ;
        RECT 36.300 27.535 36.450 27.705 ;
        RECT 36.690 27.400 36.840 27.570 ;
        RECT 38.420 27.400 38.570 27.570 ;
        RECT 38.810 27.535 38.960 27.705 ;
        RECT 39.200 27.535 39.350 27.705 ;
        RECT 39.590 27.400 39.740 27.570 ;
        RECT 41.320 27.400 41.470 27.570 ;
        RECT 41.710 27.535 41.860 27.705 ;
        RECT 42.100 27.535 42.250 27.705 ;
        RECT 42.490 27.400 42.640 27.570 ;
        RECT 44.220 27.400 44.370 27.570 ;
        RECT 44.610 27.535 44.760 27.705 ;
        RECT 45.000 27.535 45.150 27.705 ;
        RECT 45.390 27.400 45.540 27.570 ;
        RECT 47.120 27.400 47.270 27.570 ;
        RECT 47.510 27.535 47.660 27.705 ;
        RECT 47.900 27.535 48.050 27.705 ;
        RECT 48.290 27.400 48.440 27.570 ;
        RECT 50.020 27.400 50.170 27.570 ;
        RECT 50.410 27.535 50.560 27.705 ;
        RECT 50.800 27.535 50.950 27.705 ;
        RECT 51.190 27.400 51.340 27.570 ;
        RECT 52.920 27.400 53.070 27.570 ;
        RECT 53.310 27.535 53.460 27.705 ;
        RECT 53.700 27.535 53.850 27.705 ;
        RECT 54.090 27.400 54.240 27.570 ;
        RECT 55.820 27.400 55.970 27.570 ;
        RECT 56.210 27.535 56.360 27.705 ;
        RECT 56.600 27.535 56.750 27.705 ;
        RECT 56.990 27.400 57.140 27.570 ;
        RECT 58.720 27.400 58.870 27.570 ;
        RECT 59.110 27.535 59.260 27.705 ;
        RECT 59.500 27.535 59.650 27.705 ;
        RECT 59.890 27.400 60.040 27.570 ;
        RECT 61.620 27.400 61.770 27.570 ;
        RECT 62.010 27.535 62.160 27.705 ;
        RECT 62.400 27.535 62.550 27.705 ;
        RECT 62.790 27.400 62.940 27.570 ;
        RECT 64.520 27.400 64.670 27.570 ;
        RECT 64.910 27.535 65.060 27.705 ;
        RECT 65.300 27.535 65.450 27.705 ;
        RECT 65.690 27.400 65.840 27.570 ;
        RECT 67.420 27.400 67.570 27.570 ;
        RECT 67.810 27.535 67.960 27.705 ;
        RECT 68.200 27.535 68.350 27.705 ;
        RECT 68.590 27.400 68.740 27.570 ;
        RECT 70.320 27.400 70.470 27.570 ;
        RECT 70.710 27.535 70.860 27.705 ;
        RECT 71.100 27.535 71.250 27.705 ;
        RECT 71.490 27.400 71.640 27.570 ;
        RECT 73.220 27.400 73.370 27.570 ;
        RECT 73.610 27.535 73.760 27.705 ;
        RECT 74.000 27.535 74.150 27.705 ;
        RECT 74.390 27.400 74.540 27.570 ;
        RECT 76.120 27.400 76.270 27.570 ;
        RECT 76.510 27.535 76.660 27.705 ;
        RECT 76.900 27.535 77.050 27.705 ;
        RECT 77.290 27.400 77.440 27.570 ;
        RECT 79.020 27.400 79.170 27.570 ;
        RECT 79.410 27.535 79.560 27.705 ;
        RECT 79.800 27.535 79.950 27.705 ;
        RECT 80.190 27.400 80.340 27.570 ;
        RECT 81.920 27.400 82.070 27.570 ;
        RECT 82.310 27.535 82.460 27.705 ;
        RECT 82.700 27.535 82.850 27.705 ;
        RECT 83.090 27.400 83.240 27.570 ;
        RECT 84.820 27.400 84.970 27.570 ;
        RECT 85.210 27.535 85.360 27.705 ;
        RECT 85.600 27.535 85.750 27.705 ;
        RECT 85.990 27.400 86.140 27.570 ;
        RECT 87.720 27.400 87.870 27.570 ;
        RECT 88.110 27.535 88.260 27.705 ;
        RECT 88.500 27.535 88.650 27.705 ;
        RECT 88.890 27.400 89.040 27.570 ;
        RECT 90.620 27.400 90.770 27.570 ;
        RECT 91.010 27.535 91.160 27.705 ;
        RECT 91.400 27.535 91.550 27.705 ;
        RECT 91.790 27.400 91.940 27.570 ;
        RECT 0.985 27.315 1.035 27.350 ;
        POLYGON 1.035 27.350 1.070 27.315 1.035 27.315 ;
        RECT 0.985 27.190 1.070 27.315 ;
        RECT 1.690 27.190 1.775 27.350 ;
        RECT 3.885 27.315 3.935 27.350 ;
        POLYGON 3.935 27.350 3.970 27.315 3.935 27.315 ;
        RECT 3.885 27.190 3.970 27.315 ;
        RECT 4.590 27.190 4.675 27.350 ;
        RECT 6.785 27.315 6.835 27.350 ;
        POLYGON 6.835 27.350 6.870 27.315 6.835 27.315 ;
        RECT 6.785 27.190 6.870 27.315 ;
        RECT 7.490 27.190 7.575 27.350 ;
        RECT 9.685 27.315 9.735 27.350 ;
        POLYGON 9.735 27.350 9.770 27.315 9.735 27.315 ;
        RECT 9.685 27.190 9.770 27.315 ;
        RECT 10.390 27.190 10.475 27.350 ;
        RECT 12.585 27.315 12.635 27.350 ;
        POLYGON 12.635 27.350 12.670 27.315 12.635 27.315 ;
        RECT 12.585 27.190 12.670 27.315 ;
        RECT 13.290 27.190 13.375 27.350 ;
        RECT 15.485 27.315 15.535 27.350 ;
        POLYGON 15.535 27.350 15.570 27.315 15.535 27.315 ;
        RECT 15.485 27.190 15.570 27.315 ;
        RECT 16.190 27.190 16.275 27.350 ;
        RECT 18.385 27.315 18.435 27.350 ;
        POLYGON 18.435 27.350 18.470 27.315 18.435 27.315 ;
        RECT 18.385 27.190 18.470 27.315 ;
        RECT 19.090 27.190 19.175 27.350 ;
        RECT 21.285 27.315 21.335 27.350 ;
        POLYGON 21.335 27.350 21.370 27.315 21.335 27.315 ;
        RECT 21.285 27.190 21.370 27.315 ;
        RECT 21.990 27.190 22.075 27.350 ;
        RECT 24.185 27.315 24.235 27.350 ;
        POLYGON 24.235 27.350 24.270 27.315 24.235 27.315 ;
        RECT 24.185 27.190 24.270 27.315 ;
        RECT 24.890 27.190 24.975 27.350 ;
        RECT 27.085 27.315 27.135 27.350 ;
        POLYGON 27.135 27.350 27.170 27.315 27.135 27.315 ;
        RECT 27.085 27.190 27.170 27.315 ;
        RECT 27.790 27.190 27.875 27.350 ;
        RECT 29.985 27.315 30.035 27.350 ;
        POLYGON 30.035 27.350 30.070 27.315 30.035 27.315 ;
        RECT 29.985 27.190 30.070 27.315 ;
        RECT 30.690 27.190 30.775 27.350 ;
        RECT 32.885 27.315 32.935 27.350 ;
        POLYGON 32.935 27.350 32.970 27.315 32.935 27.315 ;
        RECT 32.885 27.190 32.970 27.315 ;
        RECT 33.590 27.190 33.675 27.350 ;
        RECT 35.785 27.315 35.835 27.350 ;
        POLYGON 35.835 27.350 35.870 27.315 35.835 27.315 ;
        RECT 35.785 27.190 35.870 27.315 ;
        RECT 36.490 27.190 36.575 27.350 ;
        RECT 38.685 27.315 38.735 27.350 ;
        POLYGON 38.735 27.350 38.770 27.315 38.735 27.315 ;
        RECT 38.685 27.190 38.770 27.315 ;
        RECT 39.390 27.190 39.475 27.350 ;
        RECT 41.585 27.315 41.635 27.350 ;
        POLYGON 41.635 27.350 41.670 27.315 41.635 27.315 ;
        RECT 41.585 27.190 41.670 27.315 ;
        RECT 42.290 27.190 42.375 27.350 ;
        RECT 44.485 27.315 44.535 27.350 ;
        POLYGON 44.535 27.350 44.570 27.315 44.535 27.315 ;
        RECT 44.485 27.190 44.570 27.315 ;
        RECT 45.190 27.190 45.275 27.350 ;
        RECT 47.385 27.315 47.435 27.350 ;
        POLYGON 47.435 27.350 47.470 27.315 47.435 27.315 ;
        RECT 47.385 27.190 47.470 27.315 ;
        RECT 48.090 27.190 48.175 27.350 ;
        RECT 50.285 27.315 50.335 27.350 ;
        POLYGON 50.335 27.350 50.370 27.315 50.335 27.315 ;
        RECT 50.285 27.190 50.370 27.315 ;
        RECT 50.990 27.190 51.075 27.350 ;
        RECT 53.185 27.315 53.235 27.350 ;
        POLYGON 53.235 27.350 53.270 27.315 53.235 27.315 ;
        RECT 53.185 27.190 53.270 27.315 ;
        RECT 53.890 27.190 53.975 27.350 ;
        RECT 56.085 27.315 56.135 27.350 ;
        POLYGON 56.135 27.350 56.170 27.315 56.135 27.315 ;
        RECT 56.085 27.190 56.170 27.315 ;
        RECT 56.790 27.190 56.875 27.350 ;
        RECT 58.985 27.315 59.035 27.350 ;
        POLYGON 59.035 27.350 59.070 27.315 59.035 27.315 ;
        RECT 58.985 27.190 59.070 27.315 ;
        RECT 59.690 27.190 59.775 27.350 ;
        RECT 61.885 27.315 61.935 27.350 ;
        POLYGON 61.935 27.350 61.970 27.315 61.935 27.315 ;
        RECT 61.885 27.190 61.970 27.315 ;
        RECT 62.590 27.190 62.675 27.350 ;
        RECT 64.785 27.315 64.835 27.350 ;
        POLYGON 64.835 27.350 64.870 27.315 64.835 27.315 ;
        RECT 64.785 27.190 64.870 27.315 ;
        RECT 65.490 27.190 65.575 27.350 ;
        RECT 67.685 27.315 67.735 27.350 ;
        POLYGON 67.735 27.350 67.770 27.315 67.735 27.315 ;
        RECT 67.685 27.190 67.770 27.315 ;
        RECT 68.390 27.190 68.475 27.350 ;
        RECT 70.585 27.315 70.635 27.350 ;
        POLYGON 70.635 27.350 70.670 27.315 70.635 27.315 ;
        RECT 70.585 27.190 70.670 27.315 ;
        RECT 71.290 27.190 71.375 27.350 ;
        RECT 73.485 27.315 73.535 27.350 ;
        POLYGON 73.535 27.350 73.570 27.315 73.535 27.315 ;
        RECT 73.485 27.190 73.570 27.315 ;
        RECT 74.190 27.190 74.275 27.350 ;
        RECT 76.385 27.315 76.435 27.350 ;
        POLYGON 76.435 27.350 76.470 27.315 76.435 27.315 ;
        RECT 76.385 27.190 76.470 27.315 ;
        RECT 77.090 27.190 77.175 27.350 ;
        RECT 79.285 27.315 79.335 27.350 ;
        POLYGON 79.335 27.350 79.370 27.315 79.335 27.315 ;
        RECT 79.285 27.190 79.370 27.315 ;
        RECT 79.990 27.190 80.075 27.350 ;
        RECT 82.185 27.315 82.235 27.350 ;
        POLYGON 82.235 27.350 82.270 27.315 82.235 27.315 ;
        RECT 82.185 27.190 82.270 27.315 ;
        RECT 82.890 27.190 82.975 27.350 ;
        RECT 85.085 27.315 85.135 27.350 ;
        POLYGON 85.135 27.350 85.170 27.315 85.135 27.315 ;
        RECT 85.085 27.190 85.170 27.315 ;
        RECT 85.790 27.190 85.875 27.350 ;
        RECT 87.985 27.315 88.035 27.350 ;
        POLYGON 88.035 27.350 88.070 27.315 88.035 27.315 ;
        RECT 87.985 27.190 88.070 27.315 ;
        RECT 88.690 27.190 88.775 27.350 ;
        RECT 90.885 27.315 90.935 27.350 ;
        POLYGON 90.935 27.350 90.970 27.315 90.935 27.315 ;
        RECT 90.885 27.190 90.970 27.315 ;
        RECT 91.590 27.190 91.675 27.350 ;
        RECT 0.775 26.570 0.850 26.710 ;
        RECT 0.990 26.520 1.065 26.660 ;
        RECT 1.695 26.580 1.755 26.660 ;
        POLYGON 1.695 26.580 1.755 26.580 1.755 26.520 ;
        RECT 1.910 26.570 1.985 26.710 ;
        RECT 3.675 26.570 3.750 26.710 ;
        RECT 3.890 26.520 3.965 26.660 ;
        RECT 4.595 26.580 4.655 26.660 ;
        POLYGON 4.595 26.580 4.655 26.580 4.655 26.520 ;
        RECT 4.810 26.570 4.885 26.710 ;
        RECT 6.575 26.570 6.650 26.710 ;
        RECT 6.790 26.520 6.865 26.660 ;
        RECT 7.495 26.580 7.555 26.660 ;
        POLYGON 7.495 26.580 7.555 26.580 7.555 26.520 ;
        RECT 7.710 26.570 7.785 26.710 ;
        RECT 9.475 26.570 9.550 26.710 ;
        RECT 9.690 26.520 9.765 26.660 ;
        RECT 10.395 26.580 10.455 26.660 ;
        POLYGON 10.395 26.580 10.455 26.580 10.455 26.520 ;
        RECT 10.610 26.570 10.685 26.710 ;
        RECT 12.375 26.570 12.450 26.710 ;
        RECT 12.590 26.520 12.665 26.660 ;
        RECT 13.295 26.580 13.355 26.660 ;
        POLYGON 13.295 26.580 13.355 26.580 13.355 26.520 ;
        RECT 13.510 26.570 13.585 26.710 ;
        RECT 15.275 26.570 15.350 26.710 ;
        RECT 15.490 26.520 15.565 26.660 ;
        RECT 16.195 26.580 16.255 26.660 ;
        POLYGON 16.195 26.580 16.255 26.580 16.255 26.520 ;
        RECT 16.410 26.570 16.485 26.710 ;
        RECT 18.175 26.570 18.250 26.710 ;
        RECT 18.390 26.520 18.465 26.660 ;
        RECT 19.095 26.580 19.155 26.660 ;
        POLYGON 19.095 26.580 19.155 26.580 19.155 26.520 ;
        RECT 19.310 26.570 19.385 26.710 ;
        RECT 21.075 26.570 21.150 26.710 ;
        RECT 21.290 26.520 21.365 26.660 ;
        RECT 21.995 26.580 22.055 26.660 ;
        POLYGON 21.995 26.580 22.055 26.580 22.055 26.520 ;
        RECT 22.210 26.570 22.285 26.710 ;
        RECT 23.975 26.570 24.050 26.710 ;
        RECT 24.190 26.520 24.265 26.660 ;
        RECT 24.895 26.580 24.955 26.660 ;
        POLYGON 24.895 26.580 24.955 26.580 24.955 26.520 ;
        RECT 25.110 26.570 25.185 26.710 ;
        RECT 26.875 26.570 26.950 26.710 ;
        RECT 27.090 26.520 27.165 26.660 ;
        RECT 27.795 26.580 27.855 26.660 ;
        POLYGON 27.795 26.580 27.855 26.580 27.855 26.520 ;
        RECT 28.010 26.570 28.085 26.710 ;
        RECT 29.775 26.570 29.850 26.710 ;
        RECT 29.990 26.520 30.065 26.660 ;
        RECT 30.695 26.580 30.755 26.660 ;
        POLYGON 30.695 26.580 30.755 26.580 30.755 26.520 ;
        RECT 30.910 26.570 30.985 26.710 ;
        RECT 32.675 26.570 32.750 26.710 ;
        RECT 32.890 26.520 32.965 26.660 ;
        RECT 33.595 26.580 33.655 26.660 ;
        POLYGON 33.595 26.580 33.655 26.580 33.655 26.520 ;
        RECT 33.810 26.570 33.885 26.710 ;
        RECT 35.575 26.570 35.650 26.710 ;
        RECT 35.790 26.520 35.865 26.660 ;
        RECT 36.495 26.580 36.555 26.660 ;
        POLYGON 36.495 26.580 36.555 26.580 36.555 26.520 ;
        RECT 36.710 26.570 36.785 26.710 ;
        RECT 38.475 26.570 38.550 26.710 ;
        RECT 38.690 26.520 38.765 26.660 ;
        RECT 39.395 26.580 39.455 26.660 ;
        POLYGON 39.395 26.580 39.455 26.580 39.455 26.520 ;
        RECT 39.610 26.570 39.685 26.710 ;
        RECT 41.375 26.570 41.450 26.710 ;
        RECT 41.590 26.520 41.665 26.660 ;
        RECT 42.295 26.580 42.355 26.660 ;
        POLYGON 42.295 26.580 42.355 26.580 42.355 26.520 ;
        RECT 42.510 26.570 42.585 26.710 ;
        RECT 44.275 26.570 44.350 26.710 ;
        RECT 44.490 26.520 44.565 26.660 ;
        RECT 45.195 26.580 45.255 26.660 ;
        POLYGON 45.195 26.580 45.255 26.580 45.255 26.520 ;
        RECT 45.410 26.570 45.485 26.710 ;
        RECT 47.175 26.570 47.250 26.710 ;
        RECT 47.390 26.520 47.465 26.660 ;
        RECT 48.095 26.580 48.155 26.660 ;
        POLYGON 48.095 26.580 48.155 26.580 48.155 26.520 ;
        RECT 48.310 26.570 48.385 26.710 ;
        RECT 50.075 26.570 50.150 26.710 ;
        RECT 50.290 26.520 50.365 26.660 ;
        RECT 50.995 26.580 51.055 26.660 ;
        POLYGON 50.995 26.580 51.055 26.580 51.055 26.520 ;
        RECT 51.210 26.570 51.285 26.710 ;
        RECT 52.975 26.570 53.050 26.710 ;
        RECT 53.190 26.520 53.265 26.660 ;
        RECT 53.895 26.580 53.955 26.660 ;
        POLYGON 53.895 26.580 53.955 26.580 53.955 26.520 ;
        RECT 54.110 26.570 54.185 26.710 ;
        RECT 55.875 26.570 55.950 26.710 ;
        RECT 56.090 26.520 56.165 26.660 ;
        RECT 56.795 26.580 56.855 26.660 ;
        POLYGON 56.795 26.580 56.855 26.580 56.855 26.520 ;
        RECT 57.010 26.570 57.085 26.710 ;
        RECT 58.775 26.570 58.850 26.710 ;
        RECT 58.990 26.520 59.065 26.660 ;
        RECT 59.695 26.580 59.755 26.660 ;
        POLYGON 59.695 26.580 59.755 26.580 59.755 26.520 ;
        RECT 59.910 26.570 59.985 26.710 ;
        RECT 61.675 26.570 61.750 26.710 ;
        RECT 61.890 26.520 61.965 26.660 ;
        RECT 62.595 26.580 62.655 26.660 ;
        POLYGON 62.595 26.580 62.655 26.580 62.655 26.520 ;
        RECT 62.810 26.570 62.885 26.710 ;
        RECT 64.575 26.570 64.650 26.710 ;
        RECT 64.790 26.520 64.865 26.660 ;
        RECT 65.495 26.580 65.555 26.660 ;
        POLYGON 65.495 26.580 65.555 26.580 65.555 26.520 ;
        RECT 65.710 26.570 65.785 26.710 ;
        RECT 67.475 26.570 67.550 26.710 ;
        RECT 67.690 26.520 67.765 26.660 ;
        RECT 68.395 26.580 68.455 26.660 ;
        POLYGON 68.395 26.580 68.455 26.580 68.455 26.520 ;
        RECT 68.610 26.570 68.685 26.710 ;
        RECT 70.375 26.570 70.450 26.710 ;
        RECT 70.590 26.520 70.665 26.660 ;
        RECT 71.295 26.580 71.355 26.660 ;
        POLYGON 71.295 26.580 71.355 26.580 71.355 26.520 ;
        RECT 71.510 26.570 71.585 26.710 ;
        RECT 73.275 26.570 73.350 26.710 ;
        RECT 73.490 26.520 73.565 26.660 ;
        RECT 74.195 26.580 74.255 26.660 ;
        POLYGON 74.195 26.580 74.255 26.580 74.255 26.520 ;
        RECT 74.410 26.570 74.485 26.710 ;
        RECT 76.175 26.570 76.250 26.710 ;
        RECT 76.390 26.520 76.465 26.660 ;
        RECT 77.095 26.580 77.155 26.660 ;
        POLYGON 77.095 26.580 77.155 26.580 77.155 26.520 ;
        RECT 77.310 26.570 77.385 26.710 ;
        RECT 79.075 26.570 79.150 26.710 ;
        RECT 79.290 26.520 79.365 26.660 ;
        RECT 79.995 26.580 80.055 26.660 ;
        POLYGON 79.995 26.580 80.055 26.580 80.055 26.520 ;
        RECT 80.210 26.570 80.285 26.710 ;
        RECT 81.975 26.570 82.050 26.710 ;
        RECT 82.190 26.520 82.265 26.660 ;
        RECT 82.895 26.580 82.955 26.660 ;
        POLYGON 82.895 26.580 82.955 26.580 82.955 26.520 ;
        RECT 83.110 26.570 83.185 26.710 ;
        RECT 84.875 26.570 84.950 26.710 ;
        RECT 85.090 26.520 85.165 26.660 ;
        RECT 85.795 26.580 85.855 26.660 ;
        POLYGON 85.795 26.580 85.855 26.580 85.855 26.520 ;
        RECT 86.010 26.570 86.085 26.710 ;
        RECT 87.775 26.570 87.850 26.710 ;
        RECT 87.990 26.520 88.065 26.660 ;
        RECT 88.695 26.580 88.755 26.660 ;
        POLYGON 88.695 26.580 88.755 26.580 88.755 26.520 ;
        RECT 88.910 26.570 88.985 26.710 ;
        RECT 90.675 26.570 90.750 26.710 ;
        RECT 90.890 26.520 90.965 26.660 ;
        RECT 91.595 26.580 91.655 26.660 ;
        POLYGON 91.595 26.580 91.655 26.580 91.655 26.520 ;
        RECT 91.810 26.570 91.885 26.710 ;
        RECT 0.720 26.050 0.870 26.220 ;
        RECT 1.110 26.185 1.260 26.355 ;
        RECT 1.500 26.185 1.650 26.355 ;
        RECT 1.890 26.050 2.040 26.220 ;
        RECT 3.620 26.050 3.770 26.220 ;
        RECT 4.010 26.185 4.160 26.355 ;
        RECT 4.400 26.185 4.550 26.355 ;
        RECT 4.790 26.050 4.940 26.220 ;
        RECT 6.520 26.050 6.670 26.220 ;
        RECT 6.910 26.185 7.060 26.355 ;
        RECT 7.300 26.185 7.450 26.355 ;
        RECT 7.690 26.050 7.840 26.220 ;
        RECT 9.420 26.050 9.570 26.220 ;
        RECT 9.810 26.185 9.960 26.355 ;
        RECT 10.200 26.185 10.350 26.355 ;
        RECT 10.590 26.050 10.740 26.220 ;
        RECT 12.320 26.050 12.470 26.220 ;
        RECT 12.710 26.185 12.860 26.355 ;
        RECT 13.100 26.185 13.250 26.355 ;
        RECT 13.490 26.050 13.640 26.220 ;
        RECT 15.220 26.050 15.370 26.220 ;
        RECT 15.610 26.185 15.760 26.355 ;
        RECT 16.000 26.185 16.150 26.355 ;
        RECT 16.390 26.050 16.540 26.220 ;
        RECT 18.120 26.050 18.270 26.220 ;
        RECT 18.510 26.185 18.660 26.355 ;
        RECT 18.900 26.185 19.050 26.355 ;
        RECT 19.290 26.050 19.440 26.220 ;
        RECT 21.020 26.050 21.170 26.220 ;
        RECT 21.410 26.185 21.560 26.355 ;
        RECT 21.800 26.185 21.950 26.355 ;
        RECT 22.190 26.050 22.340 26.220 ;
        RECT 23.920 26.050 24.070 26.220 ;
        RECT 24.310 26.185 24.460 26.355 ;
        RECT 24.700 26.185 24.850 26.355 ;
        RECT 25.090 26.050 25.240 26.220 ;
        RECT 26.820 26.050 26.970 26.220 ;
        RECT 27.210 26.185 27.360 26.355 ;
        RECT 27.600 26.185 27.750 26.355 ;
        RECT 27.990 26.050 28.140 26.220 ;
        RECT 29.720 26.050 29.870 26.220 ;
        RECT 30.110 26.185 30.260 26.355 ;
        RECT 30.500 26.185 30.650 26.355 ;
        RECT 30.890 26.050 31.040 26.220 ;
        RECT 32.620 26.050 32.770 26.220 ;
        RECT 33.010 26.185 33.160 26.355 ;
        RECT 33.400 26.185 33.550 26.355 ;
        RECT 33.790 26.050 33.940 26.220 ;
        RECT 35.520 26.050 35.670 26.220 ;
        RECT 35.910 26.185 36.060 26.355 ;
        RECT 36.300 26.185 36.450 26.355 ;
        RECT 36.690 26.050 36.840 26.220 ;
        RECT 38.420 26.050 38.570 26.220 ;
        RECT 38.810 26.185 38.960 26.355 ;
        RECT 39.200 26.185 39.350 26.355 ;
        RECT 39.590 26.050 39.740 26.220 ;
        RECT 41.320 26.050 41.470 26.220 ;
        RECT 41.710 26.185 41.860 26.355 ;
        RECT 42.100 26.185 42.250 26.355 ;
        RECT 42.490 26.050 42.640 26.220 ;
        RECT 44.220 26.050 44.370 26.220 ;
        RECT 44.610 26.185 44.760 26.355 ;
        RECT 45.000 26.185 45.150 26.355 ;
        RECT 45.390 26.050 45.540 26.220 ;
        RECT 47.120 26.050 47.270 26.220 ;
        RECT 47.510 26.185 47.660 26.355 ;
        RECT 47.900 26.185 48.050 26.355 ;
        RECT 48.290 26.050 48.440 26.220 ;
        RECT 50.020 26.050 50.170 26.220 ;
        RECT 50.410 26.185 50.560 26.355 ;
        RECT 50.800 26.185 50.950 26.355 ;
        RECT 51.190 26.050 51.340 26.220 ;
        RECT 52.920 26.050 53.070 26.220 ;
        RECT 53.310 26.185 53.460 26.355 ;
        RECT 53.700 26.185 53.850 26.355 ;
        RECT 54.090 26.050 54.240 26.220 ;
        RECT 55.820 26.050 55.970 26.220 ;
        RECT 56.210 26.185 56.360 26.355 ;
        RECT 56.600 26.185 56.750 26.355 ;
        RECT 56.990 26.050 57.140 26.220 ;
        RECT 58.720 26.050 58.870 26.220 ;
        RECT 59.110 26.185 59.260 26.355 ;
        RECT 59.500 26.185 59.650 26.355 ;
        RECT 59.890 26.050 60.040 26.220 ;
        RECT 61.620 26.050 61.770 26.220 ;
        RECT 62.010 26.185 62.160 26.355 ;
        RECT 62.400 26.185 62.550 26.355 ;
        RECT 62.790 26.050 62.940 26.220 ;
        RECT 64.520 26.050 64.670 26.220 ;
        RECT 64.910 26.185 65.060 26.355 ;
        RECT 65.300 26.185 65.450 26.355 ;
        RECT 65.690 26.050 65.840 26.220 ;
        RECT 67.420 26.050 67.570 26.220 ;
        RECT 67.810 26.185 67.960 26.355 ;
        RECT 68.200 26.185 68.350 26.355 ;
        RECT 68.590 26.050 68.740 26.220 ;
        RECT 70.320 26.050 70.470 26.220 ;
        RECT 70.710 26.185 70.860 26.355 ;
        RECT 71.100 26.185 71.250 26.355 ;
        RECT 71.490 26.050 71.640 26.220 ;
        RECT 73.220 26.050 73.370 26.220 ;
        RECT 73.610 26.185 73.760 26.355 ;
        RECT 74.000 26.185 74.150 26.355 ;
        RECT 74.390 26.050 74.540 26.220 ;
        RECT 76.120 26.050 76.270 26.220 ;
        RECT 76.510 26.185 76.660 26.355 ;
        RECT 76.900 26.185 77.050 26.355 ;
        RECT 77.290 26.050 77.440 26.220 ;
        RECT 79.020 26.050 79.170 26.220 ;
        RECT 79.410 26.185 79.560 26.355 ;
        RECT 79.800 26.185 79.950 26.355 ;
        RECT 80.190 26.050 80.340 26.220 ;
        RECT 81.920 26.050 82.070 26.220 ;
        RECT 82.310 26.185 82.460 26.355 ;
        RECT 82.700 26.185 82.850 26.355 ;
        RECT 83.090 26.050 83.240 26.220 ;
        RECT 84.820 26.050 84.970 26.220 ;
        RECT 85.210 26.185 85.360 26.355 ;
        RECT 85.600 26.185 85.750 26.355 ;
        RECT 85.990 26.050 86.140 26.220 ;
        RECT 87.720 26.050 87.870 26.220 ;
        RECT 88.110 26.185 88.260 26.355 ;
        RECT 88.500 26.185 88.650 26.355 ;
        RECT 88.890 26.050 89.040 26.220 ;
        RECT 90.620 26.050 90.770 26.220 ;
        RECT 91.010 26.185 91.160 26.355 ;
        RECT 91.400 26.185 91.550 26.355 ;
        RECT 91.790 26.050 91.940 26.220 ;
        RECT 0.985 25.965 1.035 26.000 ;
        POLYGON 1.035 26.000 1.070 25.965 1.035 25.965 ;
        RECT 0.985 25.840 1.070 25.965 ;
        RECT 1.690 25.840 1.775 26.000 ;
        RECT 3.885 25.965 3.935 26.000 ;
        POLYGON 3.935 26.000 3.970 25.965 3.935 25.965 ;
        RECT 3.885 25.840 3.970 25.965 ;
        RECT 4.590 25.840 4.675 26.000 ;
        RECT 6.785 25.965 6.835 26.000 ;
        POLYGON 6.835 26.000 6.870 25.965 6.835 25.965 ;
        RECT 6.785 25.840 6.870 25.965 ;
        RECT 7.490 25.840 7.575 26.000 ;
        RECT 9.685 25.965 9.735 26.000 ;
        POLYGON 9.735 26.000 9.770 25.965 9.735 25.965 ;
        RECT 9.685 25.840 9.770 25.965 ;
        RECT 10.390 25.840 10.475 26.000 ;
        RECT 12.585 25.965 12.635 26.000 ;
        POLYGON 12.635 26.000 12.670 25.965 12.635 25.965 ;
        RECT 12.585 25.840 12.670 25.965 ;
        RECT 13.290 25.840 13.375 26.000 ;
        RECT 15.485 25.965 15.535 26.000 ;
        POLYGON 15.535 26.000 15.570 25.965 15.535 25.965 ;
        RECT 15.485 25.840 15.570 25.965 ;
        RECT 16.190 25.840 16.275 26.000 ;
        RECT 18.385 25.965 18.435 26.000 ;
        POLYGON 18.435 26.000 18.470 25.965 18.435 25.965 ;
        RECT 18.385 25.840 18.470 25.965 ;
        RECT 19.090 25.840 19.175 26.000 ;
        RECT 21.285 25.965 21.335 26.000 ;
        POLYGON 21.335 26.000 21.370 25.965 21.335 25.965 ;
        RECT 21.285 25.840 21.370 25.965 ;
        RECT 21.990 25.840 22.075 26.000 ;
        RECT 24.185 25.965 24.235 26.000 ;
        POLYGON 24.235 26.000 24.270 25.965 24.235 25.965 ;
        RECT 24.185 25.840 24.270 25.965 ;
        RECT 24.890 25.840 24.975 26.000 ;
        RECT 27.085 25.965 27.135 26.000 ;
        POLYGON 27.135 26.000 27.170 25.965 27.135 25.965 ;
        RECT 27.085 25.840 27.170 25.965 ;
        RECT 27.790 25.840 27.875 26.000 ;
        RECT 29.985 25.965 30.035 26.000 ;
        POLYGON 30.035 26.000 30.070 25.965 30.035 25.965 ;
        RECT 29.985 25.840 30.070 25.965 ;
        RECT 30.690 25.840 30.775 26.000 ;
        RECT 32.885 25.965 32.935 26.000 ;
        POLYGON 32.935 26.000 32.970 25.965 32.935 25.965 ;
        RECT 32.885 25.840 32.970 25.965 ;
        RECT 33.590 25.840 33.675 26.000 ;
        RECT 35.785 25.965 35.835 26.000 ;
        POLYGON 35.835 26.000 35.870 25.965 35.835 25.965 ;
        RECT 35.785 25.840 35.870 25.965 ;
        RECT 36.490 25.840 36.575 26.000 ;
        RECT 38.685 25.965 38.735 26.000 ;
        POLYGON 38.735 26.000 38.770 25.965 38.735 25.965 ;
        RECT 38.685 25.840 38.770 25.965 ;
        RECT 39.390 25.840 39.475 26.000 ;
        RECT 41.585 25.965 41.635 26.000 ;
        POLYGON 41.635 26.000 41.670 25.965 41.635 25.965 ;
        RECT 41.585 25.840 41.670 25.965 ;
        RECT 42.290 25.840 42.375 26.000 ;
        RECT 44.485 25.965 44.535 26.000 ;
        POLYGON 44.535 26.000 44.570 25.965 44.535 25.965 ;
        RECT 44.485 25.840 44.570 25.965 ;
        RECT 45.190 25.840 45.275 26.000 ;
        RECT 47.385 25.965 47.435 26.000 ;
        POLYGON 47.435 26.000 47.470 25.965 47.435 25.965 ;
        RECT 47.385 25.840 47.470 25.965 ;
        RECT 48.090 25.840 48.175 26.000 ;
        RECT 50.285 25.965 50.335 26.000 ;
        POLYGON 50.335 26.000 50.370 25.965 50.335 25.965 ;
        RECT 50.285 25.840 50.370 25.965 ;
        RECT 50.990 25.840 51.075 26.000 ;
        RECT 53.185 25.965 53.235 26.000 ;
        POLYGON 53.235 26.000 53.270 25.965 53.235 25.965 ;
        RECT 53.185 25.840 53.270 25.965 ;
        RECT 53.890 25.840 53.975 26.000 ;
        RECT 56.085 25.965 56.135 26.000 ;
        POLYGON 56.135 26.000 56.170 25.965 56.135 25.965 ;
        RECT 56.085 25.840 56.170 25.965 ;
        RECT 56.790 25.840 56.875 26.000 ;
        RECT 58.985 25.965 59.035 26.000 ;
        POLYGON 59.035 26.000 59.070 25.965 59.035 25.965 ;
        RECT 58.985 25.840 59.070 25.965 ;
        RECT 59.690 25.840 59.775 26.000 ;
        RECT 61.885 25.965 61.935 26.000 ;
        POLYGON 61.935 26.000 61.970 25.965 61.935 25.965 ;
        RECT 61.885 25.840 61.970 25.965 ;
        RECT 62.590 25.840 62.675 26.000 ;
        RECT 64.785 25.965 64.835 26.000 ;
        POLYGON 64.835 26.000 64.870 25.965 64.835 25.965 ;
        RECT 64.785 25.840 64.870 25.965 ;
        RECT 65.490 25.840 65.575 26.000 ;
        RECT 67.685 25.965 67.735 26.000 ;
        POLYGON 67.735 26.000 67.770 25.965 67.735 25.965 ;
        RECT 67.685 25.840 67.770 25.965 ;
        RECT 68.390 25.840 68.475 26.000 ;
        RECT 70.585 25.965 70.635 26.000 ;
        POLYGON 70.635 26.000 70.670 25.965 70.635 25.965 ;
        RECT 70.585 25.840 70.670 25.965 ;
        RECT 71.290 25.840 71.375 26.000 ;
        RECT 73.485 25.965 73.535 26.000 ;
        POLYGON 73.535 26.000 73.570 25.965 73.535 25.965 ;
        RECT 73.485 25.840 73.570 25.965 ;
        RECT 74.190 25.840 74.275 26.000 ;
        RECT 76.385 25.965 76.435 26.000 ;
        POLYGON 76.435 26.000 76.470 25.965 76.435 25.965 ;
        RECT 76.385 25.840 76.470 25.965 ;
        RECT 77.090 25.840 77.175 26.000 ;
        RECT 79.285 25.965 79.335 26.000 ;
        POLYGON 79.335 26.000 79.370 25.965 79.335 25.965 ;
        RECT 79.285 25.840 79.370 25.965 ;
        RECT 79.990 25.840 80.075 26.000 ;
        RECT 82.185 25.965 82.235 26.000 ;
        POLYGON 82.235 26.000 82.270 25.965 82.235 25.965 ;
        RECT 82.185 25.840 82.270 25.965 ;
        RECT 82.890 25.840 82.975 26.000 ;
        RECT 85.085 25.965 85.135 26.000 ;
        POLYGON 85.135 26.000 85.170 25.965 85.135 25.965 ;
        RECT 85.085 25.840 85.170 25.965 ;
        RECT 85.790 25.840 85.875 26.000 ;
        RECT 87.985 25.965 88.035 26.000 ;
        POLYGON 88.035 26.000 88.070 25.965 88.035 25.965 ;
        RECT 87.985 25.840 88.070 25.965 ;
        RECT 88.690 25.840 88.775 26.000 ;
        RECT 90.885 25.965 90.935 26.000 ;
        POLYGON 90.935 26.000 90.970 25.965 90.935 25.965 ;
        RECT 90.885 25.840 90.970 25.965 ;
        RECT 91.590 25.840 91.675 26.000 ;
        RECT 0.775 25.220 0.850 25.360 ;
        RECT 0.990 25.170 1.065 25.310 ;
        RECT 1.695 25.230 1.755 25.310 ;
        POLYGON 1.695 25.230 1.755 25.230 1.755 25.170 ;
        RECT 1.910 25.220 1.985 25.360 ;
        RECT 3.675 25.220 3.750 25.360 ;
        RECT 3.890 25.170 3.965 25.310 ;
        RECT 4.595 25.230 4.655 25.310 ;
        POLYGON 4.595 25.230 4.655 25.230 4.655 25.170 ;
        RECT 4.810 25.220 4.885 25.360 ;
        RECT 6.575 25.220 6.650 25.360 ;
        RECT 6.790 25.170 6.865 25.310 ;
        RECT 7.495 25.230 7.555 25.310 ;
        POLYGON 7.495 25.230 7.555 25.230 7.555 25.170 ;
        RECT 7.710 25.220 7.785 25.360 ;
        RECT 9.475 25.220 9.550 25.360 ;
        RECT 9.690 25.170 9.765 25.310 ;
        RECT 10.395 25.230 10.455 25.310 ;
        POLYGON 10.395 25.230 10.455 25.230 10.455 25.170 ;
        RECT 10.610 25.220 10.685 25.360 ;
        RECT 12.375 25.220 12.450 25.360 ;
        RECT 12.590 25.170 12.665 25.310 ;
        RECT 13.295 25.230 13.355 25.310 ;
        POLYGON 13.295 25.230 13.355 25.230 13.355 25.170 ;
        RECT 13.510 25.220 13.585 25.360 ;
        RECT 15.275 25.220 15.350 25.360 ;
        RECT 15.490 25.170 15.565 25.310 ;
        RECT 16.195 25.230 16.255 25.310 ;
        POLYGON 16.195 25.230 16.255 25.230 16.255 25.170 ;
        RECT 16.410 25.220 16.485 25.360 ;
        RECT 18.175 25.220 18.250 25.360 ;
        RECT 18.390 25.170 18.465 25.310 ;
        RECT 19.095 25.230 19.155 25.310 ;
        POLYGON 19.095 25.230 19.155 25.230 19.155 25.170 ;
        RECT 19.310 25.220 19.385 25.360 ;
        RECT 21.075 25.220 21.150 25.360 ;
        RECT 21.290 25.170 21.365 25.310 ;
        RECT 21.995 25.230 22.055 25.310 ;
        POLYGON 21.995 25.230 22.055 25.230 22.055 25.170 ;
        RECT 22.210 25.220 22.285 25.360 ;
        RECT 23.975 25.220 24.050 25.360 ;
        RECT 24.190 25.170 24.265 25.310 ;
        RECT 24.895 25.230 24.955 25.310 ;
        POLYGON 24.895 25.230 24.955 25.230 24.955 25.170 ;
        RECT 25.110 25.220 25.185 25.360 ;
        RECT 26.875 25.220 26.950 25.360 ;
        RECT 27.090 25.170 27.165 25.310 ;
        RECT 27.795 25.230 27.855 25.310 ;
        POLYGON 27.795 25.230 27.855 25.230 27.855 25.170 ;
        RECT 28.010 25.220 28.085 25.360 ;
        RECT 29.775 25.220 29.850 25.360 ;
        RECT 29.990 25.170 30.065 25.310 ;
        RECT 30.695 25.230 30.755 25.310 ;
        POLYGON 30.695 25.230 30.755 25.230 30.755 25.170 ;
        RECT 30.910 25.220 30.985 25.360 ;
        RECT 32.675 25.220 32.750 25.360 ;
        RECT 32.890 25.170 32.965 25.310 ;
        RECT 33.595 25.230 33.655 25.310 ;
        POLYGON 33.595 25.230 33.655 25.230 33.655 25.170 ;
        RECT 33.810 25.220 33.885 25.360 ;
        RECT 35.575 25.220 35.650 25.360 ;
        RECT 35.790 25.170 35.865 25.310 ;
        RECT 36.495 25.230 36.555 25.310 ;
        POLYGON 36.495 25.230 36.555 25.230 36.555 25.170 ;
        RECT 36.710 25.220 36.785 25.360 ;
        RECT 38.475 25.220 38.550 25.360 ;
        RECT 38.690 25.170 38.765 25.310 ;
        RECT 39.395 25.230 39.455 25.310 ;
        POLYGON 39.395 25.230 39.455 25.230 39.455 25.170 ;
        RECT 39.610 25.220 39.685 25.360 ;
        RECT 41.375 25.220 41.450 25.360 ;
        RECT 41.590 25.170 41.665 25.310 ;
        RECT 42.295 25.230 42.355 25.310 ;
        POLYGON 42.295 25.230 42.355 25.230 42.355 25.170 ;
        RECT 42.510 25.220 42.585 25.360 ;
        RECT 44.275 25.220 44.350 25.360 ;
        RECT 44.490 25.170 44.565 25.310 ;
        RECT 45.195 25.230 45.255 25.310 ;
        POLYGON 45.195 25.230 45.255 25.230 45.255 25.170 ;
        RECT 45.410 25.220 45.485 25.360 ;
        RECT 47.175 25.220 47.250 25.360 ;
        RECT 47.390 25.170 47.465 25.310 ;
        RECT 48.095 25.230 48.155 25.310 ;
        POLYGON 48.095 25.230 48.155 25.230 48.155 25.170 ;
        RECT 48.310 25.220 48.385 25.360 ;
        RECT 50.075 25.220 50.150 25.360 ;
        RECT 50.290 25.170 50.365 25.310 ;
        RECT 50.995 25.230 51.055 25.310 ;
        POLYGON 50.995 25.230 51.055 25.230 51.055 25.170 ;
        RECT 51.210 25.220 51.285 25.360 ;
        RECT 52.975 25.220 53.050 25.360 ;
        RECT 53.190 25.170 53.265 25.310 ;
        RECT 53.895 25.230 53.955 25.310 ;
        POLYGON 53.895 25.230 53.955 25.230 53.955 25.170 ;
        RECT 54.110 25.220 54.185 25.360 ;
        RECT 55.875 25.220 55.950 25.360 ;
        RECT 56.090 25.170 56.165 25.310 ;
        RECT 56.795 25.230 56.855 25.310 ;
        POLYGON 56.795 25.230 56.855 25.230 56.855 25.170 ;
        RECT 57.010 25.220 57.085 25.360 ;
        RECT 58.775 25.220 58.850 25.360 ;
        RECT 58.990 25.170 59.065 25.310 ;
        RECT 59.695 25.230 59.755 25.310 ;
        POLYGON 59.695 25.230 59.755 25.230 59.755 25.170 ;
        RECT 59.910 25.220 59.985 25.360 ;
        RECT 61.675 25.220 61.750 25.360 ;
        RECT 61.890 25.170 61.965 25.310 ;
        RECT 62.595 25.230 62.655 25.310 ;
        POLYGON 62.595 25.230 62.655 25.230 62.655 25.170 ;
        RECT 62.810 25.220 62.885 25.360 ;
        RECT 64.575 25.220 64.650 25.360 ;
        RECT 64.790 25.170 64.865 25.310 ;
        RECT 65.495 25.230 65.555 25.310 ;
        POLYGON 65.495 25.230 65.555 25.230 65.555 25.170 ;
        RECT 65.710 25.220 65.785 25.360 ;
        RECT 67.475 25.220 67.550 25.360 ;
        RECT 67.690 25.170 67.765 25.310 ;
        RECT 68.395 25.230 68.455 25.310 ;
        POLYGON 68.395 25.230 68.455 25.230 68.455 25.170 ;
        RECT 68.610 25.220 68.685 25.360 ;
        RECT 70.375 25.220 70.450 25.360 ;
        RECT 70.590 25.170 70.665 25.310 ;
        RECT 71.295 25.230 71.355 25.310 ;
        POLYGON 71.295 25.230 71.355 25.230 71.355 25.170 ;
        RECT 71.510 25.220 71.585 25.360 ;
        RECT 73.275 25.220 73.350 25.360 ;
        RECT 73.490 25.170 73.565 25.310 ;
        RECT 74.195 25.230 74.255 25.310 ;
        POLYGON 74.195 25.230 74.255 25.230 74.255 25.170 ;
        RECT 74.410 25.220 74.485 25.360 ;
        RECT 76.175 25.220 76.250 25.360 ;
        RECT 76.390 25.170 76.465 25.310 ;
        RECT 77.095 25.230 77.155 25.310 ;
        POLYGON 77.095 25.230 77.155 25.230 77.155 25.170 ;
        RECT 77.310 25.220 77.385 25.360 ;
        RECT 79.075 25.220 79.150 25.360 ;
        RECT 79.290 25.170 79.365 25.310 ;
        RECT 79.995 25.230 80.055 25.310 ;
        POLYGON 79.995 25.230 80.055 25.230 80.055 25.170 ;
        RECT 80.210 25.220 80.285 25.360 ;
        RECT 81.975 25.220 82.050 25.360 ;
        RECT 82.190 25.170 82.265 25.310 ;
        RECT 82.895 25.230 82.955 25.310 ;
        POLYGON 82.895 25.230 82.955 25.230 82.955 25.170 ;
        RECT 83.110 25.220 83.185 25.360 ;
        RECT 84.875 25.220 84.950 25.360 ;
        RECT 85.090 25.170 85.165 25.310 ;
        RECT 85.795 25.230 85.855 25.310 ;
        POLYGON 85.795 25.230 85.855 25.230 85.855 25.170 ;
        RECT 86.010 25.220 86.085 25.360 ;
        RECT 87.775 25.220 87.850 25.360 ;
        RECT 87.990 25.170 88.065 25.310 ;
        RECT 88.695 25.230 88.755 25.310 ;
        POLYGON 88.695 25.230 88.755 25.230 88.755 25.170 ;
        RECT 88.910 25.220 88.985 25.360 ;
        RECT 90.675 25.220 90.750 25.360 ;
        RECT 90.890 25.170 90.965 25.310 ;
        RECT 91.595 25.230 91.655 25.310 ;
        POLYGON 91.595 25.230 91.655 25.230 91.655 25.170 ;
        RECT 91.810 25.220 91.885 25.360 ;
        RECT 0.720 24.700 0.870 24.870 ;
        RECT 1.110 24.835 1.260 25.005 ;
        RECT 1.500 24.835 1.650 25.005 ;
        RECT 1.890 24.700 2.040 24.870 ;
        RECT 3.620 24.700 3.770 24.870 ;
        RECT 4.010 24.835 4.160 25.005 ;
        RECT 4.400 24.835 4.550 25.005 ;
        RECT 4.790 24.700 4.940 24.870 ;
        RECT 6.520 24.700 6.670 24.870 ;
        RECT 6.910 24.835 7.060 25.005 ;
        RECT 7.300 24.835 7.450 25.005 ;
        RECT 7.690 24.700 7.840 24.870 ;
        RECT 9.420 24.700 9.570 24.870 ;
        RECT 9.810 24.835 9.960 25.005 ;
        RECT 10.200 24.835 10.350 25.005 ;
        RECT 10.590 24.700 10.740 24.870 ;
        RECT 12.320 24.700 12.470 24.870 ;
        RECT 12.710 24.835 12.860 25.005 ;
        RECT 13.100 24.835 13.250 25.005 ;
        RECT 13.490 24.700 13.640 24.870 ;
        RECT 15.220 24.700 15.370 24.870 ;
        RECT 15.610 24.835 15.760 25.005 ;
        RECT 16.000 24.835 16.150 25.005 ;
        RECT 16.390 24.700 16.540 24.870 ;
        RECT 18.120 24.700 18.270 24.870 ;
        RECT 18.510 24.835 18.660 25.005 ;
        RECT 18.900 24.835 19.050 25.005 ;
        RECT 19.290 24.700 19.440 24.870 ;
        RECT 21.020 24.700 21.170 24.870 ;
        RECT 21.410 24.835 21.560 25.005 ;
        RECT 21.800 24.835 21.950 25.005 ;
        RECT 22.190 24.700 22.340 24.870 ;
        RECT 23.920 24.700 24.070 24.870 ;
        RECT 24.310 24.835 24.460 25.005 ;
        RECT 24.700 24.835 24.850 25.005 ;
        RECT 25.090 24.700 25.240 24.870 ;
        RECT 26.820 24.700 26.970 24.870 ;
        RECT 27.210 24.835 27.360 25.005 ;
        RECT 27.600 24.835 27.750 25.005 ;
        RECT 27.990 24.700 28.140 24.870 ;
        RECT 29.720 24.700 29.870 24.870 ;
        RECT 30.110 24.835 30.260 25.005 ;
        RECT 30.500 24.835 30.650 25.005 ;
        RECT 30.890 24.700 31.040 24.870 ;
        RECT 32.620 24.700 32.770 24.870 ;
        RECT 33.010 24.835 33.160 25.005 ;
        RECT 33.400 24.835 33.550 25.005 ;
        RECT 33.790 24.700 33.940 24.870 ;
        RECT 35.520 24.700 35.670 24.870 ;
        RECT 35.910 24.835 36.060 25.005 ;
        RECT 36.300 24.835 36.450 25.005 ;
        RECT 36.690 24.700 36.840 24.870 ;
        RECT 38.420 24.700 38.570 24.870 ;
        RECT 38.810 24.835 38.960 25.005 ;
        RECT 39.200 24.835 39.350 25.005 ;
        RECT 39.590 24.700 39.740 24.870 ;
        RECT 41.320 24.700 41.470 24.870 ;
        RECT 41.710 24.835 41.860 25.005 ;
        RECT 42.100 24.835 42.250 25.005 ;
        RECT 42.490 24.700 42.640 24.870 ;
        RECT 44.220 24.700 44.370 24.870 ;
        RECT 44.610 24.835 44.760 25.005 ;
        RECT 45.000 24.835 45.150 25.005 ;
        RECT 45.390 24.700 45.540 24.870 ;
        RECT 47.120 24.700 47.270 24.870 ;
        RECT 47.510 24.835 47.660 25.005 ;
        RECT 47.900 24.835 48.050 25.005 ;
        RECT 48.290 24.700 48.440 24.870 ;
        RECT 50.020 24.700 50.170 24.870 ;
        RECT 50.410 24.835 50.560 25.005 ;
        RECT 50.800 24.835 50.950 25.005 ;
        RECT 51.190 24.700 51.340 24.870 ;
        RECT 52.920 24.700 53.070 24.870 ;
        RECT 53.310 24.835 53.460 25.005 ;
        RECT 53.700 24.835 53.850 25.005 ;
        RECT 54.090 24.700 54.240 24.870 ;
        RECT 55.820 24.700 55.970 24.870 ;
        RECT 56.210 24.835 56.360 25.005 ;
        RECT 56.600 24.835 56.750 25.005 ;
        RECT 56.990 24.700 57.140 24.870 ;
        RECT 58.720 24.700 58.870 24.870 ;
        RECT 59.110 24.835 59.260 25.005 ;
        RECT 59.500 24.835 59.650 25.005 ;
        RECT 59.890 24.700 60.040 24.870 ;
        RECT 61.620 24.700 61.770 24.870 ;
        RECT 62.010 24.835 62.160 25.005 ;
        RECT 62.400 24.835 62.550 25.005 ;
        RECT 62.790 24.700 62.940 24.870 ;
        RECT 64.520 24.700 64.670 24.870 ;
        RECT 64.910 24.835 65.060 25.005 ;
        RECT 65.300 24.835 65.450 25.005 ;
        RECT 65.690 24.700 65.840 24.870 ;
        RECT 67.420 24.700 67.570 24.870 ;
        RECT 67.810 24.835 67.960 25.005 ;
        RECT 68.200 24.835 68.350 25.005 ;
        RECT 68.590 24.700 68.740 24.870 ;
        RECT 70.320 24.700 70.470 24.870 ;
        RECT 70.710 24.835 70.860 25.005 ;
        RECT 71.100 24.835 71.250 25.005 ;
        RECT 71.490 24.700 71.640 24.870 ;
        RECT 73.220 24.700 73.370 24.870 ;
        RECT 73.610 24.835 73.760 25.005 ;
        RECT 74.000 24.835 74.150 25.005 ;
        RECT 74.390 24.700 74.540 24.870 ;
        RECT 76.120 24.700 76.270 24.870 ;
        RECT 76.510 24.835 76.660 25.005 ;
        RECT 76.900 24.835 77.050 25.005 ;
        RECT 77.290 24.700 77.440 24.870 ;
        RECT 79.020 24.700 79.170 24.870 ;
        RECT 79.410 24.835 79.560 25.005 ;
        RECT 79.800 24.835 79.950 25.005 ;
        RECT 80.190 24.700 80.340 24.870 ;
        RECT 81.920 24.700 82.070 24.870 ;
        RECT 82.310 24.835 82.460 25.005 ;
        RECT 82.700 24.835 82.850 25.005 ;
        RECT 83.090 24.700 83.240 24.870 ;
        RECT 84.820 24.700 84.970 24.870 ;
        RECT 85.210 24.835 85.360 25.005 ;
        RECT 85.600 24.835 85.750 25.005 ;
        RECT 85.990 24.700 86.140 24.870 ;
        RECT 87.720 24.700 87.870 24.870 ;
        RECT 88.110 24.835 88.260 25.005 ;
        RECT 88.500 24.835 88.650 25.005 ;
        RECT 88.890 24.700 89.040 24.870 ;
        RECT 90.620 24.700 90.770 24.870 ;
        RECT 91.010 24.835 91.160 25.005 ;
        RECT 91.400 24.835 91.550 25.005 ;
        RECT 91.790 24.700 91.940 24.870 ;
        RECT 0.985 24.615 1.035 24.650 ;
        POLYGON 1.035 24.650 1.070 24.615 1.035 24.615 ;
        RECT 0.985 24.490 1.070 24.615 ;
        RECT 1.690 24.490 1.775 24.650 ;
        RECT 3.885 24.615 3.935 24.650 ;
        POLYGON 3.935 24.650 3.970 24.615 3.935 24.615 ;
        RECT 3.885 24.490 3.970 24.615 ;
        RECT 4.590 24.490 4.675 24.650 ;
        RECT 6.785 24.615 6.835 24.650 ;
        POLYGON 6.835 24.650 6.870 24.615 6.835 24.615 ;
        RECT 6.785 24.490 6.870 24.615 ;
        RECT 7.490 24.490 7.575 24.650 ;
        RECT 9.685 24.615 9.735 24.650 ;
        POLYGON 9.735 24.650 9.770 24.615 9.735 24.615 ;
        RECT 9.685 24.490 9.770 24.615 ;
        RECT 10.390 24.490 10.475 24.650 ;
        RECT 12.585 24.615 12.635 24.650 ;
        POLYGON 12.635 24.650 12.670 24.615 12.635 24.615 ;
        RECT 12.585 24.490 12.670 24.615 ;
        RECT 13.290 24.490 13.375 24.650 ;
        RECT 15.485 24.615 15.535 24.650 ;
        POLYGON 15.535 24.650 15.570 24.615 15.535 24.615 ;
        RECT 15.485 24.490 15.570 24.615 ;
        RECT 16.190 24.490 16.275 24.650 ;
        RECT 18.385 24.615 18.435 24.650 ;
        POLYGON 18.435 24.650 18.470 24.615 18.435 24.615 ;
        RECT 18.385 24.490 18.470 24.615 ;
        RECT 19.090 24.490 19.175 24.650 ;
        RECT 21.285 24.615 21.335 24.650 ;
        POLYGON 21.335 24.650 21.370 24.615 21.335 24.615 ;
        RECT 21.285 24.490 21.370 24.615 ;
        RECT 21.990 24.490 22.075 24.650 ;
        RECT 24.185 24.615 24.235 24.650 ;
        POLYGON 24.235 24.650 24.270 24.615 24.235 24.615 ;
        RECT 24.185 24.490 24.270 24.615 ;
        RECT 24.890 24.490 24.975 24.650 ;
        RECT 27.085 24.615 27.135 24.650 ;
        POLYGON 27.135 24.650 27.170 24.615 27.135 24.615 ;
        RECT 27.085 24.490 27.170 24.615 ;
        RECT 27.790 24.490 27.875 24.650 ;
        RECT 29.985 24.615 30.035 24.650 ;
        POLYGON 30.035 24.650 30.070 24.615 30.035 24.615 ;
        RECT 29.985 24.490 30.070 24.615 ;
        RECT 30.690 24.490 30.775 24.650 ;
        RECT 32.885 24.615 32.935 24.650 ;
        POLYGON 32.935 24.650 32.970 24.615 32.935 24.615 ;
        RECT 32.885 24.490 32.970 24.615 ;
        RECT 33.590 24.490 33.675 24.650 ;
        RECT 35.785 24.615 35.835 24.650 ;
        POLYGON 35.835 24.650 35.870 24.615 35.835 24.615 ;
        RECT 35.785 24.490 35.870 24.615 ;
        RECT 36.490 24.490 36.575 24.650 ;
        RECT 38.685 24.615 38.735 24.650 ;
        POLYGON 38.735 24.650 38.770 24.615 38.735 24.615 ;
        RECT 38.685 24.490 38.770 24.615 ;
        RECT 39.390 24.490 39.475 24.650 ;
        RECT 41.585 24.615 41.635 24.650 ;
        POLYGON 41.635 24.650 41.670 24.615 41.635 24.615 ;
        RECT 41.585 24.490 41.670 24.615 ;
        RECT 42.290 24.490 42.375 24.650 ;
        RECT 44.485 24.615 44.535 24.650 ;
        POLYGON 44.535 24.650 44.570 24.615 44.535 24.615 ;
        RECT 44.485 24.490 44.570 24.615 ;
        RECT 45.190 24.490 45.275 24.650 ;
        RECT 47.385 24.615 47.435 24.650 ;
        POLYGON 47.435 24.650 47.470 24.615 47.435 24.615 ;
        RECT 47.385 24.490 47.470 24.615 ;
        RECT 48.090 24.490 48.175 24.650 ;
        RECT 50.285 24.615 50.335 24.650 ;
        POLYGON 50.335 24.650 50.370 24.615 50.335 24.615 ;
        RECT 50.285 24.490 50.370 24.615 ;
        RECT 50.990 24.490 51.075 24.650 ;
        RECT 53.185 24.615 53.235 24.650 ;
        POLYGON 53.235 24.650 53.270 24.615 53.235 24.615 ;
        RECT 53.185 24.490 53.270 24.615 ;
        RECT 53.890 24.490 53.975 24.650 ;
        RECT 56.085 24.615 56.135 24.650 ;
        POLYGON 56.135 24.650 56.170 24.615 56.135 24.615 ;
        RECT 56.085 24.490 56.170 24.615 ;
        RECT 56.790 24.490 56.875 24.650 ;
        RECT 58.985 24.615 59.035 24.650 ;
        POLYGON 59.035 24.650 59.070 24.615 59.035 24.615 ;
        RECT 58.985 24.490 59.070 24.615 ;
        RECT 59.690 24.490 59.775 24.650 ;
        RECT 61.885 24.615 61.935 24.650 ;
        POLYGON 61.935 24.650 61.970 24.615 61.935 24.615 ;
        RECT 61.885 24.490 61.970 24.615 ;
        RECT 62.590 24.490 62.675 24.650 ;
        RECT 64.785 24.615 64.835 24.650 ;
        POLYGON 64.835 24.650 64.870 24.615 64.835 24.615 ;
        RECT 64.785 24.490 64.870 24.615 ;
        RECT 65.490 24.490 65.575 24.650 ;
        RECT 67.685 24.615 67.735 24.650 ;
        POLYGON 67.735 24.650 67.770 24.615 67.735 24.615 ;
        RECT 67.685 24.490 67.770 24.615 ;
        RECT 68.390 24.490 68.475 24.650 ;
        RECT 70.585 24.615 70.635 24.650 ;
        POLYGON 70.635 24.650 70.670 24.615 70.635 24.615 ;
        RECT 70.585 24.490 70.670 24.615 ;
        RECT 71.290 24.490 71.375 24.650 ;
        RECT 73.485 24.615 73.535 24.650 ;
        POLYGON 73.535 24.650 73.570 24.615 73.535 24.615 ;
        RECT 73.485 24.490 73.570 24.615 ;
        RECT 74.190 24.490 74.275 24.650 ;
        RECT 76.385 24.615 76.435 24.650 ;
        POLYGON 76.435 24.650 76.470 24.615 76.435 24.615 ;
        RECT 76.385 24.490 76.470 24.615 ;
        RECT 77.090 24.490 77.175 24.650 ;
        RECT 79.285 24.615 79.335 24.650 ;
        POLYGON 79.335 24.650 79.370 24.615 79.335 24.615 ;
        RECT 79.285 24.490 79.370 24.615 ;
        RECT 79.990 24.490 80.075 24.650 ;
        RECT 82.185 24.615 82.235 24.650 ;
        POLYGON 82.235 24.650 82.270 24.615 82.235 24.615 ;
        RECT 82.185 24.490 82.270 24.615 ;
        RECT 82.890 24.490 82.975 24.650 ;
        RECT 85.085 24.615 85.135 24.650 ;
        POLYGON 85.135 24.650 85.170 24.615 85.135 24.615 ;
        RECT 85.085 24.490 85.170 24.615 ;
        RECT 85.790 24.490 85.875 24.650 ;
        RECT 87.985 24.615 88.035 24.650 ;
        POLYGON 88.035 24.650 88.070 24.615 88.035 24.615 ;
        RECT 87.985 24.490 88.070 24.615 ;
        RECT 88.690 24.490 88.775 24.650 ;
        RECT 90.885 24.615 90.935 24.650 ;
        POLYGON 90.935 24.650 90.970 24.615 90.935 24.615 ;
        RECT 90.885 24.490 90.970 24.615 ;
        RECT 91.590 24.490 91.675 24.650 ;
        RECT 0.775 23.870 0.850 24.010 ;
        RECT 0.990 23.820 1.065 23.960 ;
        RECT 1.695 23.880 1.755 23.960 ;
        POLYGON 1.695 23.880 1.755 23.880 1.755 23.820 ;
        RECT 1.910 23.870 1.985 24.010 ;
        RECT 3.675 23.870 3.750 24.010 ;
        RECT 3.890 23.820 3.965 23.960 ;
        RECT 4.595 23.880 4.655 23.960 ;
        POLYGON 4.595 23.880 4.655 23.880 4.655 23.820 ;
        RECT 4.810 23.870 4.885 24.010 ;
        RECT 6.575 23.870 6.650 24.010 ;
        RECT 6.790 23.820 6.865 23.960 ;
        RECT 7.495 23.880 7.555 23.960 ;
        POLYGON 7.495 23.880 7.555 23.880 7.555 23.820 ;
        RECT 7.710 23.870 7.785 24.010 ;
        RECT 9.475 23.870 9.550 24.010 ;
        RECT 9.690 23.820 9.765 23.960 ;
        RECT 10.395 23.880 10.455 23.960 ;
        POLYGON 10.395 23.880 10.455 23.880 10.455 23.820 ;
        RECT 10.610 23.870 10.685 24.010 ;
        RECT 12.375 23.870 12.450 24.010 ;
        RECT 12.590 23.820 12.665 23.960 ;
        RECT 13.295 23.880 13.355 23.960 ;
        POLYGON 13.295 23.880 13.355 23.880 13.355 23.820 ;
        RECT 13.510 23.870 13.585 24.010 ;
        RECT 15.275 23.870 15.350 24.010 ;
        RECT 15.490 23.820 15.565 23.960 ;
        RECT 16.195 23.880 16.255 23.960 ;
        POLYGON 16.195 23.880 16.255 23.880 16.255 23.820 ;
        RECT 16.410 23.870 16.485 24.010 ;
        RECT 18.175 23.870 18.250 24.010 ;
        RECT 18.390 23.820 18.465 23.960 ;
        RECT 19.095 23.880 19.155 23.960 ;
        POLYGON 19.095 23.880 19.155 23.880 19.155 23.820 ;
        RECT 19.310 23.870 19.385 24.010 ;
        RECT 21.075 23.870 21.150 24.010 ;
        RECT 21.290 23.820 21.365 23.960 ;
        RECT 21.995 23.880 22.055 23.960 ;
        POLYGON 21.995 23.880 22.055 23.880 22.055 23.820 ;
        RECT 22.210 23.870 22.285 24.010 ;
        RECT 23.975 23.870 24.050 24.010 ;
        RECT 24.190 23.820 24.265 23.960 ;
        RECT 24.895 23.880 24.955 23.960 ;
        POLYGON 24.895 23.880 24.955 23.880 24.955 23.820 ;
        RECT 25.110 23.870 25.185 24.010 ;
        RECT 26.875 23.870 26.950 24.010 ;
        RECT 27.090 23.820 27.165 23.960 ;
        RECT 27.795 23.880 27.855 23.960 ;
        POLYGON 27.795 23.880 27.855 23.880 27.855 23.820 ;
        RECT 28.010 23.870 28.085 24.010 ;
        RECT 29.775 23.870 29.850 24.010 ;
        RECT 29.990 23.820 30.065 23.960 ;
        RECT 30.695 23.880 30.755 23.960 ;
        POLYGON 30.695 23.880 30.755 23.880 30.755 23.820 ;
        RECT 30.910 23.870 30.985 24.010 ;
        RECT 32.675 23.870 32.750 24.010 ;
        RECT 32.890 23.820 32.965 23.960 ;
        RECT 33.595 23.880 33.655 23.960 ;
        POLYGON 33.595 23.880 33.655 23.880 33.655 23.820 ;
        RECT 33.810 23.870 33.885 24.010 ;
        RECT 35.575 23.870 35.650 24.010 ;
        RECT 35.790 23.820 35.865 23.960 ;
        RECT 36.495 23.880 36.555 23.960 ;
        POLYGON 36.495 23.880 36.555 23.880 36.555 23.820 ;
        RECT 36.710 23.870 36.785 24.010 ;
        RECT 38.475 23.870 38.550 24.010 ;
        RECT 38.690 23.820 38.765 23.960 ;
        RECT 39.395 23.880 39.455 23.960 ;
        POLYGON 39.395 23.880 39.455 23.880 39.455 23.820 ;
        RECT 39.610 23.870 39.685 24.010 ;
        RECT 41.375 23.870 41.450 24.010 ;
        RECT 41.590 23.820 41.665 23.960 ;
        RECT 42.295 23.880 42.355 23.960 ;
        POLYGON 42.295 23.880 42.355 23.880 42.355 23.820 ;
        RECT 42.510 23.870 42.585 24.010 ;
        RECT 44.275 23.870 44.350 24.010 ;
        RECT 44.490 23.820 44.565 23.960 ;
        RECT 45.195 23.880 45.255 23.960 ;
        POLYGON 45.195 23.880 45.255 23.880 45.255 23.820 ;
        RECT 45.410 23.870 45.485 24.010 ;
        RECT 47.175 23.870 47.250 24.010 ;
        RECT 47.390 23.820 47.465 23.960 ;
        RECT 48.095 23.880 48.155 23.960 ;
        POLYGON 48.095 23.880 48.155 23.880 48.155 23.820 ;
        RECT 48.310 23.870 48.385 24.010 ;
        RECT 50.075 23.870 50.150 24.010 ;
        RECT 50.290 23.820 50.365 23.960 ;
        RECT 50.995 23.880 51.055 23.960 ;
        POLYGON 50.995 23.880 51.055 23.880 51.055 23.820 ;
        RECT 51.210 23.870 51.285 24.010 ;
        RECT 52.975 23.870 53.050 24.010 ;
        RECT 53.190 23.820 53.265 23.960 ;
        RECT 53.895 23.880 53.955 23.960 ;
        POLYGON 53.895 23.880 53.955 23.880 53.955 23.820 ;
        RECT 54.110 23.870 54.185 24.010 ;
        RECT 55.875 23.870 55.950 24.010 ;
        RECT 56.090 23.820 56.165 23.960 ;
        RECT 56.795 23.880 56.855 23.960 ;
        POLYGON 56.795 23.880 56.855 23.880 56.855 23.820 ;
        RECT 57.010 23.870 57.085 24.010 ;
        RECT 58.775 23.870 58.850 24.010 ;
        RECT 58.990 23.820 59.065 23.960 ;
        RECT 59.695 23.880 59.755 23.960 ;
        POLYGON 59.695 23.880 59.755 23.880 59.755 23.820 ;
        RECT 59.910 23.870 59.985 24.010 ;
        RECT 61.675 23.870 61.750 24.010 ;
        RECT 61.890 23.820 61.965 23.960 ;
        RECT 62.595 23.880 62.655 23.960 ;
        POLYGON 62.595 23.880 62.655 23.880 62.655 23.820 ;
        RECT 62.810 23.870 62.885 24.010 ;
        RECT 64.575 23.870 64.650 24.010 ;
        RECT 64.790 23.820 64.865 23.960 ;
        RECT 65.495 23.880 65.555 23.960 ;
        POLYGON 65.495 23.880 65.555 23.880 65.555 23.820 ;
        RECT 65.710 23.870 65.785 24.010 ;
        RECT 67.475 23.870 67.550 24.010 ;
        RECT 67.690 23.820 67.765 23.960 ;
        RECT 68.395 23.880 68.455 23.960 ;
        POLYGON 68.395 23.880 68.455 23.880 68.455 23.820 ;
        RECT 68.610 23.870 68.685 24.010 ;
        RECT 70.375 23.870 70.450 24.010 ;
        RECT 70.590 23.820 70.665 23.960 ;
        RECT 71.295 23.880 71.355 23.960 ;
        POLYGON 71.295 23.880 71.355 23.880 71.355 23.820 ;
        RECT 71.510 23.870 71.585 24.010 ;
        RECT 73.275 23.870 73.350 24.010 ;
        RECT 73.490 23.820 73.565 23.960 ;
        RECT 74.195 23.880 74.255 23.960 ;
        POLYGON 74.195 23.880 74.255 23.880 74.255 23.820 ;
        RECT 74.410 23.870 74.485 24.010 ;
        RECT 76.175 23.870 76.250 24.010 ;
        RECT 76.390 23.820 76.465 23.960 ;
        RECT 77.095 23.880 77.155 23.960 ;
        POLYGON 77.095 23.880 77.155 23.880 77.155 23.820 ;
        RECT 77.310 23.870 77.385 24.010 ;
        RECT 79.075 23.870 79.150 24.010 ;
        RECT 79.290 23.820 79.365 23.960 ;
        RECT 79.995 23.880 80.055 23.960 ;
        POLYGON 79.995 23.880 80.055 23.880 80.055 23.820 ;
        RECT 80.210 23.870 80.285 24.010 ;
        RECT 81.975 23.870 82.050 24.010 ;
        RECT 82.190 23.820 82.265 23.960 ;
        RECT 82.895 23.880 82.955 23.960 ;
        POLYGON 82.895 23.880 82.955 23.880 82.955 23.820 ;
        RECT 83.110 23.870 83.185 24.010 ;
        RECT 84.875 23.870 84.950 24.010 ;
        RECT 85.090 23.820 85.165 23.960 ;
        RECT 85.795 23.880 85.855 23.960 ;
        POLYGON 85.795 23.880 85.855 23.880 85.855 23.820 ;
        RECT 86.010 23.870 86.085 24.010 ;
        RECT 87.775 23.870 87.850 24.010 ;
        RECT 87.990 23.820 88.065 23.960 ;
        RECT 88.695 23.880 88.755 23.960 ;
        POLYGON 88.695 23.880 88.755 23.880 88.755 23.820 ;
        RECT 88.910 23.870 88.985 24.010 ;
        RECT 90.675 23.870 90.750 24.010 ;
        RECT 90.890 23.820 90.965 23.960 ;
        RECT 91.595 23.880 91.655 23.960 ;
        POLYGON 91.595 23.880 91.655 23.880 91.655 23.820 ;
        RECT 91.810 23.870 91.885 24.010 ;
        RECT 0.720 23.350 0.870 23.520 ;
        RECT 1.110 23.485 1.260 23.655 ;
        RECT 1.500 23.485 1.650 23.655 ;
        RECT 1.890 23.350 2.040 23.520 ;
        RECT 3.620 23.350 3.770 23.520 ;
        RECT 4.010 23.485 4.160 23.655 ;
        RECT 4.400 23.485 4.550 23.655 ;
        RECT 4.790 23.350 4.940 23.520 ;
        RECT 6.520 23.350 6.670 23.520 ;
        RECT 6.910 23.485 7.060 23.655 ;
        RECT 7.300 23.485 7.450 23.655 ;
        RECT 7.690 23.350 7.840 23.520 ;
        RECT 9.420 23.350 9.570 23.520 ;
        RECT 9.810 23.485 9.960 23.655 ;
        RECT 10.200 23.485 10.350 23.655 ;
        RECT 10.590 23.350 10.740 23.520 ;
        RECT 12.320 23.350 12.470 23.520 ;
        RECT 12.710 23.485 12.860 23.655 ;
        RECT 13.100 23.485 13.250 23.655 ;
        RECT 13.490 23.350 13.640 23.520 ;
        RECT 15.220 23.350 15.370 23.520 ;
        RECT 15.610 23.485 15.760 23.655 ;
        RECT 16.000 23.485 16.150 23.655 ;
        RECT 16.390 23.350 16.540 23.520 ;
        RECT 18.120 23.350 18.270 23.520 ;
        RECT 18.510 23.485 18.660 23.655 ;
        RECT 18.900 23.485 19.050 23.655 ;
        RECT 19.290 23.350 19.440 23.520 ;
        RECT 21.020 23.350 21.170 23.520 ;
        RECT 21.410 23.485 21.560 23.655 ;
        RECT 21.800 23.485 21.950 23.655 ;
        RECT 22.190 23.350 22.340 23.520 ;
        RECT 23.920 23.350 24.070 23.520 ;
        RECT 24.310 23.485 24.460 23.655 ;
        RECT 24.700 23.485 24.850 23.655 ;
        RECT 25.090 23.350 25.240 23.520 ;
        RECT 26.820 23.350 26.970 23.520 ;
        RECT 27.210 23.485 27.360 23.655 ;
        RECT 27.600 23.485 27.750 23.655 ;
        RECT 27.990 23.350 28.140 23.520 ;
        RECT 29.720 23.350 29.870 23.520 ;
        RECT 30.110 23.485 30.260 23.655 ;
        RECT 30.500 23.485 30.650 23.655 ;
        RECT 30.890 23.350 31.040 23.520 ;
        RECT 32.620 23.350 32.770 23.520 ;
        RECT 33.010 23.485 33.160 23.655 ;
        RECT 33.400 23.485 33.550 23.655 ;
        RECT 33.790 23.350 33.940 23.520 ;
        RECT 35.520 23.350 35.670 23.520 ;
        RECT 35.910 23.485 36.060 23.655 ;
        RECT 36.300 23.485 36.450 23.655 ;
        RECT 36.690 23.350 36.840 23.520 ;
        RECT 38.420 23.350 38.570 23.520 ;
        RECT 38.810 23.485 38.960 23.655 ;
        RECT 39.200 23.485 39.350 23.655 ;
        RECT 39.590 23.350 39.740 23.520 ;
        RECT 41.320 23.350 41.470 23.520 ;
        RECT 41.710 23.485 41.860 23.655 ;
        RECT 42.100 23.485 42.250 23.655 ;
        RECT 42.490 23.350 42.640 23.520 ;
        RECT 44.220 23.350 44.370 23.520 ;
        RECT 44.610 23.485 44.760 23.655 ;
        RECT 45.000 23.485 45.150 23.655 ;
        RECT 45.390 23.350 45.540 23.520 ;
        RECT 47.120 23.350 47.270 23.520 ;
        RECT 47.510 23.485 47.660 23.655 ;
        RECT 47.900 23.485 48.050 23.655 ;
        RECT 48.290 23.350 48.440 23.520 ;
        RECT 50.020 23.350 50.170 23.520 ;
        RECT 50.410 23.485 50.560 23.655 ;
        RECT 50.800 23.485 50.950 23.655 ;
        RECT 51.190 23.350 51.340 23.520 ;
        RECT 52.920 23.350 53.070 23.520 ;
        RECT 53.310 23.485 53.460 23.655 ;
        RECT 53.700 23.485 53.850 23.655 ;
        RECT 54.090 23.350 54.240 23.520 ;
        RECT 55.820 23.350 55.970 23.520 ;
        RECT 56.210 23.485 56.360 23.655 ;
        RECT 56.600 23.485 56.750 23.655 ;
        RECT 56.990 23.350 57.140 23.520 ;
        RECT 58.720 23.350 58.870 23.520 ;
        RECT 59.110 23.485 59.260 23.655 ;
        RECT 59.500 23.485 59.650 23.655 ;
        RECT 59.890 23.350 60.040 23.520 ;
        RECT 61.620 23.350 61.770 23.520 ;
        RECT 62.010 23.485 62.160 23.655 ;
        RECT 62.400 23.485 62.550 23.655 ;
        RECT 62.790 23.350 62.940 23.520 ;
        RECT 64.520 23.350 64.670 23.520 ;
        RECT 64.910 23.485 65.060 23.655 ;
        RECT 65.300 23.485 65.450 23.655 ;
        RECT 65.690 23.350 65.840 23.520 ;
        RECT 67.420 23.350 67.570 23.520 ;
        RECT 67.810 23.485 67.960 23.655 ;
        RECT 68.200 23.485 68.350 23.655 ;
        RECT 68.590 23.350 68.740 23.520 ;
        RECT 70.320 23.350 70.470 23.520 ;
        RECT 70.710 23.485 70.860 23.655 ;
        RECT 71.100 23.485 71.250 23.655 ;
        RECT 71.490 23.350 71.640 23.520 ;
        RECT 73.220 23.350 73.370 23.520 ;
        RECT 73.610 23.485 73.760 23.655 ;
        RECT 74.000 23.485 74.150 23.655 ;
        RECT 74.390 23.350 74.540 23.520 ;
        RECT 76.120 23.350 76.270 23.520 ;
        RECT 76.510 23.485 76.660 23.655 ;
        RECT 76.900 23.485 77.050 23.655 ;
        RECT 77.290 23.350 77.440 23.520 ;
        RECT 79.020 23.350 79.170 23.520 ;
        RECT 79.410 23.485 79.560 23.655 ;
        RECT 79.800 23.485 79.950 23.655 ;
        RECT 80.190 23.350 80.340 23.520 ;
        RECT 81.920 23.350 82.070 23.520 ;
        RECT 82.310 23.485 82.460 23.655 ;
        RECT 82.700 23.485 82.850 23.655 ;
        RECT 83.090 23.350 83.240 23.520 ;
        RECT 84.820 23.350 84.970 23.520 ;
        RECT 85.210 23.485 85.360 23.655 ;
        RECT 85.600 23.485 85.750 23.655 ;
        RECT 85.990 23.350 86.140 23.520 ;
        RECT 87.720 23.350 87.870 23.520 ;
        RECT 88.110 23.485 88.260 23.655 ;
        RECT 88.500 23.485 88.650 23.655 ;
        RECT 88.890 23.350 89.040 23.520 ;
        RECT 90.620 23.350 90.770 23.520 ;
        RECT 91.010 23.485 91.160 23.655 ;
        RECT 91.400 23.485 91.550 23.655 ;
        RECT 91.790 23.350 91.940 23.520 ;
        RECT 0.985 23.265 1.035 23.300 ;
        POLYGON 1.035 23.300 1.070 23.265 1.035 23.265 ;
        RECT 0.985 23.140 1.070 23.265 ;
        RECT 1.690 23.140 1.775 23.300 ;
        RECT 3.885 23.265 3.935 23.300 ;
        POLYGON 3.935 23.300 3.970 23.265 3.935 23.265 ;
        RECT 3.885 23.140 3.970 23.265 ;
        RECT 4.590 23.140 4.675 23.300 ;
        RECT 6.785 23.265 6.835 23.300 ;
        POLYGON 6.835 23.300 6.870 23.265 6.835 23.265 ;
        RECT 6.785 23.140 6.870 23.265 ;
        RECT 7.490 23.140 7.575 23.300 ;
        RECT 9.685 23.265 9.735 23.300 ;
        POLYGON 9.735 23.300 9.770 23.265 9.735 23.265 ;
        RECT 9.685 23.140 9.770 23.265 ;
        RECT 10.390 23.140 10.475 23.300 ;
        RECT 12.585 23.265 12.635 23.300 ;
        POLYGON 12.635 23.300 12.670 23.265 12.635 23.265 ;
        RECT 12.585 23.140 12.670 23.265 ;
        RECT 13.290 23.140 13.375 23.300 ;
        RECT 15.485 23.265 15.535 23.300 ;
        POLYGON 15.535 23.300 15.570 23.265 15.535 23.265 ;
        RECT 15.485 23.140 15.570 23.265 ;
        RECT 16.190 23.140 16.275 23.300 ;
        RECT 18.385 23.265 18.435 23.300 ;
        POLYGON 18.435 23.300 18.470 23.265 18.435 23.265 ;
        RECT 18.385 23.140 18.470 23.265 ;
        RECT 19.090 23.140 19.175 23.300 ;
        RECT 21.285 23.265 21.335 23.300 ;
        POLYGON 21.335 23.300 21.370 23.265 21.335 23.265 ;
        RECT 21.285 23.140 21.370 23.265 ;
        RECT 21.990 23.140 22.075 23.300 ;
        RECT 24.185 23.265 24.235 23.300 ;
        POLYGON 24.235 23.300 24.270 23.265 24.235 23.265 ;
        RECT 24.185 23.140 24.270 23.265 ;
        RECT 24.890 23.140 24.975 23.300 ;
        RECT 27.085 23.265 27.135 23.300 ;
        POLYGON 27.135 23.300 27.170 23.265 27.135 23.265 ;
        RECT 27.085 23.140 27.170 23.265 ;
        RECT 27.790 23.140 27.875 23.300 ;
        RECT 29.985 23.265 30.035 23.300 ;
        POLYGON 30.035 23.300 30.070 23.265 30.035 23.265 ;
        RECT 29.985 23.140 30.070 23.265 ;
        RECT 30.690 23.140 30.775 23.300 ;
        RECT 32.885 23.265 32.935 23.300 ;
        POLYGON 32.935 23.300 32.970 23.265 32.935 23.265 ;
        RECT 32.885 23.140 32.970 23.265 ;
        RECT 33.590 23.140 33.675 23.300 ;
        RECT 35.785 23.265 35.835 23.300 ;
        POLYGON 35.835 23.300 35.870 23.265 35.835 23.265 ;
        RECT 35.785 23.140 35.870 23.265 ;
        RECT 36.490 23.140 36.575 23.300 ;
        RECT 38.685 23.265 38.735 23.300 ;
        POLYGON 38.735 23.300 38.770 23.265 38.735 23.265 ;
        RECT 38.685 23.140 38.770 23.265 ;
        RECT 39.390 23.140 39.475 23.300 ;
        RECT 41.585 23.265 41.635 23.300 ;
        POLYGON 41.635 23.300 41.670 23.265 41.635 23.265 ;
        RECT 41.585 23.140 41.670 23.265 ;
        RECT 42.290 23.140 42.375 23.300 ;
        RECT 44.485 23.265 44.535 23.300 ;
        POLYGON 44.535 23.300 44.570 23.265 44.535 23.265 ;
        RECT 44.485 23.140 44.570 23.265 ;
        RECT 45.190 23.140 45.275 23.300 ;
        RECT 47.385 23.265 47.435 23.300 ;
        POLYGON 47.435 23.300 47.470 23.265 47.435 23.265 ;
        RECT 47.385 23.140 47.470 23.265 ;
        RECT 48.090 23.140 48.175 23.300 ;
        RECT 50.285 23.265 50.335 23.300 ;
        POLYGON 50.335 23.300 50.370 23.265 50.335 23.265 ;
        RECT 50.285 23.140 50.370 23.265 ;
        RECT 50.990 23.140 51.075 23.300 ;
        RECT 53.185 23.265 53.235 23.300 ;
        POLYGON 53.235 23.300 53.270 23.265 53.235 23.265 ;
        RECT 53.185 23.140 53.270 23.265 ;
        RECT 53.890 23.140 53.975 23.300 ;
        RECT 56.085 23.265 56.135 23.300 ;
        POLYGON 56.135 23.300 56.170 23.265 56.135 23.265 ;
        RECT 56.085 23.140 56.170 23.265 ;
        RECT 56.790 23.140 56.875 23.300 ;
        RECT 58.985 23.265 59.035 23.300 ;
        POLYGON 59.035 23.300 59.070 23.265 59.035 23.265 ;
        RECT 58.985 23.140 59.070 23.265 ;
        RECT 59.690 23.140 59.775 23.300 ;
        RECT 61.885 23.265 61.935 23.300 ;
        POLYGON 61.935 23.300 61.970 23.265 61.935 23.265 ;
        RECT 61.885 23.140 61.970 23.265 ;
        RECT 62.590 23.140 62.675 23.300 ;
        RECT 64.785 23.265 64.835 23.300 ;
        POLYGON 64.835 23.300 64.870 23.265 64.835 23.265 ;
        RECT 64.785 23.140 64.870 23.265 ;
        RECT 65.490 23.140 65.575 23.300 ;
        RECT 67.685 23.265 67.735 23.300 ;
        POLYGON 67.735 23.300 67.770 23.265 67.735 23.265 ;
        RECT 67.685 23.140 67.770 23.265 ;
        RECT 68.390 23.140 68.475 23.300 ;
        RECT 70.585 23.265 70.635 23.300 ;
        POLYGON 70.635 23.300 70.670 23.265 70.635 23.265 ;
        RECT 70.585 23.140 70.670 23.265 ;
        RECT 71.290 23.140 71.375 23.300 ;
        RECT 73.485 23.265 73.535 23.300 ;
        POLYGON 73.535 23.300 73.570 23.265 73.535 23.265 ;
        RECT 73.485 23.140 73.570 23.265 ;
        RECT 74.190 23.140 74.275 23.300 ;
        RECT 76.385 23.265 76.435 23.300 ;
        POLYGON 76.435 23.300 76.470 23.265 76.435 23.265 ;
        RECT 76.385 23.140 76.470 23.265 ;
        RECT 77.090 23.140 77.175 23.300 ;
        RECT 79.285 23.265 79.335 23.300 ;
        POLYGON 79.335 23.300 79.370 23.265 79.335 23.265 ;
        RECT 79.285 23.140 79.370 23.265 ;
        RECT 79.990 23.140 80.075 23.300 ;
        RECT 82.185 23.265 82.235 23.300 ;
        POLYGON 82.235 23.300 82.270 23.265 82.235 23.265 ;
        RECT 82.185 23.140 82.270 23.265 ;
        RECT 82.890 23.140 82.975 23.300 ;
        RECT 85.085 23.265 85.135 23.300 ;
        POLYGON 85.135 23.300 85.170 23.265 85.135 23.265 ;
        RECT 85.085 23.140 85.170 23.265 ;
        RECT 85.790 23.140 85.875 23.300 ;
        RECT 87.985 23.265 88.035 23.300 ;
        POLYGON 88.035 23.300 88.070 23.265 88.035 23.265 ;
        RECT 87.985 23.140 88.070 23.265 ;
        RECT 88.690 23.140 88.775 23.300 ;
        RECT 90.885 23.265 90.935 23.300 ;
        POLYGON 90.935 23.300 90.970 23.265 90.935 23.265 ;
        RECT 90.885 23.140 90.970 23.265 ;
        RECT 91.590 23.140 91.675 23.300 ;
        RECT 0.775 22.520 0.850 22.660 ;
        RECT 0.990 22.470 1.065 22.610 ;
        RECT 1.695 22.530 1.755 22.610 ;
        POLYGON 1.695 22.530 1.755 22.530 1.755 22.470 ;
        RECT 1.910 22.520 1.985 22.660 ;
        RECT 3.675 22.520 3.750 22.660 ;
        RECT 3.890 22.470 3.965 22.610 ;
        RECT 4.595 22.530 4.655 22.610 ;
        POLYGON 4.595 22.530 4.655 22.530 4.655 22.470 ;
        RECT 4.810 22.520 4.885 22.660 ;
        RECT 6.575 22.520 6.650 22.660 ;
        RECT 6.790 22.470 6.865 22.610 ;
        RECT 7.495 22.530 7.555 22.610 ;
        POLYGON 7.495 22.530 7.555 22.530 7.555 22.470 ;
        RECT 7.710 22.520 7.785 22.660 ;
        RECT 9.475 22.520 9.550 22.660 ;
        RECT 9.690 22.470 9.765 22.610 ;
        RECT 10.395 22.530 10.455 22.610 ;
        POLYGON 10.395 22.530 10.455 22.530 10.455 22.470 ;
        RECT 10.610 22.520 10.685 22.660 ;
        RECT 12.375 22.520 12.450 22.660 ;
        RECT 12.590 22.470 12.665 22.610 ;
        RECT 13.295 22.530 13.355 22.610 ;
        POLYGON 13.295 22.530 13.355 22.530 13.355 22.470 ;
        RECT 13.510 22.520 13.585 22.660 ;
        RECT 15.275 22.520 15.350 22.660 ;
        RECT 15.490 22.470 15.565 22.610 ;
        RECT 16.195 22.530 16.255 22.610 ;
        POLYGON 16.195 22.530 16.255 22.530 16.255 22.470 ;
        RECT 16.410 22.520 16.485 22.660 ;
        RECT 18.175 22.520 18.250 22.660 ;
        RECT 18.390 22.470 18.465 22.610 ;
        RECT 19.095 22.530 19.155 22.610 ;
        POLYGON 19.095 22.530 19.155 22.530 19.155 22.470 ;
        RECT 19.310 22.520 19.385 22.660 ;
        RECT 21.075 22.520 21.150 22.660 ;
        RECT 21.290 22.470 21.365 22.610 ;
        RECT 21.995 22.530 22.055 22.610 ;
        POLYGON 21.995 22.530 22.055 22.530 22.055 22.470 ;
        RECT 22.210 22.520 22.285 22.660 ;
        RECT 23.975 22.520 24.050 22.660 ;
        RECT 24.190 22.470 24.265 22.610 ;
        RECT 24.895 22.530 24.955 22.610 ;
        POLYGON 24.895 22.530 24.955 22.530 24.955 22.470 ;
        RECT 25.110 22.520 25.185 22.660 ;
        RECT 26.875 22.520 26.950 22.660 ;
        RECT 27.090 22.470 27.165 22.610 ;
        RECT 27.795 22.530 27.855 22.610 ;
        POLYGON 27.795 22.530 27.855 22.530 27.855 22.470 ;
        RECT 28.010 22.520 28.085 22.660 ;
        RECT 29.775 22.520 29.850 22.660 ;
        RECT 29.990 22.470 30.065 22.610 ;
        RECT 30.695 22.530 30.755 22.610 ;
        POLYGON 30.695 22.530 30.755 22.530 30.755 22.470 ;
        RECT 30.910 22.520 30.985 22.660 ;
        RECT 32.675 22.520 32.750 22.660 ;
        RECT 32.890 22.470 32.965 22.610 ;
        RECT 33.595 22.530 33.655 22.610 ;
        POLYGON 33.595 22.530 33.655 22.530 33.655 22.470 ;
        RECT 33.810 22.520 33.885 22.660 ;
        RECT 35.575 22.520 35.650 22.660 ;
        RECT 35.790 22.470 35.865 22.610 ;
        RECT 36.495 22.530 36.555 22.610 ;
        POLYGON 36.495 22.530 36.555 22.530 36.555 22.470 ;
        RECT 36.710 22.520 36.785 22.660 ;
        RECT 38.475 22.520 38.550 22.660 ;
        RECT 38.690 22.470 38.765 22.610 ;
        RECT 39.395 22.530 39.455 22.610 ;
        POLYGON 39.395 22.530 39.455 22.530 39.455 22.470 ;
        RECT 39.610 22.520 39.685 22.660 ;
        RECT 41.375 22.520 41.450 22.660 ;
        RECT 41.590 22.470 41.665 22.610 ;
        RECT 42.295 22.530 42.355 22.610 ;
        POLYGON 42.295 22.530 42.355 22.530 42.355 22.470 ;
        RECT 42.510 22.520 42.585 22.660 ;
        RECT 44.275 22.520 44.350 22.660 ;
        RECT 44.490 22.470 44.565 22.610 ;
        RECT 45.195 22.530 45.255 22.610 ;
        POLYGON 45.195 22.530 45.255 22.530 45.255 22.470 ;
        RECT 45.410 22.520 45.485 22.660 ;
        RECT 47.175 22.520 47.250 22.660 ;
        RECT 47.390 22.470 47.465 22.610 ;
        RECT 48.095 22.530 48.155 22.610 ;
        POLYGON 48.095 22.530 48.155 22.530 48.155 22.470 ;
        RECT 48.310 22.520 48.385 22.660 ;
        RECT 50.075 22.520 50.150 22.660 ;
        RECT 50.290 22.470 50.365 22.610 ;
        RECT 50.995 22.530 51.055 22.610 ;
        POLYGON 50.995 22.530 51.055 22.530 51.055 22.470 ;
        RECT 51.210 22.520 51.285 22.660 ;
        RECT 52.975 22.520 53.050 22.660 ;
        RECT 53.190 22.470 53.265 22.610 ;
        RECT 53.895 22.530 53.955 22.610 ;
        POLYGON 53.895 22.530 53.955 22.530 53.955 22.470 ;
        RECT 54.110 22.520 54.185 22.660 ;
        RECT 55.875 22.520 55.950 22.660 ;
        RECT 56.090 22.470 56.165 22.610 ;
        RECT 56.795 22.530 56.855 22.610 ;
        POLYGON 56.795 22.530 56.855 22.530 56.855 22.470 ;
        RECT 57.010 22.520 57.085 22.660 ;
        RECT 58.775 22.520 58.850 22.660 ;
        RECT 58.990 22.470 59.065 22.610 ;
        RECT 59.695 22.530 59.755 22.610 ;
        POLYGON 59.695 22.530 59.755 22.530 59.755 22.470 ;
        RECT 59.910 22.520 59.985 22.660 ;
        RECT 61.675 22.520 61.750 22.660 ;
        RECT 61.890 22.470 61.965 22.610 ;
        RECT 62.595 22.530 62.655 22.610 ;
        POLYGON 62.595 22.530 62.655 22.530 62.655 22.470 ;
        RECT 62.810 22.520 62.885 22.660 ;
        RECT 64.575 22.520 64.650 22.660 ;
        RECT 64.790 22.470 64.865 22.610 ;
        RECT 65.495 22.530 65.555 22.610 ;
        POLYGON 65.495 22.530 65.555 22.530 65.555 22.470 ;
        RECT 65.710 22.520 65.785 22.660 ;
        RECT 67.475 22.520 67.550 22.660 ;
        RECT 67.690 22.470 67.765 22.610 ;
        RECT 68.395 22.530 68.455 22.610 ;
        POLYGON 68.395 22.530 68.455 22.530 68.455 22.470 ;
        RECT 68.610 22.520 68.685 22.660 ;
        RECT 70.375 22.520 70.450 22.660 ;
        RECT 70.590 22.470 70.665 22.610 ;
        RECT 71.295 22.530 71.355 22.610 ;
        POLYGON 71.295 22.530 71.355 22.530 71.355 22.470 ;
        RECT 71.510 22.520 71.585 22.660 ;
        RECT 73.275 22.520 73.350 22.660 ;
        RECT 73.490 22.470 73.565 22.610 ;
        RECT 74.195 22.530 74.255 22.610 ;
        POLYGON 74.195 22.530 74.255 22.530 74.255 22.470 ;
        RECT 74.410 22.520 74.485 22.660 ;
        RECT 76.175 22.520 76.250 22.660 ;
        RECT 76.390 22.470 76.465 22.610 ;
        RECT 77.095 22.530 77.155 22.610 ;
        POLYGON 77.095 22.530 77.155 22.530 77.155 22.470 ;
        RECT 77.310 22.520 77.385 22.660 ;
        RECT 79.075 22.520 79.150 22.660 ;
        RECT 79.290 22.470 79.365 22.610 ;
        RECT 79.995 22.530 80.055 22.610 ;
        POLYGON 79.995 22.530 80.055 22.530 80.055 22.470 ;
        RECT 80.210 22.520 80.285 22.660 ;
        RECT 81.975 22.520 82.050 22.660 ;
        RECT 82.190 22.470 82.265 22.610 ;
        RECT 82.895 22.530 82.955 22.610 ;
        POLYGON 82.895 22.530 82.955 22.530 82.955 22.470 ;
        RECT 83.110 22.520 83.185 22.660 ;
        RECT 84.875 22.520 84.950 22.660 ;
        RECT 85.090 22.470 85.165 22.610 ;
        RECT 85.795 22.530 85.855 22.610 ;
        POLYGON 85.795 22.530 85.855 22.530 85.855 22.470 ;
        RECT 86.010 22.520 86.085 22.660 ;
        RECT 87.775 22.520 87.850 22.660 ;
        RECT 87.990 22.470 88.065 22.610 ;
        RECT 88.695 22.530 88.755 22.610 ;
        POLYGON 88.695 22.530 88.755 22.530 88.755 22.470 ;
        RECT 88.910 22.520 88.985 22.660 ;
        RECT 90.675 22.520 90.750 22.660 ;
        RECT 90.890 22.470 90.965 22.610 ;
        RECT 91.595 22.530 91.655 22.610 ;
        POLYGON 91.595 22.530 91.655 22.530 91.655 22.470 ;
        RECT 91.810 22.520 91.885 22.660 ;
        RECT 0.720 22.000 0.870 22.170 ;
        RECT 1.110 22.135 1.260 22.305 ;
        RECT 1.500 22.135 1.650 22.305 ;
        RECT 1.890 22.000 2.040 22.170 ;
        RECT 3.620 22.000 3.770 22.170 ;
        RECT 4.010 22.135 4.160 22.305 ;
        RECT 4.400 22.135 4.550 22.305 ;
        RECT 4.790 22.000 4.940 22.170 ;
        RECT 6.520 22.000 6.670 22.170 ;
        RECT 6.910 22.135 7.060 22.305 ;
        RECT 7.300 22.135 7.450 22.305 ;
        RECT 7.690 22.000 7.840 22.170 ;
        RECT 9.420 22.000 9.570 22.170 ;
        RECT 9.810 22.135 9.960 22.305 ;
        RECT 10.200 22.135 10.350 22.305 ;
        RECT 10.590 22.000 10.740 22.170 ;
        RECT 12.320 22.000 12.470 22.170 ;
        RECT 12.710 22.135 12.860 22.305 ;
        RECT 13.100 22.135 13.250 22.305 ;
        RECT 13.490 22.000 13.640 22.170 ;
        RECT 15.220 22.000 15.370 22.170 ;
        RECT 15.610 22.135 15.760 22.305 ;
        RECT 16.000 22.135 16.150 22.305 ;
        RECT 16.390 22.000 16.540 22.170 ;
        RECT 18.120 22.000 18.270 22.170 ;
        RECT 18.510 22.135 18.660 22.305 ;
        RECT 18.900 22.135 19.050 22.305 ;
        RECT 19.290 22.000 19.440 22.170 ;
        RECT 21.020 22.000 21.170 22.170 ;
        RECT 21.410 22.135 21.560 22.305 ;
        RECT 21.800 22.135 21.950 22.305 ;
        RECT 22.190 22.000 22.340 22.170 ;
        RECT 23.920 22.000 24.070 22.170 ;
        RECT 24.310 22.135 24.460 22.305 ;
        RECT 24.700 22.135 24.850 22.305 ;
        RECT 25.090 22.000 25.240 22.170 ;
        RECT 26.820 22.000 26.970 22.170 ;
        RECT 27.210 22.135 27.360 22.305 ;
        RECT 27.600 22.135 27.750 22.305 ;
        RECT 27.990 22.000 28.140 22.170 ;
        RECT 29.720 22.000 29.870 22.170 ;
        RECT 30.110 22.135 30.260 22.305 ;
        RECT 30.500 22.135 30.650 22.305 ;
        RECT 30.890 22.000 31.040 22.170 ;
        RECT 32.620 22.000 32.770 22.170 ;
        RECT 33.010 22.135 33.160 22.305 ;
        RECT 33.400 22.135 33.550 22.305 ;
        RECT 33.790 22.000 33.940 22.170 ;
        RECT 35.520 22.000 35.670 22.170 ;
        RECT 35.910 22.135 36.060 22.305 ;
        RECT 36.300 22.135 36.450 22.305 ;
        RECT 36.690 22.000 36.840 22.170 ;
        RECT 38.420 22.000 38.570 22.170 ;
        RECT 38.810 22.135 38.960 22.305 ;
        RECT 39.200 22.135 39.350 22.305 ;
        RECT 39.590 22.000 39.740 22.170 ;
        RECT 41.320 22.000 41.470 22.170 ;
        RECT 41.710 22.135 41.860 22.305 ;
        RECT 42.100 22.135 42.250 22.305 ;
        RECT 42.490 22.000 42.640 22.170 ;
        RECT 44.220 22.000 44.370 22.170 ;
        RECT 44.610 22.135 44.760 22.305 ;
        RECT 45.000 22.135 45.150 22.305 ;
        RECT 45.390 22.000 45.540 22.170 ;
        RECT 47.120 22.000 47.270 22.170 ;
        RECT 47.510 22.135 47.660 22.305 ;
        RECT 47.900 22.135 48.050 22.305 ;
        RECT 48.290 22.000 48.440 22.170 ;
        RECT 50.020 22.000 50.170 22.170 ;
        RECT 50.410 22.135 50.560 22.305 ;
        RECT 50.800 22.135 50.950 22.305 ;
        RECT 51.190 22.000 51.340 22.170 ;
        RECT 52.920 22.000 53.070 22.170 ;
        RECT 53.310 22.135 53.460 22.305 ;
        RECT 53.700 22.135 53.850 22.305 ;
        RECT 54.090 22.000 54.240 22.170 ;
        RECT 55.820 22.000 55.970 22.170 ;
        RECT 56.210 22.135 56.360 22.305 ;
        RECT 56.600 22.135 56.750 22.305 ;
        RECT 56.990 22.000 57.140 22.170 ;
        RECT 58.720 22.000 58.870 22.170 ;
        RECT 59.110 22.135 59.260 22.305 ;
        RECT 59.500 22.135 59.650 22.305 ;
        RECT 59.890 22.000 60.040 22.170 ;
        RECT 61.620 22.000 61.770 22.170 ;
        RECT 62.010 22.135 62.160 22.305 ;
        RECT 62.400 22.135 62.550 22.305 ;
        RECT 62.790 22.000 62.940 22.170 ;
        RECT 64.520 22.000 64.670 22.170 ;
        RECT 64.910 22.135 65.060 22.305 ;
        RECT 65.300 22.135 65.450 22.305 ;
        RECT 65.690 22.000 65.840 22.170 ;
        RECT 67.420 22.000 67.570 22.170 ;
        RECT 67.810 22.135 67.960 22.305 ;
        RECT 68.200 22.135 68.350 22.305 ;
        RECT 68.590 22.000 68.740 22.170 ;
        RECT 70.320 22.000 70.470 22.170 ;
        RECT 70.710 22.135 70.860 22.305 ;
        RECT 71.100 22.135 71.250 22.305 ;
        RECT 71.490 22.000 71.640 22.170 ;
        RECT 73.220 22.000 73.370 22.170 ;
        RECT 73.610 22.135 73.760 22.305 ;
        RECT 74.000 22.135 74.150 22.305 ;
        RECT 74.390 22.000 74.540 22.170 ;
        RECT 76.120 22.000 76.270 22.170 ;
        RECT 76.510 22.135 76.660 22.305 ;
        RECT 76.900 22.135 77.050 22.305 ;
        RECT 77.290 22.000 77.440 22.170 ;
        RECT 79.020 22.000 79.170 22.170 ;
        RECT 79.410 22.135 79.560 22.305 ;
        RECT 79.800 22.135 79.950 22.305 ;
        RECT 80.190 22.000 80.340 22.170 ;
        RECT 81.920 22.000 82.070 22.170 ;
        RECT 82.310 22.135 82.460 22.305 ;
        RECT 82.700 22.135 82.850 22.305 ;
        RECT 83.090 22.000 83.240 22.170 ;
        RECT 84.820 22.000 84.970 22.170 ;
        RECT 85.210 22.135 85.360 22.305 ;
        RECT 85.600 22.135 85.750 22.305 ;
        RECT 85.990 22.000 86.140 22.170 ;
        RECT 87.720 22.000 87.870 22.170 ;
        RECT 88.110 22.135 88.260 22.305 ;
        RECT 88.500 22.135 88.650 22.305 ;
        RECT 88.890 22.000 89.040 22.170 ;
        RECT 90.620 22.000 90.770 22.170 ;
        RECT 91.010 22.135 91.160 22.305 ;
        RECT 91.400 22.135 91.550 22.305 ;
        RECT 91.790 22.000 91.940 22.170 ;
        RECT 0.985 21.915 1.035 21.950 ;
        POLYGON 1.035 21.950 1.070 21.915 1.035 21.915 ;
        RECT 0.985 21.790 1.070 21.915 ;
        RECT 1.690 21.790 1.775 21.950 ;
        RECT 3.885 21.915 3.935 21.950 ;
        POLYGON 3.935 21.950 3.970 21.915 3.935 21.915 ;
        RECT 3.885 21.790 3.970 21.915 ;
        RECT 4.590 21.790 4.675 21.950 ;
        RECT 6.785 21.915 6.835 21.950 ;
        POLYGON 6.835 21.950 6.870 21.915 6.835 21.915 ;
        RECT 6.785 21.790 6.870 21.915 ;
        RECT 7.490 21.790 7.575 21.950 ;
        RECT 9.685 21.915 9.735 21.950 ;
        POLYGON 9.735 21.950 9.770 21.915 9.735 21.915 ;
        RECT 9.685 21.790 9.770 21.915 ;
        RECT 10.390 21.790 10.475 21.950 ;
        RECT 12.585 21.915 12.635 21.950 ;
        POLYGON 12.635 21.950 12.670 21.915 12.635 21.915 ;
        RECT 12.585 21.790 12.670 21.915 ;
        RECT 13.290 21.790 13.375 21.950 ;
        RECT 15.485 21.915 15.535 21.950 ;
        POLYGON 15.535 21.950 15.570 21.915 15.535 21.915 ;
        RECT 15.485 21.790 15.570 21.915 ;
        RECT 16.190 21.790 16.275 21.950 ;
        RECT 18.385 21.915 18.435 21.950 ;
        POLYGON 18.435 21.950 18.470 21.915 18.435 21.915 ;
        RECT 18.385 21.790 18.470 21.915 ;
        RECT 19.090 21.790 19.175 21.950 ;
        RECT 21.285 21.915 21.335 21.950 ;
        POLYGON 21.335 21.950 21.370 21.915 21.335 21.915 ;
        RECT 21.285 21.790 21.370 21.915 ;
        RECT 21.990 21.790 22.075 21.950 ;
        RECT 24.185 21.915 24.235 21.950 ;
        POLYGON 24.235 21.950 24.270 21.915 24.235 21.915 ;
        RECT 24.185 21.790 24.270 21.915 ;
        RECT 24.890 21.790 24.975 21.950 ;
        RECT 27.085 21.915 27.135 21.950 ;
        POLYGON 27.135 21.950 27.170 21.915 27.135 21.915 ;
        RECT 27.085 21.790 27.170 21.915 ;
        RECT 27.790 21.790 27.875 21.950 ;
        RECT 29.985 21.915 30.035 21.950 ;
        POLYGON 30.035 21.950 30.070 21.915 30.035 21.915 ;
        RECT 29.985 21.790 30.070 21.915 ;
        RECT 30.690 21.790 30.775 21.950 ;
        RECT 32.885 21.915 32.935 21.950 ;
        POLYGON 32.935 21.950 32.970 21.915 32.935 21.915 ;
        RECT 32.885 21.790 32.970 21.915 ;
        RECT 33.590 21.790 33.675 21.950 ;
        RECT 35.785 21.915 35.835 21.950 ;
        POLYGON 35.835 21.950 35.870 21.915 35.835 21.915 ;
        RECT 35.785 21.790 35.870 21.915 ;
        RECT 36.490 21.790 36.575 21.950 ;
        RECT 38.685 21.915 38.735 21.950 ;
        POLYGON 38.735 21.950 38.770 21.915 38.735 21.915 ;
        RECT 38.685 21.790 38.770 21.915 ;
        RECT 39.390 21.790 39.475 21.950 ;
        RECT 41.585 21.915 41.635 21.950 ;
        POLYGON 41.635 21.950 41.670 21.915 41.635 21.915 ;
        RECT 41.585 21.790 41.670 21.915 ;
        RECT 42.290 21.790 42.375 21.950 ;
        RECT 44.485 21.915 44.535 21.950 ;
        POLYGON 44.535 21.950 44.570 21.915 44.535 21.915 ;
        RECT 44.485 21.790 44.570 21.915 ;
        RECT 45.190 21.790 45.275 21.950 ;
        RECT 47.385 21.915 47.435 21.950 ;
        POLYGON 47.435 21.950 47.470 21.915 47.435 21.915 ;
        RECT 47.385 21.790 47.470 21.915 ;
        RECT 48.090 21.790 48.175 21.950 ;
        RECT 50.285 21.915 50.335 21.950 ;
        POLYGON 50.335 21.950 50.370 21.915 50.335 21.915 ;
        RECT 50.285 21.790 50.370 21.915 ;
        RECT 50.990 21.790 51.075 21.950 ;
        RECT 53.185 21.915 53.235 21.950 ;
        POLYGON 53.235 21.950 53.270 21.915 53.235 21.915 ;
        RECT 53.185 21.790 53.270 21.915 ;
        RECT 53.890 21.790 53.975 21.950 ;
        RECT 56.085 21.915 56.135 21.950 ;
        POLYGON 56.135 21.950 56.170 21.915 56.135 21.915 ;
        RECT 56.085 21.790 56.170 21.915 ;
        RECT 56.790 21.790 56.875 21.950 ;
        RECT 58.985 21.915 59.035 21.950 ;
        POLYGON 59.035 21.950 59.070 21.915 59.035 21.915 ;
        RECT 58.985 21.790 59.070 21.915 ;
        RECT 59.690 21.790 59.775 21.950 ;
        RECT 61.885 21.915 61.935 21.950 ;
        POLYGON 61.935 21.950 61.970 21.915 61.935 21.915 ;
        RECT 61.885 21.790 61.970 21.915 ;
        RECT 62.590 21.790 62.675 21.950 ;
        RECT 64.785 21.915 64.835 21.950 ;
        POLYGON 64.835 21.950 64.870 21.915 64.835 21.915 ;
        RECT 64.785 21.790 64.870 21.915 ;
        RECT 65.490 21.790 65.575 21.950 ;
        RECT 67.685 21.915 67.735 21.950 ;
        POLYGON 67.735 21.950 67.770 21.915 67.735 21.915 ;
        RECT 67.685 21.790 67.770 21.915 ;
        RECT 68.390 21.790 68.475 21.950 ;
        RECT 70.585 21.915 70.635 21.950 ;
        POLYGON 70.635 21.950 70.670 21.915 70.635 21.915 ;
        RECT 70.585 21.790 70.670 21.915 ;
        RECT 71.290 21.790 71.375 21.950 ;
        RECT 73.485 21.915 73.535 21.950 ;
        POLYGON 73.535 21.950 73.570 21.915 73.535 21.915 ;
        RECT 73.485 21.790 73.570 21.915 ;
        RECT 74.190 21.790 74.275 21.950 ;
        RECT 76.385 21.915 76.435 21.950 ;
        POLYGON 76.435 21.950 76.470 21.915 76.435 21.915 ;
        RECT 76.385 21.790 76.470 21.915 ;
        RECT 77.090 21.790 77.175 21.950 ;
        RECT 79.285 21.915 79.335 21.950 ;
        POLYGON 79.335 21.950 79.370 21.915 79.335 21.915 ;
        RECT 79.285 21.790 79.370 21.915 ;
        RECT 79.990 21.790 80.075 21.950 ;
        RECT 82.185 21.915 82.235 21.950 ;
        POLYGON 82.235 21.950 82.270 21.915 82.235 21.915 ;
        RECT 82.185 21.790 82.270 21.915 ;
        RECT 82.890 21.790 82.975 21.950 ;
        RECT 85.085 21.915 85.135 21.950 ;
        POLYGON 85.135 21.950 85.170 21.915 85.135 21.915 ;
        RECT 85.085 21.790 85.170 21.915 ;
        RECT 85.790 21.790 85.875 21.950 ;
        RECT 87.985 21.915 88.035 21.950 ;
        POLYGON 88.035 21.950 88.070 21.915 88.035 21.915 ;
        RECT 87.985 21.790 88.070 21.915 ;
        RECT 88.690 21.790 88.775 21.950 ;
        RECT 90.885 21.915 90.935 21.950 ;
        POLYGON 90.935 21.950 90.970 21.915 90.935 21.915 ;
        RECT 90.885 21.790 90.970 21.915 ;
        RECT 91.590 21.790 91.675 21.950 ;
        RECT 0.775 21.170 0.850 21.310 ;
        RECT 0.990 21.120 1.065 21.260 ;
        RECT 1.695 21.180 1.755 21.260 ;
        POLYGON 1.695 21.180 1.755 21.180 1.755 21.120 ;
        RECT 1.910 21.170 1.985 21.310 ;
        RECT 3.675 21.170 3.750 21.310 ;
        RECT 3.890 21.120 3.965 21.260 ;
        RECT 4.595 21.180 4.655 21.260 ;
        POLYGON 4.595 21.180 4.655 21.180 4.655 21.120 ;
        RECT 4.810 21.170 4.885 21.310 ;
        RECT 6.575 21.170 6.650 21.310 ;
        RECT 6.790 21.120 6.865 21.260 ;
        RECT 7.495 21.180 7.555 21.260 ;
        POLYGON 7.495 21.180 7.555 21.180 7.555 21.120 ;
        RECT 7.710 21.170 7.785 21.310 ;
        RECT 9.475 21.170 9.550 21.310 ;
        RECT 9.690 21.120 9.765 21.260 ;
        RECT 10.395 21.180 10.455 21.260 ;
        POLYGON 10.395 21.180 10.455 21.180 10.455 21.120 ;
        RECT 10.610 21.170 10.685 21.310 ;
        RECT 12.375 21.170 12.450 21.310 ;
        RECT 12.590 21.120 12.665 21.260 ;
        RECT 13.295 21.180 13.355 21.260 ;
        POLYGON 13.295 21.180 13.355 21.180 13.355 21.120 ;
        RECT 13.510 21.170 13.585 21.310 ;
        RECT 15.275 21.170 15.350 21.310 ;
        RECT 15.490 21.120 15.565 21.260 ;
        RECT 16.195 21.180 16.255 21.260 ;
        POLYGON 16.195 21.180 16.255 21.180 16.255 21.120 ;
        RECT 16.410 21.170 16.485 21.310 ;
        RECT 18.175 21.170 18.250 21.310 ;
        RECT 18.390 21.120 18.465 21.260 ;
        RECT 19.095 21.180 19.155 21.260 ;
        POLYGON 19.095 21.180 19.155 21.180 19.155 21.120 ;
        RECT 19.310 21.170 19.385 21.310 ;
        RECT 21.075 21.170 21.150 21.310 ;
        RECT 21.290 21.120 21.365 21.260 ;
        RECT 21.995 21.180 22.055 21.260 ;
        POLYGON 21.995 21.180 22.055 21.180 22.055 21.120 ;
        RECT 22.210 21.170 22.285 21.310 ;
        RECT 23.975 21.170 24.050 21.310 ;
        RECT 24.190 21.120 24.265 21.260 ;
        RECT 24.895 21.180 24.955 21.260 ;
        POLYGON 24.895 21.180 24.955 21.180 24.955 21.120 ;
        RECT 25.110 21.170 25.185 21.310 ;
        RECT 26.875 21.170 26.950 21.310 ;
        RECT 27.090 21.120 27.165 21.260 ;
        RECT 27.795 21.180 27.855 21.260 ;
        POLYGON 27.795 21.180 27.855 21.180 27.855 21.120 ;
        RECT 28.010 21.170 28.085 21.310 ;
        RECT 29.775 21.170 29.850 21.310 ;
        RECT 29.990 21.120 30.065 21.260 ;
        RECT 30.695 21.180 30.755 21.260 ;
        POLYGON 30.695 21.180 30.755 21.180 30.755 21.120 ;
        RECT 30.910 21.170 30.985 21.310 ;
        RECT 32.675 21.170 32.750 21.310 ;
        RECT 32.890 21.120 32.965 21.260 ;
        RECT 33.595 21.180 33.655 21.260 ;
        POLYGON 33.595 21.180 33.655 21.180 33.655 21.120 ;
        RECT 33.810 21.170 33.885 21.310 ;
        RECT 35.575 21.170 35.650 21.310 ;
        RECT 35.790 21.120 35.865 21.260 ;
        RECT 36.495 21.180 36.555 21.260 ;
        POLYGON 36.495 21.180 36.555 21.180 36.555 21.120 ;
        RECT 36.710 21.170 36.785 21.310 ;
        RECT 38.475 21.170 38.550 21.310 ;
        RECT 38.690 21.120 38.765 21.260 ;
        RECT 39.395 21.180 39.455 21.260 ;
        POLYGON 39.395 21.180 39.455 21.180 39.455 21.120 ;
        RECT 39.610 21.170 39.685 21.310 ;
        RECT 41.375 21.170 41.450 21.310 ;
        RECT 41.590 21.120 41.665 21.260 ;
        RECT 42.295 21.180 42.355 21.260 ;
        POLYGON 42.295 21.180 42.355 21.180 42.355 21.120 ;
        RECT 42.510 21.170 42.585 21.310 ;
        RECT 44.275 21.170 44.350 21.310 ;
        RECT 44.490 21.120 44.565 21.260 ;
        RECT 45.195 21.180 45.255 21.260 ;
        POLYGON 45.195 21.180 45.255 21.180 45.255 21.120 ;
        RECT 45.410 21.170 45.485 21.310 ;
        RECT 47.175 21.170 47.250 21.310 ;
        RECT 47.390 21.120 47.465 21.260 ;
        RECT 48.095 21.180 48.155 21.260 ;
        POLYGON 48.095 21.180 48.155 21.180 48.155 21.120 ;
        RECT 48.310 21.170 48.385 21.310 ;
        RECT 50.075 21.170 50.150 21.310 ;
        RECT 50.290 21.120 50.365 21.260 ;
        RECT 50.995 21.180 51.055 21.260 ;
        POLYGON 50.995 21.180 51.055 21.180 51.055 21.120 ;
        RECT 51.210 21.170 51.285 21.310 ;
        RECT 52.975 21.170 53.050 21.310 ;
        RECT 53.190 21.120 53.265 21.260 ;
        RECT 53.895 21.180 53.955 21.260 ;
        POLYGON 53.895 21.180 53.955 21.180 53.955 21.120 ;
        RECT 54.110 21.170 54.185 21.310 ;
        RECT 55.875 21.170 55.950 21.310 ;
        RECT 56.090 21.120 56.165 21.260 ;
        RECT 56.795 21.180 56.855 21.260 ;
        POLYGON 56.795 21.180 56.855 21.180 56.855 21.120 ;
        RECT 57.010 21.170 57.085 21.310 ;
        RECT 58.775 21.170 58.850 21.310 ;
        RECT 58.990 21.120 59.065 21.260 ;
        RECT 59.695 21.180 59.755 21.260 ;
        POLYGON 59.695 21.180 59.755 21.180 59.755 21.120 ;
        RECT 59.910 21.170 59.985 21.310 ;
        RECT 61.675 21.170 61.750 21.310 ;
        RECT 61.890 21.120 61.965 21.260 ;
        RECT 62.595 21.180 62.655 21.260 ;
        POLYGON 62.595 21.180 62.655 21.180 62.655 21.120 ;
        RECT 62.810 21.170 62.885 21.310 ;
        RECT 64.575 21.170 64.650 21.310 ;
        RECT 64.790 21.120 64.865 21.260 ;
        RECT 65.495 21.180 65.555 21.260 ;
        POLYGON 65.495 21.180 65.555 21.180 65.555 21.120 ;
        RECT 65.710 21.170 65.785 21.310 ;
        RECT 67.475 21.170 67.550 21.310 ;
        RECT 67.690 21.120 67.765 21.260 ;
        RECT 68.395 21.180 68.455 21.260 ;
        POLYGON 68.395 21.180 68.455 21.180 68.455 21.120 ;
        RECT 68.610 21.170 68.685 21.310 ;
        RECT 70.375 21.170 70.450 21.310 ;
        RECT 70.590 21.120 70.665 21.260 ;
        RECT 71.295 21.180 71.355 21.260 ;
        POLYGON 71.295 21.180 71.355 21.180 71.355 21.120 ;
        RECT 71.510 21.170 71.585 21.310 ;
        RECT 73.275 21.170 73.350 21.310 ;
        RECT 73.490 21.120 73.565 21.260 ;
        RECT 74.195 21.180 74.255 21.260 ;
        POLYGON 74.195 21.180 74.255 21.180 74.255 21.120 ;
        RECT 74.410 21.170 74.485 21.310 ;
        RECT 76.175 21.170 76.250 21.310 ;
        RECT 76.390 21.120 76.465 21.260 ;
        RECT 77.095 21.180 77.155 21.260 ;
        POLYGON 77.095 21.180 77.155 21.180 77.155 21.120 ;
        RECT 77.310 21.170 77.385 21.310 ;
        RECT 79.075 21.170 79.150 21.310 ;
        RECT 79.290 21.120 79.365 21.260 ;
        RECT 79.995 21.180 80.055 21.260 ;
        POLYGON 79.995 21.180 80.055 21.180 80.055 21.120 ;
        RECT 80.210 21.170 80.285 21.310 ;
        RECT 81.975 21.170 82.050 21.310 ;
        RECT 82.190 21.120 82.265 21.260 ;
        RECT 82.895 21.180 82.955 21.260 ;
        POLYGON 82.895 21.180 82.955 21.180 82.955 21.120 ;
        RECT 83.110 21.170 83.185 21.310 ;
        RECT 84.875 21.170 84.950 21.310 ;
        RECT 85.090 21.120 85.165 21.260 ;
        RECT 85.795 21.180 85.855 21.260 ;
        POLYGON 85.795 21.180 85.855 21.180 85.855 21.120 ;
        RECT 86.010 21.170 86.085 21.310 ;
        RECT 87.775 21.170 87.850 21.310 ;
        RECT 87.990 21.120 88.065 21.260 ;
        RECT 88.695 21.180 88.755 21.260 ;
        POLYGON 88.695 21.180 88.755 21.180 88.755 21.120 ;
        RECT 88.910 21.170 88.985 21.310 ;
        RECT 90.675 21.170 90.750 21.310 ;
        RECT 90.890 21.120 90.965 21.260 ;
        RECT 91.595 21.180 91.655 21.260 ;
        POLYGON 91.595 21.180 91.655 21.180 91.655 21.120 ;
        RECT 91.810 21.170 91.885 21.310 ;
        RECT 0.720 20.650 0.870 20.820 ;
        RECT 1.110 20.785 1.260 20.955 ;
        RECT 1.500 20.785 1.650 20.955 ;
        RECT 1.890 20.650 2.040 20.820 ;
        RECT 3.620 20.650 3.770 20.820 ;
        RECT 4.010 20.785 4.160 20.955 ;
        RECT 4.400 20.785 4.550 20.955 ;
        RECT 4.790 20.650 4.940 20.820 ;
        RECT 6.520 20.650 6.670 20.820 ;
        RECT 6.910 20.785 7.060 20.955 ;
        RECT 7.300 20.785 7.450 20.955 ;
        RECT 7.690 20.650 7.840 20.820 ;
        RECT 9.420 20.650 9.570 20.820 ;
        RECT 9.810 20.785 9.960 20.955 ;
        RECT 10.200 20.785 10.350 20.955 ;
        RECT 10.590 20.650 10.740 20.820 ;
        RECT 12.320 20.650 12.470 20.820 ;
        RECT 12.710 20.785 12.860 20.955 ;
        RECT 13.100 20.785 13.250 20.955 ;
        RECT 13.490 20.650 13.640 20.820 ;
        RECT 15.220 20.650 15.370 20.820 ;
        RECT 15.610 20.785 15.760 20.955 ;
        RECT 16.000 20.785 16.150 20.955 ;
        RECT 16.390 20.650 16.540 20.820 ;
        RECT 18.120 20.650 18.270 20.820 ;
        RECT 18.510 20.785 18.660 20.955 ;
        RECT 18.900 20.785 19.050 20.955 ;
        RECT 19.290 20.650 19.440 20.820 ;
        RECT 21.020 20.650 21.170 20.820 ;
        RECT 21.410 20.785 21.560 20.955 ;
        RECT 21.800 20.785 21.950 20.955 ;
        RECT 22.190 20.650 22.340 20.820 ;
        RECT 23.920 20.650 24.070 20.820 ;
        RECT 24.310 20.785 24.460 20.955 ;
        RECT 24.700 20.785 24.850 20.955 ;
        RECT 25.090 20.650 25.240 20.820 ;
        RECT 26.820 20.650 26.970 20.820 ;
        RECT 27.210 20.785 27.360 20.955 ;
        RECT 27.600 20.785 27.750 20.955 ;
        RECT 27.990 20.650 28.140 20.820 ;
        RECT 29.720 20.650 29.870 20.820 ;
        RECT 30.110 20.785 30.260 20.955 ;
        RECT 30.500 20.785 30.650 20.955 ;
        RECT 30.890 20.650 31.040 20.820 ;
        RECT 32.620 20.650 32.770 20.820 ;
        RECT 33.010 20.785 33.160 20.955 ;
        RECT 33.400 20.785 33.550 20.955 ;
        RECT 33.790 20.650 33.940 20.820 ;
        RECT 35.520 20.650 35.670 20.820 ;
        RECT 35.910 20.785 36.060 20.955 ;
        RECT 36.300 20.785 36.450 20.955 ;
        RECT 36.690 20.650 36.840 20.820 ;
        RECT 38.420 20.650 38.570 20.820 ;
        RECT 38.810 20.785 38.960 20.955 ;
        RECT 39.200 20.785 39.350 20.955 ;
        RECT 39.590 20.650 39.740 20.820 ;
        RECT 41.320 20.650 41.470 20.820 ;
        RECT 41.710 20.785 41.860 20.955 ;
        RECT 42.100 20.785 42.250 20.955 ;
        RECT 42.490 20.650 42.640 20.820 ;
        RECT 44.220 20.650 44.370 20.820 ;
        RECT 44.610 20.785 44.760 20.955 ;
        RECT 45.000 20.785 45.150 20.955 ;
        RECT 45.390 20.650 45.540 20.820 ;
        RECT 47.120 20.650 47.270 20.820 ;
        RECT 47.510 20.785 47.660 20.955 ;
        RECT 47.900 20.785 48.050 20.955 ;
        RECT 48.290 20.650 48.440 20.820 ;
        RECT 50.020 20.650 50.170 20.820 ;
        RECT 50.410 20.785 50.560 20.955 ;
        RECT 50.800 20.785 50.950 20.955 ;
        RECT 51.190 20.650 51.340 20.820 ;
        RECT 52.920 20.650 53.070 20.820 ;
        RECT 53.310 20.785 53.460 20.955 ;
        RECT 53.700 20.785 53.850 20.955 ;
        RECT 54.090 20.650 54.240 20.820 ;
        RECT 55.820 20.650 55.970 20.820 ;
        RECT 56.210 20.785 56.360 20.955 ;
        RECT 56.600 20.785 56.750 20.955 ;
        RECT 56.990 20.650 57.140 20.820 ;
        RECT 58.720 20.650 58.870 20.820 ;
        RECT 59.110 20.785 59.260 20.955 ;
        RECT 59.500 20.785 59.650 20.955 ;
        RECT 59.890 20.650 60.040 20.820 ;
        RECT 61.620 20.650 61.770 20.820 ;
        RECT 62.010 20.785 62.160 20.955 ;
        RECT 62.400 20.785 62.550 20.955 ;
        RECT 62.790 20.650 62.940 20.820 ;
        RECT 64.520 20.650 64.670 20.820 ;
        RECT 64.910 20.785 65.060 20.955 ;
        RECT 65.300 20.785 65.450 20.955 ;
        RECT 65.690 20.650 65.840 20.820 ;
        RECT 67.420 20.650 67.570 20.820 ;
        RECT 67.810 20.785 67.960 20.955 ;
        RECT 68.200 20.785 68.350 20.955 ;
        RECT 68.590 20.650 68.740 20.820 ;
        RECT 70.320 20.650 70.470 20.820 ;
        RECT 70.710 20.785 70.860 20.955 ;
        RECT 71.100 20.785 71.250 20.955 ;
        RECT 71.490 20.650 71.640 20.820 ;
        RECT 73.220 20.650 73.370 20.820 ;
        RECT 73.610 20.785 73.760 20.955 ;
        RECT 74.000 20.785 74.150 20.955 ;
        RECT 74.390 20.650 74.540 20.820 ;
        RECT 76.120 20.650 76.270 20.820 ;
        RECT 76.510 20.785 76.660 20.955 ;
        RECT 76.900 20.785 77.050 20.955 ;
        RECT 77.290 20.650 77.440 20.820 ;
        RECT 79.020 20.650 79.170 20.820 ;
        RECT 79.410 20.785 79.560 20.955 ;
        RECT 79.800 20.785 79.950 20.955 ;
        RECT 80.190 20.650 80.340 20.820 ;
        RECT 81.920 20.650 82.070 20.820 ;
        RECT 82.310 20.785 82.460 20.955 ;
        RECT 82.700 20.785 82.850 20.955 ;
        RECT 83.090 20.650 83.240 20.820 ;
        RECT 84.820 20.650 84.970 20.820 ;
        RECT 85.210 20.785 85.360 20.955 ;
        RECT 85.600 20.785 85.750 20.955 ;
        RECT 85.990 20.650 86.140 20.820 ;
        RECT 87.720 20.650 87.870 20.820 ;
        RECT 88.110 20.785 88.260 20.955 ;
        RECT 88.500 20.785 88.650 20.955 ;
        RECT 88.890 20.650 89.040 20.820 ;
        RECT 90.620 20.650 90.770 20.820 ;
        RECT 91.010 20.785 91.160 20.955 ;
        RECT 91.400 20.785 91.550 20.955 ;
        RECT 91.790 20.650 91.940 20.820 ;
        RECT 0.985 20.565 1.035 20.600 ;
        POLYGON 1.035 20.600 1.070 20.565 1.035 20.565 ;
        RECT 0.985 20.440 1.070 20.565 ;
        RECT 1.690 20.440 1.775 20.600 ;
        RECT 3.885 20.565 3.935 20.600 ;
        POLYGON 3.935 20.600 3.970 20.565 3.935 20.565 ;
        RECT 3.885 20.440 3.970 20.565 ;
        RECT 4.590 20.440 4.675 20.600 ;
        RECT 6.785 20.565 6.835 20.600 ;
        POLYGON 6.835 20.600 6.870 20.565 6.835 20.565 ;
        RECT 6.785 20.440 6.870 20.565 ;
        RECT 7.490 20.440 7.575 20.600 ;
        RECT 9.685 20.565 9.735 20.600 ;
        POLYGON 9.735 20.600 9.770 20.565 9.735 20.565 ;
        RECT 9.685 20.440 9.770 20.565 ;
        RECT 10.390 20.440 10.475 20.600 ;
        RECT 12.585 20.565 12.635 20.600 ;
        POLYGON 12.635 20.600 12.670 20.565 12.635 20.565 ;
        RECT 12.585 20.440 12.670 20.565 ;
        RECT 13.290 20.440 13.375 20.600 ;
        RECT 15.485 20.565 15.535 20.600 ;
        POLYGON 15.535 20.600 15.570 20.565 15.535 20.565 ;
        RECT 15.485 20.440 15.570 20.565 ;
        RECT 16.190 20.440 16.275 20.600 ;
        RECT 18.385 20.565 18.435 20.600 ;
        POLYGON 18.435 20.600 18.470 20.565 18.435 20.565 ;
        RECT 18.385 20.440 18.470 20.565 ;
        RECT 19.090 20.440 19.175 20.600 ;
        RECT 21.285 20.565 21.335 20.600 ;
        POLYGON 21.335 20.600 21.370 20.565 21.335 20.565 ;
        RECT 21.285 20.440 21.370 20.565 ;
        RECT 21.990 20.440 22.075 20.600 ;
        RECT 24.185 20.565 24.235 20.600 ;
        POLYGON 24.235 20.600 24.270 20.565 24.235 20.565 ;
        RECT 24.185 20.440 24.270 20.565 ;
        RECT 24.890 20.440 24.975 20.600 ;
        RECT 27.085 20.565 27.135 20.600 ;
        POLYGON 27.135 20.600 27.170 20.565 27.135 20.565 ;
        RECT 27.085 20.440 27.170 20.565 ;
        RECT 27.790 20.440 27.875 20.600 ;
        RECT 29.985 20.565 30.035 20.600 ;
        POLYGON 30.035 20.600 30.070 20.565 30.035 20.565 ;
        RECT 29.985 20.440 30.070 20.565 ;
        RECT 30.690 20.440 30.775 20.600 ;
        RECT 32.885 20.565 32.935 20.600 ;
        POLYGON 32.935 20.600 32.970 20.565 32.935 20.565 ;
        RECT 32.885 20.440 32.970 20.565 ;
        RECT 33.590 20.440 33.675 20.600 ;
        RECT 35.785 20.565 35.835 20.600 ;
        POLYGON 35.835 20.600 35.870 20.565 35.835 20.565 ;
        RECT 35.785 20.440 35.870 20.565 ;
        RECT 36.490 20.440 36.575 20.600 ;
        RECT 38.685 20.565 38.735 20.600 ;
        POLYGON 38.735 20.600 38.770 20.565 38.735 20.565 ;
        RECT 38.685 20.440 38.770 20.565 ;
        RECT 39.390 20.440 39.475 20.600 ;
        RECT 41.585 20.565 41.635 20.600 ;
        POLYGON 41.635 20.600 41.670 20.565 41.635 20.565 ;
        RECT 41.585 20.440 41.670 20.565 ;
        RECT 42.290 20.440 42.375 20.600 ;
        RECT 44.485 20.565 44.535 20.600 ;
        POLYGON 44.535 20.600 44.570 20.565 44.535 20.565 ;
        RECT 44.485 20.440 44.570 20.565 ;
        RECT 45.190 20.440 45.275 20.600 ;
        RECT 47.385 20.565 47.435 20.600 ;
        POLYGON 47.435 20.600 47.470 20.565 47.435 20.565 ;
        RECT 47.385 20.440 47.470 20.565 ;
        RECT 48.090 20.440 48.175 20.600 ;
        RECT 50.285 20.565 50.335 20.600 ;
        POLYGON 50.335 20.600 50.370 20.565 50.335 20.565 ;
        RECT 50.285 20.440 50.370 20.565 ;
        RECT 50.990 20.440 51.075 20.600 ;
        RECT 53.185 20.565 53.235 20.600 ;
        POLYGON 53.235 20.600 53.270 20.565 53.235 20.565 ;
        RECT 53.185 20.440 53.270 20.565 ;
        RECT 53.890 20.440 53.975 20.600 ;
        RECT 56.085 20.565 56.135 20.600 ;
        POLYGON 56.135 20.600 56.170 20.565 56.135 20.565 ;
        RECT 56.085 20.440 56.170 20.565 ;
        RECT 56.790 20.440 56.875 20.600 ;
        RECT 58.985 20.565 59.035 20.600 ;
        POLYGON 59.035 20.600 59.070 20.565 59.035 20.565 ;
        RECT 58.985 20.440 59.070 20.565 ;
        RECT 59.690 20.440 59.775 20.600 ;
        RECT 61.885 20.565 61.935 20.600 ;
        POLYGON 61.935 20.600 61.970 20.565 61.935 20.565 ;
        RECT 61.885 20.440 61.970 20.565 ;
        RECT 62.590 20.440 62.675 20.600 ;
        RECT 64.785 20.565 64.835 20.600 ;
        POLYGON 64.835 20.600 64.870 20.565 64.835 20.565 ;
        RECT 64.785 20.440 64.870 20.565 ;
        RECT 65.490 20.440 65.575 20.600 ;
        RECT 67.685 20.565 67.735 20.600 ;
        POLYGON 67.735 20.600 67.770 20.565 67.735 20.565 ;
        RECT 67.685 20.440 67.770 20.565 ;
        RECT 68.390 20.440 68.475 20.600 ;
        RECT 70.585 20.565 70.635 20.600 ;
        POLYGON 70.635 20.600 70.670 20.565 70.635 20.565 ;
        RECT 70.585 20.440 70.670 20.565 ;
        RECT 71.290 20.440 71.375 20.600 ;
        RECT 73.485 20.565 73.535 20.600 ;
        POLYGON 73.535 20.600 73.570 20.565 73.535 20.565 ;
        RECT 73.485 20.440 73.570 20.565 ;
        RECT 74.190 20.440 74.275 20.600 ;
        RECT 76.385 20.565 76.435 20.600 ;
        POLYGON 76.435 20.600 76.470 20.565 76.435 20.565 ;
        RECT 76.385 20.440 76.470 20.565 ;
        RECT 77.090 20.440 77.175 20.600 ;
        RECT 79.285 20.565 79.335 20.600 ;
        POLYGON 79.335 20.600 79.370 20.565 79.335 20.565 ;
        RECT 79.285 20.440 79.370 20.565 ;
        RECT 79.990 20.440 80.075 20.600 ;
        RECT 82.185 20.565 82.235 20.600 ;
        POLYGON 82.235 20.600 82.270 20.565 82.235 20.565 ;
        RECT 82.185 20.440 82.270 20.565 ;
        RECT 82.890 20.440 82.975 20.600 ;
        RECT 85.085 20.565 85.135 20.600 ;
        POLYGON 85.135 20.600 85.170 20.565 85.135 20.565 ;
        RECT 85.085 20.440 85.170 20.565 ;
        RECT 85.790 20.440 85.875 20.600 ;
        RECT 87.985 20.565 88.035 20.600 ;
        POLYGON 88.035 20.600 88.070 20.565 88.035 20.565 ;
        RECT 87.985 20.440 88.070 20.565 ;
        RECT 88.690 20.440 88.775 20.600 ;
        RECT 90.885 20.565 90.935 20.600 ;
        POLYGON 90.935 20.600 90.970 20.565 90.935 20.565 ;
        RECT 90.885 20.440 90.970 20.565 ;
        RECT 91.590 20.440 91.675 20.600 ;
        RECT 0.775 19.820 0.850 19.960 ;
        RECT 0.990 19.770 1.065 19.910 ;
        RECT 1.695 19.830 1.755 19.910 ;
        POLYGON 1.695 19.830 1.755 19.830 1.755 19.770 ;
        RECT 1.910 19.820 1.985 19.960 ;
        RECT 3.675 19.820 3.750 19.960 ;
        RECT 3.890 19.770 3.965 19.910 ;
        RECT 4.595 19.830 4.655 19.910 ;
        POLYGON 4.595 19.830 4.655 19.830 4.655 19.770 ;
        RECT 4.810 19.820 4.885 19.960 ;
        RECT 6.575 19.820 6.650 19.960 ;
        RECT 6.790 19.770 6.865 19.910 ;
        RECT 7.495 19.830 7.555 19.910 ;
        POLYGON 7.495 19.830 7.555 19.830 7.555 19.770 ;
        RECT 7.710 19.820 7.785 19.960 ;
        RECT 9.475 19.820 9.550 19.960 ;
        RECT 9.690 19.770 9.765 19.910 ;
        RECT 10.395 19.830 10.455 19.910 ;
        POLYGON 10.395 19.830 10.455 19.830 10.455 19.770 ;
        RECT 10.610 19.820 10.685 19.960 ;
        RECT 12.375 19.820 12.450 19.960 ;
        RECT 12.590 19.770 12.665 19.910 ;
        RECT 13.295 19.830 13.355 19.910 ;
        POLYGON 13.295 19.830 13.355 19.830 13.355 19.770 ;
        RECT 13.510 19.820 13.585 19.960 ;
        RECT 15.275 19.820 15.350 19.960 ;
        RECT 15.490 19.770 15.565 19.910 ;
        RECT 16.195 19.830 16.255 19.910 ;
        POLYGON 16.195 19.830 16.255 19.830 16.255 19.770 ;
        RECT 16.410 19.820 16.485 19.960 ;
        RECT 18.175 19.820 18.250 19.960 ;
        RECT 18.390 19.770 18.465 19.910 ;
        RECT 19.095 19.830 19.155 19.910 ;
        POLYGON 19.095 19.830 19.155 19.830 19.155 19.770 ;
        RECT 19.310 19.820 19.385 19.960 ;
        RECT 21.075 19.820 21.150 19.960 ;
        RECT 21.290 19.770 21.365 19.910 ;
        RECT 21.995 19.830 22.055 19.910 ;
        POLYGON 21.995 19.830 22.055 19.830 22.055 19.770 ;
        RECT 22.210 19.820 22.285 19.960 ;
        RECT 23.975 19.820 24.050 19.960 ;
        RECT 24.190 19.770 24.265 19.910 ;
        RECT 24.895 19.830 24.955 19.910 ;
        POLYGON 24.895 19.830 24.955 19.830 24.955 19.770 ;
        RECT 25.110 19.820 25.185 19.960 ;
        RECT 26.875 19.820 26.950 19.960 ;
        RECT 27.090 19.770 27.165 19.910 ;
        RECT 27.795 19.830 27.855 19.910 ;
        POLYGON 27.795 19.830 27.855 19.830 27.855 19.770 ;
        RECT 28.010 19.820 28.085 19.960 ;
        RECT 29.775 19.820 29.850 19.960 ;
        RECT 29.990 19.770 30.065 19.910 ;
        RECT 30.695 19.830 30.755 19.910 ;
        POLYGON 30.695 19.830 30.755 19.830 30.755 19.770 ;
        RECT 30.910 19.820 30.985 19.960 ;
        RECT 32.675 19.820 32.750 19.960 ;
        RECT 32.890 19.770 32.965 19.910 ;
        RECT 33.595 19.830 33.655 19.910 ;
        POLYGON 33.595 19.830 33.655 19.830 33.655 19.770 ;
        RECT 33.810 19.820 33.885 19.960 ;
        RECT 35.575 19.820 35.650 19.960 ;
        RECT 35.790 19.770 35.865 19.910 ;
        RECT 36.495 19.830 36.555 19.910 ;
        POLYGON 36.495 19.830 36.555 19.830 36.555 19.770 ;
        RECT 36.710 19.820 36.785 19.960 ;
        RECT 38.475 19.820 38.550 19.960 ;
        RECT 38.690 19.770 38.765 19.910 ;
        RECT 39.395 19.830 39.455 19.910 ;
        POLYGON 39.395 19.830 39.455 19.830 39.455 19.770 ;
        RECT 39.610 19.820 39.685 19.960 ;
        RECT 41.375 19.820 41.450 19.960 ;
        RECT 41.590 19.770 41.665 19.910 ;
        RECT 42.295 19.830 42.355 19.910 ;
        POLYGON 42.295 19.830 42.355 19.830 42.355 19.770 ;
        RECT 42.510 19.820 42.585 19.960 ;
        RECT 44.275 19.820 44.350 19.960 ;
        RECT 44.490 19.770 44.565 19.910 ;
        RECT 45.195 19.830 45.255 19.910 ;
        POLYGON 45.195 19.830 45.255 19.830 45.255 19.770 ;
        RECT 45.410 19.820 45.485 19.960 ;
        RECT 47.175 19.820 47.250 19.960 ;
        RECT 47.390 19.770 47.465 19.910 ;
        RECT 48.095 19.830 48.155 19.910 ;
        POLYGON 48.095 19.830 48.155 19.830 48.155 19.770 ;
        RECT 48.310 19.820 48.385 19.960 ;
        RECT 50.075 19.820 50.150 19.960 ;
        RECT 50.290 19.770 50.365 19.910 ;
        RECT 50.995 19.830 51.055 19.910 ;
        POLYGON 50.995 19.830 51.055 19.830 51.055 19.770 ;
        RECT 51.210 19.820 51.285 19.960 ;
        RECT 52.975 19.820 53.050 19.960 ;
        RECT 53.190 19.770 53.265 19.910 ;
        RECT 53.895 19.830 53.955 19.910 ;
        POLYGON 53.895 19.830 53.955 19.830 53.955 19.770 ;
        RECT 54.110 19.820 54.185 19.960 ;
        RECT 55.875 19.820 55.950 19.960 ;
        RECT 56.090 19.770 56.165 19.910 ;
        RECT 56.795 19.830 56.855 19.910 ;
        POLYGON 56.795 19.830 56.855 19.830 56.855 19.770 ;
        RECT 57.010 19.820 57.085 19.960 ;
        RECT 58.775 19.820 58.850 19.960 ;
        RECT 58.990 19.770 59.065 19.910 ;
        RECT 59.695 19.830 59.755 19.910 ;
        POLYGON 59.695 19.830 59.755 19.830 59.755 19.770 ;
        RECT 59.910 19.820 59.985 19.960 ;
        RECT 61.675 19.820 61.750 19.960 ;
        RECT 61.890 19.770 61.965 19.910 ;
        RECT 62.595 19.830 62.655 19.910 ;
        POLYGON 62.595 19.830 62.655 19.830 62.655 19.770 ;
        RECT 62.810 19.820 62.885 19.960 ;
        RECT 64.575 19.820 64.650 19.960 ;
        RECT 64.790 19.770 64.865 19.910 ;
        RECT 65.495 19.830 65.555 19.910 ;
        POLYGON 65.495 19.830 65.555 19.830 65.555 19.770 ;
        RECT 65.710 19.820 65.785 19.960 ;
        RECT 67.475 19.820 67.550 19.960 ;
        RECT 67.690 19.770 67.765 19.910 ;
        RECT 68.395 19.830 68.455 19.910 ;
        POLYGON 68.395 19.830 68.455 19.830 68.455 19.770 ;
        RECT 68.610 19.820 68.685 19.960 ;
        RECT 70.375 19.820 70.450 19.960 ;
        RECT 70.590 19.770 70.665 19.910 ;
        RECT 71.295 19.830 71.355 19.910 ;
        POLYGON 71.295 19.830 71.355 19.830 71.355 19.770 ;
        RECT 71.510 19.820 71.585 19.960 ;
        RECT 73.275 19.820 73.350 19.960 ;
        RECT 73.490 19.770 73.565 19.910 ;
        RECT 74.195 19.830 74.255 19.910 ;
        POLYGON 74.195 19.830 74.255 19.830 74.255 19.770 ;
        RECT 74.410 19.820 74.485 19.960 ;
        RECT 76.175 19.820 76.250 19.960 ;
        RECT 76.390 19.770 76.465 19.910 ;
        RECT 77.095 19.830 77.155 19.910 ;
        POLYGON 77.095 19.830 77.155 19.830 77.155 19.770 ;
        RECT 77.310 19.820 77.385 19.960 ;
        RECT 79.075 19.820 79.150 19.960 ;
        RECT 79.290 19.770 79.365 19.910 ;
        RECT 79.995 19.830 80.055 19.910 ;
        POLYGON 79.995 19.830 80.055 19.830 80.055 19.770 ;
        RECT 80.210 19.820 80.285 19.960 ;
        RECT 81.975 19.820 82.050 19.960 ;
        RECT 82.190 19.770 82.265 19.910 ;
        RECT 82.895 19.830 82.955 19.910 ;
        POLYGON 82.895 19.830 82.955 19.830 82.955 19.770 ;
        RECT 83.110 19.820 83.185 19.960 ;
        RECT 84.875 19.820 84.950 19.960 ;
        RECT 85.090 19.770 85.165 19.910 ;
        RECT 85.795 19.830 85.855 19.910 ;
        POLYGON 85.795 19.830 85.855 19.830 85.855 19.770 ;
        RECT 86.010 19.820 86.085 19.960 ;
        RECT 87.775 19.820 87.850 19.960 ;
        RECT 87.990 19.770 88.065 19.910 ;
        RECT 88.695 19.830 88.755 19.910 ;
        POLYGON 88.695 19.830 88.755 19.830 88.755 19.770 ;
        RECT 88.910 19.820 88.985 19.960 ;
        RECT 90.675 19.820 90.750 19.960 ;
        RECT 90.890 19.770 90.965 19.910 ;
        RECT 91.595 19.830 91.655 19.910 ;
        POLYGON 91.595 19.830 91.655 19.830 91.655 19.770 ;
        RECT 91.810 19.820 91.885 19.960 ;
        RECT 0.720 19.300 0.870 19.470 ;
        RECT 1.110 19.435 1.260 19.605 ;
        RECT 1.500 19.435 1.650 19.605 ;
        RECT 1.890 19.300 2.040 19.470 ;
        RECT 3.620 19.300 3.770 19.470 ;
        RECT 4.010 19.435 4.160 19.605 ;
        RECT 4.400 19.435 4.550 19.605 ;
        RECT 4.790 19.300 4.940 19.470 ;
        RECT 6.520 19.300 6.670 19.470 ;
        RECT 6.910 19.435 7.060 19.605 ;
        RECT 7.300 19.435 7.450 19.605 ;
        RECT 7.690 19.300 7.840 19.470 ;
        RECT 9.420 19.300 9.570 19.470 ;
        RECT 9.810 19.435 9.960 19.605 ;
        RECT 10.200 19.435 10.350 19.605 ;
        RECT 10.590 19.300 10.740 19.470 ;
        RECT 12.320 19.300 12.470 19.470 ;
        RECT 12.710 19.435 12.860 19.605 ;
        RECT 13.100 19.435 13.250 19.605 ;
        RECT 13.490 19.300 13.640 19.470 ;
        RECT 15.220 19.300 15.370 19.470 ;
        RECT 15.610 19.435 15.760 19.605 ;
        RECT 16.000 19.435 16.150 19.605 ;
        RECT 16.390 19.300 16.540 19.470 ;
        RECT 18.120 19.300 18.270 19.470 ;
        RECT 18.510 19.435 18.660 19.605 ;
        RECT 18.900 19.435 19.050 19.605 ;
        RECT 19.290 19.300 19.440 19.470 ;
        RECT 21.020 19.300 21.170 19.470 ;
        RECT 21.410 19.435 21.560 19.605 ;
        RECT 21.800 19.435 21.950 19.605 ;
        RECT 22.190 19.300 22.340 19.470 ;
        RECT 23.920 19.300 24.070 19.470 ;
        RECT 24.310 19.435 24.460 19.605 ;
        RECT 24.700 19.435 24.850 19.605 ;
        RECT 25.090 19.300 25.240 19.470 ;
        RECT 26.820 19.300 26.970 19.470 ;
        RECT 27.210 19.435 27.360 19.605 ;
        RECT 27.600 19.435 27.750 19.605 ;
        RECT 27.990 19.300 28.140 19.470 ;
        RECT 29.720 19.300 29.870 19.470 ;
        RECT 30.110 19.435 30.260 19.605 ;
        RECT 30.500 19.435 30.650 19.605 ;
        RECT 30.890 19.300 31.040 19.470 ;
        RECT 32.620 19.300 32.770 19.470 ;
        RECT 33.010 19.435 33.160 19.605 ;
        RECT 33.400 19.435 33.550 19.605 ;
        RECT 33.790 19.300 33.940 19.470 ;
        RECT 35.520 19.300 35.670 19.470 ;
        RECT 35.910 19.435 36.060 19.605 ;
        RECT 36.300 19.435 36.450 19.605 ;
        RECT 36.690 19.300 36.840 19.470 ;
        RECT 38.420 19.300 38.570 19.470 ;
        RECT 38.810 19.435 38.960 19.605 ;
        RECT 39.200 19.435 39.350 19.605 ;
        RECT 39.590 19.300 39.740 19.470 ;
        RECT 41.320 19.300 41.470 19.470 ;
        RECT 41.710 19.435 41.860 19.605 ;
        RECT 42.100 19.435 42.250 19.605 ;
        RECT 42.490 19.300 42.640 19.470 ;
        RECT 44.220 19.300 44.370 19.470 ;
        RECT 44.610 19.435 44.760 19.605 ;
        RECT 45.000 19.435 45.150 19.605 ;
        RECT 45.390 19.300 45.540 19.470 ;
        RECT 47.120 19.300 47.270 19.470 ;
        RECT 47.510 19.435 47.660 19.605 ;
        RECT 47.900 19.435 48.050 19.605 ;
        RECT 48.290 19.300 48.440 19.470 ;
        RECT 50.020 19.300 50.170 19.470 ;
        RECT 50.410 19.435 50.560 19.605 ;
        RECT 50.800 19.435 50.950 19.605 ;
        RECT 51.190 19.300 51.340 19.470 ;
        RECT 52.920 19.300 53.070 19.470 ;
        RECT 53.310 19.435 53.460 19.605 ;
        RECT 53.700 19.435 53.850 19.605 ;
        RECT 54.090 19.300 54.240 19.470 ;
        RECT 55.820 19.300 55.970 19.470 ;
        RECT 56.210 19.435 56.360 19.605 ;
        RECT 56.600 19.435 56.750 19.605 ;
        RECT 56.990 19.300 57.140 19.470 ;
        RECT 58.720 19.300 58.870 19.470 ;
        RECT 59.110 19.435 59.260 19.605 ;
        RECT 59.500 19.435 59.650 19.605 ;
        RECT 59.890 19.300 60.040 19.470 ;
        RECT 61.620 19.300 61.770 19.470 ;
        RECT 62.010 19.435 62.160 19.605 ;
        RECT 62.400 19.435 62.550 19.605 ;
        RECT 62.790 19.300 62.940 19.470 ;
        RECT 64.520 19.300 64.670 19.470 ;
        RECT 64.910 19.435 65.060 19.605 ;
        RECT 65.300 19.435 65.450 19.605 ;
        RECT 65.690 19.300 65.840 19.470 ;
        RECT 67.420 19.300 67.570 19.470 ;
        RECT 67.810 19.435 67.960 19.605 ;
        RECT 68.200 19.435 68.350 19.605 ;
        RECT 68.590 19.300 68.740 19.470 ;
        RECT 70.320 19.300 70.470 19.470 ;
        RECT 70.710 19.435 70.860 19.605 ;
        RECT 71.100 19.435 71.250 19.605 ;
        RECT 71.490 19.300 71.640 19.470 ;
        RECT 73.220 19.300 73.370 19.470 ;
        RECT 73.610 19.435 73.760 19.605 ;
        RECT 74.000 19.435 74.150 19.605 ;
        RECT 74.390 19.300 74.540 19.470 ;
        RECT 76.120 19.300 76.270 19.470 ;
        RECT 76.510 19.435 76.660 19.605 ;
        RECT 76.900 19.435 77.050 19.605 ;
        RECT 77.290 19.300 77.440 19.470 ;
        RECT 79.020 19.300 79.170 19.470 ;
        RECT 79.410 19.435 79.560 19.605 ;
        RECT 79.800 19.435 79.950 19.605 ;
        RECT 80.190 19.300 80.340 19.470 ;
        RECT 81.920 19.300 82.070 19.470 ;
        RECT 82.310 19.435 82.460 19.605 ;
        RECT 82.700 19.435 82.850 19.605 ;
        RECT 83.090 19.300 83.240 19.470 ;
        RECT 84.820 19.300 84.970 19.470 ;
        RECT 85.210 19.435 85.360 19.605 ;
        RECT 85.600 19.435 85.750 19.605 ;
        RECT 85.990 19.300 86.140 19.470 ;
        RECT 87.720 19.300 87.870 19.470 ;
        RECT 88.110 19.435 88.260 19.605 ;
        RECT 88.500 19.435 88.650 19.605 ;
        RECT 88.890 19.300 89.040 19.470 ;
        RECT 90.620 19.300 90.770 19.470 ;
        RECT 91.010 19.435 91.160 19.605 ;
        RECT 91.400 19.435 91.550 19.605 ;
        RECT 91.790 19.300 91.940 19.470 ;
        RECT 0.985 19.215 1.035 19.250 ;
        POLYGON 1.035 19.250 1.070 19.215 1.035 19.215 ;
        RECT 0.985 19.090 1.070 19.215 ;
        RECT 1.690 19.090 1.775 19.250 ;
        RECT 3.885 19.215 3.935 19.250 ;
        POLYGON 3.935 19.250 3.970 19.215 3.935 19.215 ;
        RECT 3.885 19.090 3.970 19.215 ;
        RECT 4.590 19.090 4.675 19.250 ;
        RECT 6.785 19.215 6.835 19.250 ;
        POLYGON 6.835 19.250 6.870 19.215 6.835 19.215 ;
        RECT 6.785 19.090 6.870 19.215 ;
        RECT 7.490 19.090 7.575 19.250 ;
        RECT 9.685 19.215 9.735 19.250 ;
        POLYGON 9.735 19.250 9.770 19.215 9.735 19.215 ;
        RECT 9.685 19.090 9.770 19.215 ;
        RECT 10.390 19.090 10.475 19.250 ;
        RECT 12.585 19.215 12.635 19.250 ;
        POLYGON 12.635 19.250 12.670 19.215 12.635 19.215 ;
        RECT 12.585 19.090 12.670 19.215 ;
        RECT 13.290 19.090 13.375 19.250 ;
        RECT 15.485 19.215 15.535 19.250 ;
        POLYGON 15.535 19.250 15.570 19.215 15.535 19.215 ;
        RECT 15.485 19.090 15.570 19.215 ;
        RECT 16.190 19.090 16.275 19.250 ;
        RECT 18.385 19.215 18.435 19.250 ;
        POLYGON 18.435 19.250 18.470 19.215 18.435 19.215 ;
        RECT 18.385 19.090 18.470 19.215 ;
        RECT 19.090 19.090 19.175 19.250 ;
        RECT 21.285 19.215 21.335 19.250 ;
        POLYGON 21.335 19.250 21.370 19.215 21.335 19.215 ;
        RECT 21.285 19.090 21.370 19.215 ;
        RECT 21.990 19.090 22.075 19.250 ;
        RECT 24.185 19.215 24.235 19.250 ;
        POLYGON 24.235 19.250 24.270 19.215 24.235 19.215 ;
        RECT 24.185 19.090 24.270 19.215 ;
        RECT 24.890 19.090 24.975 19.250 ;
        RECT 27.085 19.215 27.135 19.250 ;
        POLYGON 27.135 19.250 27.170 19.215 27.135 19.215 ;
        RECT 27.085 19.090 27.170 19.215 ;
        RECT 27.790 19.090 27.875 19.250 ;
        RECT 29.985 19.215 30.035 19.250 ;
        POLYGON 30.035 19.250 30.070 19.215 30.035 19.215 ;
        RECT 29.985 19.090 30.070 19.215 ;
        RECT 30.690 19.090 30.775 19.250 ;
        RECT 32.885 19.215 32.935 19.250 ;
        POLYGON 32.935 19.250 32.970 19.215 32.935 19.215 ;
        RECT 32.885 19.090 32.970 19.215 ;
        RECT 33.590 19.090 33.675 19.250 ;
        RECT 35.785 19.215 35.835 19.250 ;
        POLYGON 35.835 19.250 35.870 19.215 35.835 19.215 ;
        RECT 35.785 19.090 35.870 19.215 ;
        RECT 36.490 19.090 36.575 19.250 ;
        RECT 38.685 19.215 38.735 19.250 ;
        POLYGON 38.735 19.250 38.770 19.215 38.735 19.215 ;
        RECT 38.685 19.090 38.770 19.215 ;
        RECT 39.390 19.090 39.475 19.250 ;
        RECT 41.585 19.215 41.635 19.250 ;
        POLYGON 41.635 19.250 41.670 19.215 41.635 19.215 ;
        RECT 41.585 19.090 41.670 19.215 ;
        RECT 42.290 19.090 42.375 19.250 ;
        RECT 44.485 19.215 44.535 19.250 ;
        POLYGON 44.535 19.250 44.570 19.215 44.535 19.215 ;
        RECT 44.485 19.090 44.570 19.215 ;
        RECT 45.190 19.090 45.275 19.250 ;
        RECT 47.385 19.215 47.435 19.250 ;
        POLYGON 47.435 19.250 47.470 19.215 47.435 19.215 ;
        RECT 47.385 19.090 47.470 19.215 ;
        RECT 48.090 19.090 48.175 19.250 ;
        RECT 50.285 19.215 50.335 19.250 ;
        POLYGON 50.335 19.250 50.370 19.215 50.335 19.215 ;
        RECT 50.285 19.090 50.370 19.215 ;
        RECT 50.990 19.090 51.075 19.250 ;
        RECT 53.185 19.215 53.235 19.250 ;
        POLYGON 53.235 19.250 53.270 19.215 53.235 19.215 ;
        RECT 53.185 19.090 53.270 19.215 ;
        RECT 53.890 19.090 53.975 19.250 ;
        RECT 56.085 19.215 56.135 19.250 ;
        POLYGON 56.135 19.250 56.170 19.215 56.135 19.215 ;
        RECT 56.085 19.090 56.170 19.215 ;
        RECT 56.790 19.090 56.875 19.250 ;
        RECT 58.985 19.215 59.035 19.250 ;
        POLYGON 59.035 19.250 59.070 19.215 59.035 19.215 ;
        RECT 58.985 19.090 59.070 19.215 ;
        RECT 59.690 19.090 59.775 19.250 ;
        RECT 61.885 19.215 61.935 19.250 ;
        POLYGON 61.935 19.250 61.970 19.215 61.935 19.215 ;
        RECT 61.885 19.090 61.970 19.215 ;
        RECT 62.590 19.090 62.675 19.250 ;
        RECT 64.785 19.215 64.835 19.250 ;
        POLYGON 64.835 19.250 64.870 19.215 64.835 19.215 ;
        RECT 64.785 19.090 64.870 19.215 ;
        RECT 65.490 19.090 65.575 19.250 ;
        RECT 67.685 19.215 67.735 19.250 ;
        POLYGON 67.735 19.250 67.770 19.215 67.735 19.215 ;
        RECT 67.685 19.090 67.770 19.215 ;
        RECT 68.390 19.090 68.475 19.250 ;
        RECT 70.585 19.215 70.635 19.250 ;
        POLYGON 70.635 19.250 70.670 19.215 70.635 19.215 ;
        RECT 70.585 19.090 70.670 19.215 ;
        RECT 71.290 19.090 71.375 19.250 ;
        RECT 73.485 19.215 73.535 19.250 ;
        POLYGON 73.535 19.250 73.570 19.215 73.535 19.215 ;
        RECT 73.485 19.090 73.570 19.215 ;
        RECT 74.190 19.090 74.275 19.250 ;
        RECT 76.385 19.215 76.435 19.250 ;
        POLYGON 76.435 19.250 76.470 19.215 76.435 19.215 ;
        RECT 76.385 19.090 76.470 19.215 ;
        RECT 77.090 19.090 77.175 19.250 ;
        RECT 79.285 19.215 79.335 19.250 ;
        POLYGON 79.335 19.250 79.370 19.215 79.335 19.215 ;
        RECT 79.285 19.090 79.370 19.215 ;
        RECT 79.990 19.090 80.075 19.250 ;
        RECT 82.185 19.215 82.235 19.250 ;
        POLYGON 82.235 19.250 82.270 19.215 82.235 19.215 ;
        RECT 82.185 19.090 82.270 19.215 ;
        RECT 82.890 19.090 82.975 19.250 ;
        RECT 85.085 19.215 85.135 19.250 ;
        POLYGON 85.135 19.250 85.170 19.215 85.135 19.215 ;
        RECT 85.085 19.090 85.170 19.215 ;
        RECT 85.790 19.090 85.875 19.250 ;
        RECT 87.985 19.215 88.035 19.250 ;
        POLYGON 88.035 19.250 88.070 19.215 88.035 19.215 ;
        RECT 87.985 19.090 88.070 19.215 ;
        RECT 88.690 19.090 88.775 19.250 ;
        RECT 90.885 19.215 90.935 19.250 ;
        POLYGON 90.935 19.250 90.970 19.215 90.935 19.215 ;
        RECT 90.885 19.090 90.970 19.215 ;
        RECT 91.590 19.090 91.675 19.250 ;
        RECT 0.775 18.470 0.850 18.610 ;
        RECT 0.990 18.420 1.065 18.560 ;
        RECT 1.695 18.480 1.755 18.560 ;
        POLYGON 1.695 18.480 1.755 18.480 1.755 18.420 ;
        RECT 1.910 18.470 1.985 18.610 ;
        RECT 3.675 18.470 3.750 18.610 ;
        RECT 3.890 18.420 3.965 18.560 ;
        RECT 4.595 18.480 4.655 18.560 ;
        POLYGON 4.595 18.480 4.655 18.480 4.655 18.420 ;
        RECT 4.810 18.470 4.885 18.610 ;
        RECT 6.575 18.470 6.650 18.610 ;
        RECT 6.790 18.420 6.865 18.560 ;
        RECT 7.495 18.480 7.555 18.560 ;
        POLYGON 7.495 18.480 7.555 18.480 7.555 18.420 ;
        RECT 7.710 18.470 7.785 18.610 ;
        RECT 9.475 18.470 9.550 18.610 ;
        RECT 9.690 18.420 9.765 18.560 ;
        RECT 10.395 18.480 10.455 18.560 ;
        POLYGON 10.395 18.480 10.455 18.480 10.455 18.420 ;
        RECT 10.610 18.470 10.685 18.610 ;
        RECT 12.375 18.470 12.450 18.610 ;
        RECT 12.590 18.420 12.665 18.560 ;
        RECT 13.295 18.480 13.355 18.560 ;
        POLYGON 13.295 18.480 13.355 18.480 13.355 18.420 ;
        RECT 13.510 18.470 13.585 18.610 ;
        RECT 15.275 18.470 15.350 18.610 ;
        RECT 15.490 18.420 15.565 18.560 ;
        RECT 16.195 18.480 16.255 18.560 ;
        POLYGON 16.195 18.480 16.255 18.480 16.255 18.420 ;
        RECT 16.410 18.470 16.485 18.610 ;
        RECT 18.175 18.470 18.250 18.610 ;
        RECT 18.390 18.420 18.465 18.560 ;
        RECT 19.095 18.480 19.155 18.560 ;
        POLYGON 19.095 18.480 19.155 18.480 19.155 18.420 ;
        RECT 19.310 18.470 19.385 18.610 ;
        RECT 21.075 18.470 21.150 18.610 ;
        RECT 21.290 18.420 21.365 18.560 ;
        RECT 21.995 18.480 22.055 18.560 ;
        POLYGON 21.995 18.480 22.055 18.480 22.055 18.420 ;
        RECT 22.210 18.470 22.285 18.610 ;
        RECT 23.975 18.470 24.050 18.610 ;
        RECT 24.190 18.420 24.265 18.560 ;
        RECT 24.895 18.480 24.955 18.560 ;
        POLYGON 24.895 18.480 24.955 18.480 24.955 18.420 ;
        RECT 25.110 18.470 25.185 18.610 ;
        RECT 26.875 18.470 26.950 18.610 ;
        RECT 27.090 18.420 27.165 18.560 ;
        RECT 27.795 18.480 27.855 18.560 ;
        POLYGON 27.795 18.480 27.855 18.480 27.855 18.420 ;
        RECT 28.010 18.470 28.085 18.610 ;
        RECT 29.775 18.470 29.850 18.610 ;
        RECT 29.990 18.420 30.065 18.560 ;
        RECT 30.695 18.480 30.755 18.560 ;
        POLYGON 30.695 18.480 30.755 18.480 30.755 18.420 ;
        RECT 30.910 18.470 30.985 18.610 ;
        RECT 32.675 18.470 32.750 18.610 ;
        RECT 32.890 18.420 32.965 18.560 ;
        RECT 33.595 18.480 33.655 18.560 ;
        POLYGON 33.595 18.480 33.655 18.480 33.655 18.420 ;
        RECT 33.810 18.470 33.885 18.610 ;
        RECT 35.575 18.470 35.650 18.610 ;
        RECT 35.790 18.420 35.865 18.560 ;
        RECT 36.495 18.480 36.555 18.560 ;
        POLYGON 36.495 18.480 36.555 18.480 36.555 18.420 ;
        RECT 36.710 18.470 36.785 18.610 ;
        RECT 38.475 18.470 38.550 18.610 ;
        RECT 38.690 18.420 38.765 18.560 ;
        RECT 39.395 18.480 39.455 18.560 ;
        POLYGON 39.395 18.480 39.455 18.480 39.455 18.420 ;
        RECT 39.610 18.470 39.685 18.610 ;
        RECT 41.375 18.470 41.450 18.610 ;
        RECT 41.590 18.420 41.665 18.560 ;
        RECT 42.295 18.480 42.355 18.560 ;
        POLYGON 42.295 18.480 42.355 18.480 42.355 18.420 ;
        RECT 42.510 18.470 42.585 18.610 ;
        RECT 44.275 18.470 44.350 18.610 ;
        RECT 44.490 18.420 44.565 18.560 ;
        RECT 45.195 18.480 45.255 18.560 ;
        POLYGON 45.195 18.480 45.255 18.480 45.255 18.420 ;
        RECT 45.410 18.470 45.485 18.610 ;
        RECT 47.175 18.470 47.250 18.610 ;
        RECT 47.390 18.420 47.465 18.560 ;
        RECT 48.095 18.480 48.155 18.560 ;
        POLYGON 48.095 18.480 48.155 18.480 48.155 18.420 ;
        RECT 48.310 18.470 48.385 18.610 ;
        RECT 50.075 18.470 50.150 18.610 ;
        RECT 50.290 18.420 50.365 18.560 ;
        RECT 50.995 18.480 51.055 18.560 ;
        POLYGON 50.995 18.480 51.055 18.480 51.055 18.420 ;
        RECT 51.210 18.470 51.285 18.610 ;
        RECT 52.975 18.470 53.050 18.610 ;
        RECT 53.190 18.420 53.265 18.560 ;
        RECT 53.895 18.480 53.955 18.560 ;
        POLYGON 53.895 18.480 53.955 18.480 53.955 18.420 ;
        RECT 54.110 18.470 54.185 18.610 ;
        RECT 55.875 18.470 55.950 18.610 ;
        RECT 56.090 18.420 56.165 18.560 ;
        RECT 56.795 18.480 56.855 18.560 ;
        POLYGON 56.795 18.480 56.855 18.480 56.855 18.420 ;
        RECT 57.010 18.470 57.085 18.610 ;
        RECT 58.775 18.470 58.850 18.610 ;
        RECT 58.990 18.420 59.065 18.560 ;
        RECT 59.695 18.480 59.755 18.560 ;
        POLYGON 59.695 18.480 59.755 18.480 59.755 18.420 ;
        RECT 59.910 18.470 59.985 18.610 ;
        RECT 61.675 18.470 61.750 18.610 ;
        RECT 61.890 18.420 61.965 18.560 ;
        RECT 62.595 18.480 62.655 18.560 ;
        POLYGON 62.595 18.480 62.655 18.480 62.655 18.420 ;
        RECT 62.810 18.470 62.885 18.610 ;
        RECT 64.575 18.470 64.650 18.610 ;
        RECT 64.790 18.420 64.865 18.560 ;
        RECT 65.495 18.480 65.555 18.560 ;
        POLYGON 65.495 18.480 65.555 18.480 65.555 18.420 ;
        RECT 65.710 18.470 65.785 18.610 ;
        RECT 67.475 18.470 67.550 18.610 ;
        RECT 67.690 18.420 67.765 18.560 ;
        RECT 68.395 18.480 68.455 18.560 ;
        POLYGON 68.395 18.480 68.455 18.480 68.455 18.420 ;
        RECT 68.610 18.470 68.685 18.610 ;
        RECT 70.375 18.470 70.450 18.610 ;
        RECT 70.590 18.420 70.665 18.560 ;
        RECT 71.295 18.480 71.355 18.560 ;
        POLYGON 71.295 18.480 71.355 18.480 71.355 18.420 ;
        RECT 71.510 18.470 71.585 18.610 ;
        RECT 73.275 18.470 73.350 18.610 ;
        RECT 73.490 18.420 73.565 18.560 ;
        RECT 74.195 18.480 74.255 18.560 ;
        POLYGON 74.195 18.480 74.255 18.480 74.255 18.420 ;
        RECT 74.410 18.470 74.485 18.610 ;
        RECT 76.175 18.470 76.250 18.610 ;
        RECT 76.390 18.420 76.465 18.560 ;
        RECT 77.095 18.480 77.155 18.560 ;
        POLYGON 77.095 18.480 77.155 18.480 77.155 18.420 ;
        RECT 77.310 18.470 77.385 18.610 ;
        RECT 79.075 18.470 79.150 18.610 ;
        RECT 79.290 18.420 79.365 18.560 ;
        RECT 79.995 18.480 80.055 18.560 ;
        POLYGON 79.995 18.480 80.055 18.480 80.055 18.420 ;
        RECT 80.210 18.470 80.285 18.610 ;
        RECT 81.975 18.470 82.050 18.610 ;
        RECT 82.190 18.420 82.265 18.560 ;
        RECT 82.895 18.480 82.955 18.560 ;
        POLYGON 82.895 18.480 82.955 18.480 82.955 18.420 ;
        RECT 83.110 18.470 83.185 18.610 ;
        RECT 84.875 18.470 84.950 18.610 ;
        RECT 85.090 18.420 85.165 18.560 ;
        RECT 85.795 18.480 85.855 18.560 ;
        POLYGON 85.795 18.480 85.855 18.480 85.855 18.420 ;
        RECT 86.010 18.470 86.085 18.610 ;
        RECT 87.775 18.470 87.850 18.610 ;
        RECT 87.990 18.420 88.065 18.560 ;
        RECT 88.695 18.480 88.755 18.560 ;
        POLYGON 88.695 18.480 88.755 18.480 88.755 18.420 ;
        RECT 88.910 18.470 88.985 18.610 ;
        RECT 90.675 18.470 90.750 18.610 ;
        RECT 90.890 18.420 90.965 18.560 ;
        RECT 91.595 18.480 91.655 18.560 ;
        POLYGON 91.595 18.480 91.655 18.480 91.655 18.420 ;
        RECT 91.810 18.470 91.885 18.610 ;
        RECT 0.720 17.950 0.870 18.120 ;
        RECT 1.110 18.085 1.260 18.255 ;
        RECT 1.500 18.085 1.650 18.255 ;
        RECT 1.890 17.950 2.040 18.120 ;
        RECT 3.620 17.950 3.770 18.120 ;
        RECT 4.010 18.085 4.160 18.255 ;
        RECT 4.400 18.085 4.550 18.255 ;
        RECT 4.790 17.950 4.940 18.120 ;
        RECT 6.520 17.950 6.670 18.120 ;
        RECT 6.910 18.085 7.060 18.255 ;
        RECT 7.300 18.085 7.450 18.255 ;
        RECT 7.690 17.950 7.840 18.120 ;
        RECT 9.420 17.950 9.570 18.120 ;
        RECT 9.810 18.085 9.960 18.255 ;
        RECT 10.200 18.085 10.350 18.255 ;
        RECT 10.590 17.950 10.740 18.120 ;
        RECT 12.320 17.950 12.470 18.120 ;
        RECT 12.710 18.085 12.860 18.255 ;
        RECT 13.100 18.085 13.250 18.255 ;
        RECT 13.490 17.950 13.640 18.120 ;
        RECT 15.220 17.950 15.370 18.120 ;
        RECT 15.610 18.085 15.760 18.255 ;
        RECT 16.000 18.085 16.150 18.255 ;
        RECT 16.390 17.950 16.540 18.120 ;
        RECT 18.120 17.950 18.270 18.120 ;
        RECT 18.510 18.085 18.660 18.255 ;
        RECT 18.900 18.085 19.050 18.255 ;
        RECT 19.290 17.950 19.440 18.120 ;
        RECT 21.020 17.950 21.170 18.120 ;
        RECT 21.410 18.085 21.560 18.255 ;
        RECT 21.800 18.085 21.950 18.255 ;
        RECT 22.190 17.950 22.340 18.120 ;
        RECT 23.920 17.950 24.070 18.120 ;
        RECT 24.310 18.085 24.460 18.255 ;
        RECT 24.700 18.085 24.850 18.255 ;
        RECT 25.090 17.950 25.240 18.120 ;
        RECT 26.820 17.950 26.970 18.120 ;
        RECT 27.210 18.085 27.360 18.255 ;
        RECT 27.600 18.085 27.750 18.255 ;
        RECT 27.990 17.950 28.140 18.120 ;
        RECT 29.720 17.950 29.870 18.120 ;
        RECT 30.110 18.085 30.260 18.255 ;
        RECT 30.500 18.085 30.650 18.255 ;
        RECT 30.890 17.950 31.040 18.120 ;
        RECT 32.620 17.950 32.770 18.120 ;
        RECT 33.010 18.085 33.160 18.255 ;
        RECT 33.400 18.085 33.550 18.255 ;
        RECT 33.790 17.950 33.940 18.120 ;
        RECT 35.520 17.950 35.670 18.120 ;
        RECT 35.910 18.085 36.060 18.255 ;
        RECT 36.300 18.085 36.450 18.255 ;
        RECT 36.690 17.950 36.840 18.120 ;
        RECT 38.420 17.950 38.570 18.120 ;
        RECT 38.810 18.085 38.960 18.255 ;
        RECT 39.200 18.085 39.350 18.255 ;
        RECT 39.590 17.950 39.740 18.120 ;
        RECT 41.320 17.950 41.470 18.120 ;
        RECT 41.710 18.085 41.860 18.255 ;
        RECT 42.100 18.085 42.250 18.255 ;
        RECT 42.490 17.950 42.640 18.120 ;
        RECT 44.220 17.950 44.370 18.120 ;
        RECT 44.610 18.085 44.760 18.255 ;
        RECT 45.000 18.085 45.150 18.255 ;
        RECT 45.390 17.950 45.540 18.120 ;
        RECT 47.120 17.950 47.270 18.120 ;
        RECT 47.510 18.085 47.660 18.255 ;
        RECT 47.900 18.085 48.050 18.255 ;
        RECT 48.290 17.950 48.440 18.120 ;
        RECT 50.020 17.950 50.170 18.120 ;
        RECT 50.410 18.085 50.560 18.255 ;
        RECT 50.800 18.085 50.950 18.255 ;
        RECT 51.190 17.950 51.340 18.120 ;
        RECT 52.920 17.950 53.070 18.120 ;
        RECT 53.310 18.085 53.460 18.255 ;
        RECT 53.700 18.085 53.850 18.255 ;
        RECT 54.090 17.950 54.240 18.120 ;
        RECT 55.820 17.950 55.970 18.120 ;
        RECT 56.210 18.085 56.360 18.255 ;
        RECT 56.600 18.085 56.750 18.255 ;
        RECT 56.990 17.950 57.140 18.120 ;
        RECT 58.720 17.950 58.870 18.120 ;
        RECT 59.110 18.085 59.260 18.255 ;
        RECT 59.500 18.085 59.650 18.255 ;
        RECT 59.890 17.950 60.040 18.120 ;
        RECT 61.620 17.950 61.770 18.120 ;
        RECT 62.010 18.085 62.160 18.255 ;
        RECT 62.400 18.085 62.550 18.255 ;
        RECT 62.790 17.950 62.940 18.120 ;
        RECT 64.520 17.950 64.670 18.120 ;
        RECT 64.910 18.085 65.060 18.255 ;
        RECT 65.300 18.085 65.450 18.255 ;
        RECT 65.690 17.950 65.840 18.120 ;
        RECT 67.420 17.950 67.570 18.120 ;
        RECT 67.810 18.085 67.960 18.255 ;
        RECT 68.200 18.085 68.350 18.255 ;
        RECT 68.590 17.950 68.740 18.120 ;
        RECT 70.320 17.950 70.470 18.120 ;
        RECT 70.710 18.085 70.860 18.255 ;
        RECT 71.100 18.085 71.250 18.255 ;
        RECT 71.490 17.950 71.640 18.120 ;
        RECT 73.220 17.950 73.370 18.120 ;
        RECT 73.610 18.085 73.760 18.255 ;
        RECT 74.000 18.085 74.150 18.255 ;
        RECT 74.390 17.950 74.540 18.120 ;
        RECT 76.120 17.950 76.270 18.120 ;
        RECT 76.510 18.085 76.660 18.255 ;
        RECT 76.900 18.085 77.050 18.255 ;
        RECT 77.290 17.950 77.440 18.120 ;
        RECT 79.020 17.950 79.170 18.120 ;
        RECT 79.410 18.085 79.560 18.255 ;
        RECT 79.800 18.085 79.950 18.255 ;
        RECT 80.190 17.950 80.340 18.120 ;
        RECT 81.920 17.950 82.070 18.120 ;
        RECT 82.310 18.085 82.460 18.255 ;
        RECT 82.700 18.085 82.850 18.255 ;
        RECT 83.090 17.950 83.240 18.120 ;
        RECT 84.820 17.950 84.970 18.120 ;
        RECT 85.210 18.085 85.360 18.255 ;
        RECT 85.600 18.085 85.750 18.255 ;
        RECT 85.990 17.950 86.140 18.120 ;
        RECT 87.720 17.950 87.870 18.120 ;
        RECT 88.110 18.085 88.260 18.255 ;
        RECT 88.500 18.085 88.650 18.255 ;
        RECT 88.890 17.950 89.040 18.120 ;
        RECT 90.620 17.950 90.770 18.120 ;
        RECT 91.010 18.085 91.160 18.255 ;
        RECT 91.400 18.085 91.550 18.255 ;
        RECT 91.790 17.950 91.940 18.120 ;
        RECT 0.985 17.865 1.035 17.900 ;
        POLYGON 1.035 17.900 1.070 17.865 1.035 17.865 ;
        RECT 0.985 17.740 1.070 17.865 ;
        RECT 1.690 17.740 1.775 17.900 ;
        RECT 3.885 17.865 3.935 17.900 ;
        POLYGON 3.935 17.900 3.970 17.865 3.935 17.865 ;
        RECT 3.885 17.740 3.970 17.865 ;
        RECT 4.590 17.740 4.675 17.900 ;
        RECT 6.785 17.865 6.835 17.900 ;
        POLYGON 6.835 17.900 6.870 17.865 6.835 17.865 ;
        RECT 6.785 17.740 6.870 17.865 ;
        RECT 7.490 17.740 7.575 17.900 ;
        RECT 9.685 17.865 9.735 17.900 ;
        POLYGON 9.735 17.900 9.770 17.865 9.735 17.865 ;
        RECT 9.685 17.740 9.770 17.865 ;
        RECT 10.390 17.740 10.475 17.900 ;
        RECT 12.585 17.865 12.635 17.900 ;
        POLYGON 12.635 17.900 12.670 17.865 12.635 17.865 ;
        RECT 12.585 17.740 12.670 17.865 ;
        RECT 13.290 17.740 13.375 17.900 ;
        RECT 15.485 17.865 15.535 17.900 ;
        POLYGON 15.535 17.900 15.570 17.865 15.535 17.865 ;
        RECT 15.485 17.740 15.570 17.865 ;
        RECT 16.190 17.740 16.275 17.900 ;
        RECT 18.385 17.865 18.435 17.900 ;
        POLYGON 18.435 17.900 18.470 17.865 18.435 17.865 ;
        RECT 18.385 17.740 18.470 17.865 ;
        RECT 19.090 17.740 19.175 17.900 ;
        RECT 21.285 17.865 21.335 17.900 ;
        POLYGON 21.335 17.900 21.370 17.865 21.335 17.865 ;
        RECT 21.285 17.740 21.370 17.865 ;
        RECT 21.990 17.740 22.075 17.900 ;
        RECT 24.185 17.865 24.235 17.900 ;
        POLYGON 24.235 17.900 24.270 17.865 24.235 17.865 ;
        RECT 24.185 17.740 24.270 17.865 ;
        RECT 24.890 17.740 24.975 17.900 ;
        RECT 27.085 17.865 27.135 17.900 ;
        POLYGON 27.135 17.900 27.170 17.865 27.135 17.865 ;
        RECT 27.085 17.740 27.170 17.865 ;
        RECT 27.790 17.740 27.875 17.900 ;
        RECT 29.985 17.865 30.035 17.900 ;
        POLYGON 30.035 17.900 30.070 17.865 30.035 17.865 ;
        RECT 29.985 17.740 30.070 17.865 ;
        RECT 30.690 17.740 30.775 17.900 ;
        RECT 32.885 17.865 32.935 17.900 ;
        POLYGON 32.935 17.900 32.970 17.865 32.935 17.865 ;
        RECT 32.885 17.740 32.970 17.865 ;
        RECT 33.590 17.740 33.675 17.900 ;
        RECT 35.785 17.865 35.835 17.900 ;
        POLYGON 35.835 17.900 35.870 17.865 35.835 17.865 ;
        RECT 35.785 17.740 35.870 17.865 ;
        RECT 36.490 17.740 36.575 17.900 ;
        RECT 38.685 17.865 38.735 17.900 ;
        POLYGON 38.735 17.900 38.770 17.865 38.735 17.865 ;
        RECT 38.685 17.740 38.770 17.865 ;
        RECT 39.390 17.740 39.475 17.900 ;
        RECT 41.585 17.865 41.635 17.900 ;
        POLYGON 41.635 17.900 41.670 17.865 41.635 17.865 ;
        RECT 41.585 17.740 41.670 17.865 ;
        RECT 42.290 17.740 42.375 17.900 ;
        RECT 44.485 17.865 44.535 17.900 ;
        POLYGON 44.535 17.900 44.570 17.865 44.535 17.865 ;
        RECT 44.485 17.740 44.570 17.865 ;
        RECT 45.190 17.740 45.275 17.900 ;
        RECT 47.385 17.865 47.435 17.900 ;
        POLYGON 47.435 17.900 47.470 17.865 47.435 17.865 ;
        RECT 47.385 17.740 47.470 17.865 ;
        RECT 48.090 17.740 48.175 17.900 ;
        RECT 50.285 17.865 50.335 17.900 ;
        POLYGON 50.335 17.900 50.370 17.865 50.335 17.865 ;
        RECT 50.285 17.740 50.370 17.865 ;
        RECT 50.990 17.740 51.075 17.900 ;
        RECT 53.185 17.865 53.235 17.900 ;
        POLYGON 53.235 17.900 53.270 17.865 53.235 17.865 ;
        RECT 53.185 17.740 53.270 17.865 ;
        RECT 53.890 17.740 53.975 17.900 ;
        RECT 56.085 17.865 56.135 17.900 ;
        POLYGON 56.135 17.900 56.170 17.865 56.135 17.865 ;
        RECT 56.085 17.740 56.170 17.865 ;
        RECT 56.790 17.740 56.875 17.900 ;
        RECT 58.985 17.865 59.035 17.900 ;
        POLYGON 59.035 17.900 59.070 17.865 59.035 17.865 ;
        RECT 58.985 17.740 59.070 17.865 ;
        RECT 59.690 17.740 59.775 17.900 ;
        RECT 61.885 17.865 61.935 17.900 ;
        POLYGON 61.935 17.900 61.970 17.865 61.935 17.865 ;
        RECT 61.885 17.740 61.970 17.865 ;
        RECT 62.590 17.740 62.675 17.900 ;
        RECT 64.785 17.865 64.835 17.900 ;
        POLYGON 64.835 17.900 64.870 17.865 64.835 17.865 ;
        RECT 64.785 17.740 64.870 17.865 ;
        RECT 65.490 17.740 65.575 17.900 ;
        RECT 67.685 17.865 67.735 17.900 ;
        POLYGON 67.735 17.900 67.770 17.865 67.735 17.865 ;
        RECT 67.685 17.740 67.770 17.865 ;
        RECT 68.390 17.740 68.475 17.900 ;
        RECT 70.585 17.865 70.635 17.900 ;
        POLYGON 70.635 17.900 70.670 17.865 70.635 17.865 ;
        RECT 70.585 17.740 70.670 17.865 ;
        RECT 71.290 17.740 71.375 17.900 ;
        RECT 73.485 17.865 73.535 17.900 ;
        POLYGON 73.535 17.900 73.570 17.865 73.535 17.865 ;
        RECT 73.485 17.740 73.570 17.865 ;
        RECT 74.190 17.740 74.275 17.900 ;
        RECT 76.385 17.865 76.435 17.900 ;
        POLYGON 76.435 17.900 76.470 17.865 76.435 17.865 ;
        RECT 76.385 17.740 76.470 17.865 ;
        RECT 77.090 17.740 77.175 17.900 ;
        RECT 79.285 17.865 79.335 17.900 ;
        POLYGON 79.335 17.900 79.370 17.865 79.335 17.865 ;
        RECT 79.285 17.740 79.370 17.865 ;
        RECT 79.990 17.740 80.075 17.900 ;
        RECT 82.185 17.865 82.235 17.900 ;
        POLYGON 82.235 17.900 82.270 17.865 82.235 17.865 ;
        RECT 82.185 17.740 82.270 17.865 ;
        RECT 82.890 17.740 82.975 17.900 ;
        RECT 85.085 17.865 85.135 17.900 ;
        POLYGON 85.135 17.900 85.170 17.865 85.135 17.865 ;
        RECT 85.085 17.740 85.170 17.865 ;
        RECT 85.790 17.740 85.875 17.900 ;
        RECT 87.985 17.865 88.035 17.900 ;
        POLYGON 88.035 17.900 88.070 17.865 88.035 17.865 ;
        RECT 87.985 17.740 88.070 17.865 ;
        RECT 88.690 17.740 88.775 17.900 ;
        RECT 90.885 17.865 90.935 17.900 ;
        POLYGON 90.935 17.900 90.970 17.865 90.935 17.865 ;
        RECT 90.885 17.740 90.970 17.865 ;
        RECT 91.590 17.740 91.675 17.900 ;
        RECT 0.775 17.120 0.850 17.260 ;
        RECT 0.990 17.070 1.065 17.210 ;
        RECT 1.695 17.130 1.755 17.210 ;
        POLYGON 1.695 17.130 1.755 17.130 1.755 17.070 ;
        RECT 1.910 17.120 1.985 17.260 ;
        RECT 3.675 17.120 3.750 17.260 ;
        RECT 3.890 17.070 3.965 17.210 ;
        RECT 4.595 17.130 4.655 17.210 ;
        POLYGON 4.595 17.130 4.655 17.130 4.655 17.070 ;
        RECT 4.810 17.120 4.885 17.260 ;
        RECT 6.575 17.120 6.650 17.260 ;
        RECT 6.790 17.070 6.865 17.210 ;
        RECT 7.495 17.130 7.555 17.210 ;
        POLYGON 7.495 17.130 7.555 17.130 7.555 17.070 ;
        RECT 7.710 17.120 7.785 17.260 ;
        RECT 9.475 17.120 9.550 17.260 ;
        RECT 9.690 17.070 9.765 17.210 ;
        RECT 10.395 17.130 10.455 17.210 ;
        POLYGON 10.395 17.130 10.455 17.130 10.455 17.070 ;
        RECT 10.610 17.120 10.685 17.260 ;
        RECT 12.375 17.120 12.450 17.260 ;
        RECT 12.590 17.070 12.665 17.210 ;
        RECT 13.295 17.130 13.355 17.210 ;
        POLYGON 13.295 17.130 13.355 17.130 13.355 17.070 ;
        RECT 13.510 17.120 13.585 17.260 ;
        RECT 15.275 17.120 15.350 17.260 ;
        RECT 15.490 17.070 15.565 17.210 ;
        RECT 16.195 17.130 16.255 17.210 ;
        POLYGON 16.195 17.130 16.255 17.130 16.255 17.070 ;
        RECT 16.410 17.120 16.485 17.260 ;
        RECT 18.175 17.120 18.250 17.260 ;
        RECT 18.390 17.070 18.465 17.210 ;
        RECT 19.095 17.130 19.155 17.210 ;
        POLYGON 19.095 17.130 19.155 17.130 19.155 17.070 ;
        RECT 19.310 17.120 19.385 17.260 ;
        RECT 21.075 17.120 21.150 17.260 ;
        RECT 21.290 17.070 21.365 17.210 ;
        RECT 21.995 17.130 22.055 17.210 ;
        POLYGON 21.995 17.130 22.055 17.130 22.055 17.070 ;
        RECT 22.210 17.120 22.285 17.260 ;
        RECT 23.975 17.120 24.050 17.260 ;
        RECT 24.190 17.070 24.265 17.210 ;
        RECT 24.895 17.130 24.955 17.210 ;
        POLYGON 24.895 17.130 24.955 17.130 24.955 17.070 ;
        RECT 25.110 17.120 25.185 17.260 ;
        RECT 26.875 17.120 26.950 17.260 ;
        RECT 27.090 17.070 27.165 17.210 ;
        RECT 27.795 17.130 27.855 17.210 ;
        POLYGON 27.795 17.130 27.855 17.130 27.855 17.070 ;
        RECT 28.010 17.120 28.085 17.260 ;
        RECT 29.775 17.120 29.850 17.260 ;
        RECT 29.990 17.070 30.065 17.210 ;
        RECT 30.695 17.130 30.755 17.210 ;
        POLYGON 30.695 17.130 30.755 17.130 30.755 17.070 ;
        RECT 30.910 17.120 30.985 17.260 ;
        RECT 32.675 17.120 32.750 17.260 ;
        RECT 32.890 17.070 32.965 17.210 ;
        RECT 33.595 17.130 33.655 17.210 ;
        POLYGON 33.595 17.130 33.655 17.130 33.655 17.070 ;
        RECT 33.810 17.120 33.885 17.260 ;
        RECT 35.575 17.120 35.650 17.260 ;
        RECT 35.790 17.070 35.865 17.210 ;
        RECT 36.495 17.130 36.555 17.210 ;
        POLYGON 36.495 17.130 36.555 17.130 36.555 17.070 ;
        RECT 36.710 17.120 36.785 17.260 ;
        RECT 38.475 17.120 38.550 17.260 ;
        RECT 38.690 17.070 38.765 17.210 ;
        RECT 39.395 17.130 39.455 17.210 ;
        POLYGON 39.395 17.130 39.455 17.130 39.455 17.070 ;
        RECT 39.610 17.120 39.685 17.260 ;
        RECT 41.375 17.120 41.450 17.260 ;
        RECT 41.590 17.070 41.665 17.210 ;
        RECT 42.295 17.130 42.355 17.210 ;
        POLYGON 42.295 17.130 42.355 17.130 42.355 17.070 ;
        RECT 42.510 17.120 42.585 17.260 ;
        RECT 44.275 17.120 44.350 17.260 ;
        RECT 44.490 17.070 44.565 17.210 ;
        RECT 45.195 17.130 45.255 17.210 ;
        POLYGON 45.195 17.130 45.255 17.130 45.255 17.070 ;
        RECT 45.410 17.120 45.485 17.260 ;
        RECT 47.175 17.120 47.250 17.260 ;
        RECT 47.390 17.070 47.465 17.210 ;
        RECT 48.095 17.130 48.155 17.210 ;
        POLYGON 48.095 17.130 48.155 17.130 48.155 17.070 ;
        RECT 48.310 17.120 48.385 17.260 ;
        RECT 50.075 17.120 50.150 17.260 ;
        RECT 50.290 17.070 50.365 17.210 ;
        RECT 50.995 17.130 51.055 17.210 ;
        POLYGON 50.995 17.130 51.055 17.130 51.055 17.070 ;
        RECT 51.210 17.120 51.285 17.260 ;
        RECT 52.975 17.120 53.050 17.260 ;
        RECT 53.190 17.070 53.265 17.210 ;
        RECT 53.895 17.130 53.955 17.210 ;
        POLYGON 53.895 17.130 53.955 17.130 53.955 17.070 ;
        RECT 54.110 17.120 54.185 17.260 ;
        RECT 55.875 17.120 55.950 17.260 ;
        RECT 56.090 17.070 56.165 17.210 ;
        RECT 56.795 17.130 56.855 17.210 ;
        POLYGON 56.795 17.130 56.855 17.130 56.855 17.070 ;
        RECT 57.010 17.120 57.085 17.260 ;
        RECT 58.775 17.120 58.850 17.260 ;
        RECT 58.990 17.070 59.065 17.210 ;
        RECT 59.695 17.130 59.755 17.210 ;
        POLYGON 59.695 17.130 59.755 17.130 59.755 17.070 ;
        RECT 59.910 17.120 59.985 17.260 ;
        RECT 61.675 17.120 61.750 17.260 ;
        RECT 61.890 17.070 61.965 17.210 ;
        RECT 62.595 17.130 62.655 17.210 ;
        POLYGON 62.595 17.130 62.655 17.130 62.655 17.070 ;
        RECT 62.810 17.120 62.885 17.260 ;
        RECT 64.575 17.120 64.650 17.260 ;
        RECT 64.790 17.070 64.865 17.210 ;
        RECT 65.495 17.130 65.555 17.210 ;
        POLYGON 65.495 17.130 65.555 17.130 65.555 17.070 ;
        RECT 65.710 17.120 65.785 17.260 ;
        RECT 67.475 17.120 67.550 17.260 ;
        RECT 67.690 17.070 67.765 17.210 ;
        RECT 68.395 17.130 68.455 17.210 ;
        POLYGON 68.395 17.130 68.455 17.130 68.455 17.070 ;
        RECT 68.610 17.120 68.685 17.260 ;
        RECT 70.375 17.120 70.450 17.260 ;
        RECT 70.590 17.070 70.665 17.210 ;
        RECT 71.295 17.130 71.355 17.210 ;
        POLYGON 71.295 17.130 71.355 17.130 71.355 17.070 ;
        RECT 71.510 17.120 71.585 17.260 ;
        RECT 73.275 17.120 73.350 17.260 ;
        RECT 73.490 17.070 73.565 17.210 ;
        RECT 74.195 17.130 74.255 17.210 ;
        POLYGON 74.195 17.130 74.255 17.130 74.255 17.070 ;
        RECT 74.410 17.120 74.485 17.260 ;
        RECT 76.175 17.120 76.250 17.260 ;
        RECT 76.390 17.070 76.465 17.210 ;
        RECT 77.095 17.130 77.155 17.210 ;
        POLYGON 77.095 17.130 77.155 17.130 77.155 17.070 ;
        RECT 77.310 17.120 77.385 17.260 ;
        RECT 79.075 17.120 79.150 17.260 ;
        RECT 79.290 17.070 79.365 17.210 ;
        RECT 79.995 17.130 80.055 17.210 ;
        POLYGON 79.995 17.130 80.055 17.130 80.055 17.070 ;
        RECT 80.210 17.120 80.285 17.260 ;
        RECT 81.975 17.120 82.050 17.260 ;
        RECT 82.190 17.070 82.265 17.210 ;
        RECT 82.895 17.130 82.955 17.210 ;
        POLYGON 82.895 17.130 82.955 17.130 82.955 17.070 ;
        RECT 83.110 17.120 83.185 17.260 ;
        RECT 84.875 17.120 84.950 17.260 ;
        RECT 85.090 17.070 85.165 17.210 ;
        RECT 85.795 17.130 85.855 17.210 ;
        POLYGON 85.795 17.130 85.855 17.130 85.855 17.070 ;
        RECT 86.010 17.120 86.085 17.260 ;
        RECT 87.775 17.120 87.850 17.260 ;
        RECT 87.990 17.070 88.065 17.210 ;
        RECT 88.695 17.130 88.755 17.210 ;
        POLYGON 88.695 17.130 88.755 17.130 88.755 17.070 ;
        RECT 88.910 17.120 88.985 17.260 ;
        RECT 90.675 17.120 90.750 17.260 ;
        RECT 90.890 17.070 90.965 17.210 ;
        RECT 91.595 17.130 91.655 17.210 ;
        POLYGON 91.595 17.130 91.655 17.130 91.655 17.070 ;
        RECT 91.810 17.120 91.885 17.260 ;
        RECT 0.720 16.600 0.870 16.770 ;
        RECT 1.110 16.735 1.260 16.905 ;
        RECT 1.500 16.735 1.650 16.905 ;
        RECT 1.890 16.600 2.040 16.770 ;
        RECT 3.620 16.600 3.770 16.770 ;
        RECT 4.010 16.735 4.160 16.905 ;
        RECT 4.400 16.735 4.550 16.905 ;
        RECT 4.790 16.600 4.940 16.770 ;
        RECT 6.520 16.600 6.670 16.770 ;
        RECT 6.910 16.735 7.060 16.905 ;
        RECT 7.300 16.735 7.450 16.905 ;
        RECT 7.690 16.600 7.840 16.770 ;
        RECT 9.420 16.600 9.570 16.770 ;
        RECT 9.810 16.735 9.960 16.905 ;
        RECT 10.200 16.735 10.350 16.905 ;
        RECT 10.590 16.600 10.740 16.770 ;
        RECT 12.320 16.600 12.470 16.770 ;
        RECT 12.710 16.735 12.860 16.905 ;
        RECT 13.100 16.735 13.250 16.905 ;
        RECT 13.490 16.600 13.640 16.770 ;
        RECT 15.220 16.600 15.370 16.770 ;
        RECT 15.610 16.735 15.760 16.905 ;
        RECT 16.000 16.735 16.150 16.905 ;
        RECT 16.390 16.600 16.540 16.770 ;
        RECT 18.120 16.600 18.270 16.770 ;
        RECT 18.510 16.735 18.660 16.905 ;
        RECT 18.900 16.735 19.050 16.905 ;
        RECT 19.290 16.600 19.440 16.770 ;
        RECT 21.020 16.600 21.170 16.770 ;
        RECT 21.410 16.735 21.560 16.905 ;
        RECT 21.800 16.735 21.950 16.905 ;
        RECT 22.190 16.600 22.340 16.770 ;
        RECT 23.920 16.600 24.070 16.770 ;
        RECT 24.310 16.735 24.460 16.905 ;
        RECT 24.700 16.735 24.850 16.905 ;
        RECT 25.090 16.600 25.240 16.770 ;
        RECT 26.820 16.600 26.970 16.770 ;
        RECT 27.210 16.735 27.360 16.905 ;
        RECT 27.600 16.735 27.750 16.905 ;
        RECT 27.990 16.600 28.140 16.770 ;
        RECT 29.720 16.600 29.870 16.770 ;
        RECT 30.110 16.735 30.260 16.905 ;
        RECT 30.500 16.735 30.650 16.905 ;
        RECT 30.890 16.600 31.040 16.770 ;
        RECT 32.620 16.600 32.770 16.770 ;
        RECT 33.010 16.735 33.160 16.905 ;
        RECT 33.400 16.735 33.550 16.905 ;
        RECT 33.790 16.600 33.940 16.770 ;
        RECT 35.520 16.600 35.670 16.770 ;
        RECT 35.910 16.735 36.060 16.905 ;
        RECT 36.300 16.735 36.450 16.905 ;
        RECT 36.690 16.600 36.840 16.770 ;
        RECT 38.420 16.600 38.570 16.770 ;
        RECT 38.810 16.735 38.960 16.905 ;
        RECT 39.200 16.735 39.350 16.905 ;
        RECT 39.590 16.600 39.740 16.770 ;
        RECT 41.320 16.600 41.470 16.770 ;
        RECT 41.710 16.735 41.860 16.905 ;
        RECT 42.100 16.735 42.250 16.905 ;
        RECT 42.490 16.600 42.640 16.770 ;
        RECT 44.220 16.600 44.370 16.770 ;
        RECT 44.610 16.735 44.760 16.905 ;
        RECT 45.000 16.735 45.150 16.905 ;
        RECT 45.390 16.600 45.540 16.770 ;
        RECT 47.120 16.600 47.270 16.770 ;
        RECT 47.510 16.735 47.660 16.905 ;
        RECT 47.900 16.735 48.050 16.905 ;
        RECT 48.290 16.600 48.440 16.770 ;
        RECT 50.020 16.600 50.170 16.770 ;
        RECT 50.410 16.735 50.560 16.905 ;
        RECT 50.800 16.735 50.950 16.905 ;
        RECT 51.190 16.600 51.340 16.770 ;
        RECT 52.920 16.600 53.070 16.770 ;
        RECT 53.310 16.735 53.460 16.905 ;
        RECT 53.700 16.735 53.850 16.905 ;
        RECT 54.090 16.600 54.240 16.770 ;
        RECT 55.820 16.600 55.970 16.770 ;
        RECT 56.210 16.735 56.360 16.905 ;
        RECT 56.600 16.735 56.750 16.905 ;
        RECT 56.990 16.600 57.140 16.770 ;
        RECT 58.720 16.600 58.870 16.770 ;
        RECT 59.110 16.735 59.260 16.905 ;
        RECT 59.500 16.735 59.650 16.905 ;
        RECT 59.890 16.600 60.040 16.770 ;
        RECT 61.620 16.600 61.770 16.770 ;
        RECT 62.010 16.735 62.160 16.905 ;
        RECT 62.400 16.735 62.550 16.905 ;
        RECT 62.790 16.600 62.940 16.770 ;
        RECT 64.520 16.600 64.670 16.770 ;
        RECT 64.910 16.735 65.060 16.905 ;
        RECT 65.300 16.735 65.450 16.905 ;
        RECT 65.690 16.600 65.840 16.770 ;
        RECT 67.420 16.600 67.570 16.770 ;
        RECT 67.810 16.735 67.960 16.905 ;
        RECT 68.200 16.735 68.350 16.905 ;
        RECT 68.590 16.600 68.740 16.770 ;
        RECT 70.320 16.600 70.470 16.770 ;
        RECT 70.710 16.735 70.860 16.905 ;
        RECT 71.100 16.735 71.250 16.905 ;
        RECT 71.490 16.600 71.640 16.770 ;
        RECT 73.220 16.600 73.370 16.770 ;
        RECT 73.610 16.735 73.760 16.905 ;
        RECT 74.000 16.735 74.150 16.905 ;
        RECT 74.390 16.600 74.540 16.770 ;
        RECT 76.120 16.600 76.270 16.770 ;
        RECT 76.510 16.735 76.660 16.905 ;
        RECT 76.900 16.735 77.050 16.905 ;
        RECT 77.290 16.600 77.440 16.770 ;
        RECT 79.020 16.600 79.170 16.770 ;
        RECT 79.410 16.735 79.560 16.905 ;
        RECT 79.800 16.735 79.950 16.905 ;
        RECT 80.190 16.600 80.340 16.770 ;
        RECT 81.920 16.600 82.070 16.770 ;
        RECT 82.310 16.735 82.460 16.905 ;
        RECT 82.700 16.735 82.850 16.905 ;
        RECT 83.090 16.600 83.240 16.770 ;
        RECT 84.820 16.600 84.970 16.770 ;
        RECT 85.210 16.735 85.360 16.905 ;
        RECT 85.600 16.735 85.750 16.905 ;
        RECT 85.990 16.600 86.140 16.770 ;
        RECT 87.720 16.600 87.870 16.770 ;
        RECT 88.110 16.735 88.260 16.905 ;
        RECT 88.500 16.735 88.650 16.905 ;
        RECT 88.890 16.600 89.040 16.770 ;
        RECT 90.620 16.600 90.770 16.770 ;
        RECT 91.010 16.735 91.160 16.905 ;
        RECT 91.400 16.735 91.550 16.905 ;
        RECT 91.790 16.600 91.940 16.770 ;
        RECT 0.985 16.515 1.035 16.550 ;
        POLYGON 1.035 16.550 1.070 16.515 1.035 16.515 ;
        RECT 0.985 16.390 1.070 16.515 ;
        RECT 1.690 16.390 1.775 16.550 ;
        RECT 3.885 16.515 3.935 16.550 ;
        POLYGON 3.935 16.550 3.970 16.515 3.935 16.515 ;
        RECT 3.885 16.390 3.970 16.515 ;
        RECT 4.590 16.390 4.675 16.550 ;
        RECT 6.785 16.515 6.835 16.550 ;
        POLYGON 6.835 16.550 6.870 16.515 6.835 16.515 ;
        RECT 6.785 16.390 6.870 16.515 ;
        RECT 7.490 16.390 7.575 16.550 ;
        RECT 9.685 16.515 9.735 16.550 ;
        POLYGON 9.735 16.550 9.770 16.515 9.735 16.515 ;
        RECT 9.685 16.390 9.770 16.515 ;
        RECT 10.390 16.390 10.475 16.550 ;
        RECT 12.585 16.515 12.635 16.550 ;
        POLYGON 12.635 16.550 12.670 16.515 12.635 16.515 ;
        RECT 12.585 16.390 12.670 16.515 ;
        RECT 13.290 16.390 13.375 16.550 ;
        RECT 15.485 16.515 15.535 16.550 ;
        POLYGON 15.535 16.550 15.570 16.515 15.535 16.515 ;
        RECT 15.485 16.390 15.570 16.515 ;
        RECT 16.190 16.390 16.275 16.550 ;
        RECT 18.385 16.515 18.435 16.550 ;
        POLYGON 18.435 16.550 18.470 16.515 18.435 16.515 ;
        RECT 18.385 16.390 18.470 16.515 ;
        RECT 19.090 16.390 19.175 16.550 ;
        RECT 21.285 16.515 21.335 16.550 ;
        POLYGON 21.335 16.550 21.370 16.515 21.335 16.515 ;
        RECT 21.285 16.390 21.370 16.515 ;
        RECT 21.990 16.390 22.075 16.550 ;
        RECT 24.185 16.515 24.235 16.550 ;
        POLYGON 24.235 16.550 24.270 16.515 24.235 16.515 ;
        RECT 24.185 16.390 24.270 16.515 ;
        RECT 24.890 16.390 24.975 16.550 ;
        RECT 27.085 16.515 27.135 16.550 ;
        POLYGON 27.135 16.550 27.170 16.515 27.135 16.515 ;
        RECT 27.085 16.390 27.170 16.515 ;
        RECT 27.790 16.390 27.875 16.550 ;
        RECT 29.985 16.515 30.035 16.550 ;
        POLYGON 30.035 16.550 30.070 16.515 30.035 16.515 ;
        RECT 29.985 16.390 30.070 16.515 ;
        RECT 30.690 16.390 30.775 16.550 ;
        RECT 32.885 16.515 32.935 16.550 ;
        POLYGON 32.935 16.550 32.970 16.515 32.935 16.515 ;
        RECT 32.885 16.390 32.970 16.515 ;
        RECT 33.590 16.390 33.675 16.550 ;
        RECT 35.785 16.515 35.835 16.550 ;
        POLYGON 35.835 16.550 35.870 16.515 35.835 16.515 ;
        RECT 35.785 16.390 35.870 16.515 ;
        RECT 36.490 16.390 36.575 16.550 ;
        RECT 38.685 16.515 38.735 16.550 ;
        POLYGON 38.735 16.550 38.770 16.515 38.735 16.515 ;
        RECT 38.685 16.390 38.770 16.515 ;
        RECT 39.390 16.390 39.475 16.550 ;
        RECT 41.585 16.515 41.635 16.550 ;
        POLYGON 41.635 16.550 41.670 16.515 41.635 16.515 ;
        RECT 41.585 16.390 41.670 16.515 ;
        RECT 42.290 16.390 42.375 16.550 ;
        RECT 44.485 16.515 44.535 16.550 ;
        POLYGON 44.535 16.550 44.570 16.515 44.535 16.515 ;
        RECT 44.485 16.390 44.570 16.515 ;
        RECT 45.190 16.390 45.275 16.550 ;
        RECT 47.385 16.515 47.435 16.550 ;
        POLYGON 47.435 16.550 47.470 16.515 47.435 16.515 ;
        RECT 47.385 16.390 47.470 16.515 ;
        RECT 48.090 16.390 48.175 16.550 ;
        RECT 50.285 16.515 50.335 16.550 ;
        POLYGON 50.335 16.550 50.370 16.515 50.335 16.515 ;
        RECT 50.285 16.390 50.370 16.515 ;
        RECT 50.990 16.390 51.075 16.550 ;
        RECT 53.185 16.515 53.235 16.550 ;
        POLYGON 53.235 16.550 53.270 16.515 53.235 16.515 ;
        RECT 53.185 16.390 53.270 16.515 ;
        RECT 53.890 16.390 53.975 16.550 ;
        RECT 56.085 16.515 56.135 16.550 ;
        POLYGON 56.135 16.550 56.170 16.515 56.135 16.515 ;
        RECT 56.085 16.390 56.170 16.515 ;
        RECT 56.790 16.390 56.875 16.550 ;
        RECT 58.985 16.515 59.035 16.550 ;
        POLYGON 59.035 16.550 59.070 16.515 59.035 16.515 ;
        RECT 58.985 16.390 59.070 16.515 ;
        RECT 59.690 16.390 59.775 16.550 ;
        RECT 61.885 16.515 61.935 16.550 ;
        POLYGON 61.935 16.550 61.970 16.515 61.935 16.515 ;
        RECT 61.885 16.390 61.970 16.515 ;
        RECT 62.590 16.390 62.675 16.550 ;
        RECT 64.785 16.515 64.835 16.550 ;
        POLYGON 64.835 16.550 64.870 16.515 64.835 16.515 ;
        RECT 64.785 16.390 64.870 16.515 ;
        RECT 65.490 16.390 65.575 16.550 ;
        RECT 67.685 16.515 67.735 16.550 ;
        POLYGON 67.735 16.550 67.770 16.515 67.735 16.515 ;
        RECT 67.685 16.390 67.770 16.515 ;
        RECT 68.390 16.390 68.475 16.550 ;
        RECT 70.585 16.515 70.635 16.550 ;
        POLYGON 70.635 16.550 70.670 16.515 70.635 16.515 ;
        RECT 70.585 16.390 70.670 16.515 ;
        RECT 71.290 16.390 71.375 16.550 ;
        RECT 73.485 16.515 73.535 16.550 ;
        POLYGON 73.535 16.550 73.570 16.515 73.535 16.515 ;
        RECT 73.485 16.390 73.570 16.515 ;
        RECT 74.190 16.390 74.275 16.550 ;
        RECT 76.385 16.515 76.435 16.550 ;
        POLYGON 76.435 16.550 76.470 16.515 76.435 16.515 ;
        RECT 76.385 16.390 76.470 16.515 ;
        RECT 77.090 16.390 77.175 16.550 ;
        RECT 79.285 16.515 79.335 16.550 ;
        POLYGON 79.335 16.550 79.370 16.515 79.335 16.515 ;
        RECT 79.285 16.390 79.370 16.515 ;
        RECT 79.990 16.390 80.075 16.550 ;
        RECT 82.185 16.515 82.235 16.550 ;
        POLYGON 82.235 16.550 82.270 16.515 82.235 16.515 ;
        RECT 82.185 16.390 82.270 16.515 ;
        RECT 82.890 16.390 82.975 16.550 ;
        RECT 85.085 16.515 85.135 16.550 ;
        POLYGON 85.135 16.550 85.170 16.515 85.135 16.515 ;
        RECT 85.085 16.390 85.170 16.515 ;
        RECT 85.790 16.390 85.875 16.550 ;
        RECT 87.985 16.515 88.035 16.550 ;
        POLYGON 88.035 16.550 88.070 16.515 88.035 16.515 ;
        RECT 87.985 16.390 88.070 16.515 ;
        RECT 88.690 16.390 88.775 16.550 ;
        RECT 90.885 16.515 90.935 16.550 ;
        POLYGON 90.935 16.550 90.970 16.515 90.935 16.515 ;
        RECT 90.885 16.390 90.970 16.515 ;
        RECT 91.590 16.390 91.675 16.550 ;
        RECT 0.775 15.770 0.850 15.910 ;
        RECT 0.990 15.720 1.065 15.860 ;
        RECT 1.695 15.780 1.755 15.860 ;
        POLYGON 1.695 15.780 1.755 15.780 1.755 15.720 ;
        RECT 1.910 15.770 1.985 15.910 ;
        RECT 3.675 15.770 3.750 15.910 ;
        RECT 3.890 15.720 3.965 15.860 ;
        RECT 4.595 15.780 4.655 15.860 ;
        POLYGON 4.595 15.780 4.655 15.780 4.655 15.720 ;
        RECT 4.810 15.770 4.885 15.910 ;
        RECT 6.575 15.770 6.650 15.910 ;
        RECT 6.790 15.720 6.865 15.860 ;
        RECT 7.495 15.780 7.555 15.860 ;
        POLYGON 7.495 15.780 7.555 15.780 7.555 15.720 ;
        RECT 7.710 15.770 7.785 15.910 ;
        RECT 9.475 15.770 9.550 15.910 ;
        RECT 9.690 15.720 9.765 15.860 ;
        RECT 10.395 15.780 10.455 15.860 ;
        POLYGON 10.395 15.780 10.455 15.780 10.455 15.720 ;
        RECT 10.610 15.770 10.685 15.910 ;
        RECT 12.375 15.770 12.450 15.910 ;
        RECT 12.590 15.720 12.665 15.860 ;
        RECT 13.295 15.780 13.355 15.860 ;
        POLYGON 13.295 15.780 13.355 15.780 13.355 15.720 ;
        RECT 13.510 15.770 13.585 15.910 ;
        RECT 15.275 15.770 15.350 15.910 ;
        RECT 15.490 15.720 15.565 15.860 ;
        RECT 16.195 15.780 16.255 15.860 ;
        POLYGON 16.195 15.780 16.255 15.780 16.255 15.720 ;
        RECT 16.410 15.770 16.485 15.910 ;
        RECT 18.175 15.770 18.250 15.910 ;
        RECT 18.390 15.720 18.465 15.860 ;
        RECT 19.095 15.780 19.155 15.860 ;
        POLYGON 19.095 15.780 19.155 15.780 19.155 15.720 ;
        RECT 19.310 15.770 19.385 15.910 ;
        RECT 21.075 15.770 21.150 15.910 ;
        RECT 21.290 15.720 21.365 15.860 ;
        RECT 21.995 15.780 22.055 15.860 ;
        POLYGON 21.995 15.780 22.055 15.780 22.055 15.720 ;
        RECT 22.210 15.770 22.285 15.910 ;
        RECT 23.975 15.770 24.050 15.910 ;
        RECT 24.190 15.720 24.265 15.860 ;
        RECT 24.895 15.780 24.955 15.860 ;
        POLYGON 24.895 15.780 24.955 15.780 24.955 15.720 ;
        RECT 25.110 15.770 25.185 15.910 ;
        RECT 26.875 15.770 26.950 15.910 ;
        RECT 27.090 15.720 27.165 15.860 ;
        RECT 27.795 15.780 27.855 15.860 ;
        POLYGON 27.795 15.780 27.855 15.780 27.855 15.720 ;
        RECT 28.010 15.770 28.085 15.910 ;
        RECT 29.775 15.770 29.850 15.910 ;
        RECT 29.990 15.720 30.065 15.860 ;
        RECT 30.695 15.780 30.755 15.860 ;
        POLYGON 30.695 15.780 30.755 15.780 30.755 15.720 ;
        RECT 30.910 15.770 30.985 15.910 ;
        RECT 32.675 15.770 32.750 15.910 ;
        RECT 32.890 15.720 32.965 15.860 ;
        RECT 33.595 15.780 33.655 15.860 ;
        POLYGON 33.595 15.780 33.655 15.780 33.655 15.720 ;
        RECT 33.810 15.770 33.885 15.910 ;
        RECT 35.575 15.770 35.650 15.910 ;
        RECT 35.790 15.720 35.865 15.860 ;
        RECT 36.495 15.780 36.555 15.860 ;
        POLYGON 36.495 15.780 36.555 15.780 36.555 15.720 ;
        RECT 36.710 15.770 36.785 15.910 ;
        RECT 38.475 15.770 38.550 15.910 ;
        RECT 38.690 15.720 38.765 15.860 ;
        RECT 39.395 15.780 39.455 15.860 ;
        POLYGON 39.395 15.780 39.455 15.780 39.455 15.720 ;
        RECT 39.610 15.770 39.685 15.910 ;
        RECT 41.375 15.770 41.450 15.910 ;
        RECT 41.590 15.720 41.665 15.860 ;
        RECT 42.295 15.780 42.355 15.860 ;
        POLYGON 42.295 15.780 42.355 15.780 42.355 15.720 ;
        RECT 42.510 15.770 42.585 15.910 ;
        RECT 44.275 15.770 44.350 15.910 ;
        RECT 44.490 15.720 44.565 15.860 ;
        RECT 45.195 15.780 45.255 15.860 ;
        POLYGON 45.195 15.780 45.255 15.780 45.255 15.720 ;
        RECT 45.410 15.770 45.485 15.910 ;
        RECT 47.175 15.770 47.250 15.910 ;
        RECT 47.390 15.720 47.465 15.860 ;
        RECT 48.095 15.780 48.155 15.860 ;
        POLYGON 48.095 15.780 48.155 15.780 48.155 15.720 ;
        RECT 48.310 15.770 48.385 15.910 ;
        RECT 50.075 15.770 50.150 15.910 ;
        RECT 50.290 15.720 50.365 15.860 ;
        RECT 50.995 15.780 51.055 15.860 ;
        POLYGON 50.995 15.780 51.055 15.780 51.055 15.720 ;
        RECT 51.210 15.770 51.285 15.910 ;
        RECT 52.975 15.770 53.050 15.910 ;
        RECT 53.190 15.720 53.265 15.860 ;
        RECT 53.895 15.780 53.955 15.860 ;
        POLYGON 53.895 15.780 53.955 15.780 53.955 15.720 ;
        RECT 54.110 15.770 54.185 15.910 ;
        RECT 55.875 15.770 55.950 15.910 ;
        RECT 56.090 15.720 56.165 15.860 ;
        RECT 56.795 15.780 56.855 15.860 ;
        POLYGON 56.795 15.780 56.855 15.780 56.855 15.720 ;
        RECT 57.010 15.770 57.085 15.910 ;
        RECT 58.775 15.770 58.850 15.910 ;
        RECT 58.990 15.720 59.065 15.860 ;
        RECT 59.695 15.780 59.755 15.860 ;
        POLYGON 59.695 15.780 59.755 15.780 59.755 15.720 ;
        RECT 59.910 15.770 59.985 15.910 ;
        RECT 61.675 15.770 61.750 15.910 ;
        RECT 61.890 15.720 61.965 15.860 ;
        RECT 62.595 15.780 62.655 15.860 ;
        POLYGON 62.595 15.780 62.655 15.780 62.655 15.720 ;
        RECT 62.810 15.770 62.885 15.910 ;
        RECT 64.575 15.770 64.650 15.910 ;
        RECT 64.790 15.720 64.865 15.860 ;
        RECT 65.495 15.780 65.555 15.860 ;
        POLYGON 65.495 15.780 65.555 15.780 65.555 15.720 ;
        RECT 65.710 15.770 65.785 15.910 ;
        RECT 67.475 15.770 67.550 15.910 ;
        RECT 67.690 15.720 67.765 15.860 ;
        RECT 68.395 15.780 68.455 15.860 ;
        POLYGON 68.395 15.780 68.455 15.780 68.455 15.720 ;
        RECT 68.610 15.770 68.685 15.910 ;
        RECT 70.375 15.770 70.450 15.910 ;
        RECT 70.590 15.720 70.665 15.860 ;
        RECT 71.295 15.780 71.355 15.860 ;
        POLYGON 71.295 15.780 71.355 15.780 71.355 15.720 ;
        RECT 71.510 15.770 71.585 15.910 ;
        RECT 73.275 15.770 73.350 15.910 ;
        RECT 73.490 15.720 73.565 15.860 ;
        RECT 74.195 15.780 74.255 15.860 ;
        POLYGON 74.195 15.780 74.255 15.780 74.255 15.720 ;
        RECT 74.410 15.770 74.485 15.910 ;
        RECT 76.175 15.770 76.250 15.910 ;
        RECT 76.390 15.720 76.465 15.860 ;
        RECT 77.095 15.780 77.155 15.860 ;
        POLYGON 77.095 15.780 77.155 15.780 77.155 15.720 ;
        RECT 77.310 15.770 77.385 15.910 ;
        RECT 79.075 15.770 79.150 15.910 ;
        RECT 79.290 15.720 79.365 15.860 ;
        RECT 79.995 15.780 80.055 15.860 ;
        POLYGON 79.995 15.780 80.055 15.780 80.055 15.720 ;
        RECT 80.210 15.770 80.285 15.910 ;
        RECT 81.975 15.770 82.050 15.910 ;
        RECT 82.190 15.720 82.265 15.860 ;
        RECT 82.895 15.780 82.955 15.860 ;
        POLYGON 82.895 15.780 82.955 15.780 82.955 15.720 ;
        RECT 83.110 15.770 83.185 15.910 ;
        RECT 84.875 15.770 84.950 15.910 ;
        RECT 85.090 15.720 85.165 15.860 ;
        RECT 85.795 15.780 85.855 15.860 ;
        POLYGON 85.795 15.780 85.855 15.780 85.855 15.720 ;
        RECT 86.010 15.770 86.085 15.910 ;
        RECT 87.775 15.770 87.850 15.910 ;
        RECT 87.990 15.720 88.065 15.860 ;
        RECT 88.695 15.780 88.755 15.860 ;
        POLYGON 88.695 15.780 88.755 15.780 88.755 15.720 ;
        RECT 88.910 15.770 88.985 15.910 ;
        RECT 90.675 15.770 90.750 15.910 ;
        RECT 90.890 15.720 90.965 15.860 ;
        RECT 91.595 15.780 91.655 15.860 ;
        POLYGON 91.595 15.780 91.655 15.780 91.655 15.720 ;
        RECT 91.810 15.770 91.885 15.910 ;
        RECT 0.720 15.250 0.870 15.420 ;
        RECT 1.110 15.385 1.260 15.555 ;
        RECT 1.500 15.385 1.650 15.555 ;
        RECT 1.890 15.250 2.040 15.420 ;
        RECT 3.620 15.250 3.770 15.420 ;
        RECT 4.010 15.385 4.160 15.555 ;
        RECT 4.400 15.385 4.550 15.555 ;
        RECT 4.790 15.250 4.940 15.420 ;
        RECT 6.520 15.250 6.670 15.420 ;
        RECT 6.910 15.385 7.060 15.555 ;
        RECT 7.300 15.385 7.450 15.555 ;
        RECT 7.690 15.250 7.840 15.420 ;
        RECT 9.420 15.250 9.570 15.420 ;
        RECT 9.810 15.385 9.960 15.555 ;
        RECT 10.200 15.385 10.350 15.555 ;
        RECT 10.590 15.250 10.740 15.420 ;
        RECT 12.320 15.250 12.470 15.420 ;
        RECT 12.710 15.385 12.860 15.555 ;
        RECT 13.100 15.385 13.250 15.555 ;
        RECT 13.490 15.250 13.640 15.420 ;
        RECT 15.220 15.250 15.370 15.420 ;
        RECT 15.610 15.385 15.760 15.555 ;
        RECT 16.000 15.385 16.150 15.555 ;
        RECT 16.390 15.250 16.540 15.420 ;
        RECT 18.120 15.250 18.270 15.420 ;
        RECT 18.510 15.385 18.660 15.555 ;
        RECT 18.900 15.385 19.050 15.555 ;
        RECT 19.290 15.250 19.440 15.420 ;
        RECT 21.020 15.250 21.170 15.420 ;
        RECT 21.410 15.385 21.560 15.555 ;
        RECT 21.800 15.385 21.950 15.555 ;
        RECT 22.190 15.250 22.340 15.420 ;
        RECT 23.920 15.250 24.070 15.420 ;
        RECT 24.310 15.385 24.460 15.555 ;
        RECT 24.700 15.385 24.850 15.555 ;
        RECT 25.090 15.250 25.240 15.420 ;
        RECT 26.820 15.250 26.970 15.420 ;
        RECT 27.210 15.385 27.360 15.555 ;
        RECT 27.600 15.385 27.750 15.555 ;
        RECT 27.990 15.250 28.140 15.420 ;
        RECT 29.720 15.250 29.870 15.420 ;
        RECT 30.110 15.385 30.260 15.555 ;
        RECT 30.500 15.385 30.650 15.555 ;
        RECT 30.890 15.250 31.040 15.420 ;
        RECT 32.620 15.250 32.770 15.420 ;
        RECT 33.010 15.385 33.160 15.555 ;
        RECT 33.400 15.385 33.550 15.555 ;
        RECT 33.790 15.250 33.940 15.420 ;
        RECT 35.520 15.250 35.670 15.420 ;
        RECT 35.910 15.385 36.060 15.555 ;
        RECT 36.300 15.385 36.450 15.555 ;
        RECT 36.690 15.250 36.840 15.420 ;
        RECT 38.420 15.250 38.570 15.420 ;
        RECT 38.810 15.385 38.960 15.555 ;
        RECT 39.200 15.385 39.350 15.555 ;
        RECT 39.590 15.250 39.740 15.420 ;
        RECT 41.320 15.250 41.470 15.420 ;
        RECT 41.710 15.385 41.860 15.555 ;
        RECT 42.100 15.385 42.250 15.555 ;
        RECT 42.490 15.250 42.640 15.420 ;
        RECT 44.220 15.250 44.370 15.420 ;
        RECT 44.610 15.385 44.760 15.555 ;
        RECT 45.000 15.385 45.150 15.555 ;
        RECT 45.390 15.250 45.540 15.420 ;
        RECT 47.120 15.250 47.270 15.420 ;
        RECT 47.510 15.385 47.660 15.555 ;
        RECT 47.900 15.385 48.050 15.555 ;
        RECT 48.290 15.250 48.440 15.420 ;
        RECT 50.020 15.250 50.170 15.420 ;
        RECT 50.410 15.385 50.560 15.555 ;
        RECT 50.800 15.385 50.950 15.555 ;
        RECT 51.190 15.250 51.340 15.420 ;
        RECT 52.920 15.250 53.070 15.420 ;
        RECT 53.310 15.385 53.460 15.555 ;
        RECT 53.700 15.385 53.850 15.555 ;
        RECT 54.090 15.250 54.240 15.420 ;
        RECT 55.820 15.250 55.970 15.420 ;
        RECT 56.210 15.385 56.360 15.555 ;
        RECT 56.600 15.385 56.750 15.555 ;
        RECT 56.990 15.250 57.140 15.420 ;
        RECT 58.720 15.250 58.870 15.420 ;
        RECT 59.110 15.385 59.260 15.555 ;
        RECT 59.500 15.385 59.650 15.555 ;
        RECT 59.890 15.250 60.040 15.420 ;
        RECT 61.620 15.250 61.770 15.420 ;
        RECT 62.010 15.385 62.160 15.555 ;
        RECT 62.400 15.385 62.550 15.555 ;
        RECT 62.790 15.250 62.940 15.420 ;
        RECT 64.520 15.250 64.670 15.420 ;
        RECT 64.910 15.385 65.060 15.555 ;
        RECT 65.300 15.385 65.450 15.555 ;
        RECT 65.690 15.250 65.840 15.420 ;
        RECT 67.420 15.250 67.570 15.420 ;
        RECT 67.810 15.385 67.960 15.555 ;
        RECT 68.200 15.385 68.350 15.555 ;
        RECT 68.590 15.250 68.740 15.420 ;
        RECT 70.320 15.250 70.470 15.420 ;
        RECT 70.710 15.385 70.860 15.555 ;
        RECT 71.100 15.385 71.250 15.555 ;
        RECT 71.490 15.250 71.640 15.420 ;
        RECT 73.220 15.250 73.370 15.420 ;
        RECT 73.610 15.385 73.760 15.555 ;
        RECT 74.000 15.385 74.150 15.555 ;
        RECT 74.390 15.250 74.540 15.420 ;
        RECT 76.120 15.250 76.270 15.420 ;
        RECT 76.510 15.385 76.660 15.555 ;
        RECT 76.900 15.385 77.050 15.555 ;
        RECT 77.290 15.250 77.440 15.420 ;
        RECT 79.020 15.250 79.170 15.420 ;
        RECT 79.410 15.385 79.560 15.555 ;
        RECT 79.800 15.385 79.950 15.555 ;
        RECT 80.190 15.250 80.340 15.420 ;
        RECT 81.920 15.250 82.070 15.420 ;
        RECT 82.310 15.385 82.460 15.555 ;
        RECT 82.700 15.385 82.850 15.555 ;
        RECT 83.090 15.250 83.240 15.420 ;
        RECT 84.820 15.250 84.970 15.420 ;
        RECT 85.210 15.385 85.360 15.555 ;
        RECT 85.600 15.385 85.750 15.555 ;
        RECT 85.990 15.250 86.140 15.420 ;
        RECT 87.720 15.250 87.870 15.420 ;
        RECT 88.110 15.385 88.260 15.555 ;
        RECT 88.500 15.385 88.650 15.555 ;
        RECT 88.890 15.250 89.040 15.420 ;
        RECT 90.620 15.250 90.770 15.420 ;
        RECT 91.010 15.385 91.160 15.555 ;
        RECT 91.400 15.385 91.550 15.555 ;
        RECT 91.790 15.250 91.940 15.420 ;
        RECT 0.985 15.165 1.035 15.200 ;
        POLYGON 1.035 15.200 1.070 15.165 1.035 15.165 ;
        RECT 0.985 15.040 1.070 15.165 ;
        RECT 1.690 15.040 1.775 15.200 ;
        RECT 3.885 15.165 3.935 15.200 ;
        POLYGON 3.935 15.200 3.970 15.165 3.935 15.165 ;
        RECT 3.885 15.040 3.970 15.165 ;
        RECT 4.590 15.040 4.675 15.200 ;
        RECT 6.785 15.165 6.835 15.200 ;
        POLYGON 6.835 15.200 6.870 15.165 6.835 15.165 ;
        RECT 6.785 15.040 6.870 15.165 ;
        RECT 7.490 15.040 7.575 15.200 ;
        RECT 9.685 15.165 9.735 15.200 ;
        POLYGON 9.735 15.200 9.770 15.165 9.735 15.165 ;
        RECT 9.685 15.040 9.770 15.165 ;
        RECT 10.390 15.040 10.475 15.200 ;
        RECT 12.585 15.165 12.635 15.200 ;
        POLYGON 12.635 15.200 12.670 15.165 12.635 15.165 ;
        RECT 12.585 15.040 12.670 15.165 ;
        RECT 13.290 15.040 13.375 15.200 ;
        RECT 15.485 15.165 15.535 15.200 ;
        POLYGON 15.535 15.200 15.570 15.165 15.535 15.165 ;
        RECT 15.485 15.040 15.570 15.165 ;
        RECT 16.190 15.040 16.275 15.200 ;
        RECT 18.385 15.165 18.435 15.200 ;
        POLYGON 18.435 15.200 18.470 15.165 18.435 15.165 ;
        RECT 18.385 15.040 18.470 15.165 ;
        RECT 19.090 15.040 19.175 15.200 ;
        RECT 21.285 15.165 21.335 15.200 ;
        POLYGON 21.335 15.200 21.370 15.165 21.335 15.165 ;
        RECT 21.285 15.040 21.370 15.165 ;
        RECT 21.990 15.040 22.075 15.200 ;
        RECT 24.185 15.165 24.235 15.200 ;
        POLYGON 24.235 15.200 24.270 15.165 24.235 15.165 ;
        RECT 24.185 15.040 24.270 15.165 ;
        RECT 24.890 15.040 24.975 15.200 ;
        RECT 27.085 15.165 27.135 15.200 ;
        POLYGON 27.135 15.200 27.170 15.165 27.135 15.165 ;
        RECT 27.085 15.040 27.170 15.165 ;
        RECT 27.790 15.040 27.875 15.200 ;
        RECT 29.985 15.165 30.035 15.200 ;
        POLYGON 30.035 15.200 30.070 15.165 30.035 15.165 ;
        RECT 29.985 15.040 30.070 15.165 ;
        RECT 30.690 15.040 30.775 15.200 ;
        RECT 32.885 15.165 32.935 15.200 ;
        POLYGON 32.935 15.200 32.970 15.165 32.935 15.165 ;
        RECT 32.885 15.040 32.970 15.165 ;
        RECT 33.590 15.040 33.675 15.200 ;
        RECT 35.785 15.165 35.835 15.200 ;
        POLYGON 35.835 15.200 35.870 15.165 35.835 15.165 ;
        RECT 35.785 15.040 35.870 15.165 ;
        RECT 36.490 15.040 36.575 15.200 ;
        RECT 38.685 15.165 38.735 15.200 ;
        POLYGON 38.735 15.200 38.770 15.165 38.735 15.165 ;
        RECT 38.685 15.040 38.770 15.165 ;
        RECT 39.390 15.040 39.475 15.200 ;
        RECT 41.585 15.165 41.635 15.200 ;
        POLYGON 41.635 15.200 41.670 15.165 41.635 15.165 ;
        RECT 41.585 15.040 41.670 15.165 ;
        RECT 42.290 15.040 42.375 15.200 ;
        RECT 44.485 15.165 44.535 15.200 ;
        POLYGON 44.535 15.200 44.570 15.165 44.535 15.165 ;
        RECT 44.485 15.040 44.570 15.165 ;
        RECT 45.190 15.040 45.275 15.200 ;
        RECT 47.385 15.165 47.435 15.200 ;
        POLYGON 47.435 15.200 47.470 15.165 47.435 15.165 ;
        RECT 47.385 15.040 47.470 15.165 ;
        RECT 48.090 15.040 48.175 15.200 ;
        RECT 50.285 15.165 50.335 15.200 ;
        POLYGON 50.335 15.200 50.370 15.165 50.335 15.165 ;
        RECT 50.285 15.040 50.370 15.165 ;
        RECT 50.990 15.040 51.075 15.200 ;
        RECT 53.185 15.165 53.235 15.200 ;
        POLYGON 53.235 15.200 53.270 15.165 53.235 15.165 ;
        RECT 53.185 15.040 53.270 15.165 ;
        RECT 53.890 15.040 53.975 15.200 ;
        RECT 56.085 15.165 56.135 15.200 ;
        POLYGON 56.135 15.200 56.170 15.165 56.135 15.165 ;
        RECT 56.085 15.040 56.170 15.165 ;
        RECT 56.790 15.040 56.875 15.200 ;
        RECT 58.985 15.165 59.035 15.200 ;
        POLYGON 59.035 15.200 59.070 15.165 59.035 15.165 ;
        RECT 58.985 15.040 59.070 15.165 ;
        RECT 59.690 15.040 59.775 15.200 ;
        RECT 61.885 15.165 61.935 15.200 ;
        POLYGON 61.935 15.200 61.970 15.165 61.935 15.165 ;
        RECT 61.885 15.040 61.970 15.165 ;
        RECT 62.590 15.040 62.675 15.200 ;
        RECT 64.785 15.165 64.835 15.200 ;
        POLYGON 64.835 15.200 64.870 15.165 64.835 15.165 ;
        RECT 64.785 15.040 64.870 15.165 ;
        RECT 65.490 15.040 65.575 15.200 ;
        RECT 67.685 15.165 67.735 15.200 ;
        POLYGON 67.735 15.200 67.770 15.165 67.735 15.165 ;
        RECT 67.685 15.040 67.770 15.165 ;
        RECT 68.390 15.040 68.475 15.200 ;
        RECT 70.585 15.165 70.635 15.200 ;
        POLYGON 70.635 15.200 70.670 15.165 70.635 15.165 ;
        RECT 70.585 15.040 70.670 15.165 ;
        RECT 71.290 15.040 71.375 15.200 ;
        RECT 73.485 15.165 73.535 15.200 ;
        POLYGON 73.535 15.200 73.570 15.165 73.535 15.165 ;
        RECT 73.485 15.040 73.570 15.165 ;
        RECT 74.190 15.040 74.275 15.200 ;
        RECT 76.385 15.165 76.435 15.200 ;
        POLYGON 76.435 15.200 76.470 15.165 76.435 15.165 ;
        RECT 76.385 15.040 76.470 15.165 ;
        RECT 77.090 15.040 77.175 15.200 ;
        RECT 79.285 15.165 79.335 15.200 ;
        POLYGON 79.335 15.200 79.370 15.165 79.335 15.165 ;
        RECT 79.285 15.040 79.370 15.165 ;
        RECT 79.990 15.040 80.075 15.200 ;
        RECT 82.185 15.165 82.235 15.200 ;
        POLYGON 82.235 15.200 82.270 15.165 82.235 15.165 ;
        RECT 82.185 15.040 82.270 15.165 ;
        RECT 82.890 15.040 82.975 15.200 ;
        RECT 85.085 15.165 85.135 15.200 ;
        POLYGON 85.135 15.200 85.170 15.165 85.135 15.165 ;
        RECT 85.085 15.040 85.170 15.165 ;
        RECT 85.790 15.040 85.875 15.200 ;
        RECT 87.985 15.165 88.035 15.200 ;
        POLYGON 88.035 15.200 88.070 15.165 88.035 15.165 ;
        RECT 87.985 15.040 88.070 15.165 ;
        RECT 88.690 15.040 88.775 15.200 ;
        RECT 90.885 15.165 90.935 15.200 ;
        POLYGON 90.935 15.200 90.970 15.165 90.935 15.165 ;
        RECT 90.885 15.040 90.970 15.165 ;
        RECT 91.590 15.040 91.675 15.200 ;
        RECT 0.775 14.420 0.850 14.560 ;
        RECT 0.990 14.370 1.065 14.510 ;
        RECT 1.695 14.430 1.755 14.510 ;
        POLYGON 1.695 14.430 1.755 14.430 1.755 14.370 ;
        RECT 1.910 14.420 1.985 14.560 ;
        RECT 3.675 14.420 3.750 14.560 ;
        RECT 3.890 14.370 3.965 14.510 ;
        RECT 4.595 14.430 4.655 14.510 ;
        POLYGON 4.595 14.430 4.655 14.430 4.655 14.370 ;
        RECT 4.810 14.420 4.885 14.560 ;
        RECT 6.575 14.420 6.650 14.560 ;
        RECT 6.790 14.370 6.865 14.510 ;
        RECT 7.495 14.430 7.555 14.510 ;
        POLYGON 7.495 14.430 7.555 14.430 7.555 14.370 ;
        RECT 7.710 14.420 7.785 14.560 ;
        RECT 9.475 14.420 9.550 14.560 ;
        RECT 9.690 14.370 9.765 14.510 ;
        RECT 10.395 14.430 10.455 14.510 ;
        POLYGON 10.395 14.430 10.455 14.430 10.455 14.370 ;
        RECT 10.610 14.420 10.685 14.560 ;
        RECT 12.375 14.420 12.450 14.560 ;
        RECT 12.590 14.370 12.665 14.510 ;
        RECT 13.295 14.430 13.355 14.510 ;
        POLYGON 13.295 14.430 13.355 14.430 13.355 14.370 ;
        RECT 13.510 14.420 13.585 14.560 ;
        RECT 15.275 14.420 15.350 14.560 ;
        RECT 15.490 14.370 15.565 14.510 ;
        RECT 16.195 14.430 16.255 14.510 ;
        POLYGON 16.195 14.430 16.255 14.430 16.255 14.370 ;
        RECT 16.410 14.420 16.485 14.560 ;
        RECT 18.175 14.420 18.250 14.560 ;
        RECT 18.390 14.370 18.465 14.510 ;
        RECT 19.095 14.430 19.155 14.510 ;
        POLYGON 19.095 14.430 19.155 14.430 19.155 14.370 ;
        RECT 19.310 14.420 19.385 14.560 ;
        RECT 21.075 14.420 21.150 14.560 ;
        RECT 21.290 14.370 21.365 14.510 ;
        RECT 21.995 14.430 22.055 14.510 ;
        POLYGON 21.995 14.430 22.055 14.430 22.055 14.370 ;
        RECT 22.210 14.420 22.285 14.560 ;
        RECT 23.975 14.420 24.050 14.560 ;
        RECT 24.190 14.370 24.265 14.510 ;
        RECT 24.895 14.430 24.955 14.510 ;
        POLYGON 24.895 14.430 24.955 14.430 24.955 14.370 ;
        RECT 25.110 14.420 25.185 14.560 ;
        RECT 26.875 14.420 26.950 14.560 ;
        RECT 27.090 14.370 27.165 14.510 ;
        RECT 27.795 14.430 27.855 14.510 ;
        POLYGON 27.795 14.430 27.855 14.430 27.855 14.370 ;
        RECT 28.010 14.420 28.085 14.560 ;
        RECT 29.775 14.420 29.850 14.560 ;
        RECT 29.990 14.370 30.065 14.510 ;
        RECT 30.695 14.430 30.755 14.510 ;
        POLYGON 30.695 14.430 30.755 14.430 30.755 14.370 ;
        RECT 30.910 14.420 30.985 14.560 ;
        RECT 32.675 14.420 32.750 14.560 ;
        RECT 32.890 14.370 32.965 14.510 ;
        RECT 33.595 14.430 33.655 14.510 ;
        POLYGON 33.595 14.430 33.655 14.430 33.655 14.370 ;
        RECT 33.810 14.420 33.885 14.560 ;
        RECT 35.575 14.420 35.650 14.560 ;
        RECT 35.790 14.370 35.865 14.510 ;
        RECT 36.495 14.430 36.555 14.510 ;
        POLYGON 36.495 14.430 36.555 14.430 36.555 14.370 ;
        RECT 36.710 14.420 36.785 14.560 ;
        RECT 38.475 14.420 38.550 14.560 ;
        RECT 38.690 14.370 38.765 14.510 ;
        RECT 39.395 14.430 39.455 14.510 ;
        POLYGON 39.395 14.430 39.455 14.430 39.455 14.370 ;
        RECT 39.610 14.420 39.685 14.560 ;
        RECT 41.375 14.420 41.450 14.560 ;
        RECT 41.590 14.370 41.665 14.510 ;
        RECT 42.295 14.430 42.355 14.510 ;
        POLYGON 42.295 14.430 42.355 14.430 42.355 14.370 ;
        RECT 42.510 14.420 42.585 14.560 ;
        RECT 44.275 14.420 44.350 14.560 ;
        RECT 44.490 14.370 44.565 14.510 ;
        RECT 45.195 14.430 45.255 14.510 ;
        POLYGON 45.195 14.430 45.255 14.430 45.255 14.370 ;
        RECT 45.410 14.420 45.485 14.560 ;
        RECT 47.175 14.420 47.250 14.560 ;
        RECT 47.390 14.370 47.465 14.510 ;
        RECT 48.095 14.430 48.155 14.510 ;
        POLYGON 48.095 14.430 48.155 14.430 48.155 14.370 ;
        RECT 48.310 14.420 48.385 14.560 ;
        RECT 50.075 14.420 50.150 14.560 ;
        RECT 50.290 14.370 50.365 14.510 ;
        RECT 50.995 14.430 51.055 14.510 ;
        POLYGON 50.995 14.430 51.055 14.430 51.055 14.370 ;
        RECT 51.210 14.420 51.285 14.560 ;
        RECT 52.975 14.420 53.050 14.560 ;
        RECT 53.190 14.370 53.265 14.510 ;
        RECT 53.895 14.430 53.955 14.510 ;
        POLYGON 53.895 14.430 53.955 14.430 53.955 14.370 ;
        RECT 54.110 14.420 54.185 14.560 ;
        RECT 55.875 14.420 55.950 14.560 ;
        RECT 56.090 14.370 56.165 14.510 ;
        RECT 56.795 14.430 56.855 14.510 ;
        POLYGON 56.795 14.430 56.855 14.430 56.855 14.370 ;
        RECT 57.010 14.420 57.085 14.560 ;
        RECT 58.775 14.420 58.850 14.560 ;
        RECT 58.990 14.370 59.065 14.510 ;
        RECT 59.695 14.430 59.755 14.510 ;
        POLYGON 59.695 14.430 59.755 14.430 59.755 14.370 ;
        RECT 59.910 14.420 59.985 14.560 ;
        RECT 61.675 14.420 61.750 14.560 ;
        RECT 61.890 14.370 61.965 14.510 ;
        RECT 62.595 14.430 62.655 14.510 ;
        POLYGON 62.595 14.430 62.655 14.430 62.655 14.370 ;
        RECT 62.810 14.420 62.885 14.560 ;
        RECT 64.575 14.420 64.650 14.560 ;
        RECT 64.790 14.370 64.865 14.510 ;
        RECT 65.495 14.430 65.555 14.510 ;
        POLYGON 65.495 14.430 65.555 14.430 65.555 14.370 ;
        RECT 65.710 14.420 65.785 14.560 ;
        RECT 67.475 14.420 67.550 14.560 ;
        RECT 67.690 14.370 67.765 14.510 ;
        RECT 68.395 14.430 68.455 14.510 ;
        POLYGON 68.395 14.430 68.455 14.430 68.455 14.370 ;
        RECT 68.610 14.420 68.685 14.560 ;
        RECT 70.375 14.420 70.450 14.560 ;
        RECT 70.590 14.370 70.665 14.510 ;
        RECT 71.295 14.430 71.355 14.510 ;
        POLYGON 71.295 14.430 71.355 14.430 71.355 14.370 ;
        RECT 71.510 14.420 71.585 14.560 ;
        RECT 73.275 14.420 73.350 14.560 ;
        RECT 73.490 14.370 73.565 14.510 ;
        RECT 74.195 14.430 74.255 14.510 ;
        POLYGON 74.195 14.430 74.255 14.430 74.255 14.370 ;
        RECT 74.410 14.420 74.485 14.560 ;
        RECT 76.175 14.420 76.250 14.560 ;
        RECT 76.390 14.370 76.465 14.510 ;
        RECT 77.095 14.430 77.155 14.510 ;
        POLYGON 77.095 14.430 77.155 14.430 77.155 14.370 ;
        RECT 77.310 14.420 77.385 14.560 ;
        RECT 79.075 14.420 79.150 14.560 ;
        RECT 79.290 14.370 79.365 14.510 ;
        RECT 79.995 14.430 80.055 14.510 ;
        POLYGON 79.995 14.430 80.055 14.430 80.055 14.370 ;
        RECT 80.210 14.420 80.285 14.560 ;
        RECT 81.975 14.420 82.050 14.560 ;
        RECT 82.190 14.370 82.265 14.510 ;
        RECT 82.895 14.430 82.955 14.510 ;
        POLYGON 82.895 14.430 82.955 14.430 82.955 14.370 ;
        RECT 83.110 14.420 83.185 14.560 ;
        RECT 84.875 14.420 84.950 14.560 ;
        RECT 85.090 14.370 85.165 14.510 ;
        RECT 85.795 14.430 85.855 14.510 ;
        POLYGON 85.795 14.430 85.855 14.430 85.855 14.370 ;
        RECT 86.010 14.420 86.085 14.560 ;
        RECT 87.775 14.420 87.850 14.560 ;
        RECT 87.990 14.370 88.065 14.510 ;
        RECT 88.695 14.430 88.755 14.510 ;
        POLYGON 88.695 14.430 88.755 14.430 88.755 14.370 ;
        RECT 88.910 14.420 88.985 14.560 ;
        RECT 90.675 14.420 90.750 14.560 ;
        RECT 90.890 14.370 90.965 14.510 ;
        RECT 91.595 14.430 91.655 14.510 ;
        POLYGON 91.595 14.430 91.655 14.430 91.655 14.370 ;
        RECT 91.810 14.420 91.885 14.560 ;
        RECT 0.720 13.900 0.870 14.070 ;
        RECT 1.110 14.035 1.260 14.205 ;
        RECT 1.500 14.035 1.650 14.205 ;
        RECT 1.890 13.900 2.040 14.070 ;
        RECT 3.620 13.900 3.770 14.070 ;
        RECT 4.010 14.035 4.160 14.205 ;
        RECT 4.400 14.035 4.550 14.205 ;
        RECT 4.790 13.900 4.940 14.070 ;
        RECT 6.520 13.900 6.670 14.070 ;
        RECT 6.910 14.035 7.060 14.205 ;
        RECT 7.300 14.035 7.450 14.205 ;
        RECT 7.690 13.900 7.840 14.070 ;
        RECT 9.420 13.900 9.570 14.070 ;
        RECT 9.810 14.035 9.960 14.205 ;
        RECT 10.200 14.035 10.350 14.205 ;
        RECT 10.590 13.900 10.740 14.070 ;
        RECT 12.320 13.900 12.470 14.070 ;
        RECT 12.710 14.035 12.860 14.205 ;
        RECT 13.100 14.035 13.250 14.205 ;
        RECT 13.490 13.900 13.640 14.070 ;
        RECT 15.220 13.900 15.370 14.070 ;
        RECT 15.610 14.035 15.760 14.205 ;
        RECT 16.000 14.035 16.150 14.205 ;
        RECT 16.390 13.900 16.540 14.070 ;
        RECT 18.120 13.900 18.270 14.070 ;
        RECT 18.510 14.035 18.660 14.205 ;
        RECT 18.900 14.035 19.050 14.205 ;
        RECT 19.290 13.900 19.440 14.070 ;
        RECT 21.020 13.900 21.170 14.070 ;
        RECT 21.410 14.035 21.560 14.205 ;
        RECT 21.800 14.035 21.950 14.205 ;
        RECT 22.190 13.900 22.340 14.070 ;
        RECT 23.920 13.900 24.070 14.070 ;
        RECT 24.310 14.035 24.460 14.205 ;
        RECT 24.700 14.035 24.850 14.205 ;
        RECT 25.090 13.900 25.240 14.070 ;
        RECT 26.820 13.900 26.970 14.070 ;
        RECT 27.210 14.035 27.360 14.205 ;
        RECT 27.600 14.035 27.750 14.205 ;
        RECT 27.990 13.900 28.140 14.070 ;
        RECT 29.720 13.900 29.870 14.070 ;
        RECT 30.110 14.035 30.260 14.205 ;
        RECT 30.500 14.035 30.650 14.205 ;
        RECT 30.890 13.900 31.040 14.070 ;
        RECT 32.620 13.900 32.770 14.070 ;
        RECT 33.010 14.035 33.160 14.205 ;
        RECT 33.400 14.035 33.550 14.205 ;
        RECT 33.790 13.900 33.940 14.070 ;
        RECT 35.520 13.900 35.670 14.070 ;
        RECT 35.910 14.035 36.060 14.205 ;
        RECT 36.300 14.035 36.450 14.205 ;
        RECT 36.690 13.900 36.840 14.070 ;
        RECT 38.420 13.900 38.570 14.070 ;
        RECT 38.810 14.035 38.960 14.205 ;
        RECT 39.200 14.035 39.350 14.205 ;
        RECT 39.590 13.900 39.740 14.070 ;
        RECT 41.320 13.900 41.470 14.070 ;
        RECT 41.710 14.035 41.860 14.205 ;
        RECT 42.100 14.035 42.250 14.205 ;
        RECT 42.490 13.900 42.640 14.070 ;
        RECT 44.220 13.900 44.370 14.070 ;
        RECT 44.610 14.035 44.760 14.205 ;
        RECT 45.000 14.035 45.150 14.205 ;
        RECT 45.390 13.900 45.540 14.070 ;
        RECT 47.120 13.900 47.270 14.070 ;
        RECT 47.510 14.035 47.660 14.205 ;
        RECT 47.900 14.035 48.050 14.205 ;
        RECT 48.290 13.900 48.440 14.070 ;
        RECT 50.020 13.900 50.170 14.070 ;
        RECT 50.410 14.035 50.560 14.205 ;
        RECT 50.800 14.035 50.950 14.205 ;
        RECT 51.190 13.900 51.340 14.070 ;
        RECT 52.920 13.900 53.070 14.070 ;
        RECT 53.310 14.035 53.460 14.205 ;
        RECT 53.700 14.035 53.850 14.205 ;
        RECT 54.090 13.900 54.240 14.070 ;
        RECT 55.820 13.900 55.970 14.070 ;
        RECT 56.210 14.035 56.360 14.205 ;
        RECT 56.600 14.035 56.750 14.205 ;
        RECT 56.990 13.900 57.140 14.070 ;
        RECT 58.720 13.900 58.870 14.070 ;
        RECT 59.110 14.035 59.260 14.205 ;
        RECT 59.500 14.035 59.650 14.205 ;
        RECT 59.890 13.900 60.040 14.070 ;
        RECT 61.620 13.900 61.770 14.070 ;
        RECT 62.010 14.035 62.160 14.205 ;
        RECT 62.400 14.035 62.550 14.205 ;
        RECT 62.790 13.900 62.940 14.070 ;
        RECT 64.520 13.900 64.670 14.070 ;
        RECT 64.910 14.035 65.060 14.205 ;
        RECT 65.300 14.035 65.450 14.205 ;
        RECT 65.690 13.900 65.840 14.070 ;
        RECT 67.420 13.900 67.570 14.070 ;
        RECT 67.810 14.035 67.960 14.205 ;
        RECT 68.200 14.035 68.350 14.205 ;
        RECT 68.590 13.900 68.740 14.070 ;
        RECT 70.320 13.900 70.470 14.070 ;
        RECT 70.710 14.035 70.860 14.205 ;
        RECT 71.100 14.035 71.250 14.205 ;
        RECT 71.490 13.900 71.640 14.070 ;
        RECT 73.220 13.900 73.370 14.070 ;
        RECT 73.610 14.035 73.760 14.205 ;
        RECT 74.000 14.035 74.150 14.205 ;
        RECT 74.390 13.900 74.540 14.070 ;
        RECT 76.120 13.900 76.270 14.070 ;
        RECT 76.510 14.035 76.660 14.205 ;
        RECT 76.900 14.035 77.050 14.205 ;
        RECT 77.290 13.900 77.440 14.070 ;
        RECT 79.020 13.900 79.170 14.070 ;
        RECT 79.410 14.035 79.560 14.205 ;
        RECT 79.800 14.035 79.950 14.205 ;
        RECT 80.190 13.900 80.340 14.070 ;
        RECT 81.920 13.900 82.070 14.070 ;
        RECT 82.310 14.035 82.460 14.205 ;
        RECT 82.700 14.035 82.850 14.205 ;
        RECT 83.090 13.900 83.240 14.070 ;
        RECT 84.820 13.900 84.970 14.070 ;
        RECT 85.210 14.035 85.360 14.205 ;
        RECT 85.600 14.035 85.750 14.205 ;
        RECT 85.990 13.900 86.140 14.070 ;
        RECT 87.720 13.900 87.870 14.070 ;
        RECT 88.110 14.035 88.260 14.205 ;
        RECT 88.500 14.035 88.650 14.205 ;
        RECT 88.890 13.900 89.040 14.070 ;
        RECT 90.620 13.900 90.770 14.070 ;
        RECT 91.010 14.035 91.160 14.205 ;
        RECT 91.400 14.035 91.550 14.205 ;
        RECT 91.790 13.900 91.940 14.070 ;
        RECT 0.985 13.815 1.035 13.850 ;
        POLYGON 1.035 13.850 1.070 13.815 1.035 13.815 ;
        RECT 0.985 13.690 1.070 13.815 ;
        RECT 1.690 13.690 1.775 13.850 ;
        RECT 3.885 13.815 3.935 13.850 ;
        POLYGON 3.935 13.850 3.970 13.815 3.935 13.815 ;
        RECT 3.885 13.690 3.970 13.815 ;
        RECT 4.590 13.690 4.675 13.850 ;
        RECT 6.785 13.815 6.835 13.850 ;
        POLYGON 6.835 13.850 6.870 13.815 6.835 13.815 ;
        RECT 6.785 13.690 6.870 13.815 ;
        RECT 7.490 13.690 7.575 13.850 ;
        RECT 9.685 13.815 9.735 13.850 ;
        POLYGON 9.735 13.850 9.770 13.815 9.735 13.815 ;
        RECT 9.685 13.690 9.770 13.815 ;
        RECT 10.390 13.690 10.475 13.850 ;
        RECT 12.585 13.815 12.635 13.850 ;
        POLYGON 12.635 13.850 12.670 13.815 12.635 13.815 ;
        RECT 12.585 13.690 12.670 13.815 ;
        RECT 13.290 13.690 13.375 13.850 ;
        RECT 15.485 13.815 15.535 13.850 ;
        POLYGON 15.535 13.850 15.570 13.815 15.535 13.815 ;
        RECT 15.485 13.690 15.570 13.815 ;
        RECT 16.190 13.690 16.275 13.850 ;
        RECT 18.385 13.815 18.435 13.850 ;
        POLYGON 18.435 13.850 18.470 13.815 18.435 13.815 ;
        RECT 18.385 13.690 18.470 13.815 ;
        RECT 19.090 13.690 19.175 13.850 ;
        RECT 21.285 13.815 21.335 13.850 ;
        POLYGON 21.335 13.850 21.370 13.815 21.335 13.815 ;
        RECT 21.285 13.690 21.370 13.815 ;
        RECT 21.990 13.690 22.075 13.850 ;
        RECT 24.185 13.815 24.235 13.850 ;
        POLYGON 24.235 13.850 24.270 13.815 24.235 13.815 ;
        RECT 24.185 13.690 24.270 13.815 ;
        RECT 24.890 13.690 24.975 13.850 ;
        RECT 27.085 13.815 27.135 13.850 ;
        POLYGON 27.135 13.850 27.170 13.815 27.135 13.815 ;
        RECT 27.085 13.690 27.170 13.815 ;
        RECT 27.790 13.690 27.875 13.850 ;
        RECT 29.985 13.815 30.035 13.850 ;
        POLYGON 30.035 13.850 30.070 13.815 30.035 13.815 ;
        RECT 29.985 13.690 30.070 13.815 ;
        RECT 30.690 13.690 30.775 13.850 ;
        RECT 32.885 13.815 32.935 13.850 ;
        POLYGON 32.935 13.850 32.970 13.815 32.935 13.815 ;
        RECT 32.885 13.690 32.970 13.815 ;
        RECT 33.590 13.690 33.675 13.850 ;
        RECT 35.785 13.815 35.835 13.850 ;
        POLYGON 35.835 13.850 35.870 13.815 35.835 13.815 ;
        RECT 35.785 13.690 35.870 13.815 ;
        RECT 36.490 13.690 36.575 13.850 ;
        RECT 38.685 13.815 38.735 13.850 ;
        POLYGON 38.735 13.850 38.770 13.815 38.735 13.815 ;
        RECT 38.685 13.690 38.770 13.815 ;
        RECT 39.390 13.690 39.475 13.850 ;
        RECT 41.585 13.815 41.635 13.850 ;
        POLYGON 41.635 13.850 41.670 13.815 41.635 13.815 ;
        RECT 41.585 13.690 41.670 13.815 ;
        RECT 42.290 13.690 42.375 13.850 ;
        RECT 44.485 13.815 44.535 13.850 ;
        POLYGON 44.535 13.850 44.570 13.815 44.535 13.815 ;
        RECT 44.485 13.690 44.570 13.815 ;
        RECT 45.190 13.690 45.275 13.850 ;
        RECT 47.385 13.815 47.435 13.850 ;
        POLYGON 47.435 13.850 47.470 13.815 47.435 13.815 ;
        RECT 47.385 13.690 47.470 13.815 ;
        RECT 48.090 13.690 48.175 13.850 ;
        RECT 50.285 13.815 50.335 13.850 ;
        POLYGON 50.335 13.850 50.370 13.815 50.335 13.815 ;
        RECT 50.285 13.690 50.370 13.815 ;
        RECT 50.990 13.690 51.075 13.850 ;
        RECT 53.185 13.815 53.235 13.850 ;
        POLYGON 53.235 13.850 53.270 13.815 53.235 13.815 ;
        RECT 53.185 13.690 53.270 13.815 ;
        RECT 53.890 13.690 53.975 13.850 ;
        RECT 56.085 13.815 56.135 13.850 ;
        POLYGON 56.135 13.850 56.170 13.815 56.135 13.815 ;
        RECT 56.085 13.690 56.170 13.815 ;
        RECT 56.790 13.690 56.875 13.850 ;
        RECT 58.985 13.815 59.035 13.850 ;
        POLYGON 59.035 13.850 59.070 13.815 59.035 13.815 ;
        RECT 58.985 13.690 59.070 13.815 ;
        RECT 59.690 13.690 59.775 13.850 ;
        RECT 61.885 13.815 61.935 13.850 ;
        POLYGON 61.935 13.850 61.970 13.815 61.935 13.815 ;
        RECT 61.885 13.690 61.970 13.815 ;
        RECT 62.590 13.690 62.675 13.850 ;
        RECT 64.785 13.815 64.835 13.850 ;
        POLYGON 64.835 13.850 64.870 13.815 64.835 13.815 ;
        RECT 64.785 13.690 64.870 13.815 ;
        RECT 65.490 13.690 65.575 13.850 ;
        RECT 67.685 13.815 67.735 13.850 ;
        POLYGON 67.735 13.850 67.770 13.815 67.735 13.815 ;
        RECT 67.685 13.690 67.770 13.815 ;
        RECT 68.390 13.690 68.475 13.850 ;
        RECT 70.585 13.815 70.635 13.850 ;
        POLYGON 70.635 13.850 70.670 13.815 70.635 13.815 ;
        RECT 70.585 13.690 70.670 13.815 ;
        RECT 71.290 13.690 71.375 13.850 ;
        RECT 73.485 13.815 73.535 13.850 ;
        POLYGON 73.535 13.850 73.570 13.815 73.535 13.815 ;
        RECT 73.485 13.690 73.570 13.815 ;
        RECT 74.190 13.690 74.275 13.850 ;
        RECT 76.385 13.815 76.435 13.850 ;
        POLYGON 76.435 13.850 76.470 13.815 76.435 13.815 ;
        RECT 76.385 13.690 76.470 13.815 ;
        RECT 77.090 13.690 77.175 13.850 ;
        RECT 79.285 13.815 79.335 13.850 ;
        POLYGON 79.335 13.850 79.370 13.815 79.335 13.815 ;
        RECT 79.285 13.690 79.370 13.815 ;
        RECT 79.990 13.690 80.075 13.850 ;
        RECT 82.185 13.815 82.235 13.850 ;
        POLYGON 82.235 13.850 82.270 13.815 82.235 13.815 ;
        RECT 82.185 13.690 82.270 13.815 ;
        RECT 82.890 13.690 82.975 13.850 ;
        RECT 85.085 13.815 85.135 13.850 ;
        POLYGON 85.135 13.850 85.170 13.815 85.135 13.815 ;
        RECT 85.085 13.690 85.170 13.815 ;
        RECT 85.790 13.690 85.875 13.850 ;
        RECT 87.985 13.815 88.035 13.850 ;
        POLYGON 88.035 13.850 88.070 13.815 88.035 13.815 ;
        RECT 87.985 13.690 88.070 13.815 ;
        RECT 88.690 13.690 88.775 13.850 ;
        RECT 90.885 13.815 90.935 13.850 ;
        POLYGON 90.935 13.850 90.970 13.815 90.935 13.815 ;
        RECT 90.885 13.690 90.970 13.815 ;
        RECT 91.590 13.690 91.675 13.850 ;
        RECT 0.775 13.070 0.850 13.210 ;
        RECT 0.990 13.020 1.065 13.160 ;
        RECT 1.695 13.080 1.755 13.160 ;
        POLYGON 1.695 13.080 1.755 13.080 1.755 13.020 ;
        RECT 1.910 13.070 1.985 13.210 ;
        RECT 3.675 13.070 3.750 13.210 ;
        RECT 3.890 13.020 3.965 13.160 ;
        RECT 4.595 13.080 4.655 13.160 ;
        POLYGON 4.595 13.080 4.655 13.080 4.655 13.020 ;
        RECT 4.810 13.070 4.885 13.210 ;
        RECT 6.575 13.070 6.650 13.210 ;
        RECT 6.790 13.020 6.865 13.160 ;
        RECT 7.495 13.080 7.555 13.160 ;
        POLYGON 7.495 13.080 7.555 13.080 7.555 13.020 ;
        RECT 7.710 13.070 7.785 13.210 ;
        RECT 9.475 13.070 9.550 13.210 ;
        RECT 9.690 13.020 9.765 13.160 ;
        RECT 10.395 13.080 10.455 13.160 ;
        POLYGON 10.395 13.080 10.455 13.080 10.455 13.020 ;
        RECT 10.610 13.070 10.685 13.210 ;
        RECT 12.375 13.070 12.450 13.210 ;
        RECT 12.590 13.020 12.665 13.160 ;
        RECT 13.295 13.080 13.355 13.160 ;
        POLYGON 13.295 13.080 13.355 13.080 13.355 13.020 ;
        RECT 13.510 13.070 13.585 13.210 ;
        RECT 15.275 13.070 15.350 13.210 ;
        RECT 15.490 13.020 15.565 13.160 ;
        RECT 16.195 13.080 16.255 13.160 ;
        POLYGON 16.195 13.080 16.255 13.080 16.255 13.020 ;
        RECT 16.410 13.070 16.485 13.210 ;
        RECT 18.175 13.070 18.250 13.210 ;
        RECT 18.390 13.020 18.465 13.160 ;
        RECT 19.095 13.080 19.155 13.160 ;
        POLYGON 19.095 13.080 19.155 13.080 19.155 13.020 ;
        RECT 19.310 13.070 19.385 13.210 ;
        RECT 21.075 13.070 21.150 13.210 ;
        RECT 21.290 13.020 21.365 13.160 ;
        RECT 21.995 13.080 22.055 13.160 ;
        POLYGON 21.995 13.080 22.055 13.080 22.055 13.020 ;
        RECT 22.210 13.070 22.285 13.210 ;
        RECT 23.975 13.070 24.050 13.210 ;
        RECT 24.190 13.020 24.265 13.160 ;
        RECT 24.895 13.080 24.955 13.160 ;
        POLYGON 24.895 13.080 24.955 13.080 24.955 13.020 ;
        RECT 25.110 13.070 25.185 13.210 ;
        RECT 26.875 13.070 26.950 13.210 ;
        RECT 27.090 13.020 27.165 13.160 ;
        RECT 27.795 13.080 27.855 13.160 ;
        POLYGON 27.795 13.080 27.855 13.080 27.855 13.020 ;
        RECT 28.010 13.070 28.085 13.210 ;
        RECT 29.775 13.070 29.850 13.210 ;
        RECT 29.990 13.020 30.065 13.160 ;
        RECT 30.695 13.080 30.755 13.160 ;
        POLYGON 30.695 13.080 30.755 13.080 30.755 13.020 ;
        RECT 30.910 13.070 30.985 13.210 ;
        RECT 32.675 13.070 32.750 13.210 ;
        RECT 32.890 13.020 32.965 13.160 ;
        RECT 33.595 13.080 33.655 13.160 ;
        POLYGON 33.595 13.080 33.655 13.080 33.655 13.020 ;
        RECT 33.810 13.070 33.885 13.210 ;
        RECT 35.575 13.070 35.650 13.210 ;
        RECT 35.790 13.020 35.865 13.160 ;
        RECT 36.495 13.080 36.555 13.160 ;
        POLYGON 36.495 13.080 36.555 13.080 36.555 13.020 ;
        RECT 36.710 13.070 36.785 13.210 ;
        RECT 38.475 13.070 38.550 13.210 ;
        RECT 38.690 13.020 38.765 13.160 ;
        RECT 39.395 13.080 39.455 13.160 ;
        POLYGON 39.395 13.080 39.455 13.080 39.455 13.020 ;
        RECT 39.610 13.070 39.685 13.210 ;
        RECT 41.375 13.070 41.450 13.210 ;
        RECT 41.590 13.020 41.665 13.160 ;
        RECT 42.295 13.080 42.355 13.160 ;
        POLYGON 42.295 13.080 42.355 13.080 42.355 13.020 ;
        RECT 42.510 13.070 42.585 13.210 ;
        RECT 44.275 13.070 44.350 13.210 ;
        RECT 44.490 13.020 44.565 13.160 ;
        RECT 45.195 13.080 45.255 13.160 ;
        POLYGON 45.195 13.080 45.255 13.080 45.255 13.020 ;
        RECT 45.410 13.070 45.485 13.210 ;
        RECT 47.175 13.070 47.250 13.210 ;
        RECT 47.390 13.020 47.465 13.160 ;
        RECT 48.095 13.080 48.155 13.160 ;
        POLYGON 48.095 13.080 48.155 13.080 48.155 13.020 ;
        RECT 48.310 13.070 48.385 13.210 ;
        RECT 50.075 13.070 50.150 13.210 ;
        RECT 50.290 13.020 50.365 13.160 ;
        RECT 50.995 13.080 51.055 13.160 ;
        POLYGON 50.995 13.080 51.055 13.080 51.055 13.020 ;
        RECT 51.210 13.070 51.285 13.210 ;
        RECT 52.975 13.070 53.050 13.210 ;
        RECT 53.190 13.020 53.265 13.160 ;
        RECT 53.895 13.080 53.955 13.160 ;
        POLYGON 53.895 13.080 53.955 13.080 53.955 13.020 ;
        RECT 54.110 13.070 54.185 13.210 ;
        RECT 55.875 13.070 55.950 13.210 ;
        RECT 56.090 13.020 56.165 13.160 ;
        RECT 56.795 13.080 56.855 13.160 ;
        POLYGON 56.795 13.080 56.855 13.080 56.855 13.020 ;
        RECT 57.010 13.070 57.085 13.210 ;
        RECT 58.775 13.070 58.850 13.210 ;
        RECT 58.990 13.020 59.065 13.160 ;
        RECT 59.695 13.080 59.755 13.160 ;
        POLYGON 59.695 13.080 59.755 13.080 59.755 13.020 ;
        RECT 59.910 13.070 59.985 13.210 ;
        RECT 61.675 13.070 61.750 13.210 ;
        RECT 61.890 13.020 61.965 13.160 ;
        RECT 62.595 13.080 62.655 13.160 ;
        POLYGON 62.595 13.080 62.655 13.080 62.655 13.020 ;
        RECT 62.810 13.070 62.885 13.210 ;
        RECT 64.575 13.070 64.650 13.210 ;
        RECT 64.790 13.020 64.865 13.160 ;
        RECT 65.495 13.080 65.555 13.160 ;
        POLYGON 65.495 13.080 65.555 13.080 65.555 13.020 ;
        RECT 65.710 13.070 65.785 13.210 ;
        RECT 67.475 13.070 67.550 13.210 ;
        RECT 67.690 13.020 67.765 13.160 ;
        RECT 68.395 13.080 68.455 13.160 ;
        POLYGON 68.395 13.080 68.455 13.080 68.455 13.020 ;
        RECT 68.610 13.070 68.685 13.210 ;
        RECT 70.375 13.070 70.450 13.210 ;
        RECT 70.590 13.020 70.665 13.160 ;
        RECT 71.295 13.080 71.355 13.160 ;
        POLYGON 71.295 13.080 71.355 13.080 71.355 13.020 ;
        RECT 71.510 13.070 71.585 13.210 ;
        RECT 73.275 13.070 73.350 13.210 ;
        RECT 73.490 13.020 73.565 13.160 ;
        RECT 74.195 13.080 74.255 13.160 ;
        POLYGON 74.195 13.080 74.255 13.080 74.255 13.020 ;
        RECT 74.410 13.070 74.485 13.210 ;
        RECT 76.175 13.070 76.250 13.210 ;
        RECT 76.390 13.020 76.465 13.160 ;
        RECT 77.095 13.080 77.155 13.160 ;
        POLYGON 77.095 13.080 77.155 13.080 77.155 13.020 ;
        RECT 77.310 13.070 77.385 13.210 ;
        RECT 79.075 13.070 79.150 13.210 ;
        RECT 79.290 13.020 79.365 13.160 ;
        RECT 79.995 13.080 80.055 13.160 ;
        POLYGON 79.995 13.080 80.055 13.080 80.055 13.020 ;
        RECT 80.210 13.070 80.285 13.210 ;
        RECT 81.975 13.070 82.050 13.210 ;
        RECT 82.190 13.020 82.265 13.160 ;
        RECT 82.895 13.080 82.955 13.160 ;
        POLYGON 82.895 13.080 82.955 13.080 82.955 13.020 ;
        RECT 83.110 13.070 83.185 13.210 ;
        RECT 84.875 13.070 84.950 13.210 ;
        RECT 85.090 13.020 85.165 13.160 ;
        RECT 85.795 13.080 85.855 13.160 ;
        POLYGON 85.795 13.080 85.855 13.080 85.855 13.020 ;
        RECT 86.010 13.070 86.085 13.210 ;
        RECT 87.775 13.070 87.850 13.210 ;
        RECT 87.990 13.020 88.065 13.160 ;
        RECT 88.695 13.080 88.755 13.160 ;
        POLYGON 88.695 13.080 88.755 13.080 88.755 13.020 ;
        RECT 88.910 13.070 88.985 13.210 ;
        RECT 90.675 13.070 90.750 13.210 ;
        RECT 90.890 13.020 90.965 13.160 ;
        RECT 91.595 13.080 91.655 13.160 ;
        POLYGON 91.595 13.080 91.655 13.080 91.655 13.020 ;
        RECT 91.810 13.070 91.885 13.210 ;
        RECT 0.720 12.550 0.870 12.720 ;
        RECT 1.110 12.685 1.260 12.855 ;
        RECT 1.500 12.685 1.650 12.855 ;
        RECT 1.890 12.550 2.040 12.720 ;
        RECT 3.620 12.550 3.770 12.720 ;
        RECT 4.010 12.685 4.160 12.855 ;
        RECT 4.400 12.685 4.550 12.855 ;
        RECT 4.790 12.550 4.940 12.720 ;
        RECT 6.520 12.550 6.670 12.720 ;
        RECT 6.910 12.685 7.060 12.855 ;
        RECT 7.300 12.685 7.450 12.855 ;
        RECT 7.690 12.550 7.840 12.720 ;
        RECT 9.420 12.550 9.570 12.720 ;
        RECT 9.810 12.685 9.960 12.855 ;
        RECT 10.200 12.685 10.350 12.855 ;
        RECT 10.590 12.550 10.740 12.720 ;
        RECT 12.320 12.550 12.470 12.720 ;
        RECT 12.710 12.685 12.860 12.855 ;
        RECT 13.100 12.685 13.250 12.855 ;
        RECT 13.490 12.550 13.640 12.720 ;
        RECT 15.220 12.550 15.370 12.720 ;
        RECT 15.610 12.685 15.760 12.855 ;
        RECT 16.000 12.685 16.150 12.855 ;
        RECT 16.390 12.550 16.540 12.720 ;
        RECT 18.120 12.550 18.270 12.720 ;
        RECT 18.510 12.685 18.660 12.855 ;
        RECT 18.900 12.685 19.050 12.855 ;
        RECT 19.290 12.550 19.440 12.720 ;
        RECT 21.020 12.550 21.170 12.720 ;
        RECT 21.410 12.685 21.560 12.855 ;
        RECT 21.800 12.685 21.950 12.855 ;
        RECT 22.190 12.550 22.340 12.720 ;
        RECT 23.920 12.550 24.070 12.720 ;
        RECT 24.310 12.685 24.460 12.855 ;
        RECT 24.700 12.685 24.850 12.855 ;
        RECT 25.090 12.550 25.240 12.720 ;
        RECT 26.820 12.550 26.970 12.720 ;
        RECT 27.210 12.685 27.360 12.855 ;
        RECT 27.600 12.685 27.750 12.855 ;
        RECT 27.990 12.550 28.140 12.720 ;
        RECT 29.720 12.550 29.870 12.720 ;
        RECT 30.110 12.685 30.260 12.855 ;
        RECT 30.500 12.685 30.650 12.855 ;
        RECT 30.890 12.550 31.040 12.720 ;
        RECT 32.620 12.550 32.770 12.720 ;
        RECT 33.010 12.685 33.160 12.855 ;
        RECT 33.400 12.685 33.550 12.855 ;
        RECT 33.790 12.550 33.940 12.720 ;
        RECT 35.520 12.550 35.670 12.720 ;
        RECT 35.910 12.685 36.060 12.855 ;
        RECT 36.300 12.685 36.450 12.855 ;
        RECT 36.690 12.550 36.840 12.720 ;
        RECT 38.420 12.550 38.570 12.720 ;
        RECT 38.810 12.685 38.960 12.855 ;
        RECT 39.200 12.685 39.350 12.855 ;
        RECT 39.590 12.550 39.740 12.720 ;
        RECT 41.320 12.550 41.470 12.720 ;
        RECT 41.710 12.685 41.860 12.855 ;
        RECT 42.100 12.685 42.250 12.855 ;
        RECT 42.490 12.550 42.640 12.720 ;
        RECT 44.220 12.550 44.370 12.720 ;
        RECT 44.610 12.685 44.760 12.855 ;
        RECT 45.000 12.685 45.150 12.855 ;
        RECT 45.390 12.550 45.540 12.720 ;
        RECT 47.120 12.550 47.270 12.720 ;
        RECT 47.510 12.685 47.660 12.855 ;
        RECT 47.900 12.685 48.050 12.855 ;
        RECT 48.290 12.550 48.440 12.720 ;
        RECT 50.020 12.550 50.170 12.720 ;
        RECT 50.410 12.685 50.560 12.855 ;
        RECT 50.800 12.685 50.950 12.855 ;
        RECT 51.190 12.550 51.340 12.720 ;
        RECT 52.920 12.550 53.070 12.720 ;
        RECT 53.310 12.685 53.460 12.855 ;
        RECT 53.700 12.685 53.850 12.855 ;
        RECT 54.090 12.550 54.240 12.720 ;
        RECT 55.820 12.550 55.970 12.720 ;
        RECT 56.210 12.685 56.360 12.855 ;
        RECT 56.600 12.685 56.750 12.855 ;
        RECT 56.990 12.550 57.140 12.720 ;
        RECT 58.720 12.550 58.870 12.720 ;
        RECT 59.110 12.685 59.260 12.855 ;
        RECT 59.500 12.685 59.650 12.855 ;
        RECT 59.890 12.550 60.040 12.720 ;
        RECT 61.620 12.550 61.770 12.720 ;
        RECT 62.010 12.685 62.160 12.855 ;
        RECT 62.400 12.685 62.550 12.855 ;
        RECT 62.790 12.550 62.940 12.720 ;
        RECT 64.520 12.550 64.670 12.720 ;
        RECT 64.910 12.685 65.060 12.855 ;
        RECT 65.300 12.685 65.450 12.855 ;
        RECT 65.690 12.550 65.840 12.720 ;
        RECT 67.420 12.550 67.570 12.720 ;
        RECT 67.810 12.685 67.960 12.855 ;
        RECT 68.200 12.685 68.350 12.855 ;
        RECT 68.590 12.550 68.740 12.720 ;
        RECT 70.320 12.550 70.470 12.720 ;
        RECT 70.710 12.685 70.860 12.855 ;
        RECT 71.100 12.685 71.250 12.855 ;
        RECT 71.490 12.550 71.640 12.720 ;
        RECT 73.220 12.550 73.370 12.720 ;
        RECT 73.610 12.685 73.760 12.855 ;
        RECT 74.000 12.685 74.150 12.855 ;
        RECT 74.390 12.550 74.540 12.720 ;
        RECT 76.120 12.550 76.270 12.720 ;
        RECT 76.510 12.685 76.660 12.855 ;
        RECT 76.900 12.685 77.050 12.855 ;
        RECT 77.290 12.550 77.440 12.720 ;
        RECT 79.020 12.550 79.170 12.720 ;
        RECT 79.410 12.685 79.560 12.855 ;
        RECT 79.800 12.685 79.950 12.855 ;
        RECT 80.190 12.550 80.340 12.720 ;
        RECT 81.920 12.550 82.070 12.720 ;
        RECT 82.310 12.685 82.460 12.855 ;
        RECT 82.700 12.685 82.850 12.855 ;
        RECT 83.090 12.550 83.240 12.720 ;
        RECT 84.820 12.550 84.970 12.720 ;
        RECT 85.210 12.685 85.360 12.855 ;
        RECT 85.600 12.685 85.750 12.855 ;
        RECT 85.990 12.550 86.140 12.720 ;
        RECT 87.720 12.550 87.870 12.720 ;
        RECT 88.110 12.685 88.260 12.855 ;
        RECT 88.500 12.685 88.650 12.855 ;
        RECT 88.890 12.550 89.040 12.720 ;
        RECT 90.620 12.550 90.770 12.720 ;
        RECT 91.010 12.685 91.160 12.855 ;
        RECT 91.400 12.685 91.550 12.855 ;
        RECT 91.790 12.550 91.940 12.720 ;
        RECT 0.985 12.465 1.035 12.500 ;
        POLYGON 1.035 12.500 1.070 12.465 1.035 12.465 ;
        RECT 0.985 12.340 1.070 12.465 ;
        RECT 1.690 12.340 1.775 12.500 ;
        RECT 3.885 12.465 3.935 12.500 ;
        POLYGON 3.935 12.500 3.970 12.465 3.935 12.465 ;
        RECT 3.885 12.340 3.970 12.465 ;
        RECT 4.590 12.340 4.675 12.500 ;
        RECT 6.785 12.465 6.835 12.500 ;
        POLYGON 6.835 12.500 6.870 12.465 6.835 12.465 ;
        RECT 6.785 12.340 6.870 12.465 ;
        RECT 7.490 12.340 7.575 12.500 ;
        RECT 9.685 12.465 9.735 12.500 ;
        POLYGON 9.735 12.500 9.770 12.465 9.735 12.465 ;
        RECT 9.685 12.340 9.770 12.465 ;
        RECT 10.390 12.340 10.475 12.500 ;
        RECT 12.585 12.465 12.635 12.500 ;
        POLYGON 12.635 12.500 12.670 12.465 12.635 12.465 ;
        RECT 12.585 12.340 12.670 12.465 ;
        RECT 13.290 12.340 13.375 12.500 ;
        RECT 15.485 12.465 15.535 12.500 ;
        POLYGON 15.535 12.500 15.570 12.465 15.535 12.465 ;
        RECT 15.485 12.340 15.570 12.465 ;
        RECT 16.190 12.340 16.275 12.500 ;
        RECT 18.385 12.465 18.435 12.500 ;
        POLYGON 18.435 12.500 18.470 12.465 18.435 12.465 ;
        RECT 18.385 12.340 18.470 12.465 ;
        RECT 19.090 12.340 19.175 12.500 ;
        RECT 21.285 12.465 21.335 12.500 ;
        POLYGON 21.335 12.500 21.370 12.465 21.335 12.465 ;
        RECT 21.285 12.340 21.370 12.465 ;
        RECT 21.990 12.340 22.075 12.500 ;
        RECT 24.185 12.465 24.235 12.500 ;
        POLYGON 24.235 12.500 24.270 12.465 24.235 12.465 ;
        RECT 24.185 12.340 24.270 12.465 ;
        RECT 24.890 12.340 24.975 12.500 ;
        RECT 27.085 12.465 27.135 12.500 ;
        POLYGON 27.135 12.500 27.170 12.465 27.135 12.465 ;
        RECT 27.085 12.340 27.170 12.465 ;
        RECT 27.790 12.340 27.875 12.500 ;
        RECT 29.985 12.465 30.035 12.500 ;
        POLYGON 30.035 12.500 30.070 12.465 30.035 12.465 ;
        RECT 29.985 12.340 30.070 12.465 ;
        RECT 30.690 12.340 30.775 12.500 ;
        RECT 32.885 12.465 32.935 12.500 ;
        POLYGON 32.935 12.500 32.970 12.465 32.935 12.465 ;
        RECT 32.885 12.340 32.970 12.465 ;
        RECT 33.590 12.340 33.675 12.500 ;
        RECT 35.785 12.465 35.835 12.500 ;
        POLYGON 35.835 12.500 35.870 12.465 35.835 12.465 ;
        RECT 35.785 12.340 35.870 12.465 ;
        RECT 36.490 12.340 36.575 12.500 ;
        RECT 38.685 12.465 38.735 12.500 ;
        POLYGON 38.735 12.500 38.770 12.465 38.735 12.465 ;
        RECT 38.685 12.340 38.770 12.465 ;
        RECT 39.390 12.340 39.475 12.500 ;
        RECT 41.585 12.465 41.635 12.500 ;
        POLYGON 41.635 12.500 41.670 12.465 41.635 12.465 ;
        RECT 41.585 12.340 41.670 12.465 ;
        RECT 42.290 12.340 42.375 12.500 ;
        RECT 44.485 12.465 44.535 12.500 ;
        POLYGON 44.535 12.500 44.570 12.465 44.535 12.465 ;
        RECT 44.485 12.340 44.570 12.465 ;
        RECT 45.190 12.340 45.275 12.500 ;
        RECT 47.385 12.465 47.435 12.500 ;
        POLYGON 47.435 12.500 47.470 12.465 47.435 12.465 ;
        RECT 47.385 12.340 47.470 12.465 ;
        RECT 48.090 12.340 48.175 12.500 ;
        RECT 50.285 12.465 50.335 12.500 ;
        POLYGON 50.335 12.500 50.370 12.465 50.335 12.465 ;
        RECT 50.285 12.340 50.370 12.465 ;
        RECT 50.990 12.340 51.075 12.500 ;
        RECT 53.185 12.465 53.235 12.500 ;
        POLYGON 53.235 12.500 53.270 12.465 53.235 12.465 ;
        RECT 53.185 12.340 53.270 12.465 ;
        RECT 53.890 12.340 53.975 12.500 ;
        RECT 56.085 12.465 56.135 12.500 ;
        POLYGON 56.135 12.500 56.170 12.465 56.135 12.465 ;
        RECT 56.085 12.340 56.170 12.465 ;
        RECT 56.790 12.340 56.875 12.500 ;
        RECT 58.985 12.465 59.035 12.500 ;
        POLYGON 59.035 12.500 59.070 12.465 59.035 12.465 ;
        RECT 58.985 12.340 59.070 12.465 ;
        RECT 59.690 12.340 59.775 12.500 ;
        RECT 61.885 12.465 61.935 12.500 ;
        POLYGON 61.935 12.500 61.970 12.465 61.935 12.465 ;
        RECT 61.885 12.340 61.970 12.465 ;
        RECT 62.590 12.340 62.675 12.500 ;
        RECT 64.785 12.465 64.835 12.500 ;
        POLYGON 64.835 12.500 64.870 12.465 64.835 12.465 ;
        RECT 64.785 12.340 64.870 12.465 ;
        RECT 65.490 12.340 65.575 12.500 ;
        RECT 67.685 12.465 67.735 12.500 ;
        POLYGON 67.735 12.500 67.770 12.465 67.735 12.465 ;
        RECT 67.685 12.340 67.770 12.465 ;
        RECT 68.390 12.340 68.475 12.500 ;
        RECT 70.585 12.465 70.635 12.500 ;
        POLYGON 70.635 12.500 70.670 12.465 70.635 12.465 ;
        RECT 70.585 12.340 70.670 12.465 ;
        RECT 71.290 12.340 71.375 12.500 ;
        RECT 73.485 12.465 73.535 12.500 ;
        POLYGON 73.535 12.500 73.570 12.465 73.535 12.465 ;
        RECT 73.485 12.340 73.570 12.465 ;
        RECT 74.190 12.340 74.275 12.500 ;
        RECT 76.385 12.465 76.435 12.500 ;
        POLYGON 76.435 12.500 76.470 12.465 76.435 12.465 ;
        RECT 76.385 12.340 76.470 12.465 ;
        RECT 77.090 12.340 77.175 12.500 ;
        RECT 79.285 12.465 79.335 12.500 ;
        POLYGON 79.335 12.500 79.370 12.465 79.335 12.465 ;
        RECT 79.285 12.340 79.370 12.465 ;
        RECT 79.990 12.340 80.075 12.500 ;
        RECT 82.185 12.465 82.235 12.500 ;
        POLYGON 82.235 12.500 82.270 12.465 82.235 12.465 ;
        RECT 82.185 12.340 82.270 12.465 ;
        RECT 82.890 12.340 82.975 12.500 ;
        RECT 85.085 12.465 85.135 12.500 ;
        POLYGON 85.135 12.500 85.170 12.465 85.135 12.465 ;
        RECT 85.085 12.340 85.170 12.465 ;
        RECT 85.790 12.340 85.875 12.500 ;
        RECT 87.985 12.465 88.035 12.500 ;
        POLYGON 88.035 12.500 88.070 12.465 88.035 12.465 ;
        RECT 87.985 12.340 88.070 12.465 ;
        RECT 88.690 12.340 88.775 12.500 ;
        RECT 90.885 12.465 90.935 12.500 ;
        POLYGON 90.935 12.500 90.970 12.465 90.935 12.465 ;
        RECT 90.885 12.340 90.970 12.465 ;
        RECT 91.590 12.340 91.675 12.500 ;
        RECT 0.775 11.720 0.850 11.860 ;
        RECT 0.990 11.670 1.065 11.810 ;
        RECT 1.695 11.730 1.755 11.810 ;
        POLYGON 1.695 11.730 1.755 11.730 1.755 11.670 ;
        RECT 1.910 11.720 1.985 11.860 ;
        RECT 3.675 11.720 3.750 11.860 ;
        RECT 3.890 11.670 3.965 11.810 ;
        RECT 4.595 11.730 4.655 11.810 ;
        POLYGON 4.595 11.730 4.655 11.730 4.655 11.670 ;
        RECT 4.810 11.720 4.885 11.860 ;
        RECT 6.575 11.720 6.650 11.860 ;
        RECT 6.790 11.670 6.865 11.810 ;
        RECT 7.495 11.730 7.555 11.810 ;
        POLYGON 7.495 11.730 7.555 11.730 7.555 11.670 ;
        RECT 7.710 11.720 7.785 11.860 ;
        RECT 9.475 11.720 9.550 11.860 ;
        RECT 9.690 11.670 9.765 11.810 ;
        RECT 10.395 11.730 10.455 11.810 ;
        POLYGON 10.395 11.730 10.455 11.730 10.455 11.670 ;
        RECT 10.610 11.720 10.685 11.860 ;
        RECT 12.375 11.720 12.450 11.860 ;
        RECT 12.590 11.670 12.665 11.810 ;
        RECT 13.295 11.730 13.355 11.810 ;
        POLYGON 13.295 11.730 13.355 11.730 13.355 11.670 ;
        RECT 13.510 11.720 13.585 11.860 ;
        RECT 15.275 11.720 15.350 11.860 ;
        RECT 15.490 11.670 15.565 11.810 ;
        RECT 16.195 11.730 16.255 11.810 ;
        POLYGON 16.195 11.730 16.255 11.730 16.255 11.670 ;
        RECT 16.410 11.720 16.485 11.860 ;
        RECT 18.175 11.720 18.250 11.860 ;
        RECT 18.390 11.670 18.465 11.810 ;
        RECT 19.095 11.730 19.155 11.810 ;
        POLYGON 19.095 11.730 19.155 11.730 19.155 11.670 ;
        RECT 19.310 11.720 19.385 11.860 ;
        RECT 21.075 11.720 21.150 11.860 ;
        RECT 21.290 11.670 21.365 11.810 ;
        RECT 21.995 11.730 22.055 11.810 ;
        POLYGON 21.995 11.730 22.055 11.730 22.055 11.670 ;
        RECT 22.210 11.720 22.285 11.860 ;
        RECT 23.975 11.720 24.050 11.860 ;
        RECT 24.190 11.670 24.265 11.810 ;
        RECT 24.895 11.730 24.955 11.810 ;
        POLYGON 24.895 11.730 24.955 11.730 24.955 11.670 ;
        RECT 25.110 11.720 25.185 11.860 ;
        RECT 26.875 11.720 26.950 11.860 ;
        RECT 27.090 11.670 27.165 11.810 ;
        RECT 27.795 11.730 27.855 11.810 ;
        POLYGON 27.795 11.730 27.855 11.730 27.855 11.670 ;
        RECT 28.010 11.720 28.085 11.860 ;
        RECT 29.775 11.720 29.850 11.860 ;
        RECT 29.990 11.670 30.065 11.810 ;
        RECT 30.695 11.730 30.755 11.810 ;
        POLYGON 30.695 11.730 30.755 11.730 30.755 11.670 ;
        RECT 30.910 11.720 30.985 11.860 ;
        RECT 32.675 11.720 32.750 11.860 ;
        RECT 32.890 11.670 32.965 11.810 ;
        RECT 33.595 11.730 33.655 11.810 ;
        POLYGON 33.595 11.730 33.655 11.730 33.655 11.670 ;
        RECT 33.810 11.720 33.885 11.860 ;
        RECT 35.575 11.720 35.650 11.860 ;
        RECT 35.790 11.670 35.865 11.810 ;
        RECT 36.495 11.730 36.555 11.810 ;
        POLYGON 36.495 11.730 36.555 11.730 36.555 11.670 ;
        RECT 36.710 11.720 36.785 11.860 ;
        RECT 38.475 11.720 38.550 11.860 ;
        RECT 38.690 11.670 38.765 11.810 ;
        RECT 39.395 11.730 39.455 11.810 ;
        POLYGON 39.395 11.730 39.455 11.730 39.455 11.670 ;
        RECT 39.610 11.720 39.685 11.860 ;
        RECT 41.375 11.720 41.450 11.860 ;
        RECT 41.590 11.670 41.665 11.810 ;
        RECT 42.295 11.730 42.355 11.810 ;
        POLYGON 42.295 11.730 42.355 11.730 42.355 11.670 ;
        RECT 42.510 11.720 42.585 11.860 ;
        RECT 44.275 11.720 44.350 11.860 ;
        RECT 44.490 11.670 44.565 11.810 ;
        RECT 45.195 11.730 45.255 11.810 ;
        POLYGON 45.195 11.730 45.255 11.730 45.255 11.670 ;
        RECT 45.410 11.720 45.485 11.860 ;
        RECT 47.175 11.720 47.250 11.860 ;
        RECT 47.390 11.670 47.465 11.810 ;
        RECT 48.095 11.730 48.155 11.810 ;
        POLYGON 48.095 11.730 48.155 11.730 48.155 11.670 ;
        RECT 48.310 11.720 48.385 11.860 ;
        RECT 50.075 11.720 50.150 11.860 ;
        RECT 50.290 11.670 50.365 11.810 ;
        RECT 50.995 11.730 51.055 11.810 ;
        POLYGON 50.995 11.730 51.055 11.730 51.055 11.670 ;
        RECT 51.210 11.720 51.285 11.860 ;
        RECT 52.975 11.720 53.050 11.860 ;
        RECT 53.190 11.670 53.265 11.810 ;
        RECT 53.895 11.730 53.955 11.810 ;
        POLYGON 53.895 11.730 53.955 11.730 53.955 11.670 ;
        RECT 54.110 11.720 54.185 11.860 ;
        RECT 55.875 11.720 55.950 11.860 ;
        RECT 56.090 11.670 56.165 11.810 ;
        RECT 56.795 11.730 56.855 11.810 ;
        POLYGON 56.795 11.730 56.855 11.730 56.855 11.670 ;
        RECT 57.010 11.720 57.085 11.860 ;
        RECT 58.775 11.720 58.850 11.860 ;
        RECT 58.990 11.670 59.065 11.810 ;
        RECT 59.695 11.730 59.755 11.810 ;
        POLYGON 59.695 11.730 59.755 11.730 59.755 11.670 ;
        RECT 59.910 11.720 59.985 11.860 ;
        RECT 61.675 11.720 61.750 11.860 ;
        RECT 61.890 11.670 61.965 11.810 ;
        RECT 62.595 11.730 62.655 11.810 ;
        POLYGON 62.595 11.730 62.655 11.730 62.655 11.670 ;
        RECT 62.810 11.720 62.885 11.860 ;
        RECT 64.575 11.720 64.650 11.860 ;
        RECT 64.790 11.670 64.865 11.810 ;
        RECT 65.495 11.730 65.555 11.810 ;
        POLYGON 65.495 11.730 65.555 11.730 65.555 11.670 ;
        RECT 65.710 11.720 65.785 11.860 ;
        RECT 67.475 11.720 67.550 11.860 ;
        RECT 67.690 11.670 67.765 11.810 ;
        RECT 68.395 11.730 68.455 11.810 ;
        POLYGON 68.395 11.730 68.455 11.730 68.455 11.670 ;
        RECT 68.610 11.720 68.685 11.860 ;
        RECT 70.375 11.720 70.450 11.860 ;
        RECT 70.590 11.670 70.665 11.810 ;
        RECT 71.295 11.730 71.355 11.810 ;
        POLYGON 71.295 11.730 71.355 11.730 71.355 11.670 ;
        RECT 71.510 11.720 71.585 11.860 ;
        RECT 73.275 11.720 73.350 11.860 ;
        RECT 73.490 11.670 73.565 11.810 ;
        RECT 74.195 11.730 74.255 11.810 ;
        POLYGON 74.195 11.730 74.255 11.730 74.255 11.670 ;
        RECT 74.410 11.720 74.485 11.860 ;
        RECT 76.175 11.720 76.250 11.860 ;
        RECT 76.390 11.670 76.465 11.810 ;
        RECT 77.095 11.730 77.155 11.810 ;
        POLYGON 77.095 11.730 77.155 11.730 77.155 11.670 ;
        RECT 77.310 11.720 77.385 11.860 ;
        RECT 79.075 11.720 79.150 11.860 ;
        RECT 79.290 11.670 79.365 11.810 ;
        RECT 79.995 11.730 80.055 11.810 ;
        POLYGON 79.995 11.730 80.055 11.730 80.055 11.670 ;
        RECT 80.210 11.720 80.285 11.860 ;
        RECT 81.975 11.720 82.050 11.860 ;
        RECT 82.190 11.670 82.265 11.810 ;
        RECT 82.895 11.730 82.955 11.810 ;
        POLYGON 82.895 11.730 82.955 11.730 82.955 11.670 ;
        RECT 83.110 11.720 83.185 11.860 ;
        RECT 84.875 11.720 84.950 11.860 ;
        RECT 85.090 11.670 85.165 11.810 ;
        RECT 85.795 11.730 85.855 11.810 ;
        POLYGON 85.795 11.730 85.855 11.730 85.855 11.670 ;
        RECT 86.010 11.720 86.085 11.860 ;
        RECT 87.775 11.720 87.850 11.860 ;
        RECT 87.990 11.670 88.065 11.810 ;
        RECT 88.695 11.730 88.755 11.810 ;
        POLYGON 88.695 11.730 88.755 11.730 88.755 11.670 ;
        RECT 88.910 11.720 88.985 11.860 ;
        RECT 90.675 11.720 90.750 11.860 ;
        RECT 90.890 11.670 90.965 11.810 ;
        RECT 91.595 11.730 91.655 11.810 ;
        POLYGON 91.595 11.730 91.655 11.730 91.655 11.670 ;
        RECT 91.810 11.720 91.885 11.860 ;
        RECT 0.720 11.200 0.870 11.370 ;
        RECT 1.110 11.335 1.260 11.505 ;
        RECT 1.500 11.335 1.650 11.505 ;
        RECT 1.890 11.200 2.040 11.370 ;
        RECT 3.620 11.200 3.770 11.370 ;
        RECT 4.010 11.335 4.160 11.505 ;
        RECT 4.400 11.335 4.550 11.505 ;
        RECT 4.790 11.200 4.940 11.370 ;
        RECT 6.520 11.200 6.670 11.370 ;
        RECT 6.910 11.335 7.060 11.505 ;
        RECT 7.300 11.335 7.450 11.505 ;
        RECT 7.690 11.200 7.840 11.370 ;
        RECT 9.420 11.200 9.570 11.370 ;
        RECT 9.810 11.335 9.960 11.505 ;
        RECT 10.200 11.335 10.350 11.505 ;
        RECT 10.590 11.200 10.740 11.370 ;
        RECT 12.320 11.200 12.470 11.370 ;
        RECT 12.710 11.335 12.860 11.505 ;
        RECT 13.100 11.335 13.250 11.505 ;
        RECT 13.490 11.200 13.640 11.370 ;
        RECT 15.220 11.200 15.370 11.370 ;
        RECT 15.610 11.335 15.760 11.505 ;
        RECT 16.000 11.335 16.150 11.505 ;
        RECT 16.390 11.200 16.540 11.370 ;
        RECT 18.120 11.200 18.270 11.370 ;
        RECT 18.510 11.335 18.660 11.505 ;
        RECT 18.900 11.335 19.050 11.505 ;
        RECT 19.290 11.200 19.440 11.370 ;
        RECT 21.020 11.200 21.170 11.370 ;
        RECT 21.410 11.335 21.560 11.505 ;
        RECT 21.800 11.335 21.950 11.505 ;
        RECT 22.190 11.200 22.340 11.370 ;
        RECT 23.920 11.200 24.070 11.370 ;
        RECT 24.310 11.335 24.460 11.505 ;
        RECT 24.700 11.335 24.850 11.505 ;
        RECT 25.090 11.200 25.240 11.370 ;
        RECT 26.820 11.200 26.970 11.370 ;
        RECT 27.210 11.335 27.360 11.505 ;
        RECT 27.600 11.335 27.750 11.505 ;
        RECT 27.990 11.200 28.140 11.370 ;
        RECT 29.720 11.200 29.870 11.370 ;
        RECT 30.110 11.335 30.260 11.505 ;
        RECT 30.500 11.335 30.650 11.505 ;
        RECT 30.890 11.200 31.040 11.370 ;
        RECT 32.620 11.200 32.770 11.370 ;
        RECT 33.010 11.335 33.160 11.505 ;
        RECT 33.400 11.335 33.550 11.505 ;
        RECT 33.790 11.200 33.940 11.370 ;
        RECT 35.520 11.200 35.670 11.370 ;
        RECT 35.910 11.335 36.060 11.505 ;
        RECT 36.300 11.335 36.450 11.505 ;
        RECT 36.690 11.200 36.840 11.370 ;
        RECT 38.420 11.200 38.570 11.370 ;
        RECT 38.810 11.335 38.960 11.505 ;
        RECT 39.200 11.335 39.350 11.505 ;
        RECT 39.590 11.200 39.740 11.370 ;
        RECT 41.320 11.200 41.470 11.370 ;
        RECT 41.710 11.335 41.860 11.505 ;
        RECT 42.100 11.335 42.250 11.505 ;
        RECT 42.490 11.200 42.640 11.370 ;
        RECT 44.220 11.200 44.370 11.370 ;
        RECT 44.610 11.335 44.760 11.505 ;
        RECT 45.000 11.335 45.150 11.505 ;
        RECT 45.390 11.200 45.540 11.370 ;
        RECT 47.120 11.200 47.270 11.370 ;
        RECT 47.510 11.335 47.660 11.505 ;
        RECT 47.900 11.335 48.050 11.505 ;
        RECT 48.290 11.200 48.440 11.370 ;
        RECT 50.020 11.200 50.170 11.370 ;
        RECT 50.410 11.335 50.560 11.505 ;
        RECT 50.800 11.335 50.950 11.505 ;
        RECT 51.190 11.200 51.340 11.370 ;
        RECT 52.920 11.200 53.070 11.370 ;
        RECT 53.310 11.335 53.460 11.505 ;
        RECT 53.700 11.335 53.850 11.505 ;
        RECT 54.090 11.200 54.240 11.370 ;
        RECT 55.820 11.200 55.970 11.370 ;
        RECT 56.210 11.335 56.360 11.505 ;
        RECT 56.600 11.335 56.750 11.505 ;
        RECT 56.990 11.200 57.140 11.370 ;
        RECT 58.720 11.200 58.870 11.370 ;
        RECT 59.110 11.335 59.260 11.505 ;
        RECT 59.500 11.335 59.650 11.505 ;
        RECT 59.890 11.200 60.040 11.370 ;
        RECT 61.620 11.200 61.770 11.370 ;
        RECT 62.010 11.335 62.160 11.505 ;
        RECT 62.400 11.335 62.550 11.505 ;
        RECT 62.790 11.200 62.940 11.370 ;
        RECT 64.520 11.200 64.670 11.370 ;
        RECT 64.910 11.335 65.060 11.505 ;
        RECT 65.300 11.335 65.450 11.505 ;
        RECT 65.690 11.200 65.840 11.370 ;
        RECT 67.420 11.200 67.570 11.370 ;
        RECT 67.810 11.335 67.960 11.505 ;
        RECT 68.200 11.335 68.350 11.505 ;
        RECT 68.590 11.200 68.740 11.370 ;
        RECT 70.320 11.200 70.470 11.370 ;
        RECT 70.710 11.335 70.860 11.505 ;
        RECT 71.100 11.335 71.250 11.505 ;
        RECT 71.490 11.200 71.640 11.370 ;
        RECT 73.220 11.200 73.370 11.370 ;
        RECT 73.610 11.335 73.760 11.505 ;
        RECT 74.000 11.335 74.150 11.505 ;
        RECT 74.390 11.200 74.540 11.370 ;
        RECT 76.120 11.200 76.270 11.370 ;
        RECT 76.510 11.335 76.660 11.505 ;
        RECT 76.900 11.335 77.050 11.505 ;
        RECT 77.290 11.200 77.440 11.370 ;
        RECT 79.020 11.200 79.170 11.370 ;
        RECT 79.410 11.335 79.560 11.505 ;
        RECT 79.800 11.335 79.950 11.505 ;
        RECT 80.190 11.200 80.340 11.370 ;
        RECT 81.920 11.200 82.070 11.370 ;
        RECT 82.310 11.335 82.460 11.505 ;
        RECT 82.700 11.335 82.850 11.505 ;
        RECT 83.090 11.200 83.240 11.370 ;
        RECT 84.820 11.200 84.970 11.370 ;
        RECT 85.210 11.335 85.360 11.505 ;
        RECT 85.600 11.335 85.750 11.505 ;
        RECT 85.990 11.200 86.140 11.370 ;
        RECT 87.720 11.200 87.870 11.370 ;
        RECT 88.110 11.335 88.260 11.505 ;
        RECT 88.500 11.335 88.650 11.505 ;
        RECT 88.890 11.200 89.040 11.370 ;
        RECT 90.620 11.200 90.770 11.370 ;
        RECT 91.010 11.335 91.160 11.505 ;
        RECT 91.400 11.335 91.550 11.505 ;
        RECT 91.790 11.200 91.940 11.370 ;
        RECT 0.985 11.115 1.035 11.150 ;
        POLYGON 1.035 11.150 1.070 11.115 1.035 11.115 ;
        RECT 0.985 10.990 1.070 11.115 ;
        RECT 1.690 10.990 1.775 11.150 ;
        RECT 3.885 11.115 3.935 11.150 ;
        POLYGON 3.935 11.150 3.970 11.115 3.935 11.115 ;
        RECT 3.885 10.990 3.970 11.115 ;
        RECT 4.590 10.990 4.675 11.150 ;
        RECT 6.785 11.115 6.835 11.150 ;
        POLYGON 6.835 11.150 6.870 11.115 6.835 11.115 ;
        RECT 6.785 10.990 6.870 11.115 ;
        RECT 7.490 10.990 7.575 11.150 ;
        RECT 9.685 11.115 9.735 11.150 ;
        POLYGON 9.735 11.150 9.770 11.115 9.735 11.115 ;
        RECT 9.685 10.990 9.770 11.115 ;
        RECT 10.390 10.990 10.475 11.150 ;
        RECT 12.585 11.115 12.635 11.150 ;
        POLYGON 12.635 11.150 12.670 11.115 12.635 11.115 ;
        RECT 12.585 10.990 12.670 11.115 ;
        RECT 13.290 10.990 13.375 11.150 ;
        RECT 15.485 11.115 15.535 11.150 ;
        POLYGON 15.535 11.150 15.570 11.115 15.535 11.115 ;
        RECT 15.485 10.990 15.570 11.115 ;
        RECT 16.190 10.990 16.275 11.150 ;
        RECT 18.385 11.115 18.435 11.150 ;
        POLYGON 18.435 11.150 18.470 11.115 18.435 11.115 ;
        RECT 18.385 10.990 18.470 11.115 ;
        RECT 19.090 10.990 19.175 11.150 ;
        RECT 21.285 11.115 21.335 11.150 ;
        POLYGON 21.335 11.150 21.370 11.115 21.335 11.115 ;
        RECT 21.285 10.990 21.370 11.115 ;
        RECT 21.990 10.990 22.075 11.150 ;
        RECT 24.185 11.115 24.235 11.150 ;
        POLYGON 24.235 11.150 24.270 11.115 24.235 11.115 ;
        RECT 24.185 10.990 24.270 11.115 ;
        RECT 24.890 10.990 24.975 11.150 ;
        RECT 27.085 11.115 27.135 11.150 ;
        POLYGON 27.135 11.150 27.170 11.115 27.135 11.115 ;
        RECT 27.085 10.990 27.170 11.115 ;
        RECT 27.790 10.990 27.875 11.150 ;
        RECT 29.985 11.115 30.035 11.150 ;
        POLYGON 30.035 11.150 30.070 11.115 30.035 11.115 ;
        RECT 29.985 10.990 30.070 11.115 ;
        RECT 30.690 10.990 30.775 11.150 ;
        RECT 32.885 11.115 32.935 11.150 ;
        POLYGON 32.935 11.150 32.970 11.115 32.935 11.115 ;
        RECT 32.885 10.990 32.970 11.115 ;
        RECT 33.590 10.990 33.675 11.150 ;
        RECT 35.785 11.115 35.835 11.150 ;
        POLYGON 35.835 11.150 35.870 11.115 35.835 11.115 ;
        RECT 35.785 10.990 35.870 11.115 ;
        RECT 36.490 10.990 36.575 11.150 ;
        RECT 38.685 11.115 38.735 11.150 ;
        POLYGON 38.735 11.150 38.770 11.115 38.735 11.115 ;
        RECT 38.685 10.990 38.770 11.115 ;
        RECT 39.390 10.990 39.475 11.150 ;
        RECT 41.585 11.115 41.635 11.150 ;
        POLYGON 41.635 11.150 41.670 11.115 41.635 11.115 ;
        RECT 41.585 10.990 41.670 11.115 ;
        RECT 42.290 10.990 42.375 11.150 ;
        RECT 44.485 11.115 44.535 11.150 ;
        POLYGON 44.535 11.150 44.570 11.115 44.535 11.115 ;
        RECT 44.485 10.990 44.570 11.115 ;
        RECT 45.190 10.990 45.275 11.150 ;
        RECT 47.385 11.115 47.435 11.150 ;
        POLYGON 47.435 11.150 47.470 11.115 47.435 11.115 ;
        RECT 47.385 10.990 47.470 11.115 ;
        RECT 48.090 10.990 48.175 11.150 ;
        RECT 50.285 11.115 50.335 11.150 ;
        POLYGON 50.335 11.150 50.370 11.115 50.335 11.115 ;
        RECT 50.285 10.990 50.370 11.115 ;
        RECT 50.990 10.990 51.075 11.150 ;
        RECT 53.185 11.115 53.235 11.150 ;
        POLYGON 53.235 11.150 53.270 11.115 53.235 11.115 ;
        RECT 53.185 10.990 53.270 11.115 ;
        RECT 53.890 10.990 53.975 11.150 ;
        RECT 56.085 11.115 56.135 11.150 ;
        POLYGON 56.135 11.150 56.170 11.115 56.135 11.115 ;
        RECT 56.085 10.990 56.170 11.115 ;
        RECT 56.790 10.990 56.875 11.150 ;
        RECT 58.985 11.115 59.035 11.150 ;
        POLYGON 59.035 11.150 59.070 11.115 59.035 11.115 ;
        RECT 58.985 10.990 59.070 11.115 ;
        RECT 59.690 10.990 59.775 11.150 ;
        RECT 61.885 11.115 61.935 11.150 ;
        POLYGON 61.935 11.150 61.970 11.115 61.935 11.115 ;
        RECT 61.885 10.990 61.970 11.115 ;
        RECT 62.590 10.990 62.675 11.150 ;
        RECT 64.785 11.115 64.835 11.150 ;
        POLYGON 64.835 11.150 64.870 11.115 64.835 11.115 ;
        RECT 64.785 10.990 64.870 11.115 ;
        RECT 65.490 10.990 65.575 11.150 ;
        RECT 67.685 11.115 67.735 11.150 ;
        POLYGON 67.735 11.150 67.770 11.115 67.735 11.115 ;
        RECT 67.685 10.990 67.770 11.115 ;
        RECT 68.390 10.990 68.475 11.150 ;
        RECT 70.585 11.115 70.635 11.150 ;
        POLYGON 70.635 11.150 70.670 11.115 70.635 11.115 ;
        RECT 70.585 10.990 70.670 11.115 ;
        RECT 71.290 10.990 71.375 11.150 ;
        RECT 73.485 11.115 73.535 11.150 ;
        POLYGON 73.535 11.150 73.570 11.115 73.535 11.115 ;
        RECT 73.485 10.990 73.570 11.115 ;
        RECT 74.190 10.990 74.275 11.150 ;
        RECT 76.385 11.115 76.435 11.150 ;
        POLYGON 76.435 11.150 76.470 11.115 76.435 11.115 ;
        RECT 76.385 10.990 76.470 11.115 ;
        RECT 77.090 10.990 77.175 11.150 ;
        RECT 79.285 11.115 79.335 11.150 ;
        POLYGON 79.335 11.150 79.370 11.115 79.335 11.115 ;
        RECT 79.285 10.990 79.370 11.115 ;
        RECT 79.990 10.990 80.075 11.150 ;
        RECT 82.185 11.115 82.235 11.150 ;
        POLYGON 82.235 11.150 82.270 11.115 82.235 11.115 ;
        RECT 82.185 10.990 82.270 11.115 ;
        RECT 82.890 10.990 82.975 11.150 ;
        RECT 85.085 11.115 85.135 11.150 ;
        POLYGON 85.135 11.150 85.170 11.115 85.135 11.115 ;
        RECT 85.085 10.990 85.170 11.115 ;
        RECT 85.790 10.990 85.875 11.150 ;
        RECT 87.985 11.115 88.035 11.150 ;
        POLYGON 88.035 11.150 88.070 11.115 88.035 11.115 ;
        RECT 87.985 10.990 88.070 11.115 ;
        RECT 88.690 10.990 88.775 11.150 ;
        RECT 90.885 11.115 90.935 11.150 ;
        POLYGON 90.935 11.150 90.970 11.115 90.935 11.115 ;
        RECT 90.885 10.990 90.970 11.115 ;
        RECT 91.590 10.990 91.675 11.150 ;
        RECT 0.775 10.370 0.850 10.510 ;
        RECT 0.990 10.320 1.065 10.460 ;
        RECT 1.695 10.380 1.755 10.460 ;
        POLYGON 1.695 10.380 1.755 10.380 1.755 10.320 ;
        RECT 1.910 10.370 1.985 10.510 ;
        RECT 3.675 10.370 3.750 10.510 ;
        RECT 3.890 10.320 3.965 10.460 ;
        RECT 4.595 10.380 4.655 10.460 ;
        POLYGON 4.595 10.380 4.655 10.380 4.655 10.320 ;
        RECT 4.810 10.370 4.885 10.510 ;
        RECT 6.575 10.370 6.650 10.510 ;
        RECT 6.790 10.320 6.865 10.460 ;
        RECT 7.495 10.380 7.555 10.460 ;
        POLYGON 7.495 10.380 7.555 10.380 7.555 10.320 ;
        RECT 7.710 10.370 7.785 10.510 ;
        RECT 9.475 10.370 9.550 10.510 ;
        RECT 9.690 10.320 9.765 10.460 ;
        RECT 10.395 10.380 10.455 10.460 ;
        POLYGON 10.395 10.380 10.455 10.380 10.455 10.320 ;
        RECT 10.610 10.370 10.685 10.510 ;
        RECT 12.375 10.370 12.450 10.510 ;
        RECT 12.590 10.320 12.665 10.460 ;
        RECT 13.295 10.380 13.355 10.460 ;
        POLYGON 13.295 10.380 13.355 10.380 13.355 10.320 ;
        RECT 13.510 10.370 13.585 10.510 ;
        RECT 15.275 10.370 15.350 10.510 ;
        RECT 15.490 10.320 15.565 10.460 ;
        RECT 16.195 10.380 16.255 10.460 ;
        POLYGON 16.195 10.380 16.255 10.380 16.255 10.320 ;
        RECT 16.410 10.370 16.485 10.510 ;
        RECT 18.175 10.370 18.250 10.510 ;
        RECT 18.390 10.320 18.465 10.460 ;
        RECT 19.095 10.380 19.155 10.460 ;
        POLYGON 19.095 10.380 19.155 10.380 19.155 10.320 ;
        RECT 19.310 10.370 19.385 10.510 ;
        RECT 21.075 10.370 21.150 10.510 ;
        RECT 21.290 10.320 21.365 10.460 ;
        RECT 21.995 10.380 22.055 10.460 ;
        POLYGON 21.995 10.380 22.055 10.380 22.055 10.320 ;
        RECT 22.210 10.370 22.285 10.510 ;
        RECT 23.975 10.370 24.050 10.510 ;
        RECT 24.190 10.320 24.265 10.460 ;
        RECT 24.895 10.380 24.955 10.460 ;
        POLYGON 24.895 10.380 24.955 10.380 24.955 10.320 ;
        RECT 25.110 10.370 25.185 10.510 ;
        RECT 26.875 10.370 26.950 10.510 ;
        RECT 27.090 10.320 27.165 10.460 ;
        RECT 27.795 10.380 27.855 10.460 ;
        POLYGON 27.795 10.380 27.855 10.380 27.855 10.320 ;
        RECT 28.010 10.370 28.085 10.510 ;
        RECT 29.775 10.370 29.850 10.510 ;
        RECT 29.990 10.320 30.065 10.460 ;
        RECT 30.695 10.380 30.755 10.460 ;
        POLYGON 30.695 10.380 30.755 10.380 30.755 10.320 ;
        RECT 30.910 10.370 30.985 10.510 ;
        RECT 32.675 10.370 32.750 10.510 ;
        RECT 32.890 10.320 32.965 10.460 ;
        RECT 33.595 10.380 33.655 10.460 ;
        POLYGON 33.595 10.380 33.655 10.380 33.655 10.320 ;
        RECT 33.810 10.370 33.885 10.510 ;
        RECT 35.575 10.370 35.650 10.510 ;
        RECT 35.790 10.320 35.865 10.460 ;
        RECT 36.495 10.380 36.555 10.460 ;
        POLYGON 36.495 10.380 36.555 10.380 36.555 10.320 ;
        RECT 36.710 10.370 36.785 10.510 ;
        RECT 38.475 10.370 38.550 10.510 ;
        RECT 38.690 10.320 38.765 10.460 ;
        RECT 39.395 10.380 39.455 10.460 ;
        POLYGON 39.395 10.380 39.455 10.380 39.455 10.320 ;
        RECT 39.610 10.370 39.685 10.510 ;
        RECT 41.375 10.370 41.450 10.510 ;
        RECT 41.590 10.320 41.665 10.460 ;
        RECT 42.295 10.380 42.355 10.460 ;
        POLYGON 42.295 10.380 42.355 10.380 42.355 10.320 ;
        RECT 42.510 10.370 42.585 10.510 ;
        RECT 44.275 10.370 44.350 10.510 ;
        RECT 44.490 10.320 44.565 10.460 ;
        RECT 45.195 10.380 45.255 10.460 ;
        POLYGON 45.195 10.380 45.255 10.380 45.255 10.320 ;
        RECT 45.410 10.370 45.485 10.510 ;
        RECT 47.175 10.370 47.250 10.510 ;
        RECT 47.390 10.320 47.465 10.460 ;
        RECT 48.095 10.380 48.155 10.460 ;
        POLYGON 48.095 10.380 48.155 10.380 48.155 10.320 ;
        RECT 48.310 10.370 48.385 10.510 ;
        RECT 50.075 10.370 50.150 10.510 ;
        RECT 50.290 10.320 50.365 10.460 ;
        RECT 50.995 10.380 51.055 10.460 ;
        POLYGON 50.995 10.380 51.055 10.380 51.055 10.320 ;
        RECT 51.210 10.370 51.285 10.510 ;
        RECT 52.975 10.370 53.050 10.510 ;
        RECT 53.190 10.320 53.265 10.460 ;
        RECT 53.895 10.380 53.955 10.460 ;
        POLYGON 53.895 10.380 53.955 10.380 53.955 10.320 ;
        RECT 54.110 10.370 54.185 10.510 ;
        RECT 55.875 10.370 55.950 10.510 ;
        RECT 56.090 10.320 56.165 10.460 ;
        RECT 56.795 10.380 56.855 10.460 ;
        POLYGON 56.795 10.380 56.855 10.380 56.855 10.320 ;
        RECT 57.010 10.370 57.085 10.510 ;
        RECT 58.775 10.370 58.850 10.510 ;
        RECT 58.990 10.320 59.065 10.460 ;
        RECT 59.695 10.380 59.755 10.460 ;
        POLYGON 59.695 10.380 59.755 10.380 59.755 10.320 ;
        RECT 59.910 10.370 59.985 10.510 ;
        RECT 61.675 10.370 61.750 10.510 ;
        RECT 61.890 10.320 61.965 10.460 ;
        RECT 62.595 10.380 62.655 10.460 ;
        POLYGON 62.595 10.380 62.655 10.380 62.655 10.320 ;
        RECT 62.810 10.370 62.885 10.510 ;
        RECT 64.575 10.370 64.650 10.510 ;
        RECT 64.790 10.320 64.865 10.460 ;
        RECT 65.495 10.380 65.555 10.460 ;
        POLYGON 65.495 10.380 65.555 10.380 65.555 10.320 ;
        RECT 65.710 10.370 65.785 10.510 ;
        RECT 67.475 10.370 67.550 10.510 ;
        RECT 67.690 10.320 67.765 10.460 ;
        RECT 68.395 10.380 68.455 10.460 ;
        POLYGON 68.395 10.380 68.455 10.380 68.455 10.320 ;
        RECT 68.610 10.370 68.685 10.510 ;
        RECT 70.375 10.370 70.450 10.510 ;
        RECT 70.590 10.320 70.665 10.460 ;
        RECT 71.295 10.380 71.355 10.460 ;
        POLYGON 71.295 10.380 71.355 10.380 71.355 10.320 ;
        RECT 71.510 10.370 71.585 10.510 ;
        RECT 73.275 10.370 73.350 10.510 ;
        RECT 73.490 10.320 73.565 10.460 ;
        RECT 74.195 10.380 74.255 10.460 ;
        POLYGON 74.195 10.380 74.255 10.380 74.255 10.320 ;
        RECT 74.410 10.370 74.485 10.510 ;
        RECT 76.175 10.370 76.250 10.510 ;
        RECT 76.390 10.320 76.465 10.460 ;
        RECT 77.095 10.380 77.155 10.460 ;
        POLYGON 77.095 10.380 77.155 10.380 77.155 10.320 ;
        RECT 77.310 10.370 77.385 10.510 ;
        RECT 79.075 10.370 79.150 10.510 ;
        RECT 79.290 10.320 79.365 10.460 ;
        RECT 79.995 10.380 80.055 10.460 ;
        POLYGON 79.995 10.380 80.055 10.380 80.055 10.320 ;
        RECT 80.210 10.370 80.285 10.510 ;
        RECT 81.975 10.370 82.050 10.510 ;
        RECT 82.190 10.320 82.265 10.460 ;
        RECT 82.895 10.380 82.955 10.460 ;
        POLYGON 82.895 10.380 82.955 10.380 82.955 10.320 ;
        RECT 83.110 10.370 83.185 10.510 ;
        RECT 84.875 10.370 84.950 10.510 ;
        RECT 85.090 10.320 85.165 10.460 ;
        RECT 85.795 10.380 85.855 10.460 ;
        POLYGON 85.795 10.380 85.855 10.380 85.855 10.320 ;
        RECT 86.010 10.370 86.085 10.510 ;
        RECT 87.775 10.370 87.850 10.510 ;
        RECT 87.990 10.320 88.065 10.460 ;
        RECT 88.695 10.380 88.755 10.460 ;
        POLYGON 88.695 10.380 88.755 10.380 88.755 10.320 ;
        RECT 88.910 10.370 88.985 10.510 ;
        RECT 90.675 10.370 90.750 10.510 ;
        RECT 90.890 10.320 90.965 10.460 ;
        RECT 91.595 10.380 91.655 10.460 ;
        POLYGON 91.595 10.380 91.655 10.380 91.655 10.320 ;
        RECT 91.810 10.370 91.885 10.510 ;
        RECT 0.720 9.850 0.870 10.020 ;
        RECT 1.110 9.985 1.260 10.155 ;
        RECT 1.500 9.985 1.650 10.155 ;
        RECT 1.890 9.850 2.040 10.020 ;
        RECT 3.620 9.850 3.770 10.020 ;
        RECT 4.010 9.985 4.160 10.155 ;
        RECT 4.400 9.985 4.550 10.155 ;
        RECT 4.790 9.850 4.940 10.020 ;
        RECT 6.520 9.850 6.670 10.020 ;
        RECT 6.910 9.985 7.060 10.155 ;
        RECT 7.300 9.985 7.450 10.155 ;
        RECT 7.690 9.850 7.840 10.020 ;
        RECT 9.420 9.850 9.570 10.020 ;
        RECT 9.810 9.985 9.960 10.155 ;
        RECT 10.200 9.985 10.350 10.155 ;
        RECT 10.590 9.850 10.740 10.020 ;
        RECT 12.320 9.850 12.470 10.020 ;
        RECT 12.710 9.985 12.860 10.155 ;
        RECT 13.100 9.985 13.250 10.155 ;
        RECT 13.490 9.850 13.640 10.020 ;
        RECT 15.220 9.850 15.370 10.020 ;
        RECT 15.610 9.985 15.760 10.155 ;
        RECT 16.000 9.985 16.150 10.155 ;
        RECT 16.390 9.850 16.540 10.020 ;
        RECT 18.120 9.850 18.270 10.020 ;
        RECT 18.510 9.985 18.660 10.155 ;
        RECT 18.900 9.985 19.050 10.155 ;
        RECT 19.290 9.850 19.440 10.020 ;
        RECT 21.020 9.850 21.170 10.020 ;
        RECT 21.410 9.985 21.560 10.155 ;
        RECT 21.800 9.985 21.950 10.155 ;
        RECT 22.190 9.850 22.340 10.020 ;
        RECT 23.920 9.850 24.070 10.020 ;
        RECT 24.310 9.985 24.460 10.155 ;
        RECT 24.700 9.985 24.850 10.155 ;
        RECT 25.090 9.850 25.240 10.020 ;
        RECT 26.820 9.850 26.970 10.020 ;
        RECT 27.210 9.985 27.360 10.155 ;
        RECT 27.600 9.985 27.750 10.155 ;
        RECT 27.990 9.850 28.140 10.020 ;
        RECT 29.720 9.850 29.870 10.020 ;
        RECT 30.110 9.985 30.260 10.155 ;
        RECT 30.500 9.985 30.650 10.155 ;
        RECT 30.890 9.850 31.040 10.020 ;
        RECT 32.620 9.850 32.770 10.020 ;
        RECT 33.010 9.985 33.160 10.155 ;
        RECT 33.400 9.985 33.550 10.155 ;
        RECT 33.790 9.850 33.940 10.020 ;
        RECT 35.520 9.850 35.670 10.020 ;
        RECT 35.910 9.985 36.060 10.155 ;
        RECT 36.300 9.985 36.450 10.155 ;
        RECT 36.690 9.850 36.840 10.020 ;
        RECT 38.420 9.850 38.570 10.020 ;
        RECT 38.810 9.985 38.960 10.155 ;
        RECT 39.200 9.985 39.350 10.155 ;
        RECT 39.590 9.850 39.740 10.020 ;
        RECT 41.320 9.850 41.470 10.020 ;
        RECT 41.710 9.985 41.860 10.155 ;
        RECT 42.100 9.985 42.250 10.155 ;
        RECT 42.490 9.850 42.640 10.020 ;
        RECT 44.220 9.850 44.370 10.020 ;
        RECT 44.610 9.985 44.760 10.155 ;
        RECT 45.000 9.985 45.150 10.155 ;
        RECT 45.390 9.850 45.540 10.020 ;
        RECT 47.120 9.850 47.270 10.020 ;
        RECT 47.510 9.985 47.660 10.155 ;
        RECT 47.900 9.985 48.050 10.155 ;
        RECT 48.290 9.850 48.440 10.020 ;
        RECT 50.020 9.850 50.170 10.020 ;
        RECT 50.410 9.985 50.560 10.155 ;
        RECT 50.800 9.985 50.950 10.155 ;
        RECT 51.190 9.850 51.340 10.020 ;
        RECT 52.920 9.850 53.070 10.020 ;
        RECT 53.310 9.985 53.460 10.155 ;
        RECT 53.700 9.985 53.850 10.155 ;
        RECT 54.090 9.850 54.240 10.020 ;
        RECT 55.820 9.850 55.970 10.020 ;
        RECT 56.210 9.985 56.360 10.155 ;
        RECT 56.600 9.985 56.750 10.155 ;
        RECT 56.990 9.850 57.140 10.020 ;
        RECT 58.720 9.850 58.870 10.020 ;
        RECT 59.110 9.985 59.260 10.155 ;
        RECT 59.500 9.985 59.650 10.155 ;
        RECT 59.890 9.850 60.040 10.020 ;
        RECT 61.620 9.850 61.770 10.020 ;
        RECT 62.010 9.985 62.160 10.155 ;
        RECT 62.400 9.985 62.550 10.155 ;
        RECT 62.790 9.850 62.940 10.020 ;
        RECT 64.520 9.850 64.670 10.020 ;
        RECT 64.910 9.985 65.060 10.155 ;
        RECT 65.300 9.985 65.450 10.155 ;
        RECT 65.690 9.850 65.840 10.020 ;
        RECT 67.420 9.850 67.570 10.020 ;
        RECT 67.810 9.985 67.960 10.155 ;
        RECT 68.200 9.985 68.350 10.155 ;
        RECT 68.590 9.850 68.740 10.020 ;
        RECT 70.320 9.850 70.470 10.020 ;
        RECT 70.710 9.985 70.860 10.155 ;
        RECT 71.100 9.985 71.250 10.155 ;
        RECT 71.490 9.850 71.640 10.020 ;
        RECT 73.220 9.850 73.370 10.020 ;
        RECT 73.610 9.985 73.760 10.155 ;
        RECT 74.000 9.985 74.150 10.155 ;
        RECT 74.390 9.850 74.540 10.020 ;
        RECT 76.120 9.850 76.270 10.020 ;
        RECT 76.510 9.985 76.660 10.155 ;
        RECT 76.900 9.985 77.050 10.155 ;
        RECT 77.290 9.850 77.440 10.020 ;
        RECT 79.020 9.850 79.170 10.020 ;
        RECT 79.410 9.985 79.560 10.155 ;
        RECT 79.800 9.985 79.950 10.155 ;
        RECT 80.190 9.850 80.340 10.020 ;
        RECT 81.920 9.850 82.070 10.020 ;
        RECT 82.310 9.985 82.460 10.155 ;
        RECT 82.700 9.985 82.850 10.155 ;
        RECT 83.090 9.850 83.240 10.020 ;
        RECT 84.820 9.850 84.970 10.020 ;
        RECT 85.210 9.985 85.360 10.155 ;
        RECT 85.600 9.985 85.750 10.155 ;
        RECT 85.990 9.850 86.140 10.020 ;
        RECT 87.720 9.850 87.870 10.020 ;
        RECT 88.110 9.985 88.260 10.155 ;
        RECT 88.500 9.985 88.650 10.155 ;
        RECT 88.890 9.850 89.040 10.020 ;
        RECT 90.620 9.850 90.770 10.020 ;
        RECT 91.010 9.985 91.160 10.155 ;
        RECT 91.400 9.985 91.550 10.155 ;
        RECT 91.790 9.850 91.940 10.020 ;
        RECT 0.985 9.765 1.035 9.800 ;
        POLYGON 1.035 9.800 1.070 9.765 1.035 9.765 ;
        RECT 0.985 9.640 1.070 9.765 ;
        RECT 1.690 9.640 1.775 9.800 ;
        RECT 3.885 9.765 3.935 9.800 ;
        POLYGON 3.935 9.800 3.970 9.765 3.935 9.765 ;
        RECT 3.885 9.640 3.970 9.765 ;
        RECT 4.590 9.640 4.675 9.800 ;
        RECT 6.785 9.765 6.835 9.800 ;
        POLYGON 6.835 9.800 6.870 9.765 6.835 9.765 ;
        RECT 6.785 9.640 6.870 9.765 ;
        RECT 7.490 9.640 7.575 9.800 ;
        RECT 9.685 9.765 9.735 9.800 ;
        POLYGON 9.735 9.800 9.770 9.765 9.735 9.765 ;
        RECT 9.685 9.640 9.770 9.765 ;
        RECT 10.390 9.640 10.475 9.800 ;
        RECT 12.585 9.765 12.635 9.800 ;
        POLYGON 12.635 9.800 12.670 9.765 12.635 9.765 ;
        RECT 12.585 9.640 12.670 9.765 ;
        RECT 13.290 9.640 13.375 9.800 ;
        RECT 15.485 9.765 15.535 9.800 ;
        POLYGON 15.535 9.800 15.570 9.765 15.535 9.765 ;
        RECT 15.485 9.640 15.570 9.765 ;
        RECT 16.190 9.640 16.275 9.800 ;
        RECT 18.385 9.765 18.435 9.800 ;
        POLYGON 18.435 9.800 18.470 9.765 18.435 9.765 ;
        RECT 18.385 9.640 18.470 9.765 ;
        RECT 19.090 9.640 19.175 9.800 ;
        RECT 21.285 9.765 21.335 9.800 ;
        POLYGON 21.335 9.800 21.370 9.765 21.335 9.765 ;
        RECT 21.285 9.640 21.370 9.765 ;
        RECT 21.990 9.640 22.075 9.800 ;
        RECT 24.185 9.765 24.235 9.800 ;
        POLYGON 24.235 9.800 24.270 9.765 24.235 9.765 ;
        RECT 24.185 9.640 24.270 9.765 ;
        RECT 24.890 9.640 24.975 9.800 ;
        RECT 27.085 9.765 27.135 9.800 ;
        POLYGON 27.135 9.800 27.170 9.765 27.135 9.765 ;
        RECT 27.085 9.640 27.170 9.765 ;
        RECT 27.790 9.640 27.875 9.800 ;
        RECT 29.985 9.765 30.035 9.800 ;
        POLYGON 30.035 9.800 30.070 9.765 30.035 9.765 ;
        RECT 29.985 9.640 30.070 9.765 ;
        RECT 30.690 9.640 30.775 9.800 ;
        RECT 32.885 9.765 32.935 9.800 ;
        POLYGON 32.935 9.800 32.970 9.765 32.935 9.765 ;
        RECT 32.885 9.640 32.970 9.765 ;
        RECT 33.590 9.640 33.675 9.800 ;
        RECT 35.785 9.765 35.835 9.800 ;
        POLYGON 35.835 9.800 35.870 9.765 35.835 9.765 ;
        RECT 35.785 9.640 35.870 9.765 ;
        RECT 36.490 9.640 36.575 9.800 ;
        RECT 38.685 9.765 38.735 9.800 ;
        POLYGON 38.735 9.800 38.770 9.765 38.735 9.765 ;
        RECT 38.685 9.640 38.770 9.765 ;
        RECT 39.390 9.640 39.475 9.800 ;
        RECT 41.585 9.765 41.635 9.800 ;
        POLYGON 41.635 9.800 41.670 9.765 41.635 9.765 ;
        RECT 41.585 9.640 41.670 9.765 ;
        RECT 42.290 9.640 42.375 9.800 ;
        RECT 44.485 9.765 44.535 9.800 ;
        POLYGON 44.535 9.800 44.570 9.765 44.535 9.765 ;
        RECT 44.485 9.640 44.570 9.765 ;
        RECT 45.190 9.640 45.275 9.800 ;
        RECT 47.385 9.765 47.435 9.800 ;
        POLYGON 47.435 9.800 47.470 9.765 47.435 9.765 ;
        RECT 47.385 9.640 47.470 9.765 ;
        RECT 48.090 9.640 48.175 9.800 ;
        RECT 50.285 9.765 50.335 9.800 ;
        POLYGON 50.335 9.800 50.370 9.765 50.335 9.765 ;
        RECT 50.285 9.640 50.370 9.765 ;
        RECT 50.990 9.640 51.075 9.800 ;
        RECT 53.185 9.765 53.235 9.800 ;
        POLYGON 53.235 9.800 53.270 9.765 53.235 9.765 ;
        RECT 53.185 9.640 53.270 9.765 ;
        RECT 53.890 9.640 53.975 9.800 ;
        RECT 56.085 9.765 56.135 9.800 ;
        POLYGON 56.135 9.800 56.170 9.765 56.135 9.765 ;
        RECT 56.085 9.640 56.170 9.765 ;
        RECT 56.790 9.640 56.875 9.800 ;
        RECT 58.985 9.765 59.035 9.800 ;
        POLYGON 59.035 9.800 59.070 9.765 59.035 9.765 ;
        RECT 58.985 9.640 59.070 9.765 ;
        RECT 59.690 9.640 59.775 9.800 ;
        RECT 61.885 9.765 61.935 9.800 ;
        POLYGON 61.935 9.800 61.970 9.765 61.935 9.765 ;
        RECT 61.885 9.640 61.970 9.765 ;
        RECT 62.590 9.640 62.675 9.800 ;
        RECT 64.785 9.765 64.835 9.800 ;
        POLYGON 64.835 9.800 64.870 9.765 64.835 9.765 ;
        RECT 64.785 9.640 64.870 9.765 ;
        RECT 65.490 9.640 65.575 9.800 ;
        RECT 67.685 9.765 67.735 9.800 ;
        POLYGON 67.735 9.800 67.770 9.765 67.735 9.765 ;
        RECT 67.685 9.640 67.770 9.765 ;
        RECT 68.390 9.640 68.475 9.800 ;
        RECT 70.585 9.765 70.635 9.800 ;
        POLYGON 70.635 9.800 70.670 9.765 70.635 9.765 ;
        RECT 70.585 9.640 70.670 9.765 ;
        RECT 71.290 9.640 71.375 9.800 ;
        RECT 73.485 9.765 73.535 9.800 ;
        POLYGON 73.535 9.800 73.570 9.765 73.535 9.765 ;
        RECT 73.485 9.640 73.570 9.765 ;
        RECT 74.190 9.640 74.275 9.800 ;
        RECT 76.385 9.765 76.435 9.800 ;
        POLYGON 76.435 9.800 76.470 9.765 76.435 9.765 ;
        RECT 76.385 9.640 76.470 9.765 ;
        RECT 77.090 9.640 77.175 9.800 ;
        RECT 79.285 9.765 79.335 9.800 ;
        POLYGON 79.335 9.800 79.370 9.765 79.335 9.765 ;
        RECT 79.285 9.640 79.370 9.765 ;
        RECT 79.990 9.640 80.075 9.800 ;
        RECT 82.185 9.765 82.235 9.800 ;
        POLYGON 82.235 9.800 82.270 9.765 82.235 9.765 ;
        RECT 82.185 9.640 82.270 9.765 ;
        RECT 82.890 9.640 82.975 9.800 ;
        RECT 85.085 9.765 85.135 9.800 ;
        POLYGON 85.135 9.800 85.170 9.765 85.135 9.765 ;
        RECT 85.085 9.640 85.170 9.765 ;
        RECT 85.790 9.640 85.875 9.800 ;
        RECT 87.985 9.765 88.035 9.800 ;
        POLYGON 88.035 9.800 88.070 9.765 88.035 9.765 ;
        RECT 87.985 9.640 88.070 9.765 ;
        RECT 88.690 9.640 88.775 9.800 ;
        RECT 90.885 9.765 90.935 9.800 ;
        POLYGON 90.935 9.800 90.970 9.765 90.935 9.765 ;
        RECT 90.885 9.640 90.970 9.765 ;
        RECT 91.590 9.640 91.675 9.800 ;
        RECT 0.775 9.020 0.850 9.160 ;
        RECT 0.990 8.970 1.065 9.110 ;
        RECT 1.695 9.030 1.755 9.110 ;
        POLYGON 1.695 9.030 1.755 9.030 1.755 8.970 ;
        RECT 1.910 9.020 1.985 9.160 ;
        RECT 3.675 9.020 3.750 9.160 ;
        RECT 3.890 8.970 3.965 9.110 ;
        RECT 4.595 9.030 4.655 9.110 ;
        POLYGON 4.595 9.030 4.655 9.030 4.655 8.970 ;
        RECT 4.810 9.020 4.885 9.160 ;
        RECT 6.575 9.020 6.650 9.160 ;
        RECT 6.790 8.970 6.865 9.110 ;
        RECT 7.495 9.030 7.555 9.110 ;
        POLYGON 7.495 9.030 7.555 9.030 7.555 8.970 ;
        RECT 7.710 9.020 7.785 9.160 ;
        RECT 9.475 9.020 9.550 9.160 ;
        RECT 9.690 8.970 9.765 9.110 ;
        RECT 10.395 9.030 10.455 9.110 ;
        POLYGON 10.395 9.030 10.455 9.030 10.455 8.970 ;
        RECT 10.610 9.020 10.685 9.160 ;
        RECT 12.375 9.020 12.450 9.160 ;
        RECT 12.590 8.970 12.665 9.110 ;
        RECT 13.295 9.030 13.355 9.110 ;
        POLYGON 13.295 9.030 13.355 9.030 13.355 8.970 ;
        RECT 13.510 9.020 13.585 9.160 ;
        RECT 15.275 9.020 15.350 9.160 ;
        RECT 15.490 8.970 15.565 9.110 ;
        RECT 16.195 9.030 16.255 9.110 ;
        POLYGON 16.195 9.030 16.255 9.030 16.255 8.970 ;
        RECT 16.410 9.020 16.485 9.160 ;
        RECT 18.175 9.020 18.250 9.160 ;
        RECT 18.390 8.970 18.465 9.110 ;
        RECT 19.095 9.030 19.155 9.110 ;
        POLYGON 19.095 9.030 19.155 9.030 19.155 8.970 ;
        RECT 19.310 9.020 19.385 9.160 ;
        RECT 21.075 9.020 21.150 9.160 ;
        RECT 21.290 8.970 21.365 9.110 ;
        RECT 21.995 9.030 22.055 9.110 ;
        POLYGON 21.995 9.030 22.055 9.030 22.055 8.970 ;
        RECT 22.210 9.020 22.285 9.160 ;
        RECT 23.975 9.020 24.050 9.160 ;
        RECT 24.190 8.970 24.265 9.110 ;
        RECT 24.895 9.030 24.955 9.110 ;
        POLYGON 24.895 9.030 24.955 9.030 24.955 8.970 ;
        RECT 25.110 9.020 25.185 9.160 ;
        RECT 26.875 9.020 26.950 9.160 ;
        RECT 27.090 8.970 27.165 9.110 ;
        RECT 27.795 9.030 27.855 9.110 ;
        POLYGON 27.795 9.030 27.855 9.030 27.855 8.970 ;
        RECT 28.010 9.020 28.085 9.160 ;
        RECT 29.775 9.020 29.850 9.160 ;
        RECT 29.990 8.970 30.065 9.110 ;
        RECT 30.695 9.030 30.755 9.110 ;
        POLYGON 30.695 9.030 30.755 9.030 30.755 8.970 ;
        RECT 30.910 9.020 30.985 9.160 ;
        RECT 32.675 9.020 32.750 9.160 ;
        RECT 32.890 8.970 32.965 9.110 ;
        RECT 33.595 9.030 33.655 9.110 ;
        POLYGON 33.595 9.030 33.655 9.030 33.655 8.970 ;
        RECT 33.810 9.020 33.885 9.160 ;
        RECT 35.575 9.020 35.650 9.160 ;
        RECT 35.790 8.970 35.865 9.110 ;
        RECT 36.495 9.030 36.555 9.110 ;
        POLYGON 36.495 9.030 36.555 9.030 36.555 8.970 ;
        RECT 36.710 9.020 36.785 9.160 ;
        RECT 38.475 9.020 38.550 9.160 ;
        RECT 38.690 8.970 38.765 9.110 ;
        RECT 39.395 9.030 39.455 9.110 ;
        POLYGON 39.395 9.030 39.455 9.030 39.455 8.970 ;
        RECT 39.610 9.020 39.685 9.160 ;
        RECT 41.375 9.020 41.450 9.160 ;
        RECT 41.590 8.970 41.665 9.110 ;
        RECT 42.295 9.030 42.355 9.110 ;
        POLYGON 42.295 9.030 42.355 9.030 42.355 8.970 ;
        RECT 42.510 9.020 42.585 9.160 ;
        RECT 44.275 9.020 44.350 9.160 ;
        RECT 44.490 8.970 44.565 9.110 ;
        RECT 45.195 9.030 45.255 9.110 ;
        POLYGON 45.195 9.030 45.255 9.030 45.255 8.970 ;
        RECT 45.410 9.020 45.485 9.160 ;
        RECT 47.175 9.020 47.250 9.160 ;
        RECT 47.390 8.970 47.465 9.110 ;
        RECT 48.095 9.030 48.155 9.110 ;
        POLYGON 48.095 9.030 48.155 9.030 48.155 8.970 ;
        RECT 48.310 9.020 48.385 9.160 ;
        RECT 50.075 9.020 50.150 9.160 ;
        RECT 50.290 8.970 50.365 9.110 ;
        RECT 50.995 9.030 51.055 9.110 ;
        POLYGON 50.995 9.030 51.055 9.030 51.055 8.970 ;
        RECT 51.210 9.020 51.285 9.160 ;
        RECT 52.975 9.020 53.050 9.160 ;
        RECT 53.190 8.970 53.265 9.110 ;
        RECT 53.895 9.030 53.955 9.110 ;
        POLYGON 53.895 9.030 53.955 9.030 53.955 8.970 ;
        RECT 54.110 9.020 54.185 9.160 ;
        RECT 55.875 9.020 55.950 9.160 ;
        RECT 56.090 8.970 56.165 9.110 ;
        RECT 56.795 9.030 56.855 9.110 ;
        POLYGON 56.795 9.030 56.855 9.030 56.855 8.970 ;
        RECT 57.010 9.020 57.085 9.160 ;
        RECT 58.775 9.020 58.850 9.160 ;
        RECT 58.990 8.970 59.065 9.110 ;
        RECT 59.695 9.030 59.755 9.110 ;
        POLYGON 59.695 9.030 59.755 9.030 59.755 8.970 ;
        RECT 59.910 9.020 59.985 9.160 ;
        RECT 61.675 9.020 61.750 9.160 ;
        RECT 61.890 8.970 61.965 9.110 ;
        RECT 62.595 9.030 62.655 9.110 ;
        POLYGON 62.595 9.030 62.655 9.030 62.655 8.970 ;
        RECT 62.810 9.020 62.885 9.160 ;
        RECT 64.575 9.020 64.650 9.160 ;
        RECT 64.790 8.970 64.865 9.110 ;
        RECT 65.495 9.030 65.555 9.110 ;
        POLYGON 65.495 9.030 65.555 9.030 65.555 8.970 ;
        RECT 65.710 9.020 65.785 9.160 ;
        RECT 67.475 9.020 67.550 9.160 ;
        RECT 67.690 8.970 67.765 9.110 ;
        RECT 68.395 9.030 68.455 9.110 ;
        POLYGON 68.395 9.030 68.455 9.030 68.455 8.970 ;
        RECT 68.610 9.020 68.685 9.160 ;
        RECT 70.375 9.020 70.450 9.160 ;
        RECT 70.590 8.970 70.665 9.110 ;
        RECT 71.295 9.030 71.355 9.110 ;
        POLYGON 71.295 9.030 71.355 9.030 71.355 8.970 ;
        RECT 71.510 9.020 71.585 9.160 ;
        RECT 73.275 9.020 73.350 9.160 ;
        RECT 73.490 8.970 73.565 9.110 ;
        RECT 74.195 9.030 74.255 9.110 ;
        POLYGON 74.195 9.030 74.255 9.030 74.255 8.970 ;
        RECT 74.410 9.020 74.485 9.160 ;
        RECT 76.175 9.020 76.250 9.160 ;
        RECT 76.390 8.970 76.465 9.110 ;
        RECT 77.095 9.030 77.155 9.110 ;
        POLYGON 77.095 9.030 77.155 9.030 77.155 8.970 ;
        RECT 77.310 9.020 77.385 9.160 ;
        RECT 79.075 9.020 79.150 9.160 ;
        RECT 79.290 8.970 79.365 9.110 ;
        RECT 79.995 9.030 80.055 9.110 ;
        POLYGON 79.995 9.030 80.055 9.030 80.055 8.970 ;
        RECT 80.210 9.020 80.285 9.160 ;
        RECT 81.975 9.020 82.050 9.160 ;
        RECT 82.190 8.970 82.265 9.110 ;
        RECT 82.895 9.030 82.955 9.110 ;
        POLYGON 82.895 9.030 82.955 9.030 82.955 8.970 ;
        RECT 83.110 9.020 83.185 9.160 ;
        RECT 84.875 9.020 84.950 9.160 ;
        RECT 85.090 8.970 85.165 9.110 ;
        RECT 85.795 9.030 85.855 9.110 ;
        POLYGON 85.795 9.030 85.855 9.030 85.855 8.970 ;
        RECT 86.010 9.020 86.085 9.160 ;
        RECT 87.775 9.020 87.850 9.160 ;
        RECT 87.990 8.970 88.065 9.110 ;
        RECT 88.695 9.030 88.755 9.110 ;
        POLYGON 88.695 9.030 88.755 9.030 88.755 8.970 ;
        RECT 88.910 9.020 88.985 9.160 ;
        RECT 90.675 9.020 90.750 9.160 ;
        RECT 90.890 8.970 90.965 9.110 ;
        RECT 91.595 9.030 91.655 9.110 ;
        POLYGON 91.595 9.030 91.655 9.030 91.655 8.970 ;
        RECT 91.810 9.020 91.885 9.160 ;
        RECT 0.720 8.500 0.870 8.670 ;
        RECT 1.110 8.635 1.260 8.805 ;
        RECT 1.500 8.635 1.650 8.805 ;
        RECT 1.890 8.500 2.040 8.670 ;
        RECT 3.620 8.500 3.770 8.670 ;
        RECT 4.010 8.635 4.160 8.805 ;
        RECT 4.400 8.635 4.550 8.805 ;
        RECT 4.790 8.500 4.940 8.670 ;
        RECT 6.520 8.500 6.670 8.670 ;
        RECT 6.910 8.635 7.060 8.805 ;
        RECT 7.300 8.635 7.450 8.805 ;
        RECT 7.690 8.500 7.840 8.670 ;
        RECT 9.420 8.500 9.570 8.670 ;
        RECT 9.810 8.635 9.960 8.805 ;
        RECT 10.200 8.635 10.350 8.805 ;
        RECT 10.590 8.500 10.740 8.670 ;
        RECT 12.320 8.500 12.470 8.670 ;
        RECT 12.710 8.635 12.860 8.805 ;
        RECT 13.100 8.635 13.250 8.805 ;
        RECT 13.490 8.500 13.640 8.670 ;
        RECT 15.220 8.500 15.370 8.670 ;
        RECT 15.610 8.635 15.760 8.805 ;
        RECT 16.000 8.635 16.150 8.805 ;
        RECT 16.390 8.500 16.540 8.670 ;
        RECT 18.120 8.500 18.270 8.670 ;
        RECT 18.510 8.635 18.660 8.805 ;
        RECT 18.900 8.635 19.050 8.805 ;
        RECT 19.290 8.500 19.440 8.670 ;
        RECT 21.020 8.500 21.170 8.670 ;
        RECT 21.410 8.635 21.560 8.805 ;
        RECT 21.800 8.635 21.950 8.805 ;
        RECT 22.190 8.500 22.340 8.670 ;
        RECT 23.920 8.500 24.070 8.670 ;
        RECT 24.310 8.635 24.460 8.805 ;
        RECT 24.700 8.635 24.850 8.805 ;
        RECT 25.090 8.500 25.240 8.670 ;
        RECT 26.820 8.500 26.970 8.670 ;
        RECT 27.210 8.635 27.360 8.805 ;
        RECT 27.600 8.635 27.750 8.805 ;
        RECT 27.990 8.500 28.140 8.670 ;
        RECT 29.720 8.500 29.870 8.670 ;
        RECT 30.110 8.635 30.260 8.805 ;
        RECT 30.500 8.635 30.650 8.805 ;
        RECT 30.890 8.500 31.040 8.670 ;
        RECT 32.620 8.500 32.770 8.670 ;
        RECT 33.010 8.635 33.160 8.805 ;
        RECT 33.400 8.635 33.550 8.805 ;
        RECT 33.790 8.500 33.940 8.670 ;
        RECT 35.520 8.500 35.670 8.670 ;
        RECT 35.910 8.635 36.060 8.805 ;
        RECT 36.300 8.635 36.450 8.805 ;
        RECT 36.690 8.500 36.840 8.670 ;
        RECT 38.420 8.500 38.570 8.670 ;
        RECT 38.810 8.635 38.960 8.805 ;
        RECT 39.200 8.635 39.350 8.805 ;
        RECT 39.590 8.500 39.740 8.670 ;
        RECT 41.320 8.500 41.470 8.670 ;
        RECT 41.710 8.635 41.860 8.805 ;
        RECT 42.100 8.635 42.250 8.805 ;
        RECT 42.490 8.500 42.640 8.670 ;
        RECT 44.220 8.500 44.370 8.670 ;
        RECT 44.610 8.635 44.760 8.805 ;
        RECT 45.000 8.635 45.150 8.805 ;
        RECT 45.390 8.500 45.540 8.670 ;
        RECT 47.120 8.500 47.270 8.670 ;
        RECT 47.510 8.635 47.660 8.805 ;
        RECT 47.900 8.635 48.050 8.805 ;
        RECT 48.290 8.500 48.440 8.670 ;
        RECT 50.020 8.500 50.170 8.670 ;
        RECT 50.410 8.635 50.560 8.805 ;
        RECT 50.800 8.635 50.950 8.805 ;
        RECT 51.190 8.500 51.340 8.670 ;
        RECT 52.920 8.500 53.070 8.670 ;
        RECT 53.310 8.635 53.460 8.805 ;
        RECT 53.700 8.635 53.850 8.805 ;
        RECT 54.090 8.500 54.240 8.670 ;
        RECT 55.820 8.500 55.970 8.670 ;
        RECT 56.210 8.635 56.360 8.805 ;
        RECT 56.600 8.635 56.750 8.805 ;
        RECT 56.990 8.500 57.140 8.670 ;
        RECT 58.720 8.500 58.870 8.670 ;
        RECT 59.110 8.635 59.260 8.805 ;
        RECT 59.500 8.635 59.650 8.805 ;
        RECT 59.890 8.500 60.040 8.670 ;
        RECT 61.620 8.500 61.770 8.670 ;
        RECT 62.010 8.635 62.160 8.805 ;
        RECT 62.400 8.635 62.550 8.805 ;
        RECT 62.790 8.500 62.940 8.670 ;
        RECT 64.520 8.500 64.670 8.670 ;
        RECT 64.910 8.635 65.060 8.805 ;
        RECT 65.300 8.635 65.450 8.805 ;
        RECT 65.690 8.500 65.840 8.670 ;
        RECT 67.420 8.500 67.570 8.670 ;
        RECT 67.810 8.635 67.960 8.805 ;
        RECT 68.200 8.635 68.350 8.805 ;
        RECT 68.590 8.500 68.740 8.670 ;
        RECT 70.320 8.500 70.470 8.670 ;
        RECT 70.710 8.635 70.860 8.805 ;
        RECT 71.100 8.635 71.250 8.805 ;
        RECT 71.490 8.500 71.640 8.670 ;
        RECT 73.220 8.500 73.370 8.670 ;
        RECT 73.610 8.635 73.760 8.805 ;
        RECT 74.000 8.635 74.150 8.805 ;
        RECT 74.390 8.500 74.540 8.670 ;
        RECT 76.120 8.500 76.270 8.670 ;
        RECT 76.510 8.635 76.660 8.805 ;
        RECT 76.900 8.635 77.050 8.805 ;
        RECT 77.290 8.500 77.440 8.670 ;
        RECT 79.020 8.500 79.170 8.670 ;
        RECT 79.410 8.635 79.560 8.805 ;
        RECT 79.800 8.635 79.950 8.805 ;
        RECT 80.190 8.500 80.340 8.670 ;
        RECT 81.920 8.500 82.070 8.670 ;
        RECT 82.310 8.635 82.460 8.805 ;
        RECT 82.700 8.635 82.850 8.805 ;
        RECT 83.090 8.500 83.240 8.670 ;
        RECT 84.820 8.500 84.970 8.670 ;
        RECT 85.210 8.635 85.360 8.805 ;
        RECT 85.600 8.635 85.750 8.805 ;
        RECT 85.990 8.500 86.140 8.670 ;
        RECT 87.720 8.500 87.870 8.670 ;
        RECT 88.110 8.635 88.260 8.805 ;
        RECT 88.500 8.635 88.650 8.805 ;
        RECT 88.890 8.500 89.040 8.670 ;
        RECT 90.620 8.500 90.770 8.670 ;
        RECT 91.010 8.635 91.160 8.805 ;
        RECT 91.400 8.635 91.550 8.805 ;
        RECT 91.790 8.500 91.940 8.670 ;
        RECT 0.985 8.415 1.035 8.450 ;
        POLYGON 1.035 8.450 1.070 8.415 1.035 8.415 ;
        RECT 0.985 8.290 1.070 8.415 ;
        RECT 1.690 8.290 1.775 8.450 ;
        RECT 3.885 8.415 3.935 8.450 ;
        POLYGON 3.935 8.450 3.970 8.415 3.935 8.415 ;
        RECT 3.885 8.290 3.970 8.415 ;
        RECT 4.590 8.290 4.675 8.450 ;
        RECT 6.785 8.415 6.835 8.450 ;
        POLYGON 6.835 8.450 6.870 8.415 6.835 8.415 ;
        RECT 6.785 8.290 6.870 8.415 ;
        RECT 7.490 8.290 7.575 8.450 ;
        RECT 9.685 8.415 9.735 8.450 ;
        POLYGON 9.735 8.450 9.770 8.415 9.735 8.415 ;
        RECT 9.685 8.290 9.770 8.415 ;
        RECT 10.390 8.290 10.475 8.450 ;
        RECT 12.585 8.415 12.635 8.450 ;
        POLYGON 12.635 8.450 12.670 8.415 12.635 8.415 ;
        RECT 12.585 8.290 12.670 8.415 ;
        RECT 13.290 8.290 13.375 8.450 ;
        RECT 15.485 8.415 15.535 8.450 ;
        POLYGON 15.535 8.450 15.570 8.415 15.535 8.415 ;
        RECT 15.485 8.290 15.570 8.415 ;
        RECT 16.190 8.290 16.275 8.450 ;
        RECT 18.385 8.415 18.435 8.450 ;
        POLYGON 18.435 8.450 18.470 8.415 18.435 8.415 ;
        RECT 18.385 8.290 18.470 8.415 ;
        RECT 19.090 8.290 19.175 8.450 ;
        RECT 21.285 8.415 21.335 8.450 ;
        POLYGON 21.335 8.450 21.370 8.415 21.335 8.415 ;
        RECT 21.285 8.290 21.370 8.415 ;
        RECT 21.990 8.290 22.075 8.450 ;
        RECT 24.185 8.415 24.235 8.450 ;
        POLYGON 24.235 8.450 24.270 8.415 24.235 8.415 ;
        RECT 24.185 8.290 24.270 8.415 ;
        RECT 24.890 8.290 24.975 8.450 ;
        RECT 27.085 8.415 27.135 8.450 ;
        POLYGON 27.135 8.450 27.170 8.415 27.135 8.415 ;
        RECT 27.085 8.290 27.170 8.415 ;
        RECT 27.790 8.290 27.875 8.450 ;
        RECT 29.985 8.415 30.035 8.450 ;
        POLYGON 30.035 8.450 30.070 8.415 30.035 8.415 ;
        RECT 29.985 8.290 30.070 8.415 ;
        RECT 30.690 8.290 30.775 8.450 ;
        RECT 32.885 8.415 32.935 8.450 ;
        POLYGON 32.935 8.450 32.970 8.415 32.935 8.415 ;
        RECT 32.885 8.290 32.970 8.415 ;
        RECT 33.590 8.290 33.675 8.450 ;
        RECT 35.785 8.415 35.835 8.450 ;
        POLYGON 35.835 8.450 35.870 8.415 35.835 8.415 ;
        RECT 35.785 8.290 35.870 8.415 ;
        RECT 36.490 8.290 36.575 8.450 ;
        RECT 38.685 8.415 38.735 8.450 ;
        POLYGON 38.735 8.450 38.770 8.415 38.735 8.415 ;
        RECT 38.685 8.290 38.770 8.415 ;
        RECT 39.390 8.290 39.475 8.450 ;
        RECT 41.585 8.415 41.635 8.450 ;
        POLYGON 41.635 8.450 41.670 8.415 41.635 8.415 ;
        RECT 41.585 8.290 41.670 8.415 ;
        RECT 42.290 8.290 42.375 8.450 ;
        RECT 44.485 8.415 44.535 8.450 ;
        POLYGON 44.535 8.450 44.570 8.415 44.535 8.415 ;
        RECT 44.485 8.290 44.570 8.415 ;
        RECT 45.190 8.290 45.275 8.450 ;
        RECT 47.385 8.415 47.435 8.450 ;
        POLYGON 47.435 8.450 47.470 8.415 47.435 8.415 ;
        RECT 47.385 8.290 47.470 8.415 ;
        RECT 48.090 8.290 48.175 8.450 ;
        RECT 50.285 8.415 50.335 8.450 ;
        POLYGON 50.335 8.450 50.370 8.415 50.335 8.415 ;
        RECT 50.285 8.290 50.370 8.415 ;
        RECT 50.990 8.290 51.075 8.450 ;
        RECT 53.185 8.415 53.235 8.450 ;
        POLYGON 53.235 8.450 53.270 8.415 53.235 8.415 ;
        RECT 53.185 8.290 53.270 8.415 ;
        RECT 53.890 8.290 53.975 8.450 ;
        RECT 56.085 8.415 56.135 8.450 ;
        POLYGON 56.135 8.450 56.170 8.415 56.135 8.415 ;
        RECT 56.085 8.290 56.170 8.415 ;
        RECT 56.790 8.290 56.875 8.450 ;
        RECT 58.985 8.415 59.035 8.450 ;
        POLYGON 59.035 8.450 59.070 8.415 59.035 8.415 ;
        RECT 58.985 8.290 59.070 8.415 ;
        RECT 59.690 8.290 59.775 8.450 ;
        RECT 61.885 8.415 61.935 8.450 ;
        POLYGON 61.935 8.450 61.970 8.415 61.935 8.415 ;
        RECT 61.885 8.290 61.970 8.415 ;
        RECT 62.590 8.290 62.675 8.450 ;
        RECT 64.785 8.415 64.835 8.450 ;
        POLYGON 64.835 8.450 64.870 8.415 64.835 8.415 ;
        RECT 64.785 8.290 64.870 8.415 ;
        RECT 65.490 8.290 65.575 8.450 ;
        RECT 67.685 8.415 67.735 8.450 ;
        POLYGON 67.735 8.450 67.770 8.415 67.735 8.415 ;
        RECT 67.685 8.290 67.770 8.415 ;
        RECT 68.390 8.290 68.475 8.450 ;
        RECT 70.585 8.415 70.635 8.450 ;
        POLYGON 70.635 8.450 70.670 8.415 70.635 8.415 ;
        RECT 70.585 8.290 70.670 8.415 ;
        RECT 71.290 8.290 71.375 8.450 ;
        RECT 73.485 8.415 73.535 8.450 ;
        POLYGON 73.535 8.450 73.570 8.415 73.535 8.415 ;
        RECT 73.485 8.290 73.570 8.415 ;
        RECT 74.190 8.290 74.275 8.450 ;
        RECT 76.385 8.415 76.435 8.450 ;
        POLYGON 76.435 8.450 76.470 8.415 76.435 8.415 ;
        RECT 76.385 8.290 76.470 8.415 ;
        RECT 77.090 8.290 77.175 8.450 ;
        RECT 79.285 8.415 79.335 8.450 ;
        POLYGON 79.335 8.450 79.370 8.415 79.335 8.415 ;
        RECT 79.285 8.290 79.370 8.415 ;
        RECT 79.990 8.290 80.075 8.450 ;
        RECT 82.185 8.415 82.235 8.450 ;
        POLYGON 82.235 8.450 82.270 8.415 82.235 8.415 ;
        RECT 82.185 8.290 82.270 8.415 ;
        RECT 82.890 8.290 82.975 8.450 ;
        RECT 85.085 8.415 85.135 8.450 ;
        POLYGON 85.135 8.450 85.170 8.415 85.135 8.415 ;
        RECT 85.085 8.290 85.170 8.415 ;
        RECT 85.790 8.290 85.875 8.450 ;
        RECT 87.985 8.415 88.035 8.450 ;
        POLYGON 88.035 8.450 88.070 8.415 88.035 8.415 ;
        RECT 87.985 8.290 88.070 8.415 ;
        RECT 88.690 8.290 88.775 8.450 ;
        RECT 90.885 8.415 90.935 8.450 ;
        POLYGON 90.935 8.450 90.970 8.415 90.935 8.415 ;
        RECT 90.885 8.290 90.970 8.415 ;
        RECT 91.590 8.290 91.675 8.450 ;
        RECT 0.775 7.670 0.850 7.810 ;
        RECT 0.990 7.620 1.065 7.760 ;
        RECT 1.695 7.680 1.755 7.760 ;
        POLYGON 1.695 7.680 1.755 7.680 1.755 7.620 ;
        RECT 1.910 7.670 1.985 7.810 ;
        RECT 3.675 7.670 3.750 7.810 ;
        RECT 3.890 7.620 3.965 7.760 ;
        RECT 4.595 7.680 4.655 7.760 ;
        POLYGON 4.595 7.680 4.655 7.680 4.655 7.620 ;
        RECT 4.810 7.670 4.885 7.810 ;
        RECT 6.575 7.670 6.650 7.810 ;
        RECT 6.790 7.620 6.865 7.760 ;
        RECT 7.495 7.680 7.555 7.760 ;
        POLYGON 7.495 7.680 7.555 7.680 7.555 7.620 ;
        RECT 7.710 7.670 7.785 7.810 ;
        RECT 9.475 7.670 9.550 7.810 ;
        RECT 9.690 7.620 9.765 7.760 ;
        RECT 10.395 7.680 10.455 7.760 ;
        POLYGON 10.395 7.680 10.455 7.680 10.455 7.620 ;
        RECT 10.610 7.670 10.685 7.810 ;
        RECT 12.375 7.670 12.450 7.810 ;
        RECT 12.590 7.620 12.665 7.760 ;
        RECT 13.295 7.680 13.355 7.760 ;
        POLYGON 13.295 7.680 13.355 7.680 13.355 7.620 ;
        RECT 13.510 7.670 13.585 7.810 ;
        RECT 15.275 7.670 15.350 7.810 ;
        RECT 15.490 7.620 15.565 7.760 ;
        RECT 16.195 7.680 16.255 7.760 ;
        POLYGON 16.195 7.680 16.255 7.680 16.255 7.620 ;
        RECT 16.410 7.670 16.485 7.810 ;
        RECT 18.175 7.670 18.250 7.810 ;
        RECT 18.390 7.620 18.465 7.760 ;
        RECT 19.095 7.680 19.155 7.760 ;
        POLYGON 19.095 7.680 19.155 7.680 19.155 7.620 ;
        RECT 19.310 7.670 19.385 7.810 ;
        RECT 21.075 7.670 21.150 7.810 ;
        RECT 21.290 7.620 21.365 7.760 ;
        RECT 21.995 7.680 22.055 7.760 ;
        POLYGON 21.995 7.680 22.055 7.680 22.055 7.620 ;
        RECT 22.210 7.670 22.285 7.810 ;
        RECT 23.975 7.670 24.050 7.810 ;
        RECT 24.190 7.620 24.265 7.760 ;
        RECT 24.895 7.680 24.955 7.760 ;
        POLYGON 24.895 7.680 24.955 7.680 24.955 7.620 ;
        RECT 25.110 7.670 25.185 7.810 ;
        RECT 26.875 7.670 26.950 7.810 ;
        RECT 27.090 7.620 27.165 7.760 ;
        RECT 27.795 7.680 27.855 7.760 ;
        POLYGON 27.795 7.680 27.855 7.680 27.855 7.620 ;
        RECT 28.010 7.670 28.085 7.810 ;
        RECT 29.775 7.670 29.850 7.810 ;
        RECT 29.990 7.620 30.065 7.760 ;
        RECT 30.695 7.680 30.755 7.760 ;
        POLYGON 30.695 7.680 30.755 7.680 30.755 7.620 ;
        RECT 30.910 7.670 30.985 7.810 ;
        RECT 32.675 7.670 32.750 7.810 ;
        RECT 32.890 7.620 32.965 7.760 ;
        RECT 33.595 7.680 33.655 7.760 ;
        POLYGON 33.595 7.680 33.655 7.680 33.655 7.620 ;
        RECT 33.810 7.670 33.885 7.810 ;
        RECT 35.575 7.670 35.650 7.810 ;
        RECT 35.790 7.620 35.865 7.760 ;
        RECT 36.495 7.680 36.555 7.760 ;
        POLYGON 36.495 7.680 36.555 7.680 36.555 7.620 ;
        RECT 36.710 7.670 36.785 7.810 ;
        RECT 38.475 7.670 38.550 7.810 ;
        RECT 38.690 7.620 38.765 7.760 ;
        RECT 39.395 7.680 39.455 7.760 ;
        POLYGON 39.395 7.680 39.455 7.680 39.455 7.620 ;
        RECT 39.610 7.670 39.685 7.810 ;
        RECT 41.375 7.670 41.450 7.810 ;
        RECT 41.590 7.620 41.665 7.760 ;
        RECT 42.295 7.680 42.355 7.760 ;
        POLYGON 42.295 7.680 42.355 7.680 42.355 7.620 ;
        RECT 42.510 7.670 42.585 7.810 ;
        RECT 44.275 7.670 44.350 7.810 ;
        RECT 44.490 7.620 44.565 7.760 ;
        RECT 45.195 7.680 45.255 7.760 ;
        POLYGON 45.195 7.680 45.255 7.680 45.255 7.620 ;
        RECT 45.410 7.670 45.485 7.810 ;
        RECT 47.175 7.670 47.250 7.810 ;
        RECT 47.390 7.620 47.465 7.760 ;
        RECT 48.095 7.680 48.155 7.760 ;
        POLYGON 48.095 7.680 48.155 7.680 48.155 7.620 ;
        RECT 48.310 7.670 48.385 7.810 ;
        RECT 50.075 7.670 50.150 7.810 ;
        RECT 50.290 7.620 50.365 7.760 ;
        RECT 50.995 7.680 51.055 7.760 ;
        POLYGON 50.995 7.680 51.055 7.680 51.055 7.620 ;
        RECT 51.210 7.670 51.285 7.810 ;
        RECT 52.975 7.670 53.050 7.810 ;
        RECT 53.190 7.620 53.265 7.760 ;
        RECT 53.895 7.680 53.955 7.760 ;
        POLYGON 53.895 7.680 53.955 7.680 53.955 7.620 ;
        RECT 54.110 7.670 54.185 7.810 ;
        RECT 55.875 7.670 55.950 7.810 ;
        RECT 56.090 7.620 56.165 7.760 ;
        RECT 56.795 7.680 56.855 7.760 ;
        POLYGON 56.795 7.680 56.855 7.680 56.855 7.620 ;
        RECT 57.010 7.670 57.085 7.810 ;
        RECT 58.775 7.670 58.850 7.810 ;
        RECT 58.990 7.620 59.065 7.760 ;
        RECT 59.695 7.680 59.755 7.760 ;
        POLYGON 59.695 7.680 59.755 7.680 59.755 7.620 ;
        RECT 59.910 7.670 59.985 7.810 ;
        RECT 61.675 7.670 61.750 7.810 ;
        RECT 61.890 7.620 61.965 7.760 ;
        RECT 62.595 7.680 62.655 7.760 ;
        POLYGON 62.595 7.680 62.655 7.680 62.655 7.620 ;
        RECT 62.810 7.670 62.885 7.810 ;
        RECT 64.575 7.670 64.650 7.810 ;
        RECT 64.790 7.620 64.865 7.760 ;
        RECT 65.495 7.680 65.555 7.760 ;
        POLYGON 65.495 7.680 65.555 7.680 65.555 7.620 ;
        RECT 65.710 7.670 65.785 7.810 ;
        RECT 67.475 7.670 67.550 7.810 ;
        RECT 67.690 7.620 67.765 7.760 ;
        RECT 68.395 7.680 68.455 7.760 ;
        POLYGON 68.395 7.680 68.455 7.680 68.455 7.620 ;
        RECT 68.610 7.670 68.685 7.810 ;
        RECT 70.375 7.670 70.450 7.810 ;
        RECT 70.590 7.620 70.665 7.760 ;
        RECT 71.295 7.680 71.355 7.760 ;
        POLYGON 71.295 7.680 71.355 7.680 71.355 7.620 ;
        RECT 71.510 7.670 71.585 7.810 ;
        RECT 73.275 7.670 73.350 7.810 ;
        RECT 73.490 7.620 73.565 7.760 ;
        RECT 74.195 7.680 74.255 7.760 ;
        POLYGON 74.195 7.680 74.255 7.680 74.255 7.620 ;
        RECT 74.410 7.670 74.485 7.810 ;
        RECT 76.175 7.670 76.250 7.810 ;
        RECT 76.390 7.620 76.465 7.760 ;
        RECT 77.095 7.680 77.155 7.760 ;
        POLYGON 77.095 7.680 77.155 7.680 77.155 7.620 ;
        RECT 77.310 7.670 77.385 7.810 ;
        RECT 79.075 7.670 79.150 7.810 ;
        RECT 79.290 7.620 79.365 7.760 ;
        RECT 79.995 7.680 80.055 7.760 ;
        POLYGON 79.995 7.680 80.055 7.680 80.055 7.620 ;
        RECT 80.210 7.670 80.285 7.810 ;
        RECT 81.975 7.670 82.050 7.810 ;
        RECT 82.190 7.620 82.265 7.760 ;
        RECT 82.895 7.680 82.955 7.760 ;
        POLYGON 82.895 7.680 82.955 7.680 82.955 7.620 ;
        RECT 83.110 7.670 83.185 7.810 ;
        RECT 84.875 7.670 84.950 7.810 ;
        RECT 85.090 7.620 85.165 7.760 ;
        RECT 85.795 7.680 85.855 7.760 ;
        POLYGON 85.795 7.680 85.855 7.680 85.855 7.620 ;
        RECT 86.010 7.670 86.085 7.810 ;
        RECT 87.775 7.670 87.850 7.810 ;
        RECT 87.990 7.620 88.065 7.760 ;
        RECT 88.695 7.680 88.755 7.760 ;
        POLYGON 88.695 7.680 88.755 7.680 88.755 7.620 ;
        RECT 88.910 7.670 88.985 7.810 ;
        RECT 90.675 7.670 90.750 7.810 ;
        RECT 90.890 7.620 90.965 7.760 ;
        RECT 91.595 7.680 91.655 7.760 ;
        POLYGON 91.595 7.680 91.655 7.680 91.655 7.620 ;
        RECT 91.810 7.670 91.885 7.810 ;
        RECT 0.720 7.150 0.870 7.320 ;
        RECT 1.110 7.285 1.260 7.455 ;
        RECT 1.500 7.285 1.650 7.455 ;
        RECT 1.890 7.150 2.040 7.320 ;
        RECT 3.620 7.150 3.770 7.320 ;
        RECT 4.010 7.285 4.160 7.455 ;
        RECT 4.400 7.285 4.550 7.455 ;
        RECT 4.790 7.150 4.940 7.320 ;
        RECT 6.520 7.150 6.670 7.320 ;
        RECT 6.910 7.285 7.060 7.455 ;
        RECT 7.300 7.285 7.450 7.455 ;
        RECT 7.690 7.150 7.840 7.320 ;
        RECT 9.420 7.150 9.570 7.320 ;
        RECT 9.810 7.285 9.960 7.455 ;
        RECT 10.200 7.285 10.350 7.455 ;
        RECT 10.590 7.150 10.740 7.320 ;
        RECT 12.320 7.150 12.470 7.320 ;
        RECT 12.710 7.285 12.860 7.455 ;
        RECT 13.100 7.285 13.250 7.455 ;
        RECT 13.490 7.150 13.640 7.320 ;
        RECT 15.220 7.150 15.370 7.320 ;
        RECT 15.610 7.285 15.760 7.455 ;
        RECT 16.000 7.285 16.150 7.455 ;
        RECT 16.390 7.150 16.540 7.320 ;
        RECT 18.120 7.150 18.270 7.320 ;
        RECT 18.510 7.285 18.660 7.455 ;
        RECT 18.900 7.285 19.050 7.455 ;
        RECT 19.290 7.150 19.440 7.320 ;
        RECT 21.020 7.150 21.170 7.320 ;
        RECT 21.410 7.285 21.560 7.455 ;
        RECT 21.800 7.285 21.950 7.455 ;
        RECT 22.190 7.150 22.340 7.320 ;
        RECT 23.920 7.150 24.070 7.320 ;
        RECT 24.310 7.285 24.460 7.455 ;
        RECT 24.700 7.285 24.850 7.455 ;
        RECT 25.090 7.150 25.240 7.320 ;
        RECT 26.820 7.150 26.970 7.320 ;
        RECT 27.210 7.285 27.360 7.455 ;
        RECT 27.600 7.285 27.750 7.455 ;
        RECT 27.990 7.150 28.140 7.320 ;
        RECT 29.720 7.150 29.870 7.320 ;
        RECT 30.110 7.285 30.260 7.455 ;
        RECT 30.500 7.285 30.650 7.455 ;
        RECT 30.890 7.150 31.040 7.320 ;
        RECT 32.620 7.150 32.770 7.320 ;
        RECT 33.010 7.285 33.160 7.455 ;
        RECT 33.400 7.285 33.550 7.455 ;
        RECT 33.790 7.150 33.940 7.320 ;
        RECT 35.520 7.150 35.670 7.320 ;
        RECT 35.910 7.285 36.060 7.455 ;
        RECT 36.300 7.285 36.450 7.455 ;
        RECT 36.690 7.150 36.840 7.320 ;
        RECT 38.420 7.150 38.570 7.320 ;
        RECT 38.810 7.285 38.960 7.455 ;
        RECT 39.200 7.285 39.350 7.455 ;
        RECT 39.590 7.150 39.740 7.320 ;
        RECT 41.320 7.150 41.470 7.320 ;
        RECT 41.710 7.285 41.860 7.455 ;
        RECT 42.100 7.285 42.250 7.455 ;
        RECT 42.490 7.150 42.640 7.320 ;
        RECT 44.220 7.150 44.370 7.320 ;
        RECT 44.610 7.285 44.760 7.455 ;
        RECT 45.000 7.285 45.150 7.455 ;
        RECT 45.390 7.150 45.540 7.320 ;
        RECT 47.120 7.150 47.270 7.320 ;
        RECT 47.510 7.285 47.660 7.455 ;
        RECT 47.900 7.285 48.050 7.455 ;
        RECT 48.290 7.150 48.440 7.320 ;
        RECT 50.020 7.150 50.170 7.320 ;
        RECT 50.410 7.285 50.560 7.455 ;
        RECT 50.800 7.285 50.950 7.455 ;
        RECT 51.190 7.150 51.340 7.320 ;
        RECT 52.920 7.150 53.070 7.320 ;
        RECT 53.310 7.285 53.460 7.455 ;
        RECT 53.700 7.285 53.850 7.455 ;
        RECT 54.090 7.150 54.240 7.320 ;
        RECT 55.820 7.150 55.970 7.320 ;
        RECT 56.210 7.285 56.360 7.455 ;
        RECT 56.600 7.285 56.750 7.455 ;
        RECT 56.990 7.150 57.140 7.320 ;
        RECT 58.720 7.150 58.870 7.320 ;
        RECT 59.110 7.285 59.260 7.455 ;
        RECT 59.500 7.285 59.650 7.455 ;
        RECT 59.890 7.150 60.040 7.320 ;
        RECT 61.620 7.150 61.770 7.320 ;
        RECT 62.010 7.285 62.160 7.455 ;
        RECT 62.400 7.285 62.550 7.455 ;
        RECT 62.790 7.150 62.940 7.320 ;
        RECT 64.520 7.150 64.670 7.320 ;
        RECT 64.910 7.285 65.060 7.455 ;
        RECT 65.300 7.285 65.450 7.455 ;
        RECT 65.690 7.150 65.840 7.320 ;
        RECT 67.420 7.150 67.570 7.320 ;
        RECT 67.810 7.285 67.960 7.455 ;
        RECT 68.200 7.285 68.350 7.455 ;
        RECT 68.590 7.150 68.740 7.320 ;
        RECT 70.320 7.150 70.470 7.320 ;
        RECT 70.710 7.285 70.860 7.455 ;
        RECT 71.100 7.285 71.250 7.455 ;
        RECT 71.490 7.150 71.640 7.320 ;
        RECT 73.220 7.150 73.370 7.320 ;
        RECT 73.610 7.285 73.760 7.455 ;
        RECT 74.000 7.285 74.150 7.455 ;
        RECT 74.390 7.150 74.540 7.320 ;
        RECT 76.120 7.150 76.270 7.320 ;
        RECT 76.510 7.285 76.660 7.455 ;
        RECT 76.900 7.285 77.050 7.455 ;
        RECT 77.290 7.150 77.440 7.320 ;
        RECT 79.020 7.150 79.170 7.320 ;
        RECT 79.410 7.285 79.560 7.455 ;
        RECT 79.800 7.285 79.950 7.455 ;
        RECT 80.190 7.150 80.340 7.320 ;
        RECT 81.920 7.150 82.070 7.320 ;
        RECT 82.310 7.285 82.460 7.455 ;
        RECT 82.700 7.285 82.850 7.455 ;
        RECT 83.090 7.150 83.240 7.320 ;
        RECT 84.820 7.150 84.970 7.320 ;
        RECT 85.210 7.285 85.360 7.455 ;
        RECT 85.600 7.285 85.750 7.455 ;
        RECT 85.990 7.150 86.140 7.320 ;
        RECT 87.720 7.150 87.870 7.320 ;
        RECT 88.110 7.285 88.260 7.455 ;
        RECT 88.500 7.285 88.650 7.455 ;
        RECT 88.890 7.150 89.040 7.320 ;
        RECT 90.620 7.150 90.770 7.320 ;
        RECT 91.010 7.285 91.160 7.455 ;
        RECT 91.400 7.285 91.550 7.455 ;
        RECT 91.790 7.150 91.940 7.320 ;
        RECT 0.985 7.065 1.035 7.100 ;
        POLYGON 1.035 7.100 1.070 7.065 1.035 7.065 ;
        RECT 0.985 6.940 1.070 7.065 ;
        RECT 1.690 6.940 1.775 7.100 ;
        RECT 3.885 7.065 3.935 7.100 ;
        POLYGON 3.935 7.100 3.970 7.065 3.935 7.065 ;
        RECT 3.885 6.940 3.970 7.065 ;
        RECT 4.590 6.940 4.675 7.100 ;
        RECT 6.785 7.065 6.835 7.100 ;
        POLYGON 6.835 7.100 6.870 7.065 6.835 7.065 ;
        RECT 6.785 6.940 6.870 7.065 ;
        RECT 7.490 6.940 7.575 7.100 ;
        RECT 9.685 7.065 9.735 7.100 ;
        POLYGON 9.735 7.100 9.770 7.065 9.735 7.065 ;
        RECT 9.685 6.940 9.770 7.065 ;
        RECT 10.390 6.940 10.475 7.100 ;
        RECT 12.585 7.065 12.635 7.100 ;
        POLYGON 12.635 7.100 12.670 7.065 12.635 7.065 ;
        RECT 12.585 6.940 12.670 7.065 ;
        RECT 13.290 6.940 13.375 7.100 ;
        RECT 15.485 7.065 15.535 7.100 ;
        POLYGON 15.535 7.100 15.570 7.065 15.535 7.065 ;
        RECT 15.485 6.940 15.570 7.065 ;
        RECT 16.190 6.940 16.275 7.100 ;
        RECT 18.385 7.065 18.435 7.100 ;
        POLYGON 18.435 7.100 18.470 7.065 18.435 7.065 ;
        RECT 18.385 6.940 18.470 7.065 ;
        RECT 19.090 6.940 19.175 7.100 ;
        RECT 21.285 7.065 21.335 7.100 ;
        POLYGON 21.335 7.100 21.370 7.065 21.335 7.065 ;
        RECT 21.285 6.940 21.370 7.065 ;
        RECT 21.990 6.940 22.075 7.100 ;
        RECT 24.185 7.065 24.235 7.100 ;
        POLYGON 24.235 7.100 24.270 7.065 24.235 7.065 ;
        RECT 24.185 6.940 24.270 7.065 ;
        RECT 24.890 6.940 24.975 7.100 ;
        RECT 27.085 7.065 27.135 7.100 ;
        POLYGON 27.135 7.100 27.170 7.065 27.135 7.065 ;
        RECT 27.085 6.940 27.170 7.065 ;
        RECT 27.790 6.940 27.875 7.100 ;
        RECT 29.985 7.065 30.035 7.100 ;
        POLYGON 30.035 7.100 30.070 7.065 30.035 7.065 ;
        RECT 29.985 6.940 30.070 7.065 ;
        RECT 30.690 6.940 30.775 7.100 ;
        RECT 32.885 7.065 32.935 7.100 ;
        POLYGON 32.935 7.100 32.970 7.065 32.935 7.065 ;
        RECT 32.885 6.940 32.970 7.065 ;
        RECT 33.590 6.940 33.675 7.100 ;
        RECT 35.785 7.065 35.835 7.100 ;
        POLYGON 35.835 7.100 35.870 7.065 35.835 7.065 ;
        RECT 35.785 6.940 35.870 7.065 ;
        RECT 36.490 6.940 36.575 7.100 ;
        RECT 38.685 7.065 38.735 7.100 ;
        POLYGON 38.735 7.100 38.770 7.065 38.735 7.065 ;
        RECT 38.685 6.940 38.770 7.065 ;
        RECT 39.390 6.940 39.475 7.100 ;
        RECT 41.585 7.065 41.635 7.100 ;
        POLYGON 41.635 7.100 41.670 7.065 41.635 7.065 ;
        RECT 41.585 6.940 41.670 7.065 ;
        RECT 42.290 6.940 42.375 7.100 ;
        RECT 44.485 7.065 44.535 7.100 ;
        POLYGON 44.535 7.100 44.570 7.065 44.535 7.065 ;
        RECT 44.485 6.940 44.570 7.065 ;
        RECT 45.190 6.940 45.275 7.100 ;
        RECT 47.385 7.065 47.435 7.100 ;
        POLYGON 47.435 7.100 47.470 7.065 47.435 7.065 ;
        RECT 47.385 6.940 47.470 7.065 ;
        RECT 48.090 6.940 48.175 7.100 ;
        RECT 50.285 7.065 50.335 7.100 ;
        POLYGON 50.335 7.100 50.370 7.065 50.335 7.065 ;
        RECT 50.285 6.940 50.370 7.065 ;
        RECT 50.990 6.940 51.075 7.100 ;
        RECT 53.185 7.065 53.235 7.100 ;
        POLYGON 53.235 7.100 53.270 7.065 53.235 7.065 ;
        RECT 53.185 6.940 53.270 7.065 ;
        RECT 53.890 6.940 53.975 7.100 ;
        RECT 56.085 7.065 56.135 7.100 ;
        POLYGON 56.135 7.100 56.170 7.065 56.135 7.065 ;
        RECT 56.085 6.940 56.170 7.065 ;
        RECT 56.790 6.940 56.875 7.100 ;
        RECT 58.985 7.065 59.035 7.100 ;
        POLYGON 59.035 7.100 59.070 7.065 59.035 7.065 ;
        RECT 58.985 6.940 59.070 7.065 ;
        RECT 59.690 6.940 59.775 7.100 ;
        RECT 61.885 7.065 61.935 7.100 ;
        POLYGON 61.935 7.100 61.970 7.065 61.935 7.065 ;
        RECT 61.885 6.940 61.970 7.065 ;
        RECT 62.590 6.940 62.675 7.100 ;
        RECT 64.785 7.065 64.835 7.100 ;
        POLYGON 64.835 7.100 64.870 7.065 64.835 7.065 ;
        RECT 64.785 6.940 64.870 7.065 ;
        RECT 65.490 6.940 65.575 7.100 ;
        RECT 67.685 7.065 67.735 7.100 ;
        POLYGON 67.735 7.100 67.770 7.065 67.735 7.065 ;
        RECT 67.685 6.940 67.770 7.065 ;
        RECT 68.390 6.940 68.475 7.100 ;
        RECT 70.585 7.065 70.635 7.100 ;
        POLYGON 70.635 7.100 70.670 7.065 70.635 7.065 ;
        RECT 70.585 6.940 70.670 7.065 ;
        RECT 71.290 6.940 71.375 7.100 ;
        RECT 73.485 7.065 73.535 7.100 ;
        POLYGON 73.535 7.100 73.570 7.065 73.535 7.065 ;
        RECT 73.485 6.940 73.570 7.065 ;
        RECT 74.190 6.940 74.275 7.100 ;
        RECT 76.385 7.065 76.435 7.100 ;
        POLYGON 76.435 7.100 76.470 7.065 76.435 7.065 ;
        RECT 76.385 6.940 76.470 7.065 ;
        RECT 77.090 6.940 77.175 7.100 ;
        RECT 79.285 7.065 79.335 7.100 ;
        POLYGON 79.335 7.100 79.370 7.065 79.335 7.065 ;
        RECT 79.285 6.940 79.370 7.065 ;
        RECT 79.990 6.940 80.075 7.100 ;
        RECT 82.185 7.065 82.235 7.100 ;
        POLYGON 82.235 7.100 82.270 7.065 82.235 7.065 ;
        RECT 82.185 6.940 82.270 7.065 ;
        RECT 82.890 6.940 82.975 7.100 ;
        RECT 85.085 7.065 85.135 7.100 ;
        POLYGON 85.135 7.100 85.170 7.065 85.135 7.065 ;
        RECT 85.085 6.940 85.170 7.065 ;
        RECT 85.790 6.940 85.875 7.100 ;
        RECT 87.985 7.065 88.035 7.100 ;
        POLYGON 88.035 7.100 88.070 7.065 88.035 7.065 ;
        RECT 87.985 6.940 88.070 7.065 ;
        RECT 88.690 6.940 88.775 7.100 ;
        RECT 90.885 7.065 90.935 7.100 ;
        POLYGON 90.935 7.100 90.970 7.065 90.935 7.065 ;
        RECT 90.885 6.940 90.970 7.065 ;
        RECT 91.590 6.940 91.675 7.100 ;
        RECT 0.775 6.320 0.850 6.460 ;
        RECT 0.990 6.270 1.065 6.410 ;
        RECT 1.695 6.330 1.755 6.410 ;
        POLYGON 1.695 6.330 1.755 6.330 1.755 6.270 ;
        RECT 1.910 6.320 1.985 6.460 ;
        RECT 3.675 6.320 3.750 6.460 ;
        RECT 3.890 6.270 3.965 6.410 ;
        RECT 4.595 6.330 4.655 6.410 ;
        POLYGON 4.595 6.330 4.655 6.330 4.655 6.270 ;
        RECT 4.810 6.320 4.885 6.460 ;
        RECT 6.575 6.320 6.650 6.460 ;
        RECT 6.790 6.270 6.865 6.410 ;
        RECT 7.495 6.330 7.555 6.410 ;
        POLYGON 7.495 6.330 7.555 6.330 7.555 6.270 ;
        RECT 7.710 6.320 7.785 6.460 ;
        RECT 9.475 6.320 9.550 6.460 ;
        RECT 9.690 6.270 9.765 6.410 ;
        RECT 10.395 6.330 10.455 6.410 ;
        POLYGON 10.395 6.330 10.455 6.330 10.455 6.270 ;
        RECT 10.610 6.320 10.685 6.460 ;
        RECT 12.375 6.320 12.450 6.460 ;
        RECT 12.590 6.270 12.665 6.410 ;
        RECT 13.295 6.330 13.355 6.410 ;
        POLYGON 13.295 6.330 13.355 6.330 13.355 6.270 ;
        RECT 13.510 6.320 13.585 6.460 ;
        RECT 15.275 6.320 15.350 6.460 ;
        RECT 15.490 6.270 15.565 6.410 ;
        RECT 16.195 6.330 16.255 6.410 ;
        POLYGON 16.195 6.330 16.255 6.330 16.255 6.270 ;
        RECT 16.410 6.320 16.485 6.460 ;
        RECT 18.175 6.320 18.250 6.460 ;
        RECT 18.390 6.270 18.465 6.410 ;
        RECT 19.095 6.330 19.155 6.410 ;
        POLYGON 19.095 6.330 19.155 6.330 19.155 6.270 ;
        RECT 19.310 6.320 19.385 6.460 ;
        RECT 21.075 6.320 21.150 6.460 ;
        RECT 21.290 6.270 21.365 6.410 ;
        RECT 21.995 6.330 22.055 6.410 ;
        POLYGON 21.995 6.330 22.055 6.330 22.055 6.270 ;
        RECT 22.210 6.320 22.285 6.460 ;
        RECT 23.975 6.320 24.050 6.460 ;
        RECT 24.190 6.270 24.265 6.410 ;
        RECT 24.895 6.330 24.955 6.410 ;
        POLYGON 24.895 6.330 24.955 6.330 24.955 6.270 ;
        RECT 25.110 6.320 25.185 6.460 ;
        RECT 26.875 6.320 26.950 6.460 ;
        RECT 27.090 6.270 27.165 6.410 ;
        RECT 27.795 6.330 27.855 6.410 ;
        POLYGON 27.795 6.330 27.855 6.330 27.855 6.270 ;
        RECT 28.010 6.320 28.085 6.460 ;
        RECT 29.775 6.320 29.850 6.460 ;
        RECT 29.990 6.270 30.065 6.410 ;
        RECT 30.695 6.330 30.755 6.410 ;
        POLYGON 30.695 6.330 30.755 6.330 30.755 6.270 ;
        RECT 30.910 6.320 30.985 6.460 ;
        RECT 32.675 6.320 32.750 6.460 ;
        RECT 32.890 6.270 32.965 6.410 ;
        RECT 33.595 6.330 33.655 6.410 ;
        POLYGON 33.595 6.330 33.655 6.330 33.655 6.270 ;
        RECT 33.810 6.320 33.885 6.460 ;
        RECT 35.575 6.320 35.650 6.460 ;
        RECT 35.790 6.270 35.865 6.410 ;
        RECT 36.495 6.330 36.555 6.410 ;
        POLYGON 36.495 6.330 36.555 6.330 36.555 6.270 ;
        RECT 36.710 6.320 36.785 6.460 ;
        RECT 38.475 6.320 38.550 6.460 ;
        RECT 38.690 6.270 38.765 6.410 ;
        RECT 39.395 6.330 39.455 6.410 ;
        POLYGON 39.395 6.330 39.455 6.330 39.455 6.270 ;
        RECT 39.610 6.320 39.685 6.460 ;
        RECT 41.375 6.320 41.450 6.460 ;
        RECT 41.590 6.270 41.665 6.410 ;
        RECT 42.295 6.330 42.355 6.410 ;
        POLYGON 42.295 6.330 42.355 6.330 42.355 6.270 ;
        RECT 42.510 6.320 42.585 6.460 ;
        RECT 44.275 6.320 44.350 6.460 ;
        RECT 44.490 6.270 44.565 6.410 ;
        RECT 45.195 6.330 45.255 6.410 ;
        POLYGON 45.195 6.330 45.255 6.330 45.255 6.270 ;
        RECT 45.410 6.320 45.485 6.460 ;
        RECT 47.175 6.320 47.250 6.460 ;
        RECT 47.390 6.270 47.465 6.410 ;
        RECT 48.095 6.330 48.155 6.410 ;
        POLYGON 48.095 6.330 48.155 6.330 48.155 6.270 ;
        RECT 48.310 6.320 48.385 6.460 ;
        RECT 50.075 6.320 50.150 6.460 ;
        RECT 50.290 6.270 50.365 6.410 ;
        RECT 50.995 6.330 51.055 6.410 ;
        POLYGON 50.995 6.330 51.055 6.330 51.055 6.270 ;
        RECT 51.210 6.320 51.285 6.460 ;
        RECT 52.975 6.320 53.050 6.460 ;
        RECT 53.190 6.270 53.265 6.410 ;
        RECT 53.895 6.330 53.955 6.410 ;
        POLYGON 53.895 6.330 53.955 6.330 53.955 6.270 ;
        RECT 54.110 6.320 54.185 6.460 ;
        RECT 55.875 6.320 55.950 6.460 ;
        RECT 56.090 6.270 56.165 6.410 ;
        RECT 56.795 6.330 56.855 6.410 ;
        POLYGON 56.795 6.330 56.855 6.330 56.855 6.270 ;
        RECT 57.010 6.320 57.085 6.460 ;
        RECT 58.775 6.320 58.850 6.460 ;
        RECT 58.990 6.270 59.065 6.410 ;
        RECT 59.695 6.330 59.755 6.410 ;
        POLYGON 59.695 6.330 59.755 6.330 59.755 6.270 ;
        RECT 59.910 6.320 59.985 6.460 ;
        RECT 61.675 6.320 61.750 6.460 ;
        RECT 61.890 6.270 61.965 6.410 ;
        RECT 62.595 6.330 62.655 6.410 ;
        POLYGON 62.595 6.330 62.655 6.330 62.655 6.270 ;
        RECT 62.810 6.320 62.885 6.460 ;
        RECT 64.575 6.320 64.650 6.460 ;
        RECT 64.790 6.270 64.865 6.410 ;
        RECT 65.495 6.330 65.555 6.410 ;
        POLYGON 65.495 6.330 65.555 6.330 65.555 6.270 ;
        RECT 65.710 6.320 65.785 6.460 ;
        RECT 67.475 6.320 67.550 6.460 ;
        RECT 67.690 6.270 67.765 6.410 ;
        RECT 68.395 6.330 68.455 6.410 ;
        POLYGON 68.395 6.330 68.455 6.330 68.455 6.270 ;
        RECT 68.610 6.320 68.685 6.460 ;
        RECT 70.375 6.320 70.450 6.460 ;
        RECT 70.590 6.270 70.665 6.410 ;
        RECT 71.295 6.330 71.355 6.410 ;
        POLYGON 71.295 6.330 71.355 6.330 71.355 6.270 ;
        RECT 71.510 6.320 71.585 6.460 ;
        RECT 73.275 6.320 73.350 6.460 ;
        RECT 73.490 6.270 73.565 6.410 ;
        RECT 74.195 6.330 74.255 6.410 ;
        POLYGON 74.195 6.330 74.255 6.330 74.255 6.270 ;
        RECT 74.410 6.320 74.485 6.460 ;
        RECT 76.175 6.320 76.250 6.460 ;
        RECT 76.390 6.270 76.465 6.410 ;
        RECT 77.095 6.330 77.155 6.410 ;
        POLYGON 77.095 6.330 77.155 6.330 77.155 6.270 ;
        RECT 77.310 6.320 77.385 6.460 ;
        RECT 79.075 6.320 79.150 6.460 ;
        RECT 79.290 6.270 79.365 6.410 ;
        RECT 79.995 6.330 80.055 6.410 ;
        POLYGON 79.995 6.330 80.055 6.330 80.055 6.270 ;
        RECT 80.210 6.320 80.285 6.460 ;
        RECT 81.975 6.320 82.050 6.460 ;
        RECT 82.190 6.270 82.265 6.410 ;
        RECT 82.895 6.330 82.955 6.410 ;
        POLYGON 82.895 6.330 82.955 6.330 82.955 6.270 ;
        RECT 83.110 6.320 83.185 6.460 ;
        RECT 84.875 6.320 84.950 6.460 ;
        RECT 85.090 6.270 85.165 6.410 ;
        RECT 85.795 6.330 85.855 6.410 ;
        POLYGON 85.795 6.330 85.855 6.330 85.855 6.270 ;
        RECT 86.010 6.320 86.085 6.460 ;
        RECT 87.775 6.320 87.850 6.460 ;
        RECT 87.990 6.270 88.065 6.410 ;
        RECT 88.695 6.330 88.755 6.410 ;
        POLYGON 88.695 6.330 88.755 6.330 88.755 6.270 ;
        RECT 88.910 6.320 88.985 6.460 ;
        RECT 90.675 6.320 90.750 6.460 ;
        RECT 90.890 6.270 90.965 6.410 ;
        RECT 91.595 6.330 91.655 6.410 ;
        POLYGON 91.595 6.330 91.655 6.330 91.655 6.270 ;
        RECT 91.810 6.320 91.885 6.460 ;
        RECT 0.720 5.800 0.870 5.970 ;
        RECT 1.110 5.935 1.260 6.105 ;
        RECT 1.500 5.935 1.650 6.105 ;
        RECT 1.890 5.800 2.040 5.970 ;
        RECT 3.620 5.800 3.770 5.970 ;
        RECT 4.010 5.935 4.160 6.105 ;
        RECT 4.400 5.935 4.550 6.105 ;
        RECT 4.790 5.800 4.940 5.970 ;
        RECT 6.520 5.800 6.670 5.970 ;
        RECT 6.910 5.935 7.060 6.105 ;
        RECT 7.300 5.935 7.450 6.105 ;
        RECT 7.690 5.800 7.840 5.970 ;
        RECT 9.420 5.800 9.570 5.970 ;
        RECT 9.810 5.935 9.960 6.105 ;
        RECT 10.200 5.935 10.350 6.105 ;
        RECT 10.590 5.800 10.740 5.970 ;
        RECT 12.320 5.800 12.470 5.970 ;
        RECT 12.710 5.935 12.860 6.105 ;
        RECT 13.100 5.935 13.250 6.105 ;
        RECT 13.490 5.800 13.640 5.970 ;
        RECT 15.220 5.800 15.370 5.970 ;
        RECT 15.610 5.935 15.760 6.105 ;
        RECT 16.000 5.935 16.150 6.105 ;
        RECT 16.390 5.800 16.540 5.970 ;
        RECT 18.120 5.800 18.270 5.970 ;
        RECT 18.510 5.935 18.660 6.105 ;
        RECT 18.900 5.935 19.050 6.105 ;
        RECT 19.290 5.800 19.440 5.970 ;
        RECT 21.020 5.800 21.170 5.970 ;
        RECT 21.410 5.935 21.560 6.105 ;
        RECT 21.800 5.935 21.950 6.105 ;
        RECT 22.190 5.800 22.340 5.970 ;
        RECT 23.920 5.800 24.070 5.970 ;
        RECT 24.310 5.935 24.460 6.105 ;
        RECT 24.700 5.935 24.850 6.105 ;
        RECT 25.090 5.800 25.240 5.970 ;
        RECT 26.820 5.800 26.970 5.970 ;
        RECT 27.210 5.935 27.360 6.105 ;
        RECT 27.600 5.935 27.750 6.105 ;
        RECT 27.990 5.800 28.140 5.970 ;
        RECT 29.720 5.800 29.870 5.970 ;
        RECT 30.110 5.935 30.260 6.105 ;
        RECT 30.500 5.935 30.650 6.105 ;
        RECT 30.890 5.800 31.040 5.970 ;
        RECT 32.620 5.800 32.770 5.970 ;
        RECT 33.010 5.935 33.160 6.105 ;
        RECT 33.400 5.935 33.550 6.105 ;
        RECT 33.790 5.800 33.940 5.970 ;
        RECT 35.520 5.800 35.670 5.970 ;
        RECT 35.910 5.935 36.060 6.105 ;
        RECT 36.300 5.935 36.450 6.105 ;
        RECT 36.690 5.800 36.840 5.970 ;
        RECT 38.420 5.800 38.570 5.970 ;
        RECT 38.810 5.935 38.960 6.105 ;
        RECT 39.200 5.935 39.350 6.105 ;
        RECT 39.590 5.800 39.740 5.970 ;
        RECT 41.320 5.800 41.470 5.970 ;
        RECT 41.710 5.935 41.860 6.105 ;
        RECT 42.100 5.935 42.250 6.105 ;
        RECT 42.490 5.800 42.640 5.970 ;
        RECT 44.220 5.800 44.370 5.970 ;
        RECT 44.610 5.935 44.760 6.105 ;
        RECT 45.000 5.935 45.150 6.105 ;
        RECT 45.390 5.800 45.540 5.970 ;
        RECT 47.120 5.800 47.270 5.970 ;
        RECT 47.510 5.935 47.660 6.105 ;
        RECT 47.900 5.935 48.050 6.105 ;
        RECT 48.290 5.800 48.440 5.970 ;
        RECT 50.020 5.800 50.170 5.970 ;
        RECT 50.410 5.935 50.560 6.105 ;
        RECT 50.800 5.935 50.950 6.105 ;
        RECT 51.190 5.800 51.340 5.970 ;
        RECT 52.920 5.800 53.070 5.970 ;
        RECT 53.310 5.935 53.460 6.105 ;
        RECT 53.700 5.935 53.850 6.105 ;
        RECT 54.090 5.800 54.240 5.970 ;
        RECT 55.820 5.800 55.970 5.970 ;
        RECT 56.210 5.935 56.360 6.105 ;
        RECT 56.600 5.935 56.750 6.105 ;
        RECT 56.990 5.800 57.140 5.970 ;
        RECT 58.720 5.800 58.870 5.970 ;
        RECT 59.110 5.935 59.260 6.105 ;
        RECT 59.500 5.935 59.650 6.105 ;
        RECT 59.890 5.800 60.040 5.970 ;
        RECT 61.620 5.800 61.770 5.970 ;
        RECT 62.010 5.935 62.160 6.105 ;
        RECT 62.400 5.935 62.550 6.105 ;
        RECT 62.790 5.800 62.940 5.970 ;
        RECT 64.520 5.800 64.670 5.970 ;
        RECT 64.910 5.935 65.060 6.105 ;
        RECT 65.300 5.935 65.450 6.105 ;
        RECT 65.690 5.800 65.840 5.970 ;
        RECT 67.420 5.800 67.570 5.970 ;
        RECT 67.810 5.935 67.960 6.105 ;
        RECT 68.200 5.935 68.350 6.105 ;
        RECT 68.590 5.800 68.740 5.970 ;
        RECT 70.320 5.800 70.470 5.970 ;
        RECT 70.710 5.935 70.860 6.105 ;
        RECT 71.100 5.935 71.250 6.105 ;
        RECT 71.490 5.800 71.640 5.970 ;
        RECT 73.220 5.800 73.370 5.970 ;
        RECT 73.610 5.935 73.760 6.105 ;
        RECT 74.000 5.935 74.150 6.105 ;
        RECT 74.390 5.800 74.540 5.970 ;
        RECT 76.120 5.800 76.270 5.970 ;
        RECT 76.510 5.935 76.660 6.105 ;
        RECT 76.900 5.935 77.050 6.105 ;
        RECT 77.290 5.800 77.440 5.970 ;
        RECT 79.020 5.800 79.170 5.970 ;
        RECT 79.410 5.935 79.560 6.105 ;
        RECT 79.800 5.935 79.950 6.105 ;
        RECT 80.190 5.800 80.340 5.970 ;
        RECT 81.920 5.800 82.070 5.970 ;
        RECT 82.310 5.935 82.460 6.105 ;
        RECT 82.700 5.935 82.850 6.105 ;
        RECT 83.090 5.800 83.240 5.970 ;
        RECT 84.820 5.800 84.970 5.970 ;
        RECT 85.210 5.935 85.360 6.105 ;
        RECT 85.600 5.935 85.750 6.105 ;
        RECT 85.990 5.800 86.140 5.970 ;
        RECT 87.720 5.800 87.870 5.970 ;
        RECT 88.110 5.935 88.260 6.105 ;
        RECT 88.500 5.935 88.650 6.105 ;
        RECT 88.890 5.800 89.040 5.970 ;
        RECT 90.620 5.800 90.770 5.970 ;
        RECT 91.010 5.935 91.160 6.105 ;
        RECT 91.400 5.935 91.550 6.105 ;
        RECT 91.790 5.800 91.940 5.970 ;
        RECT 0.985 5.715 1.035 5.750 ;
        POLYGON 1.035 5.750 1.070 5.715 1.035 5.715 ;
        RECT 0.985 5.590 1.070 5.715 ;
        RECT 1.690 5.590 1.775 5.750 ;
        RECT 3.885 5.715 3.935 5.750 ;
        POLYGON 3.935 5.750 3.970 5.715 3.935 5.715 ;
        RECT 3.885 5.590 3.970 5.715 ;
        RECT 4.590 5.590 4.675 5.750 ;
        RECT 6.785 5.715 6.835 5.750 ;
        POLYGON 6.835 5.750 6.870 5.715 6.835 5.715 ;
        RECT 6.785 5.590 6.870 5.715 ;
        RECT 7.490 5.590 7.575 5.750 ;
        RECT 9.685 5.715 9.735 5.750 ;
        POLYGON 9.735 5.750 9.770 5.715 9.735 5.715 ;
        RECT 9.685 5.590 9.770 5.715 ;
        RECT 10.390 5.590 10.475 5.750 ;
        RECT 12.585 5.715 12.635 5.750 ;
        POLYGON 12.635 5.750 12.670 5.715 12.635 5.715 ;
        RECT 12.585 5.590 12.670 5.715 ;
        RECT 13.290 5.590 13.375 5.750 ;
        RECT 15.485 5.715 15.535 5.750 ;
        POLYGON 15.535 5.750 15.570 5.715 15.535 5.715 ;
        RECT 15.485 5.590 15.570 5.715 ;
        RECT 16.190 5.590 16.275 5.750 ;
        RECT 18.385 5.715 18.435 5.750 ;
        POLYGON 18.435 5.750 18.470 5.715 18.435 5.715 ;
        RECT 18.385 5.590 18.470 5.715 ;
        RECT 19.090 5.590 19.175 5.750 ;
        RECT 21.285 5.715 21.335 5.750 ;
        POLYGON 21.335 5.750 21.370 5.715 21.335 5.715 ;
        RECT 21.285 5.590 21.370 5.715 ;
        RECT 21.990 5.590 22.075 5.750 ;
        RECT 24.185 5.715 24.235 5.750 ;
        POLYGON 24.235 5.750 24.270 5.715 24.235 5.715 ;
        RECT 24.185 5.590 24.270 5.715 ;
        RECT 24.890 5.590 24.975 5.750 ;
        RECT 27.085 5.715 27.135 5.750 ;
        POLYGON 27.135 5.750 27.170 5.715 27.135 5.715 ;
        RECT 27.085 5.590 27.170 5.715 ;
        RECT 27.790 5.590 27.875 5.750 ;
        RECT 29.985 5.715 30.035 5.750 ;
        POLYGON 30.035 5.750 30.070 5.715 30.035 5.715 ;
        RECT 29.985 5.590 30.070 5.715 ;
        RECT 30.690 5.590 30.775 5.750 ;
        RECT 32.885 5.715 32.935 5.750 ;
        POLYGON 32.935 5.750 32.970 5.715 32.935 5.715 ;
        RECT 32.885 5.590 32.970 5.715 ;
        RECT 33.590 5.590 33.675 5.750 ;
        RECT 35.785 5.715 35.835 5.750 ;
        POLYGON 35.835 5.750 35.870 5.715 35.835 5.715 ;
        RECT 35.785 5.590 35.870 5.715 ;
        RECT 36.490 5.590 36.575 5.750 ;
        RECT 38.685 5.715 38.735 5.750 ;
        POLYGON 38.735 5.750 38.770 5.715 38.735 5.715 ;
        RECT 38.685 5.590 38.770 5.715 ;
        RECT 39.390 5.590 39.475 5.750 ;
        RECT 41.585 5.715 41.635 5.750 ;
        POLYGON 41.635 5.750 41.670 5.715 41.635 5.715 ;
        RECT 41.585 5.590 41.670 5.715 ;
        RECT 42.290 5.590 42.375 5.750 ;
        RECT 44.485 5.715 44.535 5.750 ;
        POLYGON 44.535 5.750 44.570 5.715 44.535 5.715 ;
        RECT 44.485 5.590 44.570 5.715 ;
        RECT 45.190 5.590 45.275 5.750 ;
        RECT 47.385 5.715 47.435 5.750 ;
        POLYGON 47.435 5.750 47.470 5.715 47.435 5.715 ;
        RECT 47.385 5.590 47.470 5.715 ;
        RECT 48.090 5.590 48.175 5.750 ;
        RECT 50.285 5.715 50.335 5.750 ;
        POLYGON 50.335 5.750 50.370 5.715 50.335 5.715 ;
        RECT 50.285 5.590 50.370 5.715 ;
        RECT 50.990 5.590 51.075 5.750 ;
        RECT 53.185 5.715 53.235 5.750 ;
        POLYGON 53.235 5.750 53.270 5.715 53.235 5.715 ;
        RECT 53.185 5.590 53.270 5.715 ;
        RECT 53.890 5.590 53.975 5.750 ;
        RECT 56.085 5.715 56.135 5.750 ;
        POLYGON 56.135 5.750 56.170 5.715 56.135 5.715 ;
        RECT 56.085 5.590 56.170 5.715 ;
        RECT 56.790 5.590 56.875 5.750 ;
        RECT 58.985 5.715 59.035 5.750 ;
        POLYGON 59.035 5.750 59.070 5.715 59.035 5.715 ;
        RECT 58.985 5.590 59.070 5.715 ;
        RECT 59.690 5.590 59.775 5.750 ;
        RECT 61.885 5.715 61.935 5.750 ;
        POLYGON 61.935 5.750 61.970 5.715 61.935 5.715 ;
        RECT 61.885 5.590 61.970 5.715 ;
        RECT 62.590 5.590 62.675 5.750 ;
        RECT 64.785 5.715 64.835 5.750 ;
        POLYGON 64.835 5.750 64.870 5.715 64.835 5.715 ;
        RECT 64.785 5.590 64.870 5.715 ;
        RECT 65.490 5.590 65.575 5.750 ;
        RECT 67.685 5.715 67.735 5.750 ;
        POLYGON 67.735 5.750 67.770 5.715 67.735 5.715 ;
        RECT 67.685 5.590 67.770 5.715 ;
        RECT 68.390 5.590 68.475 5.750 ;
        RECT 70.585 5.715 70.635 5.750 ;
        POLYGON 70.635 5.750 70.670 5.715 70.635 5.715 ;
        RECT 70.585 5.590 70.670 5.715 ;
        RECT 71.290 5.590 71.375 5.750 ;
        RECT 73.485 5.715 73.535 5.750 ;
        POLYGON 73.535 5.750 73.570 5.715 73.535 5.715 ;
        RECT 73.485 5.590 73.570 5.715 ;
        RECT 74.190 5.590 74.275 5.750 ;
        RECT 76.385 5.715 76.435 5.750 ;
        POLYGON 76.435 5.750 76.470 5.715 76.435 5.715 ;
        RECT 76.385 5.590 76.470 5.715 ;
        RECT 77.090 5.590 77.175 5.750 ;
        RECT 79.285 5.715 79.335 5.750 ;
        POLYGON 79.335 5.750 79.370 5.715 79.335 5.715 ;
        RECT 79.285 5.590 79.370 5.715 ;
        RECT 79.990 5.590 80.075 5.750 ;
        RECT 82.185 5.715 82.235 5.750 ;
        POLYGON 82.235 5.750 82.270 5.715 82.235 5.715 ;
        RECT 82.185 5.590 82.270 5.715 ;
        RECT 82.890 5.590 82.975 5.750 ;
        RECT 85.085 5.715 85.135 5.750 ;
        POLYGON 85.135 5.750 85.170 5.715 85.135 5.715 ;
        RECT 85.085 5.590 85.170 5.715 ;
        RECT 85.790 5.590 85.875 5.750 ;
        RECT 87.985 5.715 88.035 5.750 ;
        POLYGON 88.035 5.750 88.070 5.715 88.035 5.715 ;
        RECT 87.985 5.590 88.070 5.715 ;
        RECT 88.690 5.590 88.775 5.750 ;
        RECT 90.885 5.715 90.935 5.750 ;
        POLYGON 90.935 5.750 90.970 5.715 90.935 5.715 ;
        RECT 90.885 5.590 90.970 5.715 ;
        RECT 91.590 5.590 91.675 5.750 ;
        RECT 0.775 4.970 0.850 5.110 ;
        RECT 0.990 4.920 1.065 5.060 ;
        RECT 1.695 4.980 1.755 5.060 ;
        POLYGON 1.695 4.980 1.755 4.980 1.755 4.920 ;
        RECT 1.910 4.970 1.985 5.110 ;
        RECT 3.675 4.970 3.750 5.110 ;
        RECT 3.890 4.920 3.965 5.060 ;
        RECT 4.595 4.980 4.655 5.060 ;
        POLYGON 4.595 4.980 4.655 4.980 4.655 4.920 ;
        RECT 4.810 4.970 4.885 5.110 ;
        RECT 6.575 4.970 6.650 5.110 ;
        RECT 6.790 4.920 6.865 5.060 ;
        RECT 7.495 4.980 7.555 5.060 ;
        POLYGON 7.495 4.980 7.555 4.980 7.555 4.920 ;
        RECT 7.710 4.970 7.785 5.110 ;
        RECT 9.475 4.970 9.550 5.110 ;
        RECT 9.690 4.920 9.765 5.060 ;
        RECT 10.395 4.980 10.455 5.060 ;
        POLYGON 10.395 4.980 10.455 4.980 10.455 4.920 ;
        RECT 10.610 4.970 10.685 5.110 ;
        RECT 12.375 4.970 12.450 5.110 ;
        RECT 12.590 4.920 12.665 5.060 ;
        RECT 13.295 4.980 13.355 5.060 ;
        POLYGON 13.295 4.980 13.355 4.980 13.355 4.920 ;
        RECT 13.510 4.970 13.585 5.110 ;
        RECT 15.275 4.970 15.350 5.110 ;
        RECT 15.490 4.920 15.565 5.060 ;
        RECT 16.195 4.980 16.255 5.060 ;
        POLYGON 16.195 4.980 16.255 4.980 16.255 4.920 ;
        RECT 16.410 4.970 16.485 5.110 ;
        RECT 18.175 4.970 18.250 5.110 ;
        RECT 18.390 4.920 18.465 5.060 ;
        RECT 19.095 4.980 19.155 5.060 ;
        POLYGON 19.095 4.980 19.155 4.980 19.155 4.920 ;
        RECT 19.310 4.970 19.385 5.110 ;
        RECT 21.075 4.970 21.150 5.110 ;
        RECT 21.290 4.920 21.365 5.060 ;
        RECT 21.995 4.980 22.055 5.060 ;
        POLYGON 21.995 4.980 22.055 4.980 22.055 4.920 ;
        RECT 22.210 4.970 22.285 5.110 ;
        RECT 23.975 4.970 24.050 5.110 ;
        RECT 24.190 4.920 24.265 5.060 ;
        RECT 24.895 4.980 24.955 5.060 ;
        POLYGON 24.895 4.980 24.955 4.980 24.955 4.920 ;
        RECT 25.110 4.970 25.185 5.110 ;
        RECT 26.875 4.970 26.950 5.110 ;
        RECT 27.090 4.920 27.165 5.060 ;
        RECT 27.795 4.980 27.855 5.060 ;
        POLYGON 27.795 4.980 27.855 4.980 27.855 4.920 ;
        RECT 28.010 4.970 28.085 5.110 ;
        RECT 29.775 4.970 29.850 5.110 ;
        RECT 29.990 4.920 30.065 5.060 ;
        RECT 30.695 4.980 30.755 5.060 ;
        POLYGON 30.695 4.980 30.755 4.980 30.755 4.920 ;
        RECT 30.910 4.970 30.985 5.110 ;
        RECT 32.675 4.970 32.750 5.110 ;
        RECT 32.890 4.920 32.965 5.060 ;
        RECT 33.595 4.980 33.655 5.060 ;
        POLYGON 33.595 4.980 33.655 4.980 33.655 4.920 ;
        RECT 33.810 4.970 33.885 5.110 ;
        RECT 35.575 4.970 35.650 5.110 ;
        RECT 35.790 4.920 35.865 5.060 ;
        RECT 36.495 4.980 36.555 5.060 ;
        POLYGON 36.495 4.980 36.555 4.980 36.555 4.920 ;
        RECT 36.710 4.970 36.785 5.110 ;
        RECT 38.475 4.970 38.550 5.110 ;
        RECT 38.690 4.920 38.765 5.060 ;
        RECT 39.395 4.980 39.455 5.060 ;
        POLYGON 39.395 4.980 39.455 4.980 39.455 4.920 ;
        RECT 39.610 4.970 39.685 5.110 ;
        RECT 41.375 4.970 41.450 5.110 ;
        RECT 41.590 4.920 41.665 5.060 ;
        RECT 42.295 4.980 42.355 5.060 ;
        POLYGON 42.295 4.980 42.355 4.980 42.355 4.920 ;
        RECT 42.510 4.970 42.585 5.110 ;
        RECT 44.275 4.970 44.350 5.110 ;
        RECT 44.490 4.920 44.565 5.060 ;
        RECT 45.195 4.980 45.255 5.060 ;
        POLYGON 45.195 4.980 45.255 4.980 45.255 4.920 ;
        RECT 45.410 4.970 45.485 5.110 ;
        RECT 47.175 4.970 47.250 5.110 ;
        RECT 47.390 4.920 47.465 5.060 ;
        RECT 48.095 4.980 48.155 5.060 ;
        POLYGON 48.095 4.980 48.155 4.980 48.155 4.920 ;
        RECT 48.310 4.970 48.385 5.110 ;
        RECT 50.075 4.970 50.150 5.110 ;
        RECT 50.290 4.920 50.365 5.060 ;
        RECT 50.995 4.980 51.055 5.060 ;
        POLYGON 50.995 4.980 51.055 4.980 51.055 4.920 ;
        RECT 51.210 4.970 51.285 5.110 ;
        RECT 52.975 4.970 53.050 5.110 ;
        RECT 53.190 4.920 53.265 5.060 ;
        RECT 53.895 4.980 53.955 5.060 ;
        POLYGON 53.895 4.980 53.955 4.980 53.955 4.920 ;
        RECT 54.110 4.970 54.185 5.110 ;
        RECT 55.875 4.970 55.950 5.110 ;
        RECT 56.090 4.920 56.165 5.060 ;
        RECT 56.795 4.980 56.855 5.060 ;
        POLYGON 56.795 4.980 56.855 4.980 56.855 4.920 ;
        RECT 57.010 4.970 57.085 5.110 ;
        RECT 58.775 4.970 58.850 5.110 ;
        RECT 58.990 4.920 59.065 5.060 ;
        RECT 59.695 4.980 59.755 5.060 ;
        POLYGON 59.695 4.980 59.755 4.980 59.755 4.920 ;
        RECT 59.910 4.970 59.985 5.110 ;
        RECT 61.675 4.970 61.750 5.110 ;
        RECT 61.890 4.920 61.965 5.060 ;
        RECT 62.595 4.980 62.655 5.060 ;
        POLYGON 62.595 4.980 62.655 4.980 62.655 4.920 ;
        RECT 62.810 4.970 62.885 5.110 ;
        RECT 64.575 4.970 64.650 5.110 ;
        RECT 64.790 4.920 64.865 5.060 ;
        RECT 65.495 4.980 65.555 5.060 ;
        POLYGON 65.495 4.980 65.555 4.980 65.555 4.920 ;
        RECT 65.710 4.970 65.785 5.110 ;
        RECT 67.475 4.970 67.550 5.110 ;
        RECT 67.690 4.920 67.765 5.060 ;
        RECT 68.395 4.980 68.455 5.060 ;
        POLYGON 68.395 4.980 68.455 4.980 68.455 4.920 ;
        RECT 68.610 4.970 68.685 5.110 ;
        RECT 70.375 4.970 70.450 5.110 ;
        RECT 70.590 4.920 70.665 5.060 ;
        RECT 71.295 4.980 71.355 5.060 ;
        POLYGON 71.295 4.980 71.355 4.980 71.355 4.920 ;
        RECT 71.510 4.970 71.585 5.110 ;
        RECT 73.275 4.970 73.350 5.110 ;
        RECT 73.490 4.920 73.565 5.060 ;
        RECT 74.195 4.980 74.255 5.060 ;
        POLYGON 74.195 4.980 74.255 4.980 74.255 4.920 ;
        RECT 74.410 4.970 74.485 5.110 ;
        RECT 76.175 4.970 76.250 5.110 ;
        RECT 76.390 4.920 76.465 5.060 ;
        RECT 77.095 4.980 77.155 5.060 ;
        POLYGON 77.095 4.980 77.155 4.980 77.155 4.920 ;
        RECT 77.310 4.970 77.385 5.110 ;
        RECT 79.075 4.970 79.150 5.110 ;
        RECT 79.290 4.920 79.365 5.060 ;
        RECT 79.995 4.980 80.055 5.060 ;
        POLYGON 79.995 4.980 80.055 4.980 80.055 4.920 ;
        RECT 80.210 4.970 80.285 5.110 ;
        RECT 81.975 4.970 82.050 5.110 ;
        RECT 82.190 4.920 82.265 5.060 ;
        RECT 82.895 4.980 82.955 5.060 ;
        POLYGON 82.895 4.980 82.955 4.980 82.955 4.920 ;
        RECT 83.110 4.970 83.185 5.110 ;
        RECT 84.875 4.970 84.950 5.110 ;
        RECT 85.090 4.920 85.165 5.060 ;
        RECT 85.795 4.980 85.855 5.060 ;
        POLYGON 85.795 4.980 85.855 4.980 85.855 4.920 ;
        RECT 86.010 4.970 86.085 5.110 ;
        RECT 87.775 4.970 87.850 5.110 ;
        RECT 87.990 4.920 88.065 5.060 ;
        RECT 88.695 4.980 88.755 5.060 ;
        POLYGON 88.695 4.980 88.755 4.980 88.755 4.920 ;
        RECT 88.910 4.970 88.985 5.110 ;
        RECT 90.675 4.970 90.750 5.110 ;
        RECT 90.890 4.920 90.965 5.060 ;
        RECT 91.595 4.980 91.655 5.060 ;
        POLYGON 91.595 4.980 91.655 4.980 91.655 4.920 ;
        RECT 91.810 4.970 91.885 5.110 ;
        RECT 0.720 4.450 0.870 4.620 ;
        RECT 1.110 4.585 1.260 4.755 ;
        RECT 1.500 4.585 1.650 4.755 ;
        RECT 1.890 4.450 2.040 4.620 ;
        RECT 3.620 4.450 3.770 4.620 ;
        RECT 4.010 4.585 4.160 4.755 ;
        RECT 4.400 4.585 4.550 4.755 ;
        RECT 4.790 4.450 4.940 4.620 ;
        RECT 6.520 4.450 6.670 4.620 ;
        RECT 6.910 4.585 7.060 4.755 ;
        RECT 7.300 4.585 7.450 4.755 ;
        RECT 7.690 4.450 7.840 4.620 ;
        RECT 9.420 4.450 9.570 4.620 ;
        RECT 9.810 4.585 9.960 4.755 ;
        RECT 10.200 4.585 10.350 4.755 ;
        RECT 10.590 4.450 10.740 4.620 ;
        RECT 12.320 4.450 12.470 4.620 ;
        RECT 12.710 4.585 12.860 4.755 ;
        RECT 13.100 4.585 13.250 4.755 ;
        RECT 13.490 4.450 13.640 4.620 ;
        RECT 15.220 4.450 15.370 4.620 ;
        RECT 15.610 4.585 15.760 4.755 ;
        RECT 16.000 4.585 16.150 4.755 ;
        RECT 16.390 4.450 16.540 4.620 ;
        RECT 18.120 4.450 18.270 4.620 ;
        RECT 18.510 4.585 18.660 4.755 ;
        RECT 18.900 4.585 19.050 4.755 ;
        RECT 19.290 4.450 19.440 4.620 ;
        RECT 21.020 4.450 21.170 4.620 ;
        RECT 21.410 4.585 21.560 4.755 ;
        RECT 21.800 4.585 21.950 4.755 ;
        RECT 22.190 4.450 22.340 4.620 ;
        RECT 23.920 4.450 24.070 4.620 ;
        RECT 24.310 4.585 24.460 4.755 ;
        RECT 24.700 4.585 24.850 4.755 ;
        RECT 25.090 4.450 25.240 4.620 ;
        RECT 26.820 4.450 26.970 4.620 ;
        RECT 27.210 4.585 27.360 4.755 ;
        RECT 27.600 4.585 27.750 4.755 ;
        RECT 27.990 4.450 28.140 4.620 ;
        RECT 29.720 4.450 29.870 4.620 ;
        RECT 30.110 4.585 30.260 4.755 ;
        RECT 30.500 4.585 30.650 4.755 ;
        RECT 30.890 4.450 31.040 4.620 ;
        RECT 32.620 4.450 32.770 4.620 ;
        RECT 33.010 4.585 33.160 4.755 ;
        RECT 33.400 4.585 33.550 4.755 ;
        RECT 33.790 4.450 33.940 4.620 ;
        RECT 35.520 4.450 35.670 4.620 ;
        RECT 35.910 4.585 36.060 4.755 ;
        RECT 36.300 4.585 36.450 4.755 ;
        RECT 36.690 4.450 36.840 4.620 ;
        RECT 38.420 4.450 38.570 4.620 ;
        RECT 38.810 4.585 38.960 4.755 ;
        RECT 39.200 4.585 39.350 4.755 ;
        RECT 39.590 4.450 39.740 4.620 ;
        RECT 41.320 4.450 41.470 4.620 ;
        RECT 41.710 4.585 41.860 4.755 ;
        RECT 42.100 4.585 42.250 4.755 ;
        RECT 42.490 4.450 42.640 4.620 ;
        RECT 44.220 4.450 44.370 4.620 ;
        RECT 44.610 4.585 44.760 4.755 ;
        RECT 45.000 4.585 45.150 4.755 ;
        RECT 45.390 4.450 45.540 4.620 ;
        RECT 47.120 4.450 47.270 4.620 ;
        RECT 47.510 4.585 47.660 4.755 ;
        RECT 47.900 4.585 48.050 4.755 ;
        RECT 48.290 4.450 48.440 4.620 ;
        RECT 50.020 4.450 50.170 4.620 ;
        RECT 50.410 4.585 50.560 4.755 ;
        RECT 50.800 4.585 50.950 4.755 ;
        RECT 51.190 4.450 51.340 4.620 ;
        RECT 52.920 4.450 53.070 4.620 ;
        RECT 53.310 4.585 53.460 4.755 ;
        RECT 53.700 4.585 53.850 4.755 ;
        RECT 54.090 4.450 54.240 4.620 ;
        RECT 55.820 4.450 55.970 4.620 ;
        RECT 56.210 4.585 56.360 4.755 ;
        RECT 56.600 4.585 56.750 4.755 ;
        RECT 56.990 4.450 57.140 4.620 ;
        RECT 58.720 4.450 58.870 4.620 ;
        RECT 59.110 4.585 59.260 4.755 ;
        RECT 59.500 4.585 59.650 4.755 ;
        RECT 59.890 4.450 60.040 4.620 ;
        RECT 61.620 4.450 61.770 4.620 ;
        RECT 62.010 4.585 62.160 4.755 ;
        RECT 62.400 4.585 62.550 4.755 ;
        RECT 62.790 4.450 62.940 4.620 ;
        RECT 64.520 4.450 64.670 4.620 ;
        RECT 64.910 4.585 65.060 4.755 ;
        RECT 65.300 4.585 65.450 4.755 ;
        RECT 65.690 4.450 65.840 4.620 ;
        RECT 67.420 4.450 67.570 4.620 ;
        RECT 67.810 4.585 67.960 4.755 ;
        RECT 68.200 4.585 68.350 4.755 ;
        RECT 68.590 4.450 68.740 4.620 ;
        RECT 70.320 4.450 70.470 4.620 ;
        RECT 70.710 4.585 70.860 4.755 ;
        RECT 71.100 4.585 71.250 4.755 ;
        RECT 71.490 4.450 71.640 4.620 ;
        RECT 73.220 4.450 73.370 4.620 ;
        RECT 73.610 4.585 73.760 4.755 ;
        RECT 74.000 4.585 74.150 4.755 ;
        RECT 74.390 4.450 74.540 4.620 ;
        RECT 76.120 4.450 76.270 4.620 ;
        RECT 76.510 4.585 76.660 4.755 ;
        RECT 76.900 4.585 77.050 4.755 ;
        RECT 77.290 4.450 77.440 4.620 ;
        RECT 79.020 4.450 79.170 4.620 ;
        RECT 79.410 4.585 79.560 4.755 ;
        RECT 79.800 4.585 79.950 4.755 ;
        RECT 80.190 4.450 80.340 4.620 ;
        RECT 81.920 4.450 82.070 4.620 ;
        RECT 82.310 4.585 82.460 4.755 ;
        RECT 82.700 4.585 82.850 4.755 ;
        RECT 83.090 4.450 83.240 4.620 ;
        RECT 84.820 4.450 84.970 4.620 ;
        RECT 85.210 4.585 85.360 4.755 ;
        RECT 85.600 4.585 85.750 4.755 ;
        RECT 85.990 4.450 86.140 4.620 ;
        RECT 87.720 4.450 87.870 4.620 ;
        RECT 88.110 4.585 88.260 4.755 ;
        RECT 88.500 4.585 88.650 4.755 ;
        RECT 88.890 4.450 89.040 4.620 ;
        RECT 90.620 4.450 90.770 4.620 ;
        RECT 91.010 4.585 91.160 4.755 ;
        RECT 91.400 4.585 91.550 4.755 ;
        RECT 91.790 4.450 91.940 4.620 ;
        RECT 0.985 4.365 1.035 4.400 ;
        POLYGON 1.035 4.400 1.070 4.365 1.035 4.365 ;
        RECT 0.985 4.240 1.070 4.365 ;
        RECT 1.690 4.240 1.775 4.400 ;
        RECT 3.885 4.365 3.935 4.400 ;
        POLYGON 3.935 4.400 3.970 4.365 3.935 4.365 ;
        RECT 3.885 4.240 3.970 4.365 ;
        RECT 4.590 4.240 4.675 4.400 ;
        RECT 6.785 4.365 6.835 4.400 ;
        POLYGON 6.835 4.400 6.870 4.365 6.835 4.365 ;
        RECT 6.785 4.240 6.870 4.365 ;
        RECT 7.490 4.240 7.575 4.400 ;
        RECT 9.685 4.365 9.735 4.400 ;
        POLYGON 9.735 4.400 9.770 4.365 9.735 4.365 ;
        RECT 9.685 4.240 9.770 4.365 ;
        RECT 10.390 4.240 10.475 4.400 ;
        RECT 12.585 4.365 12.635 4.400 ;
        POLYGON 12.635 4.400 12.670 4.365 12.635 4.365 ;
        RECT 12.585 4.240 12.670 4.365 ;
        RECT 13.290 4.240 13.375 4.400 ;
        RECT 15.485 4.365 15.535 4.400 ;
        POLYGON 15.535 4.400 15.570 4.365 15.535 4.365 ;
        RECT 15.485 4.240 15.570 4.365 ;
        RECT 16.190 4.240 16.275 4.400 ;
        RECT 18.385 4.365 18.435 4.400 ;
        POLYGON 18.435 4.400 18.470 4.365 18.435 4.365 ;
        RECT 18.385 4.240 18.470 4.365 ;
        RECT 19.090 4.240 19.175 4.400 ;
        RECT 21.285 4.365 21.335 4.400 ;
        POLYGON 21.335 4.400 21.370 4.365 21.335 4.365 ;
        RECT 21.285 4.240 21.370 4.365 ;
        RECT 21.990 4.240 22.075 4.400 ;
        RECT 24.185 4.365 24.235 4.400 ;
        POLYGON 24.235 4.400 24.270 4.365 24.235 4.365 ;
        RECT 24.185 4.240 24.270 4.365 ;
        RECT 24.890 4.240 24.975 4.400 ;
        RECT 27.085 4.365 27.135 4.400 ;
        POLYGON 27.135 4.400 27.170 4.365 27.135 4.365 ;
        RECT 27.085 4.240 27.170 4.365 ;
        RECT 27.790 4.240 27.875 4.400 ;
        RECT 29.985 4.365 30.035 4.400 ;
        POLYGON 30.035 4.400 30.070 4.365 30.035 4.365 ;
        RECT 29.985 4.240 30.070 4.365 ;
        RECT 30.690 4.240 30.775 4.400 ;
        RECT 32.885 4.365 32.935 4.400 ;
        POLYGON 32.935 4.400 32.970 4.365 32.935 4.365 ;
        RECT 32.885 4.240 32.970 4.365 ;
        RECT 33.590 4.240 33.675 4.400 ;
        RECT 35.785 4.365 35.835 4.400 ;
        POLYGON 35.835 4.400 35.870 4.365 35.835 4.365 ;
        RECT 35.785 4.240 35.870 4.365 ;
        RECT 36.490 4.240 36.575 4.400 ;
        RECT 38.685 4.365 38.735 4.400 ;
        POLYGON 38.735 4.400 38.770 4.365 38.735 4.365 ;
        RECT 38.685 4.240 38.770 4.365 ;
        RECT 39.390 4.240 39.475 4.400 ;
        RECT 41.585 4.365 41.635 4.400 ;
        POLYGON 41.635 4.400 41.670 4.365 41.635 4.365 ;
        RECT 41.585 4.240 41.670 4.365 ;
        RECT 42.290 4.240 42.375 4.400 ;
        RECT 44.485 4.365 44.535 4.400 ;
        POLYGON 44.535 4.400 44.570 4.365 44.535 4.365 ;
        RECT 44.485 4.240 44.570 4.365 ;
        RECT 45.190 4.240 45.275 4.400 ;
        RECT 47.385 4.365 47.435 4.400 ;
        POLYGON 47.435 4.400 47.470 4.365 47.435 4.365 ;
        RECT 47.385 4.240 47.470 4.365 ;
        RECT 48.090 4.240 48.175 4.400 ;
        RECT 50.285 4.365 50.335 4.400 ;
        POLYGON 50.335 4.400 50.370 4.365 50.335 4.365 ;
        RECT 50.285 4.240 50.370 4.365 ;
        RECT 50.990 4.240 51.075 4.400 ;
        RECT 53.185 4.365 53.235 4.400 ;
        POLYGON 53.235 4.400 53.270 4.365 53.235 4.365 ;
        RECT 53.185 4.240 53.270 4.365 ;
        RECT 53.890 4.240 53.975 4.400 ;
        RECT 56.085 4.365 56.135 4.400 ;
        POLYGON 56.135 4.400 56.170 4.365 56.135 4.365 ;
        RECT 56.085 4.240 56.170 4.365 ;
        RECT 56.790 4.240 56.875 4.400 ;
        RECT 58.985 4.365 59.035 4.400 ;
        POLYGON 59.035 4.400 59.070 4.365 59.035 4.365 ;
        RECT 58.985 4.240 59.070 4.365 ;
        RECT 59.690 4.240 59.775 4.400 ;
        RECT 61.885 4.365 61.935 4.400 ;
        POLYGON 61.935 4.400 61.970 4.365 61.935 4.365 ;
        RECT 61.885 4.240 61.970 4.365 ;
        RECT 62.590 4.240 62.675 4.400 ;
        RECT 64.785 4.365 64.835 4.400 ;
        POLYGON 64.835 4.400 64.870 4.365 64.835 4.365 ;
        RECT 64.785 4.240 64.870 4.365 ;
        RECT 65.490 4.240 65.575 4.400 ;
        RECT 67.685 4.365 67.735 4.400 ;
        POLYGON 67.735 4.400 67.770 4.365 67.735 4.365 ;
        RECT 67.685 4.240 67.770 4.365 ;
        RECT 68.390 4.240 68.475 4.400 ;
        RECT 70.585 4.365 70.635 4.400 ;
        POLYGON 70.635 4.400 70.670 4.365 70.635 4.365 ;
        RECT 70.585 4.240 70.670 4.365 ;
        RECT 71.290 4.240 71.375 4.400 ;
        RECT 73.485 4.365 73.535 4.400 ;
        POLYGON 73.535 4.400 73.570 4.365 73.535 4.365 ;
        RECT 73.485 4.240 73.570 4.365 ;
        RECT 74.190 4.240 74.275 4.400 ;
        RECT 76.385 4.365 76.435 4.400 ;
        POLYGON 76.435 4.400 76.470 4.365 76.435 4.365 ;
        RECT 76.385 4.240 76.470 4.365 ;
        RECT 77.090 4.240 77.175 4.400 ;
        RECT 79.285 4.365 79.335 4.400 ;
        POLYGON 79.335 4.400 79.370 4.365 79.335 4.365 ;
        RECT 79.285 4.240 79.370 4.365 ;
        RECT 79.990 4.240 80.075 4.400 ;
        RECT 82.185 4.365 82.235 4.400 ;
        POLYGON 82.235 4.400 82.270 4.365 82.235 4.365 ;
        RECT 82.185 4.240 82.270 4.365 ;
        RECT 82.890 4.240 82.975 4.400 ;
        RECT 85.085 4.365 85.135 4.400 ;
        POLYGON 85.135 4.400 85.170 4.365 85.135 4.365 ;
        RECT 85.085 4.240 85.170 4.365 ;
        RECT 85.790 4.240 85.875 4.400 ;
        RECT 87.985 4.365 88.035 4.400 ;
        POLYGON 88.035 4.400 88.070 4.365 88.035 4.365 ;
        RECT 87.985 4.240 88.070 4.365 ;
        RECT 88.690 4.240 88.775 4.400 ;
        RECT 90.885 4.365 90.935 4.400 ;
        POLYGON 90.935 4.400 90.970 4.365 90.935 4.365 ;
        RECT 90.885 4.240 90.970 4.365 ;
        RECT 91.590 4.240 91.675 4.400 ;
        RECT 0.775 3.620 0.850 3.760 ;
        RECT 0.990 3.570 1.065 3.710 ;
        RECT 1.695 3.630 1.755 3.710 ;
        POLYGON 1.695 3.630 1.755 3.630 1.755 3.570 ;
        RECT 1.910 3.620 1.985 3.760 ;
        RECT 3.675 3.620 3.750 3.760 ;
        RECT 3.890 3.570 3.965 3.710 ;
        RECT 4.595 3.630 4.655 3.710 ;
        POLYGON 4.595 3.630 4.655 3.630 4.655 3.570 ;
        RECT 4.810 3.620 4.885 3.760 ;
        RECT 6.575 3.620 6.650 3.760 ;
        RECT 6.790 3.570 6.865 3.710 ;
        RECT 7.495 3.630 7.555 3.710 ;
        POLYGON 7.495 3.630 7.555 3.630 7.555 3.570 ;
        RECT 7.710 3.620 7.785 3.760 ;
        RECT 9.475 3.620 9.550 3.760 ;
        RECT 9.690 3.570 9.765 3.710 ;
        RECT 10.395 3.630 10.455 3.710 ;
        POLYGON 10.395 3.630 10.455 3.630 10.455 3.570 ;
        RECT 10.610 3.620 10.685 3.760 ;
        RECT 12.375 3.620 12.450 3.760 ;
        RECT 12.590 3.570 12.665 3.710 ;
        RECT 13.295 3.630 13.355 3.710 ;
        POLYGON 13.295 3.630 13.355 3.630 13.355 3.570 ;
        RECT 13.510 3.620 13.585 3.760 ;
        RECT 15.275 3.620 15.350 3.760 ;
        RECT 15.490 3.570 15.565 3.710 ;
        RECT 16.195 3.630 16.255 3.710 ;
        POLYGON 16.195 3.630 16.255 3.630 16.255 3.570 ;
        RECT 16.410 3.620 16.485 3.760 ;
        RECT 18.175 3.620 18.250 3.760 ;
        RECT 18.390 3.570 18.465 3.710 ;
        RECT 19.095 3.630 19.155 3.710 ;
        POLYGON 19.095 3.630 19.155 3.630 19.155 3.570 ;
        RECT 19.310 3.620 19.385 3.760 ;
        RECT 21.075 3.620 21.150 3.760 ;
        RECT 21.290 3.570 21.365 3.710 ;
        RECT 21.995 3.630 22.055 3.710 ;
        POLYGON 21.995 3.630 22.055 3.630 22.055 3.570 ;
        RECT 22.210 3.620 22.285 3.760 ;
        RECT 23.975 3.620 24.050 3.760 ;
        RECT 24.190 3.570 24.265 3.710 ;
        RECT 24.895 3.630 24.955 3.710 ;
        POLYGON 24.895 3.630 24.955 3.630 24.955 3.570 ;
        RECT 25.110 3.620 25.185 3.760 ;
        RECT 26.875 3.620 26.950 3.760 ;
        RECT 27.090 3.570 27.165 3.710 ;
        RECT 27.795 3.630 27.855 3.710 ;
        POLYGON 27.795 3.630 27.855 3.630 27.855 3.570 ;
        RECT 28.010 3.620 28.085 3.760 ;
        RECT 29.775 3.620 29.850 3.760 ;
        RECT 29.990 3.570 30.065 3.710 ;
        RECT 30.695 3.630 30.755 3.710 ;
        POLYGON 30.695 3.630 30.755 3.630 30.755 3.570 ;
        RECT 30.910 3.620 30.985 3.760 ;
        RECT 32.675 3.620 32.750 3.760 ;
        RECT 32.890 3.570 32.965 3.710 ;
        RECT 33.595 3.630 33.655 3.710 ;
        POLYGON 33.595 3.630 33.655 3.630 33.655 3.570 ;
        RECT 33.810 3.620 33.885 3.760 ;
        RECT 35.575 3.620 35.650 3.760 ;
        RECT 35.790 3.570 35.865 3.710 ;
        RECT 36.495 3.630 36.555 3.710 ;
        POLYGON 36.495 3.630 36.555 3.630 36.555 3.570 ;
        RECT 36.710 3.620 36.785 3.760 ;
        RECT 38.475 3.620 38.550 3.760 ;
        RECT 38.690 3.570 38.765 3.710 ;
        RECT 39.395 3.630 39.455 3.710 ;
        POLYGON 39.395 3.630 39.455 3.630 39.455 3.570 ;
        RECT 39.610 3.620 39.685 3.760 ;
        RECT 41.375 3.620 41.450 3.760 ;
        RECT 41.590 3.570 41.665 3.710 ;
        RECT 42.295 3.630 42.355 3.710 ;
        POLYGON 42.295 3.630 42.355 3.630 42.355 3.570 ;
        RECT 42.510 3.620 42.585 3.760 ;
        RECT 44.275 3.620 44.350 3.760 ;
        RECT 44.490 3.570 44.565 3.710 ;
        RECT 45.195 3.630 45.255 3.710 ;
        POLYGON 45.195 3.630 45.255 3.630 45.255 3.570 ;
        RECT 45.410 3.620 45.485 3.760 ;
        RECT 47.175 3.620 47.250 3.760 ;
        RECT 47.390 3.570 47.465 3.710 ;
        RECT 48.095 3.630 48.155 3.710 ;
        POLYGON 48.095 3.630 48.155 3.630 48.155 3.570 ;
        RECT 48.310 3.620 48.385 3.760 ;
        RECT 50.075 3.620 50.150 3.760 ;
        RECT 50.290 3.570 50.365 3.710 ;
        RECT 50.995 3.630 51.055 3.710 ;
        POLYGON 50.995 3.630 51.055 3.630 51.055 3.570 ;
        RECT 51.210 3.620 51.285 3.760 ;
        RECT 52.975 3.620 53.050 3.760 ;
        RECT 53.190 3.570 53.265 3.710 ;
        RECT 53.895 3.630 53.955 3.710 ;
        POLYGON 53.895 3.630 53.955 3.630 53.955 3.570 ;
        RECT 54.110 3.620 54.185 3.760 ;
        RECT 55.875 3.620 55.950 3.760 ;
        RECT 56.090 3.570 56.165 3.710 ;
        RECT 56.795 3.630 56.855 3.710 ;
        POLYGON 56.795 3.630 56.855 3.630 56.855 3.570 ;
        RECT 57.010 3.620 57.085 3.760 ;
        RECT 58.775 3.620 58.850 3.760 ;
        RECT 58.990 3.570 59.065 3.710 ;
        RECT 59.695 3.630 59.755 3.710 ;
        POLYGON 59.695 3.630 59.755 3.630 59.755 3.570 ;
        RECT 59.910 3.620 59.985 3.760 ;
        RECT 61.675 3.620 61.750 3.760 ;
        RECT 61.890 3.570 61.965 3.710 ;
        RECT 62.595 3.630 62.655 3.710 ;
        POLYGON 62.595 3.630 62.655 3.630 62.655 3.570 ;
        RECT 62.810 3.620 62.885 3.760 ;
        RECT 64.575 3.620 64.650 3.760 ;
        RECT 64.790 3.570 64.865 3.710 ;
        RECT 65.495 3.630 65.555 3.710 ;
        POLYGON 65.495 3.630 65.555 3.630 65.555 3.570 ;
        RECT 65.710 3.620 65.785 3.760 ;
        RECT 67.475 3.620 67.550 3.760 ;
        RECT 67.690 3.570 67.765 3.710 ;
        RECT 68.395 3.630 68.455 3.710 ;
        POLYGON 68.395 3.630 68.455 3.630 68.455 3.570 ;
        RECT 68.610 3.620 68.685 3.760 ;
        RECT 70.375 3.620 70.450 3.760 ;
        RECT 70.590 3.570 70.665 3.710 ;
        RECT 71.295 3.630 71.355 3.710 ;
        POLYGON 71.295 3.630 71.355 3.630 71.355 3.570 ;
        RECT 71.510 3.620 71.585 3.760 ;
        RECT 73.275 3.620 73.350 3.760 ;
        RECT 73.490 3.570 73.565 3.710 ;
        RECT 74.195 3.630 74.255 3.710 ;
        POLYGON 74.195 3.630 74.255 3.630 74.255 3.570 ;
        RECT 74.410 3.620 74.485 3.760 ;
        RECT 76.175 3.620 76.250 3.760 ;
        RECT 76.390 3.570 76.465 3.710 ;
        RECT 77.095 3.630 77.155 3.710 ;
        POLYGON 77.095 3.630 77.155 3.630 77.155 3.570 ;
        RECT 77.310 3.620 77.385 3.760 ;
        RECT 79.075 3.620 79.150 3.760 ;
        RECT 79.290 3.570 79.365 3.710 ;
        RECT 79.995 3.630 80.055 3.710 ;
        POLYGON 79.995 3.630 80.055 3.630 80.055 3.570 ;
        RECT 80.210 3.620 80.285 3.760 ;
        RECT 81.975 3.620 82.050 3.760 ;
        RECT 82.190 3.570 82.265 3.710 ;
        RECT 82.895 3.630 82.955 3.710 ;
        POLYGON 82.895 3.630 82.955 3.630 82.955 3.570 ;
        RECT 83.110 3.620 83.185 3.760 ;
        RECT 84.875 3.620 84.950 3.760 ;
        RECT 85.090 3.570 85.165 3.710 ;
        RECT 85.795 3.630 85.855 3.710 ;
        POLYGON 85.795 3.630 85.855 3.630 85.855 3.570 ;
        RECT 86.010 3.620 86.085 3.760 ;
        RECT 87.775 3.620 87.850 3.760 ;
        RECT 87.990 3.570 88.065 3.710 ;
        RECT 88.695 3.630 88.755 3.710 ;
        POLYGON 88.695 3.630 88.755 3.630 88.755 3.570 ;
        RECT 88.910 3.620 88.985 3.760 ;
        RECT 90.675 3.620 90.750 3.760 ;
        RECT 90.890 3.570 90.965 3.710 ;
        RECT 91.595 3.630 91.655 3.710 ;
        POLYGON 91.595 3.630 91.655 3.630 91.655 3.570 ;
        RECT 91.810 3.620 91.885 3.760 ;
        RECT 0.720 3.100 0.870 3.270 ;
        RECT 1.110 3.235 1.260 3.405 ;
        RECT 1.500 3.235 1.650 3.405 ;
        RECT 1.890 3.100 2.040 3.270 ;
        RECT 3.620 3.100 3.770 3.270 ;
        RECT 4.010 3.235 4.160 3.405 ;
        RECT 4.400 3.235 4.550 3.405 ;
        RECT 4.790 3.100 4.940 3.270 ;
        RECT 6.520 3.100 6.670 3.270 ;
        RECT 6.910 3.235 7.060 3.405 ;
        RECT 7.300 3.235 7.450 3.405 ;
        RECT 7.690 3.100 7.840 3.270 ;
        RECT 9.420 3.100 9.570 3.270 ;
        RECT 9.810 3.235 9.960 3.405 ;
        RECT 10.200 3.235 10.350 3.405 ;
        RECT 10.590 3.100 10.740 3.270 ;
        RECT 12.320 3.100 12.470 3.270 ;
        RECT 12.710 3.235 12.860 3.405 ;
        RECT 13.100 3.235 13.250 3.405 ;
        RECT 13.490 3.100 13.640 3.270 ;
        RECT 15.220 3.100 15.370 3.270 ;
        RECT 15.610 3.235 15.760 3.405 ;
        RECT 16.000 3.235 16.150 3.405 ;
        RECT 16.390 3.100 16.540 3.270 ;
        RECT 18.120 3.100 18.270 3.270 ;
        RECT 18.510 3.235 18.660 3.405 ;
        RECT 18.900 3.235 19.050 3.405 ;
        RECT 19.290 3.100 19.440 3.270 ;
        RECT 21.020 3.100 21.170 3.270 ;
        RECT 21.410 3.235 21.560 3.405 ;
        RECT 21.800 3.235 21.950 3.405 ;
        RECT 22.190 3.100 22.340 3.270 ;
        RECT 23.920 3.100 24.070 3.270 ;
        RECT 24.310 3.235 24.460 3.405 ;
        RECT 24.700 3.235 24.850 3.405 ;
        RECT 25.090 3.100 25.240 3.270 ;
        RECT 26.820 3.100 26.970 3.270 ;
        RECT 27.210 3.235 27.360 3.405 ;
        RECT 27.600 3.235 27.750 3.405 ;
        RECT 27.990 3.100 28.140 3.270 ;
        RECT 29.720 3.100 29.870 3.270 ;
        RECT 30.110 3.235 30.260 3.405 ;
        RECT 30.500 3.235 30.650 3.405 ;
        RECT 30.890 3.100 31.040 3.270 ;
        RECT 32.620 3.100 32.770 3.270 ;
        RECT 33.010 3.235 33.160 3.405 ;
        RECT 33.400 3.235 33.550 3.405 ;
        RECT 33.790 3.100 33.940 3.270 ;
        RECT 35.520 3.100 35.670 3.270 ;
        RECT 35.910 3.235 36.060 3.405 ;
        RECT 36.300 3.235 36.450 3.405 ;
        RECT 36.690 3.100 36.840 3.270 ;
        RECT 38.420 3.100 38.570 3.270 ;
        RECT 38.810 3.235 38.960 3.405 ;
        RECT 39.200 3.235 39.350 3.405 ;
        RECT 39.590 3.100 39.740 3.270 ;
        RECT 41.320 3.100 41.470 3.270 ;
        RECT 41.710 3.235 41.860 3.405 ;
        RECT 42.100 3.235 42.250 3.405 ;
        RECT 42.490 3.100 42.640 3.270 ;
        RECT 44.220 3.100 44.370 3.270 ;
        RECT 44.610 3.235 44.760 3.405 ;
        RECT 45.000 3.235 45.150 3.405 ;
        RECT 45.390 3.100 45.540 3.270 ;
        RECT 47.120 3.100 47.270 3.270 ;
        RECT 47.510 3.235 47.660 3.405 ;
        RECT 47.900 3.235 48.050 3.405 ;
        RECT 48.290 3.100 48.440 3.270 ;
        RECT 50.020 3.100 50.170 3.270 ;
        RECT 50.410 3.235 50.560 3.405 ;
        RECT 50.800 3.235 50.950 3.405 ;
        RECT 51.190 3.100 51.340 3.270 ;
        RECT 52.920 3.100 53.070 3.270 ;
        RECT 53.310 3.235 53.460 3.405 ;
        RECT 53.700 3.235 53.850 3.405 ;
        RECT 54.090 3.100 54.240 3.270 ;
        RECT 55.820 3.100 55.970 3.270 ;
        RECT 56.210 3.235 56.360 3.405 ;
        RECT 56.600 3.235 56.750 3.405 ;
        RECT 56.990 3.100 57.140 3.270 ;
        RECT 58.720 3.100 58.870 3.270 ;
        RECT 59.110 3.235 59.260 3.405 ;
        RECT 59.500 3.235 59.650 3.405 ;
        RECT 59.890 3.100 60.040 3.270 ;
        RECT 61.620 3.100 61.770 3.270 ;
        RECT 62.010 3.235 62.160 3.405 ;
        RECT 62.400 3.235 62.550 3.405 ;
        RECT 62.790 3.100 62.940 3.270 ;
        RECT 64.520 3.100 64.670 3.270 ;
        RECT 64.910 3.235 65.060 3.405 ;
        RECT 65.300 3.235 65.450 3.405 ;
        RECT 65.690 3.100 65.840 3.270 ;
        RECT 67.420 3.100 67.570 3.270 ;
        RECT 67.810 3.235 67.960 3.405 ;
        RECT 68.200 3.235 68.350 3.405 ;
        RECT 68.590 3.100 68.740 3.270 ;
        RECT 70.320 3.100 70.470 3.270 ;
        RECT 70.710 3.235 70.860 3.405 ;
        RECT 71.100 3.235 71.250 3.405 ;
        RECT 71.490 3.100 71.640 3.270 ;
        RECT 73.220 3.100 73.370 3.270 ;
        RECT 73.610 3.235 73.760 3.405 ;
        RECT 74.000 3.235 74.150 3.405 ;
        RECT 74.390 3.100 74.540 3.270 ;
        RECT 76.120 3.100 76.270 3.270 ;
        RECT 76.510 3.235 76.660 3.405 ;
        RECT 76.900 3.235 77.050 3.405 ;
        RECT 77.290 3.100 77.440 3.270 ;
        RECT 79.020 3.100 79.170 3.270 ;
        RECT 79.410 3.235 79.560 3.405 ;
        RECT 79.800 3.235 79.950 3.405 ;
        RECT 80.190 3.100 80.340 3.270 ;
        RECT 81.920 3.100 82.070 3.270 ;
        RECT 82.310 3.235 82.460 3.405 ;
        RECT 82.700 3.235 82.850 3.405 ;
        RECT 83.090 3.100 83.240 3.270 ;
        RECT 84.820 3.100 84.970 3.270 ;
        RECT 85.210 3.235 85.360 3.405 ;
        RECT 85.600 3.235 85.750 3.405 ;
        RECT 85.990 3.100 86.140 3.270 ;
        RECT 87.720 3.100 87.870 3.270 ;
        RECT 88.110 3.235 88.260 3.405 ;
        RECT 88.500 3.235 88.650 3.405 ;
        RECT 88.890 3.100 89.040 3.270 ;
        RECT 90.620 3.100 90.770 3.270 ;
        RECT 91.010 3.235 91.160 3.405 ;
        RECT 91.400 3.235 91.550 3.405 ;
        RECT 91.790 3.100 91.940 3.270 ;
        RECT 0.985 3.015 1.035 3.050 ;
        POLYGON 1.035 3.050 1.070 3.015 1.035 3.015 ;
        RECT 0.985 2.890 1.070 3.015 ;
        RECT 1.690 2.890 1.775 3.050 ;
        RECT 3.885 3.015 3.935 3.050 ;
        POLYGON 3.935 3.050 3.970 3.015 3.935 3.015 ;
        RECT 3.885 2.890 3.970 3.015 ;
        RECT 4.590 2.890 4.675 3.050 ;
        RECT 6.785 3.015 6.835 3.050 ;
        POLYGON 6.835 3.050 6.870 3.015 6.835 3.015 ;
        RECT 6.785 2.890 6.870 3.015 ;
        RECT 7.490 2.890 7.575 3.050 ;
        RECT 9.685 3.015 9.735 3.050 ;
        POLYGON 9.735 3.050 9.770 3.015 9.735 3.015 ;
        RECT 9.685 2.890 9.770 3.015 ;
        RECT 10.390 2.890 10.475 3.050 ;
        RECT 12.585 3.015 12.635 3.050 ;
        POLYGON 12.635 3.050 12.670 3.015 12.635 3.015 ;
        RECT 12.585 2.890 12.670 3.015 ;
        RECT 13.290 2.890 13.375 3.050 ;
        RECT 15.485 3.015 15.535 3.050 ;
        POLYGON 15.535 3.050 15.570 3.015 15.535 3.015 ;
        RECT 15.485 2.890 15.570 3.015 ;
        RECT 16.190 2.890 16.275 3.050 ;
        RECT 18.385 3.015 18.435 3.050 ;
        POLYGON 18.435 3.050 18.470 3.015 18.435 3.015 ;
        RECT 18.385 2.890 18.470 3.015 ;
        RECT 19.090 2.890 19.175 3.050 ;
        RECT 21.285 3.015 21.335 3.050 ;
        POLYGON 21.335 3.050 21.370 3.015 21.335 3.015 ;
        RECT 21.285 2.890 21.370 3.015 ;
        RECT 21.990 2.890 22.075 3.050 ;
        RECT 24.185 3.015 24.235 3.050 ;
        POLYGON 24.235 3.050 24.270 3.015 24.235 3.015 ;
        RECT 24.185 2.890 24.270 3.015 ;
        RECT 24.890 2.890 24.975 3.050 ;
        RECT 27.085 3.015 27.135 3.050 ;
        POLYGON 27.135 3.050 27.170 3.015 27.135 3.015 ;
        RECT 27.085 2.890 27.170 3.015 ;
        RECT 27.790 2.890 27.875 3.050 ;
        RECT 29.985 3.015 30.035 3.050 ;
        POLYGON 30.035 3.050 30.070 3.015 30.035 3.015 ;
        RECT 29.985 2.890 30.070 3.015 ;
        RECT 30.690 2.890 30.775 3.050 ;
        RECT 32.885 3.015 32.935 3.050 ;
        POLYGON 32.935 3.050 32.970 3.015 32.935 3.015 ;
        RECT 32.885 2.890 32.970 3.015 ;
        RECT 33.590 2.890 33.675 3.050 ;
        RECT 35.785 3.015 35.835 3.050 ;
        POLYGON 35.835 3.050 35.870 3.015 35.835 3.015 ;
        RECT 35.785 2.890 35.870 3.015 ;
        RECT 36.490 2.890 36.575 3.050 ;
        RECT 38.685 3.015 38.735 3.050 ;
        POLYGON 38.735 3.050 38.770 3.015 38.735 3.015 ;
        RECT 38.685 2.890 38.770 3.015 ;
        RECT 39.390 2.890 39.475 3.050 ;
        RECT 41.585 3.015 41.635 3.050 ;
        POLYGON 41.635 3.050 41.670 3.015 41.635 3.015 ;
        RECT 41.585 2.890 41.670 3.015 ;
        RECT 42.290 2.890 42.375 3.050 ;
        RECT 44.485 3.015 44.535 3.050 ;
        POLYGON 44.535 3.050 44.570 3.015 44.535 3.015 ;
        RECT 44.485 2.890 44.570 3.015 ;
        RECT 45.190 2.890 45.275 3.050 ;
        RECT 47.385 3.015 47.435 3.050 ;
        POLYGON 47.435 3.050 47.470 3.015 47.435 3.015 ;
        RECT 47.385 2.890 47.470 3.015 ;
        RECT 48.090 2.890 48.175 3.050 ;
        RECT 50.285 3.015 50.335 3.050 ;
        POLYGON 50.335 3.050 50.370 3.015 50.335 3.015 ;
        RECT 50.285 2.890 50.370 3.015 ;
        RECT 50.990 2.890 51.075 3.050 ;
        RECT 53.185 3.015 53.235 3.050 ;
        POLYGON 53.235 3.050 53.270 3.015 53.235 3.015 ;
        RECT 53.185 2.890 53.270 3.015 ;
        RECT 53.890 2.890 53.975 3.050 ;
        RECT 56.085 3.015 56.135 3.050 ;
        POLYGON 56.135 3.050 56.170 3.015 56.135 3.015 ;
        RECT 56.085 2.890 56.170 3.015 ;
        RECT 56.790 2.890 56.875 3.050 ;
        RECT 58.985 3.015 59.035 3.050 ;
        POLYGON 59.035 3.050 59.070 3.015 59.035 3.015 ;
        RECT 58.985 2.890 59.070 3.015 ;
        RECT 59.690 2.890 59.775 3.050 ;
        RECT 61.885 3.015 61.935 3.050 ;
        POLYGON 61.935 3.050 61.970 3.015 61.935 3.015 ;
        RECT 61.885 2.890 61.970 3.015 ;
        RECT 62.590 2.890 62.675 3.050 ;
        RECT 64.785 3.015 64.835 3.050 ;
        POLYGON 64.835 3.050 64.870 3.015 64.835 3.015 ;
        RECT 64.785 2.890 64.870 3.015 ;
        RECT 65.490 2.890 65.575 3.050 ;
        RECT 67.685 3.015 67.735 3.050 ;
        POLYGON 67.735 3.050 67.770 3.015 67.735 3.015 ;
        RECT 67.685 2.890 67.770 3.015 ;
        RECT 68.390 2.890 68.475 3.050 ;
        RECT 70.585 3.015 70.635 3.050 ;
        POLYGON 70.635 3.050 70.670 3.015 70.635 3.015 ;
        RECT 70.585 2.890 70.670 3.015 ;
        RECT 71.290 2.890 71.375 3.050 ;
        RECT 73.485 3.015 73.535 3.050 ;
        POLYGON 73.535 3.050 73.570 3.015 73.535 3.015 ;
        RECT 73.485 2.890 73.570 3.015 ;
        RECT 74.190 2.890 74.275 3.050 ;
        RECT 76.385 3.015 76.435 3.050 ;
        POLYGON 76.435 3.050 76.470 3.015 76.435 3.015 ;
        RECT 76.385 2.890 76.470 3.015 ;
        RECT 77.090 2.890 77.175 3.050 ;
        RECT 79.285 3.015 79.335 3.050 ;
        POLYGON 79.335 3.050 79.370 3.015 79.335 3.015 ;
        RECT 79.285 2.890 79.370 3.015 ;
        RECT 79.990 2.890 80.075 3.050 ;
        RECT 82.185 3.015 82.235 3.050 ;
        POLYGON 82.235 3.050 82.270 3.015 82.235 3.015 ;
        RECT 82.185 2.890 82.270 3.015 ;
        RECT 82.890 2.890 82.975 3.050 ;
        RECT 85.085 3.015 85.135 3.050 ;
        POLYGON 85.135 3.050 85.170 3.015 85.135 3.015 ;
        RECT 85.085 2.890 85.170 3.015 ;
        RECT 85.790 2.890 85.875 3.050 ;
        RECT 87.985 3.015 88.035 3.050 ;
        POLYGON 88.035 3.050 88.070 3.015 88.035 3.015 ;
        RECT 87.985 2.890 88.070 3.015 ;
        RECT 88.690 2.890 88.775 3.050 ;
        RECT 90.885 3.015 90.935 3.050 ;
        POLYGON 90.935 3.050 90.970 3.015 90.935 3.015 ;
        RECT 90.885 2.890 90.970 3.015 ;
        RECT 91.590 2.890 91.675 3.050 ;
        RECT 0.775 2.270 0.850 2.410 ;
        RECT 0.990 2.220 1.065 2.360 ;
        RECT 1.695 2.280 1.755 2.360 ;
        POLYGON 1.695 2.280 1.755 2.280 1.755 2.220 ;
        RECT 1.910 2.270 1.985 2.410 ;
        RECT 3.675 2.270 3.750 2.410 ;
        RECT 3.890 2.220 3.965 2.360 ;
        RECT 4.595 2.280 4.655 2.360 ;
        POLYGON 4.595 2.280 4.655 2.280 4.655 2.220 ;
        RECT 4.810 2.270 4.885 2.410 ;
        RECT 6.575 2.270 6.650 2.410 ;
        RECT 6.790 2.220 6.865 2.360 ;
        RECT 7.495 2.280 7.555 2.360 ;
        POLYGON 7.495 2.280 7.555 2.280 7.555 2.220 ;
        RECT 7.710 2.270 7.785 2.410 ;
        RECT 9.475 2.270 9.550 2.410 ;
        RECT 9.690 2.220 9.765 2.360 ;
        RECT 10.395 2.280 10.455 2.360 ;
        POLYGON 10.395 2.280 10.455 2.280 10.455 2.220 ;
        RECT 10.610 2.270 10.685 2.410 ;
        RECT 12.375 2.270 12.450 2.410 ;
        RECT 12.590 2.220 12.665 2.360 ;
        RECT 13.295 2.280 13.355 2.360 ;
        POLYGON 13.295 2.280 13.355 2.280 13.355 2.220 ;
        RECT 13.510 2.270 13.585 2.410 ;
        RECT 15.275 2.270 15.350 2.410 ;
        RECT 15.490 2.220 15.565 2.360 ;
        RECT 16.195 2.280 16.255 2.360 ;
        POLYGON 16.195 2.280 16.255 2.280 16.255 2.220 ;
        RECT 16.410 2.270 16.485 2.410 ;
        RECT 18.175 2.270 18.250 2.410 ;
        RECT 18.390 2.220 18.465 2.360 ;
        RECT 19.095 2.280 19.155 2.360 ;
        POLYGON 19.095 2.280 19.155 2.280 19.155 2.220 ;
        RECT 19.310 2.270 19.385 2.410 ;
        RECT 21.075 2.270 21.150 2.410 ;
        RECT 21.290 2.220 21.365 2.360 ;
        RECT 21.995 2.280 22.055 2.360 ;
        POLYGON 21.995 2.280 22.055 2.280 22.055 2.220 ;
        RECT 22.210 2.270 22.285 2.410 ;
        RECT 23.975 2.275 24.050 2.415 ;
        RECT 24.190 2.225 24.265 2.365 ;
        RECT 24.895 2.285 24.955 2.365 ;
        POLYGON 24.895 2.285 24.955 2.285 24.955 2.225 ;
        RECT 25.110 2.275 25.185 2.415 ;
        RECT 26.875 2.275 26.950 2.415 ;
        RECT 27.090 2.225 27.165 2.365 ;
        RECT 27.795 2.285 27.855 2.365 ;
        POLYGON 27.795 2.285 27.855 2.285 27.855 2.225 ;
        RECT 28.010 2.275 28.085 2.415 ;
        RECT 29.775 2.275 29.850 2.415 ;
        RECT 29.990 2.225 30.065 2.365 ;
        RECT 30.695 2.285 30.755 2.365 ;
        POLYGON 30.695 2.285 30.755 2.285 30.755 2.225 ;
        RECT 30.910 2.275 30.985 2.415 ;
        RECT 32.675 2.275 32.750 2.415 ;
        RECT 32.890 2.225 32.965 2.365 ;
        RECT 33.595 2.285 33.655 2.365 ;
        POLYGON 33.595 2.285 33.655 2.285 33.655 2.225 ;
        RECT 33.810 2.275 33.885 2.415 ;
        RECT 35.575 2.275 35.650 2.415 ;
        RECT 35.790 2.225 35.865 2.365 ;
        RECT 36.495 2.285 36.555 2.365 ;
        POLYGON 36.495 2.285 36.555 2.285 36.555 2.225 ;
        RECT 36.710 2.275 36.785 2.415 ;
        RECT 38.475 2.275 38.550 2.415 ;
        RECT 38.690 2.225 38.765 2.365 ;
        RECT 39.395 2.285 39.455 2.365 ;
        POLYGON 39.395 2.285 39.455 2.285 39.455 2.225 ;
        RECT 39.610 2.275 39.685 2.415 ;
        RECT 41.375 2.275 41.450 2.415 ;
        RECT 41.590 2.225 41.665 2.365 ;
        RECT 42.295 2.285 42.355 2.365 ;
        POLYGON 42.295 2.285 42.355 2.285 42.355 2.225 ;
        RECT 42.510 2.275 42.585 2.415 ;
        RECT 44.275 2.275 44.350 2.415 ;
        RECT 44.490 2.225 44.565 2.365 ;
        RECT 45.195 2.285 45.255 2.365 ;
        POLYGON 45.195 2.285 45.255 2.285 45.255 2.225 ;
        RECT 45.410 2.275 45.485 2.415 ;
        RECT 47.175 2.275 47.250 2.415 ;
        RECT 47.390 2.225 47.465 2.365 ;
        RECT 48.095 2.285 48.155 2.365 ;
        POLYGON 48.095 2.285 48.155 2.285 48.155 2.225 ;
        RECT 48.310 2.275 48.385 2.415 ;
        RECT 50.075 2.275 50.150 2.415 ;
        RECT 50.290 2.225 50.365 2.365 ;
        RECT 50.995 2.285 51.055 2.365 ;
        POLYGON 50.995 2.285 51.055 2.285 51.055 2.225 ;
        RECT 51.210 2.275 51.285 2.415 ;
        RECT 52.975 2.275 53.050 2.415 ;
        RECT 53.190 2.225 53.265 2.365 ;
        RECT 53.895 2.285 53.955 2.365 ;
        POLYGON 53.895 2.285 53.955 2.285 53.955 2.225 ;
        RECT 54.110 2.275 54.185 2.415 ;
        RECT 55.875 2.275 55.950 2.415 ;
        RECT 56.090 2.225 56.165 2.365 ;
        RECT 56.795 2.285 56.855 2.365 ;
        POLYGON 56.795 2.285 56.855 2.285 56.855 2.225 ;
        RECT 57.010 2.275 57.085 2.415 ;
        RECT 58.775 2.275 58.850 2.415 ;
        RECT 58.990 2.225 59.065 2.365 ;
        RECT 59.695 2.285 59.755 2.365 ;
        POLYGON 59.695 2.285 59.755 2.285 59.755 2.225 ;
        RECT 59.910 2.275 59.985 2.415 ;
        RECT 61.675 2.275 61.750 2.415 ;
        RECT 61.890 2.225 61.965 2.365 ;
        RECT 62.595 2.285 62.655 2.365 ;
        POLYGON 62.595 2.285 62.655 2.285 62.655 2.225 ;
        RECT 62.810 2.275 62.885 2.415 ;
        RECT 64.575 2.275 64.650 2.415 ;
        RECT 64.790 2.225 64.865 2.365 ;
        RECT 65.495 2.285 65.555 2.365 ;
        POLYGON 65.495 2.285 65.555 2.285 65.555 2.225 ;
        RECT 65.710 2.275 65.785 2.415 ;
        RECT 67.475 2.275 67.550 2.415 ;
        RECT 67.690 2.225 67.765 2.365 ;
        RECT 68.395 2.285 68.455 2.365 ;
        POLYGON 68.395 2.285 68.455 2.285 68.455 2.225 ;
        RECT 68.610 2.275 68.685 2.415 ;
        RECT 70.375 2.275 70.450 2.415 ;
        RECT 70.590 2.225 70.665 2.365 ;
        RECT 71.295 2.285 71.355 2.365 ;
        POLYGON 71.295 2.285 71.355 2.285 71.355 2.225 ;
        RECT 71.510 2.275 71.585 2.415 ;
        RECT 73.275 2.275 73.350 2.415 ;
        RECT 73.490 2.225 73.565 2.365 ;
        RECT 74.195 2.285 74.255 2.365 ;
        POLYGON 74.195 2.285 74.255 2.285 74.255 2.225 ;
        RECT 74.410 2.275 74.485 2.415 ;
        RECT 76.175 2.275 76.250 2.415 ;
        RECT 76.390 2.225 76.465 2.365 ;
        RECT 77.095 2.285 77.155 2.365 ;
        POLYGON 77.095 2.285 77.155 2.285 77.155 2.225 ;
        RECT 77.310 2.275 77.385 2.415 ;
        RECT 79.075 2.275 79.150 2.415 ;
        RECT 79.290 2.225 79.365 2.365 ;
        RECT 79.995 2.285 80.055 2.365 ;
        POLYGON 79.995 2.285 80.055 2.285 80.055 2.225 ;
        RECT 80.210 2.275 80.285 2.415 ;
        RECT 81.975 2.275 82.050 2.415 ;
        RECT 82.190 2.225 82.265 2.365 ;
        RECT 82.895 2.285 82.955 2.365 ;
        POLYGON 82.895 2.285 82.955 2.285 82.955 2.225 ;
        RECT 83.110 2.275 83.185 2.415 ;
        RECT 84.875 2.275 84.950 2.415 ;
        RECT 85.090 2.225 85.165 2.365 ;
        RECT 85.795 2.285 85.855 2.365 ;
        POLYGON 85.795 2.285 85.855 2.285 85.855 2.225 ;
        RECT 86.010 2.275 86.085 2.415 ;
        RECT 87.775 2.275 87.850 2.415 ;
        RECT 87.990 2.225 88.065 2.365 ;
        RECT 88.695 2.285 88.755 2.365 ;
        POLYGON 88.695 2.285 88.755 2.285 88.755 2.225 ;
        RECT 88.910 2.275 88.985 2.415 ;
        RECT 90.675 2.275 90.750 2.415 ;
        RECT 90.890 2.225 90.965 2.365 ;
        RECT 91.595 2.285 91.655 2.365 ;
        POLYGON 91.595 2.285 91.655 2.285 91.655 2.225 ;
        RECT 91.810 2.275 91.885 2.415 ;
        RECT 0.720 1.750 0.870 1.920 ;
        RECT 1.110 1.885 1.260 2.055 ;
        RECT 1.500 1.885 1.650 2.055 ;
        RECT 1.890 1.750 2.040 1.920 ;
        RECT 3.620 1.750 3.770 1.920 ;
        RECT 4.010 1.885 4.160 2.055 ;
        RECT 4.400 1.885 4.550 2.055 ;
        RECT 4.790 1.750 4.940 1.920 ;
        RECT 6.520 1.750 6.670 1.920 ;
        RECT 6.910 1.885 7.060 2.055 ;
        RECT 7.300 1.885 7.450 2.055 ;
        RECT 7.690 1.750 7.840 1.920 ;
        RECT 9.420 1.750 9.570 1.920 ;
        RECT 9.810 1.885 9.960 2.055 ;
        RECT 10.200 1.885 10.350 2.055 ;
        RECT 10.590 1.750 10.740 1.920 ;
        RECT 12.320 1.750 12.470 1.920 ;
        RECT 12.710 1.885 12.860 2.055 ;
        RECT 13.100 1.885 13.250 2.055 ;
        RECT 13.490 1.750 13.640 1.920 ;
        RECT 15.220 1.750 15.370 1.920 ;
        RECT 15.610 1.885 15.760 2.055 ;
        RECT 16.000 1.885 16.150 2.055 ;
        RECT 16.390 1.750 16.540 1.920 ;
        RECT 18.120 1.750 18.270 1.920 ;
        RECT 18.510 1.885 18.660 2.055 ;
        RECT 18.900 1.885 19.050 2.055 ;
        RECT 19.290 1.750 19.440 1.920 ;
        RECT 21.020 1.750 21.170 1.920 ;
        RECT 21.410 1.885 21.560 2.055 ;
        RECT 21.800 1.885 21.950 2.055 ;
        RECT 22.190 1.750 22.340 1.920 ;
        RECT 23.920 1.755 24.070 1.925 ;
        RECT 24.310 1.890 24.460 2.060 ;
        RECT 24.700 1.890 24.850 2.060 ;
        RECT 25.090 1.755 25.240 1.925 ;
        RECT 26.820 1.755 26.970 1.925 ;
        RECT 27.210 1.890 27.360 2.060 ;
        RECT 27.600 1.890 27.750 2.060 ;
        RECT 27.990 1.755 28.140 1.925 ;
        RECT 29.720 1.755 29.870 1.925 ;
        RECT 30.110 1.890 30.260 2.060 ;
        RECT 30.500 1.890 30.650 2.060 ;
        RECT 30.890 1.755 31.040 1.925 ;
        RECT 32.620 1.755 32.770 1.925 ;
        RECT 33.010 1.890 33.160 2.060 ;
        RECT 33.400 1.890 33.550 2.060 ;
        RECT 33.790 1.755 33.940 1.925 ;
        RECT 35.520 1.755 35.670 1.925 ;
        RECT 35.910 1.890 36.060 2.060 ;
        RECT 36.300 1.890 36.450 2.060 ;
        RECT 36.690 1.755 36.840 1.925 ;
        RECT 38.420 1.755 38.570 1.925 ;
        RECT 38.810 1.890 38.960 2.060 ;
        RECT 39.200 1.890 39.350 2.060 ;
        RECT 39.590 1.755 39.740 1.925 ;
        RECT 41.320 1.755 41.470 1.925 ;
        RECT 41.710 1.890 41.860 2.060 ;
        RECT 42.100 1.890 42.250 2.060 ;
        RECT 42.490 1.755 42.640 1.925 ;
        RECT 44.220 1.755 44.370 1.925 ;
        RECT 44.610 1.890 44.760 2.060 ;
        RECT 45.000 1.890 45.150 2.060 ;
        RECT 45.390 1.755 45.540 1.925 ;
        RECT 47.120 1.755 47.270 1.925 ;
        RECT 47.510 1.890 47.660 2.060 ;
        RECT 47.900 1.890 48.050 2.060 ;
        RECT 48.290 1.755 48.440 1.925 ;
        RECT 50.020 1.755 50.170 1.925 ;
        RECT 50.410 1.890 50.560 2.060 ;
        RECT 50.800 1.890 50.950 2.060 ;
        RECT 51.190 1.755 51.340 1.925 ;
        RECT 52.920 1.755 53.070 1.925 ;
        RECT 53.310 1.890 53.460 2.060 ;
        RECT 53.700 1.890 53.850 2.060 ;
        RECT 54.090 1.755 54.240 1.925 ;
        RECT 55.820 1.755 55.970 1.925 ;
        RECT 56.210 1.890 56.360 2.060 ;
        RECT 56.600 1.890 56.750 2.060 ;
        RECT 56.990 1.755 57.140 1.925 ;
        RECT 58.720 1.755 58.870 1.925 ;
        RECT 59.110 1.890 59.260 2.060 ;
        RECT 59.500 1.890 59.650 2.060 ;
        RECT 59.890 1.755 60.040 1.925 ;
        RECT 61.620 1.755 61.770 1.925 ;
        RECT 62.010 1.890 62.160 2.060 ;
        RECT 62.400 1.890 62.550 2.060 ;
        RECT 62.790 1.755 62.940 1.925 ;
        RECT 64.520 1.755 64.670 1.925 ;
        RECT 64.910 1.890 65.060 2.060 ;
        RECT 65.300 1.890 65.450 2.060 ;
        RECT 65.690 1.755 65.840 1.925 ;
        RECT 67.420 1.755 67.570 1.925 ;
        RECT 67.810 1.890 67.960 2.060 ;
        RECT 68.200 1.890 68.350 2.060 ;
        RECT 68.590 1.755 68.740 1.925 ;
        RECT 70.320 1.755 70.470 1.925 ;
        RECT 70.710 1.890 70.860 2.060 ;
        RECT 71.100 1.890 71.250 2.060 ;
        RECT 71.490 1.755 71.640 1.925 ;
        RECT 73.220 1.755 73.370 1.925 ;
        RECT 73.610 1.890 73.760 2.060 ;
        RECT 74.000 1.890 74.150 2.060 ;
        RECT 74.390 1.755 74.540 1.925 ;
        RECT 76.120 1.755 76.270 1.925 ;
        RECT 76.510 1.890 76.660 2.060 ;
        RECT 76.900 1.890 77.050 2.060 ;
        RECT 77.290 1.755 77.440 1.925 ;
        RECT 79.020 1.755 79.170 1.925 ;
        RECT 79.410 1.890 79.560 2.060 ;
        RECT 79.800 1.890 79.950 2.060 ;
        RECT 80.190 1.755 80.340 1.925 ;
        RECT 81.920 1.755 82.070 1.925 ;
        RECT 82.310 1.890 82.460 2.060 ;
        RECT 82.700 1.890 82.850 2.060 ;
        RECT 83.090 1.755 83.240 1.925 ;
        RECT 84.820 1.755 84.970 1.925 ;
        RECT 85.210 1.890 85.360 2.060 ;
        RECT 85.600 1.890 85.750 2.060 ;
        RECT 85.990 1.755 86.140 1.925 ;
        RECT 87.720 1.755 87.870 1.925 ;
        RECT 88.110 1.890 88.260 2.060 ;
        RECT 88.500 1.890 88.650 2.060 ;
        RECT 88.890 1.755 89.040 1.925 ;
        RECT 90.620 1.755 90.770 1.925 ;
        RECT 91.010 1.890 91.160 2.060 ;
        RECT 91.400 1.890 91.550 2.060 ;
        RECT 91.790 1.755 91.940 1.925 ;
        RECT 0.985 1.665 1.035 1.700 ;
        POLYGON 1.035 1.700 1.070 1.665 1.035 1.665 ;
        RECT 0.985 1.540 1.070 1.665 ;
        RECT 1.690 1.540 1.775 1.700 ;
        RECT 3.885 1.665 3.935 1.700 ;
        POLYGON 3.935 1.700 3.970 1.665 3.935 1.665 ;
        RECT 3.885 1.540 3.970 1.665 ;
        RECT 4.590 1.540 4.675 1.700 ;
        RECT 6.785 1.665 6.835 1.700 ;
        POLYGON 6.835 1.700 6.870 1.665 6.835 1.665 ;
        RECT 6.785 1.540 6.870 1.665 ;
        RECT 7.490 1.540 7.575 1.700 ;
        RECT 9.685 1.665 9.735 1.700 ;
        POLYGON 9.735 1.700 9.770 1.665 9.735 1.665 ;
        RECT 9.685 1.540 9.770 1.665 ;
        RECT 10.390 1.540 10.475 1.700 ;
        RECT 12.585 1.665 12.635 1.700 ;
        POLYGON 12.635 1.700 12.670 1.665 12.635 1.665 ;
        RECT 12.585 1.540 12.670 1.665 ;
        RECT 13.290 1.540 13.375 1.700 ;
        RECT 15.485 1.665 15.535 1.700 ;
        POLYGON 15.535 1.700 15.570 1.665 15.535 1.665 ;
        RECT 15.485 1.540 15.570 1.665 ;
        RECT 16.190 1.540 16.275 1.700 ;
        RECT 18.385 1.665 18.435 1.700 ;
        POLYGON 18.435 1.700 18.470 1.665 18.435 1.665 ;
        RECT 18.385 1.540 18.470 1.665 ;
        RECT 19.090 1.540 19.175 1.700 ;
        RECT 21.285 1.665 21.335 1.700 ;
        POLYGON 21.335 1.700 21.370 1.665 21.335 1.665 ;
        RECT 21.285 1.540 21.370 1.665 ;
        RECT 21.990 1.540 22.075 1.700 ;
        RECT 24.185 1.670 24.235 1.705 ;
        POLYGON 24.235 1.705 24.270 1.670 24.235 1.670 ;
        RECT 24.185 1.545 24.270 1.670 ;
        RECT 24.890 1.545 24.975 1.705 ;
        RECT 27.085 1.670 27.135 1.705 ;
        POLYGON 27.135 1.705 27.170 1.670 27.135 1.670 ;
        RECT 27.085 1.545 27.170 1.670 ;
        RECT 27.790 1.545 27.875 1.705 ;
        RECT 29.985 1.670 30.035 1.705 ;
        POLYGON 30.035 1.705 30.070 1.670 30.035 1.670 ;
        RECT 29.985 1.545 30.070 1.670 ;
        RECT 30.690 1.545 30.775 1.705 ;
        RECT 32.885 1.670 32.935 1.705 ;
        POLYGON 32.935 1.705 32.970 1.670 32.935 1.670 ;
        RECT 32.885 1.545 32.970 1.670 ;
        RECT 33.590 1.545 33.675 1.705 ;
        RECT 35.785 1.670 35.835 1.705 ;
        POLYGON 35.835 1.705 35.870 1.670 35.835 1.670 ;
        RECT 35.785 1.545 35.870 1.670 ;
        RECT 36.490 1.545 36.575 1.705 ;
        RECT 38.685 1.670 38.735 1.705 ;
        POLYGON 38.735 1.705 38.770 1.670 38.735 1.670 ;
        RECT 38.685 1.545 38.770 1.670 ;
        RECT 39.390 1.545 39.475 1.705 ;
        RECT 41.585 1.670 41.635 1.705 ;
        POLYGON 41.635 1.705 41.670 1.670 41.635 1.670 ;
        RECT 41.585 1.545 41.670 1.670 ;
        RECT 42.290 1.545 42.375 1.705 ;
        RECT 44.485 1.670 44.535 1.705 ;
        POLYGON 44.535 1.705 44.570 1.670 44.535 1.670 ;
        RECT 44.485 1.545 44.570 1.670 ;
        RECT 45.190 1.545 45.275 1.705 ;
        RECT 47.385 1.670 47.435 1.705 ;
        POLYGON 47.435 1.705 47.470 1.670 47.435 1.670 ;
        RECT 47.385 1.545 47.470 1.670 ;
        RECT 48.090 1.545 48.175 1.705 ;
        RECT 50.285 1.670 50.335 1.705 ;
        POLYGON 50.335 1.705 50.370 1.670 50.335 1.670 ;
        RECT 50.285 1.545 50.370 1.670 ;
        RECT 50.990 1.545 51.075 1.705 ;
        RECT 53.185 1.670 53.235 1.705 ;
        POLYGON 53.235 1.705 53.270 1.670 53.235 1.670 ;
        RECT 53.185 1.545 53.270 1.670 ;
        RECT 53.890 1.545 53.975 1.705 ;
        RECT 56.085 1.670 56.135 1.705 ;
        POLYGON 56.135 1.705 56.170 1.670 56.135 1.670 ;
        RECT 56.085 1.545 56.170 1.670 ;
        RECT 56.790 1.545 56.875 1.705 ;
        RECT 58.985 1.670 59.035 1.705 ;
        POLYGON 59.035 1.705 59.070 1.670 59.035 1.670 ;
        RECT 58.985 1.545 59.070 1.670 ;
        RECT 59.690 1.545 59.775 1.705 ;
        RECT 61.885 1.670 61.935 1.705 ;
        POLYGON 61.935 1.705 61.970 1.670 61.935 1.670 ;
        RECT 61.885 1.545 61.970 1.670 ;
        RECT 62.590 1.545 62.675 1.705 ;
        RECT 64.785 1.670 64.835 1.705 ;
        POLYGON 64.835 1.705 64.870 1.670 64.835 1.670 ;
        RECT 64.785 1.545 64.870 1.670 ;
        RECT 65.490 1.545 65.575 1.705 ;
        RECT 67.685 1.670 67.735 1.705 ;
        POLYGON 67.735 1.705 67.770 1.670 67.735 1.670 ;
        RECT 67.685 1.545 67.770 1.670 ;
        RECT 68.390 1.545 68.475 1.705 ;
        RECT 70.585 1.670 70.635 1.705 ;
        POLYGON 70.635 1.705 70.670 1.670 70.635 1.670 ;
        RECT 70.585 1.545 70.670 1.670 ;
        RECT 71.290 1.545 71.375 1.705 ;
        RECT 73.485 1.670 73.535 1.705 ;
        POLYGON 73.535 1.705 73.570 1.670 73.535 1.670 ;
        RECT 73.485 1.545 73.570 1.670 ;
        RECT 74.190 1.545 74.275 1.705 ;
        RECT 76.385 1.670 76.435 1.705 ;
        POLYGON 76.435 1.705 76.470 1.670 76.435 1.670 ;
        RECT 76.385 1.545 76.470 1.670 ;
        RECT 77.090 1.545 77.175 1.705 ;
        RECT 79.285 1.670 79.335 1.705 ;
        POLYGON 79.335 1.705 79.370 1.670 79.335 1.670 ;
        RECT 79.285 1.545 79.370 1.670 ;
        RECT 79.990 1.545 80.075 1.705 ;
        RECT 82.185 1.670 82.235 1.705 ;
        POLYGON 82.235 1.705 82.270 1.670 82.235 1.670 ;
        RECT 82.185 1.545 82.270 1.670 ;
        RECT 82.890 1.545 82.975 1.705 ;
        RECT 85.085 1.670 85.135 1.705 ;
        POLYGON 85.135 1.705 85.170 1.670 85.135 1.670 ;
        RECT 85.085 1.545 85.170 1.670 ;
        RECT 85.790 1.545 85.875 1.705 ;
        RECT 87.985 1.670 88.035 1.705 ;
        POLYGON 88.035 1.705 88.070 1.670 88.035 1.670 ;
        RECT 87.985 1.545 88.070 1.670 ;
        RECT 88.690 1.545 88.775 1.705 ;
        RECT 90.885 1.670 90.935 1.705 ;
        POLYGON 90.935 1.705 90.970 1.670 90.935 1.670 ;
        RECT 90.885 1.545 90.970 1.670 ;
        RECT 91.590 1.545 91.675 1.705 ;
        RECT 0.775 0.920 0.850 1.060 ;
        RECT 0.990 0.870 1.065 1.010 ;
        RECT 1.695 0.930 1.755 1.010 ;
        POLYGON 1.695 0.930 1.755 0.930 1.755 0.870 ;
        RECT 1.910 0.920 1.985 1.060 ;
        RECT 3.675 0.920 3.750 1.060 ;
        RECT 3.890 0.870 3.965 1.010 ;
        RECT 4.595 0.930 4.655 1.010 ;
        POLYGON 4.595 0.930 4.655 0.930 4.655 0.870 ;
        RECT 4.810 0.920 4.885 1.060 ;
        RECT 6.575 0.920 6.650 1.060 ;
        RECT 6.790 0.870 6.865 1.010 ;
        RECT 7.495 0.930 7.555 1.010 ;
        POLYGON 7.495 0.930 7.555 0.930 7.555 0.870 ;
        RECT 7.710 0.920 7.785 1.060 ;
        RECT 9.475 0.920 9.550 1.060 ;
        RECT 9.690 0.870 9.765 1.010 ;
        RECT 10.395 0.930 10.455 1.010 ;
        POLYGON 10.395 0.930 10.455 0.930 10.455 0.870 ;
        RECT 10.610 0.920 10.685 1.060 ;
        RECT 12.375 0.920 12.450 1.060 ;
        RECT 12.590 0.870 12.665 1.010 ;
        RECT 13.295 0.930 13.355 1.010 ;
        POLYGON 13.295 0.930 13.355 0.930 13.355 0.870 ;
        RECT 13.510 0.920 13.585 1.060 ;
        RECT 15.275 0.920 15.350 1.060 ;
        RECT 15.490 0.870 15.565 1.010 ;
        RECT 16.195 0.930 16.255 1.010 ;
        POLYGON 16.195 0.930 16.255 0.930 16.255 0.870 ;
        RECT 16.410 0.920 16.485 1.060 ;
        RECT 18.175 0.920 18.250 1.060 ;
        RECT 18.390 0.870 18.465 1.010 ;
        RECT 19.095 0.930 19.155 1.010 ;
        POLYGON 19.095 0.930 19.155 0.930 19.155 0.870 ;
        RECT 19.310 0.920 19.385 1.060 ;
        RECT 21.075 0.920 21.150 1.060 ;
        RECT 21.290 0.870 21.365 1.010 ;
        RECT 21.995 0.930 22.055 1.010 ;
        POLYGON 21.995 0.930 22.055 0.930 22.055 0.870 ;
        RECT 22.210 0.920 22.285 1.060 ;
        RECT 23.975 0.925 24.050 1.065 ;
        RECT 24.190 0.875 24.265 1.015 ;
        RECT 24.895 0.935 24.955 1.015 ;
        POLYGON 24.895 0.935 24.955 0.935 24.955 0.875 ;
        RECT 25.110 0.925 25.185 1.065 ;
        RECT 26.875 0.925 26.950 1.065 ;
        RECT 27.090 0.875 27.165 1.015 ;
        RECT 27.795 0.935 27.855 1.015 ;
        POLYGON 27.795 0.935 27.855 0.935 27.855 0.875 ;
        RECT 28.010 0.925 28.085 1.065 ;
        RECT 29.775 0.925 29.850 1.065 ;
        RECT 29.990 0.875 30.065 1.015 ;
        RECT 30.695 0.935 30.755 1.015 ;
        POLYGON 30.695 0.935 30.755 0.935 30.755 0.875 ;
        RECT 30.910 0.925 30.985 1.065 ;
        RECT 32.675 0.925 32.750 1.065 ;
        RECT 32.890 0.875 32.965 1.015 ;
        RECT 33.595 0.935 33.655 1.015 ;
        POLYGON 33.595 0.935 33.655 0.935 33.655 0.875 ;
        RECT 33.810 0.925 33.885 1.065 ;
        RECT 35.575 0.925 35.650 1.065 ;
        RECT 35.790 0.875 35.865 1.015 ;
        RECT 36.495 0.935 36.555 1.015 ;
        POLYGON 36.495 0.935 36.555 0.935 36.555 0.875 ;
        RECT 36.710 0.925 36.785 1.065 ;
        RECT 38.475 0.925 38.550 1.065 ;
        RECT 38.690 0.875 38.765 1.015 ;
        RECT 39.395 0.935 39.455 1.015 ;
        POLYGON 39.395 0.935 39.455 0.935 39.455 0.875 ;
        RECT 39.610 0.925 39.685 1.065 ;
        RECT 41.375 0.925 41.450 1.065 ;
        RECT 41.590 0.875 41.665 1.015 ;
        RECT 42.295 0.935 42.355 1.015 ;
        POLYGON 42.295 0.935 42.355 0.935 42.355 0.875 ;
        RECT 42.510 0.925 42.585 1.065 ;
        RECT 44.275 0.925 44.350 1.065 ;
        RECT 44.490 0.875 44.565 1.015 ;
        RECT 45.195 0.935 45.255 1.015 ;
        POLYGON 45.195 0.935 45.255 0.935 45.255 0.875 ;
        RECT 45.410 0.925 45.485 1.065 ;
        RECT 47.175 0.925 47.250 1.065 ;
        RECT 47.390 0.875 47.465 1.015 ;
        RECT 48.095 0.935 48.155 1.015 ;
        POLYGON 48.095 0.935 48.155 0.935 48.155 0.875 ;
        RECT 48.310 0.925 48.385 1.065 ;
        RECT 50.075 0.925 50.150 1.065 ;
        RECT 50.290 0.875 50.365 1.015 ;
        RECT 50.995 0.935 51.055 1.015 ;
        POLYGON 50.995 0.935 51.055 0.935 51.055 0.875 ;
        RECT 51.210 0.925 51.285 1.065 ;
        RECT 52.975 0.925 53.050 1.065 ;
        RECT 53.190 0.875 53.265 1.015 ;
        RECT 53.895 0.935 53.955 1.015 ;
        POLYGON 53.895 0.935 53.955 0.935 53.955 0.875 ;
        RECT 54.110 0.925 54.185 1.065 ;
        RECT 55.875 0.925 55.950 1.065 ;
        RECT 56.090 0.875 56.165 1.015 ;
        RECT 56.795 0.935 56.855 1.015 ;
        POLYGON 56.795 0.935 56.855 0.935 56.855 0.875 ;
        RECT 57.010 0.925 57.085 1.065 ;
        RECT 58.775 0.925 58.850 1.065 ;
        RECT 58.990 0.875 59.065 1.015 ;
        RECT 59.695 0.935 59.755 1.015 ;
        POLYGON 59.695 0.935 59.755 0.935 59.755 0.875 ;
        RECT 59.910 0.925 59.985 1.065 ;
        RECT 61.675 0.925 61.750 1.065 ;
        RECT 61.890 0.875 61.965 1.015 ;
        RECT 62.595 0.935 62.655 1.015 ;
        POLYGON 62.595 0.935 62.655 0.935 62.655 0.875 ;
        RECT 62.810 0.925 62.885 1.065 ;
        RECT 64.575 0.925 64.650 1.065 ;
        RECT 64.790 0.875 64.865 1.015 ;
        RECT 65.495 0.935 65.555 1.015 ;
        POLYGON 65.495 0.935 65.555 0.935 65.555 0.875 ;
        RECT 65.710 0.925 65.785 1.065 ;
        RECT 67.475 0.925 67.550 1.065 ;
        RECT 67.690 0.875 67.765 1.015 ;
        RECT 68.395 0.935 68.455 1.015 ;
        POLYGON 68.395 0.935 68.455 0.935 68.455 0.875 ;
        RECT 68.610 0.925 68.685 1.065 ;
        RECT 70.375 0.925 70.450 1.065 ;
        RECT 70.590 0.875 70.665 1.015 ;
        RECT 71.295 0.935 71.355 1.015 ;
        POLYGON 71.295 0.935 71.355 0.935 71.355 0.875 ;
        RECT 71.510 0.925 71.585 1.065 ;
        RECT 73.275 0.925 73.350 1.065 ;
        RECT 73.490 0.875 73.565 1.015 ;
        RECT 74.195 0.935 74.255 1.015 ;
        POLYGON 74.195 0.935 74.255 0.935 74.255 0.875 ;
        RECT 74.410 0.925 74.485 1.065 ;
        RECT 76.175 0.925 76.250 1.065 ;
        RECT 76.390 0.875 76.465 1.015 ;
        RECT 77.095 0.935 77.155 1.015 ;
        POLYGON 77.095 0.935 77.155 0.935 77.155 0.875 ;
        RECT 77.310 0.925 77.385 1.065 ;
        RECT 79.075 0.925 79.150 1.065 ;
        RECT 79.290 0.875 79.365 1.015 ;
        RECT 79.995 0.935 80.055 1.015 ;
        POLYGON 79.995 0.935 80.055 0.935 80.055 0.875 ;
        RECT 80.210 0.925 80.285 1.065 ;
        RECT 81.975 0.925 82.050 1.065 ;
        RECT 82.190 0.875 82.265 1.015 ;
        RECT 82.895 0.935 82.955 1.015 ;
        POLYGON 82.895 0.935 82.955 0.935 82.955 0.875 ;
        RECT 83.110 0.925 83.185 1.065 ;
        RECT 84.875 0.925 84.950 1.065 ;
        RECT 85.090 0.875 85.165 1.015 ;
        RECT 85.795 0.935 85.855 1.015 ;
        POLYGON 85.795 0.935 85.855 0.935 85.855 0.875 ;
        RECT 86.010 0.925 86.085 1.065 ;
        RECT 87.775 0.925 87.850 1.065 ;
        RECT 87.990 0.875 88.065 1.015 ;
        RECT 88.695 0.935 88.755 1.015 ;
        POLYGON 88.695 0.935 88.755 0.935 88.755 0.875 ;
        RECT 88.910 0.925 88.985 1.065 ;
        RECT 90.675 0.925 90.750 1.065 ;
        RECT 90.890 0.875 90.965 1.015 ;
        RECT 91.595 0.935 91.655 1.015 ;
        POLYGON 91.595 0.935 91.655 0.935 91.655 0.875 ;
        RECT 91.810 0.925 91.885 1.065 ;
        RECT 0.720 0.400 0.870 0.570 ;
        RECT 1.110 0.535 1.260 0.705 ;
        RECT 1.500 0.535 1.650 0.705 ;
        RECT 1.890 0.400 2.040 0.570 ;
        RECT 3.620 0.400 3.770 0.570 ;
        RECT 4.010 0.535 4.160 0.705 ;
        RECT 4.400 0.535 4.550 0.705 ;
        RECT 4.790 0.400 4.940 0.570 ;
        RECT 6.520 0.400 6.670 0.570 ;
        RECT 6.910 0.535 7.060 0.705 ;
        RECT 7.300 0.535 7.450 0.705 ;
        RECT 7.690 0.400 7.840 0.570 ;
        RECT 9.420 0.400 9.570 0.570 ;
        RECT 9.810 0.535 9.960 0.705 ;
        RECT 10.200 0.535 10.350 0.705 ;
        RECT 10.590 0.400 10.740 0.570 ;
        RECT 12.320 0.400 12.470 0.570 ;
        RECT 12.710 0.535 12.860 0.705 ;
        RECT 13.100 0.535 13.250 0.705 ;
        RECT 13.490 0.400 13.640 0.570 ;
        RECT 15.220 0.400 15.370 0.570 ;
        RECT 15.610 0.535 15.760 0.705 ;
        RECT 16.000 0.535 16.150 0.705 ;
        RECT 16.390 0.400 16.540 0.570 ;
        RECT 18.120 0.400 18.270 0.570 ;
        RECT 18.510 0.535 18.660 0.705 ;
        RECT 18.900 0.535 19.050 0.705 ;
        RECT 19.290 0.400 19.440 0.570 ;
        RECT 21.020 0.400 21.170 0.570 ;
        RECT 21.410 0.535 21.560 0.705 ;
        RECT 21.800 0.535 21.950 0.705 ;
        RECT 22.190 0.400 22.340 0.570 ;
        RECT 23.920 0.405 24.070 0.575 ;
        RECT 24.310 0.540 24.460 0.710 ;
        RECT 24.700 0.540 24.850 0.710 ;
        RECT 25.090 0.405 25.240 0.575 ;
        RECT 26.820 0.405 26.970 0.575 ;
        RECT 27.210 0.540 27.360 0.710 ;
        RECT 27.600 0.540 27.750 0.710 ;
        RECT 27.990 0.405 28.140 0.575 ;
        RECT 29.720 0.405 29.870 0.575 ;
        RECT 30.110 0.540 30.260 0.710 ;
        RECT 30.500 0.540 30.650 0.710 ;
        RECT 30.890 0.405 31.040 0.575 ;
        RECT 32.620 0.405 32.770 0.575 ;
        RECT 33.010 0.540 33.160 0.710 ;
        RECT 33.400 0.540 33.550 0.710 ;
        RECT 33.790 0.405 33.940 0.575 ;
        RECT 35.520 0.405 35.670 0.575 ;
        RECT 35.910 0.540 36.060 0.710 ;
        RECT 36.300 0.540 36.450 0.710 ;
        RECT 36.690 0.405 36.840 0.575 ;
        RECT 38.420 0.405 38.570 0.575 ;
        RECT 38.810 0.540 38.960 0.710 ;
        RECT 39.200 0.540 39.350 0.710 ;
        RECT 39.590 0.405 39.740 0.575 ;
        RECT 41.320 0.405 41.470 0.575 ;
        RECT 41.710 0.540 41.860 0.710 ;
        RECT 42.100 0.540 42.250 0.710 ;
        RECT 42.490 0.405 42.640 0.575 ;
        RECT 44.220 0.405 44.370 0.575 ;
        RECT 44.610 0.540 44.760 0.710 ;
        RECT 45.000 0.540 45.150 0.710 ;
        RECT 45.390 0.405 45.540 0.575 ;
        RECT 47.120 0.405 47.270 0.575 ;
        RECT 47.510 0.540 47.660 0.710 ;
        RECT 47.900 0.540 48.050 0.710 ;
        RECT 48.290 0.405 48.440 0.575 ;
        RECT 50.020 0.405 50.170 0.575 ;
        RECT 50.410 0.540 50.560 0.710 ;
        RECT 50.800 0.540 50.950 0.710 ;
        RECT 51.190 0.405 51.340 0.575 ;
        RECT 52.920 0.405 53.070 0.575 ;
        RECT 53.310 0.540 53.460 0.710 ;
        RECT 53.700 0.540 53.850 0.710 ;
        RECT 54.090 0.405 54.240 0.575 ;
        RECT 55.820 0.405 55.970 0.575 ;
        RECT 56.210 0.540 56.360 0.710 ;
        RECT 56.600 0.540 56.750 0.710 ;
        RECT 56.990 0.405 57.140 0.575 ;
        RECT 58.720 0.405 58.870 0.575 ;
        RECT 59.110 0.540 59.260 0.710 ;
        RECT 59.500 0.540 59.650 0.710 ;
        RECT 59.890 0.405 60.040 0.575 ;
        RECT 61.620 0.405 61.770 0.575 ;
        RECT 62.010 0.540 62.160 0.710 ;
        RECT 62.400 0.540 62.550 0.710 ;
        RECT 62.790 0.405 62.940 0.575 ;
        RECT 64.520 0.405 64.670 0.575 ;
        RECT 64.910 0.540 65.060 0.710 ;
        RECT 65.300 0.540 65.450 0.710 ;
        RECT 65.690 0.405 65.840 0.575 ;
        RECT 67.420 0.405 67.570 0.575 ;
        RECT 67.810 0.540 67.960 0.710 ;
        RECT 68.200 0.540 68.350 0.710 ;
        RECT 68.590 0.405 68.740 0.575 ;
        RECT 70.320 0.405 70.470 0.575 ;
        RECT 70.710 0.540 70.860 0.710 ;
        RECT 71.100 0.540 71.250 0.710 ;
        RECT 71.490 0.405 71.640 0.575 ;
        RECT 73.220 0.405 73.370 0.575 ;
        RECT 73.610 0.540 73.760 0.710 ;
        RECT 74.000 0.540 74.150 0.710 ;
        RECT 74.390 0.405 74.540 0.575 ;
        RECT 76.120 0.405 76.270 0.575 ;
        RECT 76.510 0.540 76.660 0.710 ;
        RECT 76.900 0.540 77.050 0.710 ;
        RECT 77.290 0.405 77.440 0.575 ;
        RECT 79.020 0.405 79.170 0.575 ;
        RECT 79.410 0.540 79.560 0.710 ;
        RECT 79.800 0.540 79.950 0.710 ;
        RECT 80.190 0.405 80.340 0.575 ;
        RECT 81.920 0.405 82.070 0.575 ;
        RECT 82.310 0.540 82.460 0.710 ;
        RECT 82.700 0.540 82.850 0.710 ;
        RECT 83.090 0.405 83.240 0.575 ;
        RECT 84.820 0.405 84.970 0.575 ;
        RECT 85.210 0.540 85.360 0.710 ;
        RECT 85.600 0.540 85.750 0.710 ;
        RECT 85.990 0.405 86.140 0.575 ;
        RECT 87.720 0.405 87.870 0.575 ;
        RECT 88.110 0.540 88.260 0.710 ;
        RECT 88.500 0.540 88.650 0.710 ;
        RECT 88.890 0.405 89.040 0.575 ;
        RECT 90.620 0.405 90.770 0.575 ;
        RECT 91.010 0.540 91.160 0.710 ;
        RECT 91.400 0.540 91.550 0.710 ;
        RECT 91.790 0.405 91.940 0.575 ;
        RECT 0.985 0.315 1.035 0.350 ;
        POLYGON 1.035 0.350 1.070 0.315 1.035 0.315 ;
        RECT 0.985 0.190 1.070 0.315 ;
        RECT 1.690 0.190 1.775 0.350 ;
        RECT 3.885 0.315 3.935 0.350 ;
        POLYGON 3.935 0.350 3.970 0.315 3.935 0.315 ;
        RECT 3.885 0.190 3.970 0.315 ;
        RECT 4.590 0.190 4.675 0.350 ;
        RECT 6.785 0.315 6.835 0.350 ;
        POLYGON 6.835 0.350 6.870 0.315 6.835 0.315 ;
        RECT 6.785 0.190 6.870 0.315 ;
        RECT 7.490 0.190 7.575 0.350 ;
        RECT 9.685 0.315 9.735 0.350 ;
        POLYGON 9.735 0.350 9.770 0.315 9.735 0.315 ;
        RECT 9.685 0.190 9.770 0.315 ;
        RECT 10.390 0.190 10.475 0.350 ;
        RECT 12.585 0.315 12.635 0.350 ;
        POLYGON 12.635 0.350 12.670 0.315 12.635 0.315 ;
        RECT 12.585 0.190 12.670 0.315 ;
        RECT 13.290 0.190 13.375 0.350 ;
        RECT 15.485 0.315 15.535 0.350 ;
        POLYGON 15.535 0.350 15.570 0.315 15.535 0.315 ;
        RECT 15.485 0.190 15.570 0.315 ;
        RECT 16.190 0.190 16.275 0.350 ;
        RECT 18.385 0.315 18.435 0.350 ;
        POLYGON 18.435 0.350 18.470 0.315 18.435 0.315 ;
        RECT 18.385 0.190 18.470 0.315 ;
        RECT 19.090 0.190 19.175 0.350 ;
        RECT 21.285 0.315 21.335 0.350 ;
        POLYGON 21.335 0.350 21.370 0.315 21.335 0.315 ;
        RECT 21.285 0.190 21.370 0.315 ;
        RECT 21.990 0.190 22.075 0.350 ;
        RECT 24.185 0.320 24.235 0.355 ;
        POLYGON 24.235 0.355 24.270 0.320 24.235 0.320 ;
        RECT 24.185 0.195 24.270 0.320 ;
        RECT 24.890 0.195 24.975 0.355 ;
        RECT 27.085 0.320 27.135 0.355 ;
        POLYGON 27.135 0.355 27.170 0.320 27.135 0.320 ;
        RECT 27.085 0.195 27.170 0.320 ;
        RECT 27.790 0.195 27.875 0.355 ;
        RECT 29.985 0.320 30.035 0.355 ;
        POLYGON 30.035 0.355 30.070 0.320 30.035 0.320 ;
        RECT 29.985 0.195 30.070 0.320 ;
        RECT 30.690 0.195 30.775 0.355 ;
        RECT 32.885 0.320 32.935 0.355 ;
        POLYGON 32.935 0.355 32.970 0.320 32.935 0.320 ;
        RECT 32.885 0.195 32.970 0.320 ;
        RECT 33.590 0.195 33.675 0.355 ;
        RECT 35.785 0.320 35.835 0.355 ;
        POLYGON 35.835 0.355 35.870 0.320 35.835 0.320 ;
        RECT 35.785 0.195 35.870 0.320 ;
        RECT 36.490 0.195 36.575 0.355 ;
        RECT 38.685 0.320 38.735 0.355 ;
        POLYGON 38.735 0.355 38.770 0.320 38.735 0.320 ;
        RECT 38.685 0.195 38.770 0.320 ;
        RECT 39.390 0.195 39.475 0.355 ;
        RECT 41.585 0.320 41.635 0.355 ;
        POLYGON 41.635 0.355 41.670 0.320 41.635 0.320 ;
        RECT 41.585 0.195 41.670 0.320 ;
        RECT 42.290 0.195 42.375 0.355 ;
        RECT 44.485 0.320 44.535 0.355 ;
        POLYGON 44.535 0.355 44.570 0.320 44.535 0.320 ;
        RECT 44.485 0.195 44.570 0.320 ;
        RECT 45.190 0.195 45.275 0.355 ;
        RECT 47.385 0.320 47.435 0.355 ;
        POLYGON 47.435 0.355 47.470 0.320 47.435 0.320 ;
        RECT 47.385 0.195 47.470 0.320 ;
        RECT 48.090 0.195 48.175 0.355 ;
        RECT 50.285 0.320 50.335 0.355 ;
        POLYGON 50.335 0.355 50.370 0.320 50.335 0.320 ;
        RECT 50.285 0.195 50.370 0.320 ;
        RECT 50.990 0.195 51.075 0.355 ;
        RECT 53.185 0.320 53.235 0.355 ;
        POLYGON 53.235 0.355 53.270 0.320 53.235 0.320 ;
        RECT 53.185 0.195 53.270 0.320 ;
        RECT 53.890 0.195 53.975 0.355 ;
        RECT 56.085 0.320 56.135 0.355 ;
        POLYGON 56.135 0.355 56.170 0.320 56.135 0.320 ;
        RECT 56.085 0.195 56.170 0.320 ;
        RECT 56.790 0.195 56.875 0.355 ;
        RECT 58.985 0.320 59.035 0.355 ;
        POLYGON 59.035 0.355 59.070 0.320 59.035 0.320 ;
        RECT 58.985 0.195 59.070 0.320 ;
        RECT 59.690 0.195 59.775 0.355 ;
        RECT 61.885 0.320 61.935 0.355 ;
        POLYGON 61.935 0.355 61.970 0.320 61.935 0.320 ;
        RECT 61.885 0.195 61.970 0.320 ;
        RECT 62.590 0.195 62.675 0.355 ;
        RECT 64.785 0.320 64.835 0.355 ;
        POLYGON 64.835 0.355 64.870 0.320 64.835 0.320 ;
        RECT 64.785 0.195 64.870 0.320 ;
        RECT 65.490 0.195 65.575 0.355 ;
        RECT 67.685 0.320 67.735 0.355 ;
        POLYGON 67.735 0.355 67.770 0.320 67.735 0.320 ;
        RECT 67.685 0.195 67.770 0.320 ;
        RECT 68.390 0.195 68.475 0.355 ;
        RECT 70.585 0.320 70.635 0.355 ;
        POLYGON 70.635 0.355 70.670 0.320 70.635 0.320 ;
        RECT 70.585 0.195 70.670 0.320 ;
        RECT 71.290 0.195 71.375 0.355 ;
        RECT 73.485 0.320 73.535 0.355 ;
        POLYGON 73.535 0.355 73.570 0.320 73.535 0.320 ;
        RECT 73.485 0.195 73.570 0.320 ;
        RECT 74.190 0.195 74.275 0.355 ;
        RECT 76.385 0.320 76.435 0.355 ;
        POLYGON 76.435 0.355 76.470 0.320 76.435 0.320 ;
        RECT 76.385 0.195 76.470 0.320 ;
        RECT 77.090 0.195 77.175 0.355 ;
        RECT 79.285 0.320 79.335 0.355 ;
        POLYGON 79.335 0.355 79.370 0.320 79.335 0.320 ;
        RECT 79.285 0.195 79.370 0.320 ;
        RECT 79.990 0.195 80.075 0.355 ;
        RECT 82.185 0.320 82.235 0.355 ;
        POLYGON 82.235 0.355 82.270 0.320 82.235 0.320 ;
        RECT 82.185 0.195 82.270 0.320 ;
        RECT 82.890 0.195 82.975 0.355 ;
        RECT 85.085 0.320 85.135 0.355 ;
        POLYGON 85.135 0.355 85.170 0.320 85.135 0.320 ;
        RECT 85.085 0.195 85.170 0.320 ;
        RECT 85.790 0.195 85.875 0.355 ;
        RECT 87.985 0.320 88.035 0.355 ;
        POLYGON 88.035 0.355 88.070 0.320 88.035 0.320 ;
        RECT 87.985 0.195 88.070 0.320 ;
        RECT 88.690 0.195 88.775 0.355 ;
        RECT 90.885 0.320 90.935 0.355 ;
        POLYGON 90.935 0.355 90.970 0.320 90.935 0.320 ;
        RECT 90.885 0.195 90.970 0.320 ;
        RECT 91.590 0.195 91.675 0.355 ;
      LAYER met1 ;
        RECT 23.200 38.310 69.245 38.480 ;
        RECT 69.600 38.310 92.445 38.480 ;
  END
END 10T_32x32_magic_flattened
END LIBRARY

