magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< nwell >>
rect 0 0 720 806
<< pmos >>
rect 204 102 240 704
rect 296 102 332 704
rect 388 102 424 704
rect 480 102 516 704
<< pdiff >>
rect 148 692 204 704
rect 148 658 159 692
rect 193 658 204 692
rect 148 624 204 658
rect 148 590 159 624
rect 193 590 204 624
rect 148 556 204 590
rect 148 522 159 556
rect 193 522 204 556
rect 148 488 204 522
rect 148 454 159 488
rect 193 454 204 488
rect 148 420 204 454
rect 148 386 159 420
rect 193 386 204 420
rect 148 352 204 386
rect 148 318 159 352
rect 193 318 204 352
rect 148 284 204 318
rect 148 250 159 284
rect 193 250 204 284
rect 148 216 204 250
rect 148 182 159 216
rect 193 182 204 216
rect 148 148 204 182
rect 148 114 159 148
rect 193 114 204 148
rect 148 102 204 114
rect 240 692 296 704
rect 240 658 251 692
rect 285 658 296 692
rect 240 624 296 658
rect 240 590 251 624
rect 285 590 296 624
rect 240 556 296 590
rect 240 522 251 556
rect 285 522 296 556
rect 240 488 296 522
rect 240 454 251 488
rect 285 454 296 488
rect 240 420 296 454
rect 240 386 251 420
rect 285 386 296 420
rect 240 352 296 386
rect 240 318 251 352
rect 285 318 296 352
rect 240 284 296 318
rect 240 250 251 284
rect 285 250 296 284
rect 240 216 296 250
rect 240 182 251 216
rect 285 182 296 216
rect 240 148 296 182
rect 240 114 251 148
rect 285 114 296 148
rect 240 102 296 114
rect 332 692 388 704
rect 332 658 343 692
rect 377 658 388 692
rect 332 624 388 658
rect 332 590 343 624
rect 377 590 388 624
rect 332 556 388 590
rect 332 522 343 556
rect 377 522 388 556
rect 332 488 388 522
rect 332 454 343 488
rect 377 454 388 488
rect 332 420 388 454
rect 332 386 343 420
rect 377 386 388 420
rect 332 352 388 386
rect 332 318 343 352
rect 377 318 388 352
rect 332 284 388 318
rect 332 250 343 284
rect 377 250 388 284
rect 332 216 388 250
rect 332 182 343 216
rect 377 182 388 216
rect 332 148 388 182
rect 332 114 343 148
rect 377 114 388 148
rect 332 102 388 114
rect 424 692 480 704
rect 424 658 435 692
rect 469 658 480 692
rect 424 624 480 658
rect 424 590 435 624
rect 469 590 480 624
rect 424 556 480 590
rect 424 522 435 556
rect 469 522 480 556
rect 424 488 480 522
rect 424 454 435 488
rect 469 454 480 488
rect 424 420 480 454
rect 424 386 435 420
rect 469 386 480 420
rect 424 352 480 386
rect 424 318 435 352
rect 469 318 480 352
rect 424 284 480 318
rect 424 250 435 284
rect 469 250 480 284
rect 424 216 480 250
rect 424 182 435 216
rect 469 182 480 216
rect 424 148 480 182
rect 424 114 435 148
rect 469 114 480 148
rect 424 102 480 114
rect 516 692 572 704
rect 516 658 527 692
rect 561 658 572 692
rect 516 624 572 658
rect 516 590 527 624
rect 561 590 572 624
rect 516 556 572 590
rect 516 522 527 556
rect 561 522 572 556
rect 516 488 572 522
rect 516 454 527 488
rect 561 454 572 488
rect 516 420 572 454
rect 516 386 527 420
rect 561 386 572 420
rect 516 352 572 386
rect 516 318 527 352
rect 561 318 572 352
rect 516 284 572 318
rect 516 250 527 284
rect 561 250 572 284
rect 516 216 572 250
rect 516 182 527 216
rect 561 182 572 216
rect 516 148 572 182
rect 516 114 527 148
rect 561 114 572 148
rect 516 102 572 114
<< pdiffc >>
rect 159 658 193 692
rect 159 590 193 624
rect 159 522 193 556
rect 159 454 193 488
rect 159 386 193 420
rect 159 318 193 352
rect 159 250 193 284
rect 159 182 193 216
rect 159 114 193 148
rect 251 658 285 692
rect 251 590 285 624
rect 251 522 285 556
rect 251 454 285 488
rect 251 386 285 420
rect 251 318 285 352
rect 251 250 285 284
rect 251 182 285 216
rect 251 114 285 148
rect 343 658 377 692
rect 343 590 377 624
rect 343 522 377 556
rect 343 454 377 488
rect 343 386 377 420
rect 343 318 377 352
rect 343 250 377 284
rect 343 182 377 216
rect 343 114 377 148
rect 435 658 469 692
rect 435 590 469 624
rect 435 522 469 556
rect 435 454 469 488
rect 435 386 469 420
rect 435 318 469 352
rect 435 250 469 284
rect 435 182 469 216
rect 435 114 469 148
rect 527 658 561 692
rect 527 590 561 624
rect 527 522 561 556
rect 527 454 561 488
rect 527 386 561 420
rect 527 318 561 352
rect 527 250 561 284
rect 527 182 561 216
rect 527 114 561 148
<< nsubdiff >>
rect 36 658 94 704
rect 36 624 48 658
rect 82 624 94 658
rect 36 590 94 624
rect 36 556 48 590
rect 82 556 94 590
rect 36 522 94 556
rect 36 488 48 522
rect 82 488 94 522
rect 36 454 94 488
rect 36 420 48 454
rect 82 420 94 454
rect 36 386 94 420
rect 36 352 48 386
rect 82 352 94 386
rect 36 318 94 352
rect 36 284 48 318
rect 82 284 94 318
rect 36 250 94 284
rect 36 216 48 250
rect 82 216 94 250
rect 36 182 94 216
rect 36 148 48 182
rect 82 148 94 182
rect 36 102 94 148
rect 626 658 684 704
rect 626 624 638 658
rect 672 624 684 658
rect 626 590 684 624
rect 626 556 638 590
rect 672 556 684 590
rect 626 522 684 556
rect 626 488 638 522
rect 672 488 684 522
rect 626 454 684 488
rect 626 420 638 454
rect 672 420 684 454
rect 626 386 684 420
rect 626 352 638 386
rect 672 352 684 386
rect 626 318 684 352
rect 626 284 638 318
rect 672 284 684 318
rect 626 250 684 284
rect 626 216 638 250
rect 672 216 684 250
rect 626 182 684 216
rect 626 148 638 182
rect 672 148 684 182
rect 626 102 684 148
<< nsubdiffcont >>
rect 48 624 82 658
rect 48 556 82 590
rect 48 488 82 522
rect 48 420 82 454
rect 48 352 82 386
rect 48 284 82 318
rect 48 216 82 250
rect 48 148 82 182
rect 638 624 672 658
rect 638 556 672 590
rect 638 488 672 522
rect 638 420 672 454
rect 638 352 672 386
rect 638 284 672 318
rect 638 216 672 250
rect 638 148 672 182
<< poly >>
rect 191 786 529 806
rect 191 752 207 786
rect 241 752 275 786
rect 309 752 343 786
rect 377 752 411 786
rect 445 752 479 786
rect 513 752 529 786
rect 191 736 529 752
rect 204 704 240 736
rect 296 704 332 736
rect 388 704 424 736
rect 480 704 516 736
rect 204 70 240 102
rect 296 70 332 102
rect 388 70 424 102
rect 480 70 516 102
rect 191 54 529 70
rect 191 20 207 54
rect 241 20 275 54
rect 309 20 343 54
rect 377 20 411 54
rect 445 20 479 54
rect 513 20 529 54
rect 191 0 529 20
<< polycont >>
rect 207 752 241 786
rect 275 752 309 786
rect 343 752 377 786
rect 411 752 445 786
rect 479 752 513 786
rect 207 20 241 54
rect 275 20 309 54
rect 343 20 377 54
rect 411 20 445 54
rect 479 20 513 54
<< locali >>
rect 191 752 199 786
rect 241 752 271 786
rect 309 752 343 786
rect 377 752 411 786
rect 449 752 479 786
rect 521 752 529 786
rect 159 692 193 708
rect 48 672 82 674
rect 48 600 82 624
rect 48 528 82 556
rect 48 456 82 488
rect 48 386 82 420
rect 48 318 82 350
rect 48 250 82 278
rect 48 182 82 206
rect 48 132 82 134
rect 159 624 193 638
rect 159 556 193 566
rect 159 488 193 494
rect 159 420 193 422
rect 159 384 193 386
rect 159 312 193 318
rect 159 240 193 250
rect 159 168 193 182
rect 159 98 193 114
rect 251 692 285 708
rect 251 624 285 638
rect 251 556 285 566
rect 251 488 285 494
rect 251 420 285 422
rect 251 384 285 386
rect 251 312 285 318
rect 251 240 285 250
rect 251 168 285 182
rect 251 98 285 114
rect 343 692 377 708
rect 343 624 377 638
rect 343 556 377 566
rect 343 488 377 494
rect 343 420 377 422
rect 343 384 377 386
rect 343 312 377 318
rect 343 240 377 250
rect 343 168 377 182
rect 343 98 377 114
rect 435 692 469 708
rect 435 624 469 638
rect 435 556 469 566
rect 435 488 469 494
rect 435 420 469 422
rect 435 384 469 386
rect 435 312 469 318
rect 435 240 469 250
rect 435 168 469 182
rect 435 98 469 114
rect 527 692 561 708
rect 527 624 561 638
rect 527 556 561 566
rect 527 488 561 494
rect 527 420 561 422
rect 527 384 561 386
rect 527 312 561 318
rect 527 240 561 250
rect 527 168 561 182
rect 638 672 672 674
rect 638 600 672 624
rect 638 528 672 556
rect 638 456 672 488
rect 638 386 672 420
rect 638 318 672 350
rect 638 250 672 278
rect 638 182 672 206
rect 638 132 672 134
rect 527 98 561 114
rect 191 20 199 54
rect 241 20 271 54
rect 309 20 343 54
rect 377 20 411 54
rect 449 20 479 54
rect 521 20 529 54
<< viali >>
rect 199 752 207 786
rect 207 752 233 786
rect 271 752 275 786
rect 275 752 305 786
rect 343 752 377 786
rect 415 752 445 786
rect 445 752 449 786
rect 487 752 513 786
rect 513 752 521 786
rect 48 658 82 672
rect 48 638 82 658
rect 48 590 82 600
rect 48 566 82 590
rect 48 522 82 528
rect 48 494 82 522
rect 48 454 82 456
rect 48 422 82 454
rect 48 352 82 384
rect 48 350 82 352
rect 48 284 82 312
rect 48 278 82 284
rect 48 216 82 240
rect 48 206 82 216
rect 48 148 82 168
rect 48 134 82 148
rect 159 658 193 672
rect 159 638 193 658
rect 159 590 193 600
rect 159 566 193 590
rect 159 522 193 528
rect 159 494 193 522
rect 159 454 193 456
rect 159 422 193 454
rect 159 352 193 384
rect 159 350 193 352
rect 159 284 193 312
rect 159 278 193 284
rect 159 216 193 240
rect 159 206 193 216
rect 159 148 193 168
rect 159 134 193 148
rect 251 658 285 672
rect 251 638 285 658
rect 251 590 285 600
rect 251 566 285 590
rect 251 522 285 528
rect 251 494 285 522
rect 251 454 285 456
rect 251 422 285 454
rect 251 352 285 384
rect 251 350 285 352
rect 251 284 285 312
rect 251 278 285 284
rect 251 216 285 240
rect 251 206 285 216
rect 251 148 285 168
rect 251 134 285 148
rect 343 658 377 672
rect 343 638 377 658
rect 343 590 377 600
rect 343 566 377 590
rect 343 522 377 528
rect 343 494 377 522
rect 343 454 377 456
rect 343 422 377 454
rect 343 352 377 384
rect 343 350 377 352
rect 343 284 377 312
rect 343 278 377 284
rect 343 216 377 240
rect 343 206 377 216
rect 343 148 377 168
rect 343 134 377 148
rect 435 658 469 672
rect 435 638 469 658
rect 435 590 469 600
rect 435 566 469 590
rect 435 522 469 528
rect 435 494 469 522
rect 435 454 469 456
rect 435 422 469 454
rect 435 352 469 384
rect 435 350 469 352
rect 435 284 469 312
rect 435 278 469 284
rect 435 216 469 240
rect 435 206 469 216
rect 435 148 469 168
rect 435 134 469 148
rect 527 658 561 672
rect 527 638 561 658
rect 527 590 561 600
rect 527 566 561 590
rect 527 522 561 528
rect 527 494 561 522
rect 527 454 561 456
rect 527 422 561 454
rect 527 352 561 384
rect 527 350 561 352
rect 527 284 561 312
rect 527 278 561 284
rect 527 216 561 240
rect 527 206 561 216
rect 527 148 561 168
rect 527 134 561 148
rect 638 658 672 672
rect 638 638 672 658
rect 638 590 672 600
rect 638 566 672 590
rect 638 522 672 528
rect 638 494 672 522
rect 638 454 672 456
rect 638 422 672 454
rect 638 352 672 384
rect 638 350 672 352
rect 638 284 672 312
rect 638 278 672 284
rect 638 216 672 240
rect 638 206 672 216
rect 638 148 672 168
rect 638 134 672 148
rect 199 20 207 54
rect 207 20 233 54
rect 271 20 275 54
rect 275 20 305 54
rect 343 20 377 54
rect 415 20 445 54
rect 445 20 449 54
rect 487 20 513 54
rect 513 20 521 54
<< metal1 >>
rect 187 786 533 806
rect 187 752 199 786
rect 233 752 271 786
rect 305 752 343 786
rect 377 752 415 786
rect 449 752 487 786
rect 521 752 533 786
rect 187 740 533 752
rect 36 672 94 684
rect 36 638 48 672
rect 82 638 94 672
rect 36 600 94 638
rect 36 566 48 600
rect 82 566 94 600
rect 36 528 94 566
rect 36 494 48 528
rect 82 494 94 528
rect 36 456 94 494
rect 36 422 48 456
rect 82 422 94 456
rect 36 384 94 422
rect 36 350 48 384
rect 82 350 94 384
rect 36 312 94 350
rect 36 278 48 312
rect 82 278 94 312
rect 36 240 94 278
rect 36 206 48 240
rect 82 206 94 240
rect 36 168 94 206
rect 36 134 48 168
rect 82 134 94 168
rect 36 122 94 134
rect 150 672 202 684
rect 150 638 159 672
rect 193 638 202 672
rect 150 600 202 638
rect 150 566 159 600
rect 193 566 202 600
rect 150 528 202 566
rect 150 494 159 528
rect 193 494 202 528
rect 150 456 202 494
rect 150 422 159 456
rect 193 422 202 456
rect 150 384 202 422
rect 150 372 159 384
rect 193 372 202 384
rect 150 312 202 320
rect 150 308 159 312
rect 193 308 202 312
rect 150 244 202 256
rect 150 180 202 192
rect 150 122 202 128
rect 242 678 294 684
rect 242 614 294 626
rect 242 550 294 562
rect 242 494 251 498
rect 285 494 294 498
rect 242 486 294 494
rect 242 422 251 434
rect 285 422 294 434
rect 242 384 294 422
rect 242 350 251 384
rect 285 350 294 384
rect 242 312 294 350
rect 242 278 251 312
rect 285 278 294 312
rect 242 240 294 278
rect 242 206 251 240
rect 285 206 294 240
rect 242 168 294 206
rect 242 134 251 168
rect 285 134 294 168
rect 242 122 294 134
rect 334 672 386 684
rect 334 638 343 672
rect 377 638 386 672
rect 334 600 386 638
rect 334 566 343 600
rect 377 566 386 600
rect 334 528 386 566
rect 334 494 343 528
rect 377 494 386 528
rect 334 456 386 494
rect 334 422 343 456
rect 377 422 386 456
rect 334 384 386 422
rect 334 372 343 384
rect 377 372 386 384
rect 334 312 386 320
rect 334 308 343 312
rect 377 308 386 312
rect 334 244 386 256
rect 334 180 386 192
rect 334 122 386 128
rect 426 678 478 684
rect 426 614 478 626
rect 426 550 478 562
rect 426 494 435 498
rect 469 494 478 498
rect 426 486 478 494
rect 426 422 435 434
rect 469 422 478 434
rect 426 384 478 422
rect 426 350 435 384
rect 469 350 478 384
rect 426 312 478 350
rect 426 278 435 312
rect 469 278 478 312
rect 426 240 478 278
rect 426 206 435 240
rect 469 206 478 240
rect 426 168 478 206
rect 426 134 435 168
rect 469 134 478 168
rect 426 122 478 134
rect 518 672 570 684
rect 518 638 527 672
rect 561 638 570 672
rect 518 600 570 638
rect 518 566 527 600
rect 561 566 570 600
rect 518 528 570 566
rect 518 494 527 528
rect 561 494 570 528
rect 518 456 570 494
rect 518 422 527 456
rect 561 422 570 456
rect 518 384 570 422
rect 518 372 527 384
rect 561 372 570 384
rect 518 312 570 320
rect 518 308 527 312
rect 561 308 570 312
rect 518 244 570 256
rect 518 180 570 192
rect 518 122 570 128
rect 626 672 684 684
rect 626 638 638 672
rect 672 638 684 672
rect 626 600 684 638
rect 626 566 638 600
rect 672 566 684 600
rect 626 528 684 566
rect 626 494 638 528
rect 672 494 684 528
rect 626 456 684 494
rect 626 422 638 456
rect 672 422 684 456
rect 626 384 684 422
rect 626 350 638 384
rect 672 350 684 384
rect 626 312 684 350
rect 626 278 638 312
rect 672 278 684 312
rect 626 240 684 278
rect 626 206 638 240
rect 672 206 684 240
rect 626 168 684 206
rect 626 134 638 168
rect 672 134 684 168
rect 626 122 684 134
rect 187 54 533 66
rect 187 20 199 54
rect 233 20 271 54
rect 305 20 343 54
rect 377 20 415 54
rect 449 20 487 54
rect 521 20 533 54
rect 187 0 533 20
<< via1 >>
rect 150 350 159 372
rect 159 350 193 372
rect 193 350 202 372
rect 150 320 202 350
rect 150 278 159 308
rect 159 278 193 308
rect 193 278 202 308
rect 150 256 202 278
rect 150 240 202 244
rect 150 206 159 240
rect 159 206 193 240
rect 193 206 202 240
rect 150 192 202 206
rect 150 168 202 180
rect 150 134 159 168
rect 159 134 193 168
rect 193 134 202 168
rect 150 128 202 134
rect 242 672 294 678
rect 242 638 251 672
rect 251 638 285 672
rect 285 638 294 672
rect 242 626 294 638
rect 242 600 294 614
rect 242 566 251 600
rect 251 566 285 600
rect 285 566 294 600
rect 242 562 294 566
rect 242 528 294 550
rect 242 498 251 528
rect 251 498 285 528
rect 285 498 294 528
rect 242 456 294 486
rect 242 434 251 456
rect 251 434 285 456
rect 285 434 294 456
rect 334 350 343 372
rect 343 350 377 372
rect 377 350 386 372
rect 334 320 386 350
rect 334 278 343 308
rect 343 278 377 308
rect 377 278 386 308
rect 334 256 386 278
rect 334 240 386 244
rect 334 206 343 240
rect 343 206 377 240
rect 377 206 386 240
rect 334 192 386 206
rect 334 168 386 180
rect 334 134 343 168
rect 343 134 377 168
rect 377 134 386 168
rect 334 128 386 134
rect 426 672 478 678
rect 426 638 435 672
rect 435 638 469 672
rect 469 638 478 672
rect 426 626 478 638
rect 426 600 478 614
rect 426 566 435 600
rect 435 566 469 600
rect 469 566 478 600
rect 426 562 478 566
rect 426 528 478 550
rect 426 498 435 528
rect 435 498 469 528
rect 469 498 478 528
rect 426 456 478 486
rect 426 434 435 456
rect 435 434 469 456
rect 469 434 478 456
rect 518 350 527 372
rect 527 350 561 372
rect 561 350 570 372
rect 518 320 570 350
rect 518 278 527 308
rect 527 278 561 308
rect 561 278 570 308
rect 518 256 570 278
rect 518 240 570 244
rect 518 206 527 240
rect 527 206 561 240
rect 561 206 570 240
rect 518 192 570 206
rect 518 168 570 180
rect 518 134 527 168
rect 527 134 561 168
rect 561 134 570 168
rect 518 128 570 134
<< metal2 >>
rect 10 678 710 684
rect 10 626 242 678
rect 294 626 426 678
rect 478 626 710 678
rect 10 614 710 626
rect 10 562 242 614
rect 294 562 426 614
rect 478 562 710 614
rect 10 550 710 562
rect 10 498 242 550
rect 294 498 426 550
rect 478 498 710 550
rect 10 486 710 498
rect 10 434 242 486
rect 294 434 426 486
rect 478 434 710 486
rect 10 428 710 434
rect 10 372 710 378
rect 10 320 150 372
rect 202 320 334 372
rect 386 320 518 372
rect 570 320 710 372
rect 10 308 710 320
rect 10 256 150 308
rect 202 256 334 308
rect 386 256 518 308
rect 570 256 710 308
rect 10 244 710 256
rect 10 192 150 244
rect 202 192 334 244
rect 386 192 518 244
rect 570 192 710 244
rect 10 180 710 192
rect 10 128 150 180
rect 202 128 334 180
rect 386 128 518 180
rect 570 128 710 180
rect 10 122 710 128
<< labels >>
flabel comment s 176 403 176 403 0 FreeSans 300 0 0 0 S
flabel comment s 268 403 268 403 0 FreeSans 300 0 0 0 S
flabel comment s 360 403 360 403 0 FreeSans 300 0 0 0 S
flabel comment s 452 403 452 403 0 FreeSans 300 0 0 0 S
flabel comment s 176 403 176 403 0 FreeSans 300 0 0 0 S
flabel comment s 268 403 268 403 0 FreeSans 300 0 0 0 D
flabel comment s 360 403 360 403 0 FreeSans 300 0 0 0 S
flabel comment s 452 403 452 403 0 FreeSans 300 0 0 0 D
flabel comment s 544 403 544 403 0 FreeSans 300 0 0 0 S
flabel metal1 s 321 762 379 787 0 FreeSans 100 0 0 0 GATE
port 3 nsew
flabel metal1 s 341 22 399 47 0 FreeSans 100 0 0 0 GATE
port 3 nsew
flabel metal1 s 638 396 672 407 0 FreeSans 100 0 0 0 BULK
port 1 nsew
flabel metal1 s 49 396 83 407 0 FreeSans 100 0 0 0 BULK
port 1 nsew
flabel metal2 s 54 540 69 606 0 FreeSans 100 0 0 0 DRAIN
port 2 nsew
flabel metal2 s 56 231 70 294 0 FreeSans 100 0 0 0 SOURCE
port 4 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 9538682
string GDS_START 9523116
<< end >>
