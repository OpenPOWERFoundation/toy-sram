`timescale 1 ps / 1 ps

module sky130_fd_pr__pfet_01v8 (
    input G,
    input D
);

endmodule
