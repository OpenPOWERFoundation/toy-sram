magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< pwell >>
rect 78 371 89 386
<< obsli1 >>
rect 137 447 679 463
rect 137 413 139 447
rect 173 413 211 447
rect 245 413 283 447
rect 317 413 355 447
rect 389 413 427 447
rect 461 413 499 447
rect 533 413 571 447
rect 605 413 643 447
rect 677 413 679 447
rect 137 397 679 413
rect 47 329 81 357
rect 47 257 81 295
rect 47 185 81 223
rect 47 113 81 151
rect 47 51 81 79
rect 133 51 167 357
rect 219 329 253 357
rect 219 257 253 295
rect 219 185 253 223
rect 219 113 253 151
rect 219 51 253 79
rect 305 51 339 357
rect 391 329 425 357
rect 391 257 425 295
rect 391 185 425 223
rect 391 113 425 151
rect 391 51 425 79
rect 477 51 511 357
rect 563 329 597 357
rect 563 257 597 295
rect 563 185 597 223
rect 563 113 597 151
rect 563 51 597 79
rect 649 51 683 357
rect 735 329 769 357
rect 735 257 769 295
rect 735 185 769 223
rect 735 113 769 151
rect 735 51 769 79
<< obsli1c >>
rect 139 413 173 447
rect 211 413 245 447
rect 283 413 317 447
rect 355 413 389 447
rect 427 413 461 447
rect 499 413 533 447
rect 571 413 605 447
rect 643 413 677 447
rect 47 295 81 329
rect 47 223 81 257
rect 47 151 81 185
rect 47 79 81 113
rect 219 295 253 329
rect 219 223 253 257
rect 219 151 253 185
rect 219 79 253 113
rect 391 295 425 329
rect 391 223 425 257
rect 391 151 425 185
rect 391 79 425 113
rect 563 295 597 329
rect 563 223 597 257
rect 563 151 597 185
rect 563 79 597 113
rect 735 295 769 329
rect 735 223 769 257
rect 735 151 769 185
rect 735 79 769 113
<< metal1 >>
rect 127 447 689 459
rect 127 413 139 447
rect 173 413 211 447
rect 245 413 283 447
rect 317 413 355 447
rect 389 413 427 447
rect 461 413 499 447
rect 533 413 571 447
rect 605 413 643 447
rect 677 413 689 447
rect 127 401 689 413
rect 41 329 87 357
rect 41 295 47 329
rect 81 295 87 329
rect 41 257 87 295
rect 41 223 47 257
rect 81 223 87 257
rect 41 185 87 223
rect 41 151 47 185
rect 81 151 87 185
rect 41 113 87 151
rect 41 79 47 113
rect 81 79 87 113
rect 41 -29 87 79
rect 213 329 259 357
rect 213 295 219 329
rect 253 295 259 329
rect 213 257 259 295
rect 213 223 219 257
rect 253 223 259 257
rect 213 185 259 223
rect 213 151 219 185
rect 253 151 259 185
rect 213 113 259 151
rect 213 79 219 113
rect 253 79 259 113
rect 213 -29 259 79
rect 385 329 431 357
rect 385 295 391 329
rect 425 295 431 329
rect 385 257 431 295
rect 385 223 391 257
rect 425 223 431 257
rect 385 185 431 223
rect 385 151 391 185
rect 425 151 431 185
rect 385 113 431 151
rect 385 79 391 113
rect 425 79 431 113
rect 385 -29 431 79
rect 557 329 603 357
rect 557 295 563 329
rect 597 295 603 329
rect 557 257 603 295
rect 557 223 563 257
rect 597 223 603 257
rect 557 185 603 223
rect 557 151 563 185
rect 597 151 603 185
rect 557 113 603 151
rect 557 79 563 113
rect 597 79 603 113
rect 557 -29 603 79
rect 729 329 775 357
rect 729 295 735 329
rect 769 295 775 329
rect 729 257 775 295
rect 729 223 735 257
rect 769 223 775 257
rect 729 185 775 223
rect 729 151 735 185
rect 769 151 775 185
rect 729 113 775 151
rect 729 79 735 113
rect 769 79 775 113
rect 729 -29 775 79
rect 41 -89 775 -29
<< obsm1 >>
rect 124 51 176 357
rect 296 51 348 357
rect 468 51 520 357
rect 640 51 692 357
<< obsm2 >>
rect 117 203 183 357
rect 289 203 355 357
rect 461 203 527 357
rect 633 203 699 357
<< metal3 >>
rect 117 291 699 357
rect 117 203 183 291
rect 289 203 355 291
rect 461 203 527 291
rect 633 203 699 291
<< labels >>
rlabel metal3 s 633 203 699 291 6 DRAIN
port 1 nsew
rlabel metal3 s 461 203 527 291 6 DRAIN
port 1 nsew
rlabel metal3 s 289 203 355 291 6 DRAIN
port 1 nsew
rlabel metal3 s 117 291 699 357 6 DRAIN
port 1 nsew
rlabel metal3 s 117 203 183 291 6 DRAIN
port 1 nsew
rlabel metal1 s 127 401 689 459 6 GATE
port 2 nsew
rlabel metal1 s 729 -29 775 357 6 SOURCE
port 3 nsew
rlabel metal1 s 557 -29 603 357 6 SOURCE
port 3 nsew
rlabel metal1 s 385 -29 431 357 6 SOURCE
port 3 nsew
rlabel metal1 s 213 -29 259 357 6 SOURCE
port 3 nsew
rlabel metal1 s 41 -29 87 357 6 SOURCE
port 3 nsew
rlabel metal1 s 41 -89 775 -29 8 SOURCE
port 3 nsew
rlabel pwell s 78 371 89 386 6 SUBSTRATE
port 4 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 36 -89 780 463
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 5929566
string GDS_START 5915584
<< end >>
