magic
tech sky130A
magscale 1 2
timestamp 1658882323
<< error_s >>
rect 15 8624 28 8640
rect 83 8624 98 8638
rect 117 8626 130 8640
rect 198 8636 351 8682
rect 180 8624 372 8636
rect 451 8624 464 8640
rect 546 8624 565 8640
rect 580 8624 586 8640
rect 595 8624 608 8640
rect 663 8624 678 8638
rect 697 8626 710 8640
rect 778 8636 931 8682
rect 760 8624 952 8636
rect 1031 8624 1044 8640
rect 1126 8624 1145 8640
rect 1160 8624 1166 8640
rect 1175 8624 1188 8640
rect 1243 8624 1258 8638
rect 1277 8626 1290 8640
rect 1358 8636 1511 8682
rect 1340 8624 1532 8636
rect 1611 8624 1624 8640
rect 1706 8624 1725 8640
rect 1740 8624 1746 8640
rect 1755 8624 1768 8640
rect 1823 8624 1838 8638
rect 1857 8626 1870 8640
rect 1938 8636 2091 8682
rect 1920 8624 2112 8636
rect 2191 8624 2204 8640
rect 2286 8624 2305 8640
rect 2320 8624 2326 8640
rect 2335 8624 2348 8640
rect 2403 8624 2418 8638
rect 2437 8626 2450 8640
rect 2518 8636 2671 8682
rect 2500 8624 2692 8636
rect 2771 8624 2784 8640
rect 2866 8624 2885 8640
rect 2900 8624 2906 8640
rect 2915 8624 2928 8640
rect 2983 8624 2998 8638
rect 3017 8626 3030 8640
rect 3098 8636 3251 8682
rect 3080 8624 3272 8636
rect 3351 8624 3364 8640
rect 3446 8624 3465 8640
rect 3480 8624 3486 8640
rect 3495 8624 3508 8640
rect 3563 8624 3578 8638
rect 3597 8626 3610 8640
rect 3678 8636 3831 8682
rect 3660 8624 3852 8636
rect 3931 8624 3944 8640
rect 4026 8624 4045 8640
rect 4060 8624 4066 8640
rect 4075 8624 4088 8640
rect 4143 8624 4158 8638
rect 4177 8626 4190 8640
rect 4258 8636 4411 8682
rect 4240 8624 4432 8636
rect 4511 8624 4524 8640
rect 4606 8624 4625 8640
rect 4640 8624 4646 8640
rect 4655 8624 4668 8640
rect 4723 8624 4738 8638
rect 4757 8626 4770 8640
rect 4838 8636 4991 8682
rect 4820 8624 5012 8636
rect 5091 8624 5104 8640
rect 5186 8624 5205 8640
rect 5220 8624 5226 8640
rect 5235 8624 5248 8640
rect 5303 8624 5318 8638
rect 5337 8626 5350 8640
rect 5418 8636 5571 8682
rect 5400 8624 5592 8636
rect 5671 8624 5684 8640
rect 5766 8624 5785 8640
rect 5800 8624 5806 8640
rect 5815 8624 5828 8640
rect 5883 8624 5898 8638
rect 5917 8626 5930 8640
rect 5998 8636 6151 8682
rect 5980 8624 6172 8636
rect 6251 8624 6264 8640
rect 6346 8624 6365 8640
rect 6380 8624 6386 8640
rect 6395 8624 6408 8640
rect 6463 8624 6478 8638
rect 6497 8626 6510 8640
rect 6578 8636 6731 8682
rect 6560 8624 6752 8636
rect 6831 8624 6844 8640
rect 6926 8624 6945 8640
rect 6960 8624 6966 8640
rect 6975 8624 6988 8640
rect 7043 8624 7058 8638
rect 7077 8626 7090 8640
rect 7158 8636 7311 8682
rect 7140 8624 7332 8636
rect 7411 8624 7424 8640
rect 7506 8624 7525 8640
rect 7540 8624 7546 8640
rect 7555 8624 7568 8640
rect 7623 8624 7638 8638
rect 7657 8626 7670 8640
rect 7738 8636 7891 8682
rect 7720 8624 7912 8636
rect 7991 8624 8004 8640
rect 8086 8624 8105 8640
rect 8120 8624 8126 8640
rect 8135 8624 8148 8640
rect 8203 8624 8218 8638
rect 8237 8626 8250 8640
rect 8318 8636 8471 8682
rect 8300 8624 8492 8636
rect 8571 8624 8584 8640
rect 8666 8624 8685 8640
rect 8700 8624 8706 8640
rect 8715 8624 8728 8640
rect 8783 8624 8798 8638
rect 8817 8626 8830 8640
rect 8898 8636 9051 8682
rect 8880 8624 9072 8636
rect 9151 8624 9164 8640
rect 9246 8624 9265 8640
rect 9280 8624 9286 8640
rect 9295 8624 9308 8640
rect 9363 8624 9378 8638
rect 9397 8626 9410 8640
rect 9478 8636 9631 8682
rect 9460 8624 9652 8636
rect 9731 8624 9744 8640
rect 9826 8624 9845 8640
rect 9860 8624 9866 8640
rect 9875 8624 9888 8640
rect 9943 8624 9958 8638
rect 9977 8626 9990 8640
rect 10058 8636 10211 8682
rect 10040 8624 10232 8636
rect 10311 8624 10324 8640
rect 10406 8624 10425 8640
rect 10440 8624 10446 8640
rect 10455 8624 10468 8640
rect 10523 8624 10538 8638
rect 10557 8626 10570 8640
rect 10638 8636 10791 8682
rect 10620 8624 10812 8636
rect 10891 8624 10904 8640
rect 10986 8624 11005 8640
rect 11020 8624 11026 8640
rect 11035 8624 11048 8640
rect 11103 8624 11118 8638
rect 11137 8626 11150 8640
rect 11218 8636 11371 8682
rect 11200 8624 11392 8636
rect 11471 8624 11484 8640
rect 11566 8624 11585 8640
rect 11600 8624 11606 8640
rect 11615 8624 11628 8640
rect 11683 8624 11698 8638
rect 11717 8626 11730 8640
rect 11798 8636 11951 8682
rect 11780 8624 11972 8636
rect 12051 8624 12064 8640
rect 12146 8624 12165 8640
rect 12180 8624 12186 8640
rect 12195 8624 12208 8640
rect 12263 8624 12278 8638
rect 12297 8626 12310 8640
rect 12378 8636 12531 8682
rect 12360 8624 12552 8636
rect 12631 8624 12644 8640
rect 12726 8624 12745 8640
rect 12760 8624 12766 8640
rect 12775 8624 12788 8640
rect 12843 8624 12858 8638
rect 12877 8626 12890 8640
rect 12958 8636 13111 8682
rect 12940 8624 13132 8636
rect 13211 8624 13224 8640
rect 13306 8624 13325 8640
rect 13340 8624 13346 8640
rect 13355 8624 13368 8640
rect 13423 8624 13438 8638
rect 13457 8626 13470 8640
rect 13538 8636 13691 8682
rect 13520 8624 13712 8636
rect 13791 8624 13804 8640
rect 13886 8624 13905 8640
rect 13920 8624 13926 8640
rect 13935 8624 13948 8640
rect 14003 8624 14018 8638
rect 14037 8626 14050 8640
rect 14118 8636 14271 8682
rect 14100 8624 14292 8636
rect 14371 8624 14384 8640
rect 14466 8624 14485 8640
rect 14500 8624 14506 8640
rect 14515 8624 14528 8640
rect 14583 8624 14598 8638
rect 14617 8626 14630 8640
rect 14698 8636 14851 8682
rect 14680 8624 14872 8636
rect 14951 8624 14964 8640
rect 15046 8624 15065 8640
rect 15080 8624 15086 8640
rect 15095 8624 15108 8640
rect 15163 8624 15178 8638
rect 15197 8626 15210 8640
rect 15278 8636 15431 8682
rect 15260 8624 15452 8636
rect 15531 8624 15544 8640
rect 15626 8624 15645 8640
rect 15660 8624 15666 8640
rect 15675 8624 15688 8640
rect 15743 8624 15758 8638
rect 15777 8626 15790 8640
rect 15858 8636 16011 8682
rect 15840 8624 16032 8636
rect 16111 8624 16124 8640
rect 16206 8624 16225 8640
rect 16240 8624 16246 8640
rect 16255 8624 16268 8640
rect 16323 8624 16338 8638
rect 16357 8626 16370 8640
rect 16438 8636 16591 8682
rect 16420 8624 16612 8636
rect 16691 8624 16704 8640
rect 16786 8624 16805 8640
rect 16820 8624 16826 8640
rect 16835 8624 16848 8640
rect 16903 8624 16918 8638
rect 16937 8626 16950 8640
rect 17018 8636 17171 8682
rect 17000 8624 17192 8636
rect 17271 8624 17284 8640
rect 17366 8624 17385 8640
rect 17400 8624 17406 8640
rect 17415 8624 17428 8640
rect 17483 8624 17498 8638
rect 17517 8626 17530 8640
rect 17598 8636 17751 8682
rect 17580 8624 17772 8636
rect 17851 8624 17864 8640
rect 17946 8624 17965 8640
rect 17980 8624 17986 8640
rect 17995 8624 18008 8640
rect 18063 8624 18078 8638
rect 18097 8626 18110 8640
rect 18178 8636 18331 8682
rect 18160 8624 18352 8636
rect 18431 8624 18444 8640
rect 18532 8624 18545 8640
rect 0 8610 18545 8624
rect 15 8540 28 8610
rect 73 8584 102 8598
rect 155 8584 171 8598
rect 209 8594 215 8596
rect 222 8594 330 8610
rect 337 8594 343 8596
rect 351 8594 366 8610
rect 432 8604 451 8607
rect 73 8582 171 8584
rect 198 8582 366 8594
rect 381 8584 397 8598
rect 432 8585 454 8604
rect 464 8598 480 8599
rect 463 8596 480 8598
rect 464 8591 480 8596
rect 454 8584 460 8585
rect 463 8584 492 8591
rect 381 8583 492 8584
rect 381 8582 498 8583
rect 57 8574 108 8582
rect 155 8574 189 8582
rect 57 8562 82 8574
rect 89 8562 108 8574
rect 162 8572 189 8574
rect 198 8572 419 8582
rect 454 8579 460 8582
rect 162 8568 419 8572
rect 57 8554 108 8562
rect 155 8554 419 8568
rect 463 8574 498 8582
rect 9 8506 28 8540
rect 73 8546 102 8554
rect 73 8540 90 8546
rect 73 8538 107 8540
rect 155 8538 171 8554
rect 172 8544 380 8554
rect 381 8544 397 8554
rect 445 8550 460 8565
rect 463 8562 464 8574
rect 471 8562 498 8574
rect 463 8554 498 8562
rect 463 8553 492 8554
rect 183 8540 397 8544
rect 198 8538 397 8540
rect 432 8540 445 8550
rect 463 8540 480 8553
rect 432 8538 480 8540
rect 74 8534 107 8538
rect 70 8532 107 8534
rect 70 8531 137 8532
rect 70 8526 101 8531
rect 107 8526 137 8531
rect 70 8522 137 8526
rect 43 8519 137 8522
rect 43 8512 92 8519
rect 43 8506 73 8512
rect 92 8507 97 8512
rect 9 8490 89 8506
rect 101 8498 137 8519
rect 198 8514 387 8538
rect 432 8537 479 8538
rect 445 8532 479 8537
rect 213 8511 387 8514
rect 206 8508 387 8511
rect 415 8531 479 8532
rect 9 8488 28 8490
rect 43 8488 77 8490
rect 9 8472 89 8488
rect 9 8466 28 8472
rect -1 8450 28 8466
rect 43 8456 73 8472
rect 101 8450 107 8498
rect 110 8492 129 8498
rect 144 8492 174 8500
rect 110 8484 174 8492
rect 110 8468 190 8484
rect 206 8477 268 8508
rect 284 8477 346 8508
rect 415 8506 464 8531
rect 479 8506 509 8522
rect 378 8492 408 8500
rect 415 8498 525 8506
rect 378 8484 423 8492
rect 110 8466 129 8468
rect 144 8466 190 8468
rect 110 8450 190 8466
rect 217 8464 252 8477
rect 293 8474 330 8477
rect 293 8472 335 8474
rect 222 8461 252 8464
rect 231 8457 238 8461
rect 238 8456 239 8457
rect 197 8450 207 8456
rect -7 8442 34 8450
rect -7 8416 8 8442
rect 15 8416 34 8442
rect 98 8438 129 8450
rect 144 8438 247 8450
rect 259 8440 285 8466
rect 300 8461 330 8472
rect 362 8468 424 8484
rect 362 8466 408 8468
rect 362 8450 424 8466
rect 436 8450 442 8498
rect 445 8490 525 8498
rect 445 8488 464 8490
rect 479 8488 513 8490
rect 445 8472 525 8488
rect 445 8450 464 8472
rect 479 8456 509 8472
rect 537 8466 543 8540
rect 546 8466 565 8610
rect 580 8466 586 8610
rect 595 8540 608 8610
rect 653 8584 682 8598
rect 735 8584 751 8598
rect 789 8594 795 8596
rect 802 8594 910 8610
rect 917 8594 923 8596
rect 931 8594 946 8610
rect 1012 8604 1031 8607
rect 653 8582 751 8584
rect 778 8582 946 8594
rect 961 8584 977 8598
rect 1012 8585 1034 8604
rect 1044 8598 1060 8599
rect 1043 8596 1060 8598
rect 1044 8591 1060 8596
rect 1034 8584 1040 8585
rect 1043 8584 1072 8591
rect 961 8583 1072 8584
rect 961 8582 1078 8583
rect 637 8574 688 8582
rect 735 8574 769 8582
rect 637 8562 662 8574
rect 669 8562 688 8574
rect 742 8572 769 8574
rect 778 8572 999 8582
rect 1034 8579 1040 8582
rect 742 8568 999 8572
rect 637 8554 688 8562
rect 735 8554 999 8568
rect 1043 8574 1078 8582
rect 589 8506 608 8540
rect 653 8546 682 8554
rect 653 8540 670 8546
rect 653 8538 687 8540
rect 735 8538 751 8554
rect 752 8544 960 8554
rect 961 8544 977 8554
rect 1025 8550 1040 8565
rect 1043 8562 1044 8574
rect 1051 8562 1078 8574
rect 1043 8554 1078 8562
rect 1043 8553 1072 8554
rect 763 8540 977 8544
rect 778 8538 977 8540
rect 1012 8540 1025 8550
rect 1043 8540 1060 8553
rect 1012 8538 1060 8540
rect 654 8534 687 8538
rect 650 8532 687 8534
rect 650 8531 717 8532
rect 650 8526 681 8531
rect 687 8526 717 8531
rect 650 8522 717 8526
rect 623 8519 717 8522
rect 623 8512 672 8519
rect 623 8506 653 8512
rect 672 8507 677 8512
rect 589 8490 669 8506
rect 681 8498 717 8519
rect 778 8514 967 8538
rect 1012 8537 1059 8538
rect 1025 8532 1059 8537
rect 793 8511 967 8514
rect 786 8508 967 8511
rect 995 8531 1059 8532
rect 589 8488 608 8490
rect 623 8488 657 8490
rect 589 8472 669 8488
rect 589 8466 608 8472
rect 305 8440 408 8450
rect 259 8438 408 8440
rect 429 8438 464 8450
rect 98 8436 260 8438
rect 110 8416 129 8436
rect 144 8434 174 8436
rect -7 8408 34 8416
rect 116 8412 129 8416
rect 181 8420 260 8436
rect 292 8436 464 8438
rect 292 8420 371 8436
rect 378 8434 408 8436
rect -1 8398 28 8408
rect 43 8398 73 8412
rect 116 8398 159 8412
rect 181 8408 371 8420
rect 436 8416 442 8436
rect 166 8398 196 8408
rect 197 8398 355 8408
rect 359 8398 389 8408
rect 393 8398 423 8412
rect 451 8398 464 8436
rect 536 8450 565 8466
rect 579 8450 608 8466
rect 623 8456 653 8472
rect 681 8450 687 8498
rect 690 8492 709 8498
rect 724 8492 754 8500
rect 690 8484 754 8492
rect 690 8468 770 8484
rect 786 8477 848 8508
rect 864 8477 926 8508
rect 995 8506 1044 8531
rect 1059 8506 1089 8522
rect 958 8492 988 8500
rect 995 8498 1105 8506
rect 958 8484 1003 8492
rect 690 8466 709 8468
rect 724 8466 770 8468
rect 690 8450 770 8466
rect 797 8464 832 8477
rect 873 8474 910 8477
rect 873 8472 915 8474
rect 802 8461 832 8464
rect 811 8457 818 8461
rect 818 8456 819 8457
rect 777 8450 787 8456
rect 536 8442 571 8450
rect 536 8416 537 8442
rect 544 8416 571 8442
rect 479 8398 509 8412
rect 536 8408 571 8416
rect 573 8442 614 8450
rect 573 8416 588 8442
rect 595 8416 614 8442
rect 678 8438 709 8450
rect 724 8438 827 8450
rect 839 8440 865 8466
rect 880 8461 910 8472
rect 942 8468 1004 8484
rect 942 8466 988 8468
rect 942 8450 1004 8466
rect 1016 8450 1022 8498
rect 1025 8490 1105 8498
rect 1025 8488 1044 8490
rect 1059 8488 1093 8490
rect 1025 8472 1105 8488
rect 1025 8450 1044 8472
rect 1059 8456 1089 8472
rect 1117 8466 1123 8540
rect 1126 8466 1145 8610
rect 1160 8466 1166 8610
rect 1175 8540 1188 8610
rect 1233 8584 1262 8598
rect 1315 8584 1331 8598
rect 1369 8594 1375 8596
rect 1382 8594 1490 8610
rect 1497 8594 1503 8596
rect 1511 8594 1526 8610
rect 1592 8604 1611 8607
rect 1233 8582 1331 8584
rect 1358 8582 1526 8594
rect 1541 8584 1557 8598
rect 1592 8585 1614 8604
rect 1624 8598 1640 8599
rect 1623 8596 1640 8598
rect 1624 8591 1640 8596
rect 1614 8584 1620 8585
rect 1623 8584 1652 8591
rect 1541 8583 1652 8584
rect 1541 8582 1658 8583
rect 1217 8574 1268 8582
rect 1315 8574 1349 8582
rect 1217 8562 1242 8574
rect 1249 8562 1268 8574
rect 1322 8572 1349 8574
rect 1358 8572 1579 8582
rect 1614 8579 1620 8582
rect 1322 8568 1579 8572
rect 1217 8554 1268 8562
rect 1315 8554 1579 8568
rect 1623 8574 1658 8582
rect 1169 8506 1188 8540
rect 1233 8546 1262 8554
rect 1233 8540 1250 8546
rect 1233 8538 1267 8540
rect 1315 8538 1331 8554
rect 1332 8544 1540 8554
rect 1541 8544 1557 8554
rect 1605 8550 1620 8565
rect 1623 8562 1624 8574
rect 1631 8562 1658 8574
rect 1623 8554 1658 8562
rect 1623 8553 1652 8554
rect 1343 8540 1557 8544
rect 1358 8538 1557 8540
rect 1592 8540 1605 8550
rect 1623 8540 1640 8553
rect 1592 8538 1640 8540
rect 1234 8534 1267 8538
rect 1230 8532 1267 8534
rect 1230 8531 1297 8532
rect 1230 8526 1261 8531
rect 1267 8526 1297 8531
rect 1230 8522 1297 8526
rect 1203 8519 1297 8522
rect 1203 8512 1252 8519
rect 1203 8506 1233 8512
rect 1252 8507 1257 8512
rect 1169 8490 1249 8506
rect 1261 8498 1297 8519
rect 1358 8514 1547 8538
rect 1592 8537 1639 8538
rect 1605 8532 1639 8537
rect 1373 8511 1547 8514
rect 1366 8508 1547 8511
rect 1575 8531 1639 8532
rect 1169 8488 1188 8490
rect 1203 8488 1237 8490
rect 1169 8472 1249 8488
rect 1169 8466 1188 8472
rect 885 8440 988 8450
rect 839 8438 988 8440
rect 1009 8438 1044 8450
rect 678 8436 840 8438
rect 690 8416 709 8436
rect 724 8434 754 8436
rect 573 8408 614 8416
rect 696 8412 709 8416
rect 761 8420 840 8436
rect 872 8436 1044 8438
rect 872 8420 951 8436
rect 958 8434 988 8436
rect 536 8398 565 8408
rect 579 8398 608 8408
rect 623 8398 653 8412
rect 696 8398 739 8412
rect 761 8408 951 8420
rect 1016 8416 1022 8436
rect 746 8398 776 8408
rect 777 8398 935 8408
rect 939 8398 969 8408
rect 973 8398 1003 8412
rect 1031 8398 1044 8436
rect 1116 8450 1145 8466
rect 1159 8450 1188 8466
rect 1203 8456 1233 8472
rect 1261 8450 1267 8498
rect 1270 8492 1289 8498
rect 1304 8492 1334 8500
rect 1270 8484 1334 8492
rect 1270 8468 1350 8484
rect 1366 8477 1428 8508
rect 1444 8477 1506 8508
rect 1575 8506 1624 8531
rect 1639 8506 1669 8522
rect 1538 8492 1568 8500
rect 1575 8498 1685 8506
rect 1538 8484 1583 8492
rect 1270 8466 1289 8468
rect 1304 8466 1350 8468
rect 1270 8450 1350 8466
rect 1377 8464 1412 8477
rect 1453 8474 1490 8477
rect 1453 8472 1495 8474
rect 1382 8461 1412 8464
rect 1391 8457 1398 8461
rect 1398 8456 1399 8457
rect 1357 8450 1367 8456
rect 1116 8442 1151 8450
rect 1116 8416 1117 8442
rect 1124 8416 1151 8442
rect 1059 8398 1089 8412
rect 1116 8408 1151 8416
rect 1153 8442 1194 8450
rect 1153 8416 1168 8442
rect 1175 8416 1194 8442
rect 1258 8438 1289 8450
rect 1304 8438 1407 8450
rect 1419 8440 1445 8466
rect 1460 8461 1490 8472
rect 1522 8468 1584 8484
rect 1522 8466 1568 8468
rect 1522 8450 1584 8466
rect 1596 8450 1602 8498
rect 1605 8490 1685 8498
rect 1605 8488 1624 8490
rect 1639 8488 1673 8490
rect 1605 8472 1685 8488
rect 1605 8450 1624 8472
rect 1639 8456 1669 8472
rect 1697 8466 1703 8540
rect 1706 8466 1725 8610
rect 1740 8466 1746 8610
rect 1755 8540 1768 8610
rect 1813 8584 1842 8598
rect 1895 8584 1911 8598
rect 1949 8594 1955 8596
rect 1962 8594 2070 8610
rect 2077 8594 2083 8596
rect 2091 8594 2106 8610
rect 2172 8604 2191 8607
rect 1813 8582 1911 8584
rect 1938 8582 2106 8594
rect 2121 8584 2137 8598
rect 2172 8585 2194 8604
rect 2204 8598 2220 8599
rect 2203 8596 2220 8598
rect 2204 8591 2220 8596
rect 2194 8584 2200 8585
rect 2203 8584 2232 8591
rect 2121 8583 2232 8584
rect 2121 8582 2238 8583
rect 1797 8574 1848 8582
rect 1895 8574 1929 8582
rect 1797 8562 1822 8574
rect 1829 8562 1848 8574
rect 1902 8572 1929 8574
rect 1938 8572 2159 8582
rect 2194 8579 2200 8582
rect 1902 8568 2159 8572
rect 1797 8554 1848 8562
rect 1895 8554 2159 8568
rect 2203 8574 2238 8582
rect 1749 8506 1768 8540
rect 1813 8546 1842 8554
rect 1813 8540 1830 8546
rect 1813 8538 1847 8540
rect 1895 8538 1911 8554
rect 1912 8544 2120 8554
rect 2121 8544 2137 8554
rect 2185 8550 2200 8565
rect 2203 8562 2204 8574
rect 2211 8562 2238 8574
rect 2203 8554 2238 8562
rect 2203 8553 2232 8554
rect 1923 8540 2137 8544
rect 1938 8538 2137 8540
rect 2172 8540 2185 8550
rect 2203 8540 2220 8553
rect 2172 8538 2220 8540
rect 1814 8534 1847 8538
rect 1810 8532 1847 8534
rect 1810 8531 1877 8532
rect 1810 8526 1841 8531
rect 1847 8526 1877 8531
rect 1810 8522 1877 8526
rect 1783 8519 1877 8522
rect 1783 8512 1832 8519
rect 1783 8506 1813 8512
rect 1832 8507 1837 8512
rect 1749 8490 1829 8506
rect 1841 8498 1877 8519
rect 1938 8514 2127 8538
rect 2172 8537 2219 8538
rect 2185 8532 2219 8537
rect 1953 8511 2127 8514
rect 1946 8508 2127 8511
rect 2155 8531 2219 8532
rect 1749 8488 1768 8490
rect 1783 8488 1817 8490
rect 1749 8472 1829 8488
rect 1749 8466 1768 8472
rect 1465 8440 1568 8450
rect 1419 8438 1568 8440
rect 1589 8438 1624 8450
rect 1258 8436 1420 8438
rect 1270 8416 1289 8436
rect 1304 8434 1334 8436
rect 1153 8408 1194 8416
rect 1276 8412 1289 8416
rect 1341 8420 1420 8436
rect 1452 8436 1624 8438
rect 1452 8420 1531 8436
rect 1538 8434 1568 8436
rect 1116 8398 1145 8408
rect 1159 8398 1188 8408
rect 1203 8398 1233 8412
rect 1276 8398 1319 8412
rect 1341 8408 1531 8420
rect 1596 8416 1602 8436
rect 1326 8398 1356 8408
rect 1357 8398 1515 8408
rect 1519 8398 1549 8408
rect 1553 8398 1583 8412
rect 1611 8398 1624 8436
rect 1696 8450 1725 8466
rect 1739 8450 1768 8466
rect 1783 8456 1813 8472
rect 1841 8450 1847 8498
rect 1850 8492 1869 8498
rect 1884 8492 1914 8500
rect 1850 8484 1914 8492
rect 1850 8468 1930 8484
rect 1946 8477 2008 8508
rect 2024 8477 2086 8508
rect 2155 8506 2204 8531
rect 2219 8506 2249 8522
rect 2118 8492 2148 8500
rect 2155 8498 2265 8506
rect 2118 8484 2163 8492
rect 1850 8466 1869 8468
rect 1884 8466 1930 8468
rect 1850 8450 1930 8466
rect 1957 8464 1992 8477
rect 2033 8474 2070 8477
rect 2033 8472 2075 8474
rect 1962 8461 1992 8464
rect 1971 8457 1978 8461
rect 1978 8456 1979 8457
rect 1937 8450 1947 8456
rect 1696 8442 1731 8450
rect 1696 8416 1697 8442
rect 1704 8416 1731 8442
rect 1639 8398 1669 8412
rect 1696 8408 1731 8416
rect 1733 8442 1774 8450
rect 1733 8416 1748 8442
rect 1755 8416 1774 8442
rect 1838 8438 1869 8450
rect 1884 8438 1987 8450
rect 1999 8440 2025 8466
rect 2040 8461 2070 8472
rect 2102 8468 2164 8484
rect 2102 8466 2148 8468
rect 2102 8450 2164 8466
rect 2176 8450 2182 8498
rect 2185 8490 2265 8498
rect 2185 8488 2204 8490
rect 2219 8488 2253 8490
rect 2185 8472 2265 8488
rect 2185 8450 2204 8472
rect 2219 8456 2249 8472
rect 2277 8466 2283 8540
rect 2286 8466 2305 8610
rect 2320 8466 2326 8610
rect 2335 8540 2348 8610
rect 2393 8584 2422 8598
rect 2475 8584 2491 8598
rect 2529 8594 2535 8596
rect 2542 8594 2650 8610
rect 2657 8594 2663 8596
rect 2671 8594 2686 8610
rect 2752 8604 2771 8607
rect 2393 8582 2491 8584
rect 2518 8582 2686 8594
rect 2701 8584 2717 8598
rect 2752 8585 2774 8604
rect 2784 8598 2800 8599
rect 2783 8596 2800 8598
rect 2784 8591 2800 8596
rect 2774 8584 2780 8585
rect 2783 8584 2812 8591
rect 2701 8583 2812 8584
rect 2701 8582 2818 8583
rect 2377 8574 2428 8582
rect 2475 8574 2509 8582
rect 2377 8562 2402 8574
rect 2409 8562 2428 8574
rect 2482 8572 2509 8574
rect 2518 8572 2739 8582
rect 2774 8579 2780 8582
rect 2482 8568 2739 8572
rect 2377 8554 2428 8562
rect 2475 8554 2739 8568
rect 2783 8574 2818 8582
rect 2329 8506 2348 8540
rect 2393 8546 2422 8554
rect 2393 8540 2410 8546
rect 2393 8538 2427 8540
rect 2475 8538 2491 8554
rect 2492 8544 2700 8554
rect 2701 8544 2717 8554
rect 2765 8550 2780 8565
rect 2783 8562 2784 8574
rect 2791 8562 2818 8574
rect 2783 8554 2818 8562
rect 2783 8553 2812 8554
rect 2503 8540 2717 8544
rect 2518 8538 2717 8540
rect 2752 8540 2765 8550
rect 2783 8540 2800 8553
rect 2752 8538 2800 8540
rect 2394 8534 2427 8538
rect 2390 8532 2427 8534
rect 2390 8531 2457 8532
rect 2390 8526 2421 8531
rect 2427 8526 2457 8531
rect 2390 8522 2457 8526
rect 2363 8519 2457 8522
rect 2363 8512 2412 8519
rect 2363 8506 2393 8512
rect 2412 8507 2417 8512
rect 2329 8490 2409 8506
rect 2421 8498 2457 8519
rect 2518 8514 2707 8538
rect 2752 8537 2799 8538
rect 2765 8532 2799 8537
rect 2533 8511 2707 8514
rect 2526 8508 2707 8511
rect 2735 8531 2799 8532
rect 2329 8488 2348 8490
rect 2363 8488 2397 8490
rect 2329 8472 2409 8488
rect 2329 8466 2348 8472
rect 2045 8440 2148 8450
rect 1999 8438 2148 8440
rect 2169 8438 2204 8450
rect 1838 8436 2000 8438
rect 1850 8416 1869 8436
rect 1884 8434 1914 8436
rect 1733 8408 1774 8416
rect 1856 8412 1869 8416
rect 1921 8420 2000 8436
rect 2032 8436 2204 8438
rect 2032 8420 2111 8436
rect 2118 8434 2148 8436
rect 1696 8398 1725 8408
rect 1739 8398 1768 8408
rect 1783 8398 1813 8412
rect 1856 8398 1899 8412
rect 1921 8408 2111 8420
rect 2176 8416 2182 8436
rect 1906 8398 1936 8408
rect 1937 8398 2095 8408
rect 2099 8398 2129 8408
rect 2133 8398 2163 8412
rect 2191 8398 2204 8436
rect 2276 8450 2305 8466
rect 2319 8450 2348 8466
rect 2363 8456 2393 8472
rect 2421 8450 2427 8498
rect 2430 8492 2449 8498
rect 2464 8492 2494 8500
rect 2430 8484 2494 8492
rect 2430 8468 2510 8484
rect 2526 8477 2588 8508
rect 2604 8477 2666 8508
rect 2735 8506 2784 8531
rect 2799 8506 2829 8522
rect 2698 8492 2728 8500
rect 2735 8498 2845 8506
rect 2698 8484 2743 8492
rect 2430 8466 2449 8468
rect 2464 8466 2510 8468
rect 2430 8450 2510 8466
rect 2537 8464 2572 8477
rect 2613 8474 2650 8477
rect 2613 8472 2655 8474
rect 2542 8461 2572 8464
rect 2551 8457 2558 8461
rect 2558 8456 2559 8457
rect 2517 8450 2527 8456
rect 2276 8442 2311 8450
rect 2276 8416 2277 8442
rect 2284 8416 2311 8442
rect 2219 8398 2249 8412
rect 2276 8408 2311 8416
rect 2313 8442 2354 8450
rect 2313 8416 2328 8442
rect 2335 8416 2354 8442
rect 2418 8438 2449 8450
rect 2464 8438 2567 8450
rect 2579 8440 2605 8466
rect 2620 8461 2650 8472
rect 2682 8468 2744 8484
rect 2682 8466 2728 8468
rect 2682 8450 2744 8466
rect 2756 8450 2762 8498
rect 2765 8490 2845 8498
rect 2765 8488 2784 8490
rect 2799 8488 2833 8490
rect 2765 8472 2845 8488
rect 2765 8450 2784 8472
rect 2799 8456 2829 8472
rect 2857 8466 2863 8540
rect 2866 8466 2885 8610
rect 2900 8466 2906 8610
rect 2915 8540 2928 8610
rect 2973 8584 3002 8598
rect 3055 8584 3071 8598
rect 3109 8594 3115 8596
rect 3122 8594 3230 8610
rect 3237 8594 3243 8596
rect 3251 8594 3266 8610
rect 3332 8604 3351 8607
rect 2973 8582 3071 8584
rect 3098 8582 3266 8594
rect 3281 8584 3297 8598
rect 3332 8585 3354 8604
rect 3364 8598 3380 8599
rect 3363 8596 3380 8598
rect 3364 8591 3380 8596
rect 3354 8584 3360 8585
rect 3363 8584 3392 8591
rect 3281 8583 3392 8584
rect 3281 8582 3398 8583
rect 2957 8574 3008 8582
rect 3055 8574 3089 8582
rect 2957 8562 2982 8574
rect 2989 8562 3008 8574
rect 3062 8572 3089 8574
rect 3098 8572 3319 8582
rect 3354 8579 3360 8582
rect 3062 8568 3319 8572
rect 2957 8554 3008 8562
rect 3055 8554 3319 8568
rect 3363 8574 3398 8582
rect 2909 8506 2928 8540
rect 2973 8546 3002 8554
rect 2973 8540 2990 8546
rect 2973 8538 3007 8540
rect 3055 8538 3071 8554
rect 3072 8544 3280 8554
rect 3281 8544 3297 8554
rect 3345 8550 3360 8565
rect 3363 8562 3364 8574
rect 3371 8562 3398 8574
rect 3363 8554 3398 8562
rect 3363 8553 3392 8554
rect 3083 8540 3297 8544
rect 3098 8538 3297 8540
rect 3332 8540 3345 8550
rect 3363 8540 3380 8553
rect 3332 8538 3380 8540
rect 2974 8534 3007 8538
rect 2970 8532 3007 8534
rect 2970 8531 3037 8532
rect 2970 8526 3001 8531
rect 3007 8526 3037 8531
rect 2970 8522 3037 8526
rect 2943 8519 3037 8522
rect 2943 8512 2992 8519
rect 2943 8506 2973 8512
rect 2992 8507 2997 8512
rect 2909 8490 2989 8506
rect 3001 8498 3037 8519
rect 3098 8514 3287 8538
rect 3332 8537 3379 8538
rect 3345 8532 3379 8537
rect 3113 8511 3287 8514
rect 3106 8508 3287 8511
rect 3315 8531 3379 8532
rect 2909 8488 2928 8490
rect 2943 8488 2977 8490
rect 2909 8472 2989 8488
rect 2909 8466 2928 8472
rect 2625 8440 2728 8450
rect 2579 8438 2728 8440
rect 2749 8438 2784 8450
rect 2418 8436 2580 8438
rect 2430 8416 2449 8436
rect 2464 8434 2494 8436
rect 2313 8408 2354 8416
rect 2436 8412 2449 8416
rect 2501 8420 2580 8436
rect 2612 8436 2784 8438
rect 2612 8420 2691 8436
rect 2698 8434 2728 8436
rect 2276 8398 2305 8408
rect 2319 8398 2348 8408
rect 2363 8398 2393 8412
rect 2436 8398 2479 8412
rect 2501 8408 2691 8420
rect 2756 8416 2762 8436
rect 2486 8398 2516 8408
rect 2517 8398 2675 8408
rect 2679 8398 2709 8408
rect 2713 8398 2743 8412
rect 2771 8398 2784 8436
rect 2856 8450 2885 8466
rect 2899 8450 2928 8466
rect 2943 8456 2973 8472
rect 3001 8450 3007 8498
rect 3010 8492 3029 8498
rect 3044 8492 3074 8500
rect 3010 8484 3074 8492
rect 3010 8468 3090 8484
rect 3106 8477 3168 8508
rect 3184 8477 3246 8508
rect 3315 8506 3364 8531
rect 3379 8506 3409 8522
rect 3278 8492 3308 8500
rect 3315 8498 3425 8506
rect 3278 8484 3323 8492
rect 3010 8466 3029 8468
rect 3044 8466 3090 8468
rect 3010 8450 3090 8466
rect 3117 8464 3152 8477
rect 3193 8474 3230 8477
rect 3193 8472 3235 8474
rect 3122 8461 3152 8464
rect 3131 8457 3138 8461
rect 3138 8456 3139 8457
rect 3097 8450 3107 8456
rect 2856 8442 2891 8450
rect 2856 8416 2857 8442
rect 2864 8416 2891 8442
rect 2799 8398 2829 8412
rect 2856 8408 2891 8416
rect 2893 8442 2934 8450
rect 2893 8416 2908 8442
rect 2915 8416 2934 8442
rect 2998 8438 3029 8450
rect 3044 8438 3147 8450
rect 3159 8440 3185 8466
rect 3200 8461 3230 8472
rect 3262 8468 3324 8484
rect 3262 8466 3308 8468
rect 3262 8450 3324 8466
rect 3336 8450 3342 8498
rect 3345 8490 3425 8498
rect 3345 8488 3364 8490
rect 3379 8488 3413 8490
rect 3345 8472 3425 8488
rect 3345 8450 3364 8472
rect 3379 8456 3409 8472
rect 3437 8466 3443 8540
rect 3446 8466 3465 8610
rect 3480 8466 3486 8610
rect 3495 8540 3508 8610
rect 3553 8584 3582 8598
rect 3635 8584 3651 8598
rect 3689 8594 3695 8596
rect 3702 8594 3810 8610
rect 3817 8594 3823 8596
rect 3831 8594 3846 8610
rect 3912 8604 3931 8607
rect 3553 8582 3651 8584
rect 3678 8582 3846 8594
rect 3861 8584 3877 8598
rect 3912 8585 3934 8604
rect 3944 8598 3960 8599
rect 3943 8596 3960 8598
rect 3944 8591 3960 8596
rect 3934 8584 3940 8585
rect 3943 8584 3972 8591
rect 3861 8583 3972 8584
rect 3861 8582 3978 8583
rect 3537 8574 3588 8582
rect 3635 8574 3669 8582
rect 3537 8562 3562 8574
rect 3569 8562 3588 8574
rect 3642 8572 3669 8574
rect 3678 8572 3899 8582
rect 3934 8579 3940 8582
rect 3642 8568 3899 8572
rect 3537 8554 3588 8562
rect 3635 8554 3899 8568
rect 3943 8574 3978 8582
rect 3489 8506 3508 8540
rect 3553 8546 3582 8554
rect 3553 8540 3570 8546
rect 3553 8538 3587 8540
rect 3635 8538 3651 8554
rect 3652 8544 3860 8554
rect 3861 8544 3877 8554
rect 3925 8550 3940 8565
rect 3943 8562 3944 8574
rect 3951 8562 3978 8574
rect 3943 8554 3978 8562
rect 3943 8553 3972 8554
rect 3663 8540 3877 8544
rect 3678 8538 3877 8540
rect 3912 8540 3925 8550
rect 3943 8540 3960 8553
rect 3912 8538 3960 8540
rect 3554 8534 3587 8538
rect 3550 8532 3587 8534
rect 3550 8531 3617 8532
rect 3550 8526 3581 8531
rect 3587 8526 3617 8531
rect 3550 8522 3617 8526
rect 3523 8519 3617 8522
rect 3523 8512 3572 8519
rect 3523 8506 3553 8512
rect 3572 8507 3577 8512
rect 3489 8490 3569 8506
rect 3581 8498 3617 8519
rect 3678 8514 3867 8538
rect 3912 8537 3959 8538
rect 3925 8532 3959 8537
rect 3693 8511 3867 8514
rect 3686 8508 3867 8511
rect 3895 8531 3959 8532
rect 3489 8488 3508 8490
rect 3523 8488 3557 8490
rect 3489 8472 3569 8488
rect 3489 8466 3508 8472
rect 3205 8440 3308 8450
rect 3159 8438 3308 8440
rect 3329 8438 3364 8450
rect 2998 8436 3160 8438
rect 3010 8416 3029 8436
rect 3044 8434 3074 8436
rect 2893 8408 2934 8416
rect 3016 8412 3029 8416
rect 3081 8420 3160 8436
rect 3192 8436 3364 8438
rect 3192 8420 3271 8436
rect 3278 8434 3308 8436
rect 2856 8398 2885 8408
rect 2899 8398 2928 8408
rect 2943 8398 2973 8412
rect 3016 8398 3059 8412
rect 3081 8408 3271 8420
rect 3336 8416 3342 8436
rect 3066 8398 3096 8408
rect 3097 8398 3255 8408
rect 3259 8398 3289 8408
rect 3293 8398 3323 8412
rect 3351 8398 3364 8436
rect 3436 8450 3465 8466
rect 3479 8450 3508 8466
rect 3523 8456 3553 8472
rect 3581 8450 3587 8498
rect 3590 8492 3609 8498
rect 3624 8492 3654 8500
rect 3590 8484 3654 8492
rect 3590 8468 3670 8484
rect 3686 8477 3748 8508
rect 3764 8477 3826 8508
rect 3895 8506 3944 8531
rect 3959 8506 3989 8522
rect 3858 8492 3888 8500
rect 3895 8498 4005 8506
rect 3858 8484 3903 8492
rect 3590 8466 3609 8468
rect 3624 8466 3670 8468
rect 3590 8450 3670 8466
rect 3697 8464 3732 8477
rect 3773 8474 3810 8477
rect 3773 8472 3815 8474
rect 3702 8461 3732 8464
rect 3711 8457 3718 8461
rect 3718 8456 3719 8457
rect 3677 8450 3687 8456
rect 3436 8442 3471 8450
rect 3436 8416 3437 8442
rect 3444 8416 3471 8442
rect 3379 8398 3409 8412
rect 3436 8408 3471 8416
rect 3473 8442 3514 8450
rect 3473 8416 3488 8442
rect 3495 8416 3514 8442
rect 3578 8438 3609 8450
rect 3624 8438 3727 8450
rect 3739 8440 3765 8466
rect 3780 8461 3810 8472
rect 3842 8468 3904 8484
rect 3842 8466 3888 8468
rect 3842 8450 3904 8466
rect 3916 8450 3922 8498
rect 3925 8490 4005 8498
rect 3925 8488 3944 8490
rect 3959 8488 3993 8490
rect 3925 8472 4005 8488
rect 3925 8450 3944 8472
rect 3959 8456 3989 8472
rect 4017 8466 4023 8540
rect 4026 8466 4045 8610
rect 4060 8466 4066 8610
rect 4075 8540 4088 8610
rect 4133 8584 4162 8598
rect 4215 8584 4231 8598
rect 4269 8594 4275 8596
rect 4282 8594 4390 8610
rect 4397 8594 4403 8596
rect 4411 8594 4426 8610
rect 4492 8604 4511 8607
rect 4133 8582 4231 8584
rect 4258 8582 4426 8594
rect 4441 8584 4457 8598
rect 4492 8585 4514 8604
rect 4524 8598 4540 8599
rect 4523 8596 4540 8598
rect 4524 8591 4540 8596
rect 4514 8584 4520 8585
rect 4523 8584 4552 8591
rect 4441 8583 4552 8584
rect 4441 8582 4558 8583
rect 4117 8574 4168 8582
rect 4215 8574 4249 8582
rect 4117 8562 4142 8574
rect 4149 8562 4168 8574
rect 4222 8572 4249 8574
rect 4258 8572 4479 8582
rect 4514 8579 4520 8582
rect 4222 8568 4479 8572
rect 4117 8554 4168 8562
rect 4215 8554 4479 8568
rect 4523 8574 4558 8582
rect 4069 8506 4088 8540
rect 4133 8546 4162 8554
rect 4133 8540 4150 8546
rect 4133 8538 4167 8540
rect 4215 8538 4231 8554
rect 4232 8544 4440 8554
rect 4441 8544 4457 8554
rect 4505 8550 4520 8565
rect 4523 8562 4524 8574
rect 4531 8562 4558 8574
rect 4523 8554 4558 8562
rect 4523 8553 4552 8554
rect 4243 8540 4457 8544
rect 4258 8538 4457 8540
rect 4492 8540 4505 8550
rect 4523 8540 4540 8553
rect 4492 8538 4540 8540
rect 4134 8534 4167 8538
rect 4130 8532 4167 8534
rect 4130 8531 4197 8532
rect 4130 8526 4161 8531
rect 4167 8526 4197 8531
rect 4130 8522 4197 8526
rect 4103 8519 4197 8522
rect 4103 8512 4152 8519
rect 4103 8506 4133 8512
rect 4152 8507 4157 8512
rect 4069 8490 4149 8506
rect 4161 8498 4197 8519
rect 4258 8514 4447 8538
rect 4492 8537 4539 8538
rect 4505 8532 4539 8537
rect 4273 8511 4447 8514
rect 4266 8508 4447 8511
rect 4475 8531 4539 8532
rect 4069 8488 4088 8490
rect 4103 8488 4137 8490
rect 4069 8472 4149 8488
rect 4069 8466 4088 8472
rect 3785 8440 3888 8450
rect 3739 8438 3888 8440
rect 3909 8438 3944 8450
rect 3578 8436 3740 8438
rect 3590 8416 3609 8436
rect 3624 8434 3654 8436
rect 3473 8408 3514 8416
rect 3596 8412 3609 8416
rect 3661 8420 3740 8436
rect 3772 8436 3944 8438
rect 3772 8420 3851 8436
rect 3858 8434 3888 8436
rect 3436 8398 3465 8408
rect 3479 8398 3508 8408
rect 3523 8398 3553 8412
rect 3596 8398 3639 8412
rect 3661 8408 3851 8420
rect 3916 8416 3922 8436
rect 3646 8398 3676 8408
rect 3677 8398 3835 8408
rect 3839 8398 3869 8408
rect 3873 8398 3903 8412
rect 3931 8398 3944 8436
rect 4016 8450 4045 8466
rect 4059 8450 4088 8466
rect 4103 8456 4133 8472
rect 4161 8450 4167 8498
rect 4170 8492 4189 8498
rect 4204 8492 4234 8500
rect 4170 8484 4234 8492
rect 4170 8468 4250 8484
rect 4266 8477 4328 8508
rect 4344 8477 4406 8508
rect 4475 8506 4524 8531
rect 4539 8506 4569 8522
rect 4438 8492 4468 8500
rect 4475 8498 4585 8506
rect 4438 8484 4483 8492
rect 4170 8466 4189 8468
rect 4204 8466 4250 8468
rect 4170 8450 4250 8466
rect 4277 8464 4312 8477
rect 4353 8474 4390 8477
rect 4353 8472 4395 8474
rect 4282 8461 4312 8464
rect 4291 8457 4298 8461
rect 4298 8456 4299 8457
rect 4257 8450 4267 8456
rect 4016 8442 4051 8450
rect 4016 8416 4017 8442
rect 4024 8416 4051 8442
rect 3959 8398 3989 8412
rect 4016 8408 4051 8416
rect 4053 8442 4094 8450
rect 4053 8416 4068 8442
rect 4075 8416 4094 8442
rect 4158 8438 4189 8450
rect 4204 8438 4307 8450
rect 4319 8440 4345 8466
rect 4360 8461 4390 8472
rect 4422 8468 4484 8484
rect 4422 8466 4468 8468
rect 4422 8450 4484 8466
rect 4496 8450 4502 8498
rect 4505 8490 4585 8498
rect 4505 8488 4524 8490
rect 4539 8488 4573 8490
rect 4505 8472 4585 8488
rect 4505 8450 4524 8472
rect 4539 8456 4569 8472
rect 4597 8466 4603 8540
rect 4606 8466 4625 8610
rect 4640 8466 4646 8610
rect 4655 8540 4668 8610
rect 4713 8584 4742 8598
rect 4795 8584 4811 8598
rect 4849 8594 4855 8596
rect 4862 8594 4970 8610
rect 4977 8594 4983 8596
rect 4991 8594 5006 8610
rect 5072 8604 5091 8607
rect 4713 8582 4811 8584
rect 4838 8582 5006 8594
rect 5021 8584 5037 8598
rect 5072 8585 5094 8604
rect 5104 8598 5120 8599
rect 5103 8596 5120 8598
rect 5104 8591 5120 8596
rect 5094 8584 5100 8585
rect 5103 8584 5132 8591
rect 5021 8583 5132 8584
rect 5021 8582 5138 8583
rect 4697 8574 4748 8582
rect 4795 8574 4829 8582
rect 4697 8562 4722 8574
rect 4729 8562 4748 8574
rect 4802 8572 4829 8574
rect 4838 8572 5059 8582
rect 5094 8579 5100 8582
rect 4802 8568 5059 8572
rect 4697 8554 4748 8562
rect 4795 8554 5059 8568
rect 5103 8574 5138 8582
rect 4649 8506 4668 8540
rect 4713 8546 4742 8554
rect 4713 8540 4730 8546
rect 4713 8538 4747 8540
rect 4795 8538 4811 8554
rect 4812 8544 5020 8554
rect 5021 8544 5037 8554
rect 5085 8550 5100 8565
rect 5103 8562 5104 8574
rect 5111 8562 5138 8574
rect 5103 8554 5138 8562
rect 5103 8553 5132 8554
rect 4823 8540 5037 8544
rect 4838 8538 5037 8540
rect 5072 8540 5085 8550
rect 5103 8540 5120 8553
rect 5072 8538 5120 8540
rect 4714 8534 4747 8538
rect 4710 8532 4747 8534
rect 4710 8531 4777 8532
rect 4710 8526 4741 8531
rect 4747 8526 4777 8531
rect 4710 8522 4777 8526
rect 4683 8519 4777 8522
rect 4683 8512 4732 8519
rect 4683 8506 4713 8512
rect 4732 8507 4737 8512
rect 4649 8490 4729 8506
rect 4741 8498 4777 8519
rect 4838 8514 5027 8538
rect 5072 8537 5119 8538
rect 5085 8532 5119 8537
rect 4853 8511 5027 8514
rect 4846 8508 5027 8511
rect 5055 8531 5119 8532
rect 4649 8488 4668 8490
rect 4683 8488 4717 8490
rect 4649 8472 4729 8488
rect 4649 8466 4668 8472
rect 4365 8440 4468 8450
rect 4319 8438 4468 8440
rect 4489 8438 4524 8450
rect 4158 8436 4320 8438
rect 4170 8416 4189 8436
rect 4204 8434 4234 8436
rect 4053 8408 4094 8416
rect 4176 8412 4189 8416
rect 4241 8420 4320 8436
rect 4352 8436 4524 8438
rect 4352 8420 4431 8436
rect 4438 8434 4468 8436
rect 4016 8398 4045 8408
rect 4059 8398 4088 8408
rect 4103 8398 4133 8412
rect 4176 8398 4219 8412
rect 4241 8408 4431 8420
rect 4496 8416 4502 8436
rect 4226 8398 4256 8408
rect 4257 8398 4415 8408
rect 4419 8398 4449 8408
rect 4453 8398 4483 8412
rect 4511 8398 4524 8436
rect 4596 8450 4625 8466
rect 4639 8450 4668 8466
rect 4683 8456 4713 8472
rect 4741 8450 4747 8498
rect 4750 8492 4769 8498
rect 4784 8492 4814 8500
rect 4750 8484 4814 8492
rect 4750 8468 4830 8484
rect 4846 8477 4908 8508
rect 4924 8477 4986 8508
rect 5055 8506 5104 8531
rect 5119 8506 5149 8522
rect 5018 8492 5048 8500
rect 5055 8498 5165 8506
rect 5018 8484 5063 8492
rect 4750 8466 4769 8468
rect 4784 8466 4830 8468
rect 4750 8450 4830 8466
rect 4857 8464 4892 8477
rect 4933 8474 4970 8477
rect 4933 8472 4975 8474
rect 4862 8461 4892 8464
rect 4871 8457 4878 8461
rect 4878 8456 4879 8457
rect 4837 8450 4847 8456
rect 4596 8442 4631 8450
rect 4596 8416 4597 8442
rect 4604 8416 4631 8442
rect 4539 8398 4569 8412
rect 4596 8408 4631 8416
rect 4633 8442 4674 8450
rect 4633 8416 4648 8442
rect 4655 8416 4674 8442
rect 4738 8438 4769 8450
rect 4784 8438 4887 8450
rect 4899 8440 4925 8466
rect 4940 8461 4970 8472
rect 5002 8468 5064 8484
rect 5002 8466 5048 8468
rect 5002 8450 5064 8466
rect 5076 8450 5082 8498
rect 5085 8490 5165 8498
rect 5085 8488 5104 8490
rect 5119 8488 5153 8490
rect 5085 8472 5165 8488
rect 5085 8450 5104 8472
rect 5119 8456 5149 8472
rect 5177 8466 5183 8540
rect 5186 8466 5205 8610
rect 5220 8466 5226 8610
rect 5235 8540 5248 8610
rect 5293 8584 5322 8598
rect 5375 8584 5391 8598
rect 5429 8594 5435 8596
rect 5442 8594 5550 8610
rect 5557 8594 5563 8596
rect 5571 8594 5586 8610
rect 5652 8604 5671 8607
rect 5293 8582 5391 8584
rect 5418 8582 5586 8594
rect 5601 8584 5617 8598
rect 5652 8585 5674 8604
rect 5684 8598 5700 8599
rect 5683 8596 5700 8598
rect 5684 8591 5700 8596
rect 5674 8584 5680 8585
rect 5683 8584 5712 8591
rect 5601 8583 5712 8584
rect 5601 8582 5718 8583
rect 5277 8574 5328 8582
rect 5375 8574 5409 8582
rect 5277 8562 5302 8574
rect 5309 8562 5328 8574
rect 5382 8572 5409 8574
rect 5418 8572 5639 8582
rect 5674 8579 5680 8582
rect 5382 8568 5639 8572
rect 5277 8554 5328 8562
rect 5375 8554 5639 8568
rect 5683 8574 5718 8582
rect 5229 8506 5248 8540
rect 5293 8546 5322 8554
rect 5293 8540 5310 8546
rect 5293 8538 5327 8540
rect 5375 8538 5391 8554
rect 5392 8544 5600 8554
rect 5601 8544 5617 8554
rect 5665 8550 5680 8565
rect 5683 8562 5684 8574
rect 5691 8562 5718 8574
rect 5683 8554 5718 8562
rect 5683 8553 5712 8554
rect 5403 8540 5617 8544
rect 5418 8538 5617 8540
rect 5652 8540 5665 8550
rect 5683 8540 5700 8553
rect 5652 8538 5700 8540
rect 5294 8534 5327 8538
rect 5290 8532 5327 8534
rect 5290 8531 5357 8532
rect 5290 8526 5321 8531
rect 5327 8526 5357 8531
rect 5290 8522 5357 8526
rect 5263 8519 5357 8522
rect 5263 8512 5312 8519
rect 5263 8506 5293 8512
rect 5312 8507 5317 8512
rect 5229 8490 5309 8506
rect 5321 8498 5357 8519
rect 5418 8514 5607 8538
rect 5652 8537 5699 8538
rect 5665 8532 5699 8537
rect 5433 8511 5607 8514
rect 5426 8508 5607 8511
rect 5635 8531 5699 8532
rect 5229 8488 5248 8490
rect 5263 8488 5297 8490
rect 5229 8472 5309 8488
rect 5229 8466 5248 8472
rect 4945 8440 5048 8450
rect 4899 8438 5048 8440
rect 5069 8438 5104 8450
rect 4738 8436 4900 8438
rect 4750 8416 4769 8436
rect 4784 8434 4814 8436
rect 4633 8408 4674 8416
rect 4756 8412 4769 8416
rect 4821 8420 4900 8436
rect 4932 8436 5104 8438
rect 4932 8420 5011 8436
rect 5018 8434 5048 8436
rect 4596 8398 4625 8408
rect 4639 8398 4668 8408
rect 4683 8398 4713 8412
rect 4756 8398 4799 8412
rect 4821 8408 5011 8420
rect 5076 8416 5082 8436
rect 4806 8398 4836 8408
rect 4837 8398 4995 8408
rect 4999 8398 5029 8408
rect 5033 8398 5063 8412
rect 5091 8398 5104 8436
rect 5176 8450 5205 8466
rect 5219 8450 5248 8466
rect 5263 8456 5293 8472
rect 5321 8450 5327 8498
rect 5330 8492 5349 8498
rect 5364 8492 5394 8500
rect 5330 8484 5394 8492
rect 5330 8468 5410 8484
rect 5426 8477 5488 8508
rect 5504 8477 5566 8508
rect 5635 8506 5684 8531
rect 5699 8506 5729 8522
rect 5598 8492 5628 8500
rect 5635 8498 5745 8506
rect 5598 8484 5643 8492
rect 5330 8466 5349 8468
rect 5364 8466 5410 8468
rect 5330 8450 5410 8466
rect 5437 8464 5472 8477
rect 5513 8474 5550 8477
rect 5513 8472 5555 8474
rect 5442 8461 5472 8464
rect 5451 8457 5458 8461
rect 5458 8456 5459 8457
rect 5417 8450 5427 8456
rect 5176 8442 5211 8450
rect 5176 8416 5177 8442
rect 5184 8416 5211 8442
rect 5119 8398 5149 8412
rect 5176 8408 5211 8416
rect 5213 8442 5254 8450
rect 5213 8416 5228 8442
rect 5235 8416 5254 8442
rect 5318 8438 5349 8450
rect 5364 8438 5467 8450
rect 5479 8440 5505 8466
rect 5520 8461 5550 8472
rect 5582 8468 5644 8484
rect 5582 8466 5628 8468
rect 5582 8450 5644 8466
rect 5656 8450 5662 8498
rect 5665 8490 5745 8498
rect 5665 8488 5684 8490
rect 5699 8488 5733 8490
rect 5665 8472 5745 8488
rect 5665 8450 5684 8472
rect 5699 8456 5729 8472
rect 5757 8466 5763 8540
rect 5766 8466 5785 8610
rect 5800 8466 5806 8610
rect 5815 8540 5828 8610
rect 5873 8584 5902 8598
rect 5955 8584 5971 8598
rect 6009 8594 6015 8596
rect 6022 8594 6130 8610
rect 6137 8594 6143 8596
rect 6151 8594 6166 8610
rect 6232 8604 6251 8607
rect 5873 8582 5971 8584
rect 5998 8582 6166 8594
rect 6181 8584 6197 8598
rect 6232 8585 6254 8604
rect 6264 8598 6280 8599
rect 6263 8596 6280 8598
rect 6264 8591 6280 8596
rect 6254 8584 6260 8585
rect 6263 8584 6292 8591
rect 6181 8583 6292 8584
rect 6181 8582 6298 8583
rect 5857 8574 5908 8582
rect 5955 8574 5989 8582
rect 5857 8562 5882 8574
rect 5889 8562 5908 8574
rect 5962 8572 5989 8574
rect 5998 8572 6219 8582
rect 6254 8579 6260 8582
rect 5962 8568 6219 8572
rect 5857 8554 5908 8562
rect 5955 8554 6219 8568
rect 6263 8574 6298 8582
rect 5809 8506 5828 8540
rect 5873 8546 5902 8554
rect 5873 8540 5890 8546
rect 5873 8538 5907 8540
rect 5955 8538 5971 8554
rect 5972 8544 6180 8554
rect 6181 8544 6197 8554
rect 6245 8550 6260 8565
rect 6263 8562 6264 8574
rect 6271 8562 6298 8574
rect 6263 8554 6298 8562
rect 6263 8553 6292 8554
rect 5983 8540 6197 8544
rect 5998 8538 6197 8540
rect 6232 8540 6245 8550
rect 6263 8540 6280 8553
rect 6232 8538 6280 8540
rect 5874 8534 5907 8538
rect 5870 8532 5907 8534
rect 5870 8531 5937 8532
rect 5870 8526 5901 8531
rect 5907 8526 5937 8531
rect 5870 8522 5937 8526
rect 5843 8519 5937 8522
rect 5843 8512 5892 8519
rect 5843 8506 5873 8512
rect 5892 8507 5897 8512
rect 5809 8490 5889 8506
rect 5901 8498 5937 8519
rect 5998 8514 6187 8538
rect 6232 8537 6279 8538
rect 6245 8532 6279 8537
rect 6013 8511 6187 8514
rect 6006 8508 6187 8511
rect 6215 8531 6279 8532
rect 5809 8488 5828 8490
rect 5843 8488 5877 8490
rect 5809 8472 5889 8488
rect 5809 8466 5828 8472
rect 5525 8440 5628 8450
rect 5479 8438 5628 8440
rect 5649 8438 5684 8450
rect 5318 8436 5480 8438
rect 5330 8416 5349 8436
rect 5364 8434 5394 8436
rect 5213 8408 5254 8416
rect 5336 8412 5349 8416
rect 5401 8420 5480 8436
rect 5512 8436 5684 8438
rect 5512 8420 5591 8436
rect 5598 8434 5628 8436
rect 5176 8398 5205 8408
rect 5219 8398 5248 8408
rect 5263 8398 5293 8412
rect 5336 8398 5379 8412
rect 5401 8408 5591 8420
rect 5656 8416 5662 8436
rect 5386 8398 5416 8408
rect 5417 8398 5575 8408
rect 5579 8398 5609 8408
rect 5613 8398 5643 8412
rect 5671 8398 5684 8436
rect 5756 8450 5785 8466
rect 5799 8450 5828 8466
rect 5843 8456 5873 8472
rect 5901 8450 5907 8498
rect 5910 8492 5929 8498
rect 5944 8492 5974 8500
rect 5910 8484 5974 8492
rect 5910 8468 5990 8484
rect 6006 8477 6068 8508
rect 6084 8477 6146 8508
rect 6215 8506 6264 8531
rect 6279 8506 6309 8522
rect 6178 8492 6208 8500
rect 6215 8498 6325 8506
rect 6178 8484 6223 8492
rect 5910 8466 5929 8468
rect 5944 8466 5990 8468
rect 5910 8450 5990 8466
rect 6017 8464 6052 8477
rect 6093 8474 6130 8477
rect 6093 8472 6135 8474
rect 6022 8461 6052 8464
rect 6031 8457 6038 8461
rect 6038 8456 6039 8457
rect 5997 8450 6007 8456
rect 5756 8442 5791 8450
rect 5756 8416 5757 8442
rect 5764 8416 5791 8442
rect 5699 8398 5729 8412
rect 5756 8408 5791 8416
rect 5793 8442 5834 8450
rect 5793 8416 5808 8442
rect 5815 8416 5834 8442
rect 5898 8438 5929 8450
rect 5944 8438 6047 8450
rect 6059 8440 6085 8466
rect 6100 8461 6130 8472
rect 6162 8468 6224 8484
rect 6162 8466 6208 8468
rect 6162 8450 6224 8466
rect 6236 8450 6242 8498
rect 6245 8490 6325 8498
rect 6245 8488 6264 8490
rect 6279 8488 6313 8490
rect 6245 8472 6325 8488
rect 6245 8450 6264 8472
rect 6279 8456 6309 8472
rect 6337 8466 6343 8540
rect 6346 8466 6365 8610
rect 6380 8466 6386 8610
rect 6395 8540 6408 8610
rect 6453 8584 6482 8598
rect 6535 8584 6551 8598
rect 6589 8594 6595 8596
rect 6602 8594 6710 8610
rect 6717 8594 6723 8596
rect 6731 8594 6746 8610
rect 6812 8604 6831 8607
rect 6453 8582 6551 8584
rect 6578 8582 6746 8594
rect 6761 8584 6777 8598
rect 6812 8585 6834 8604
rect 6844 8598 6860 8599
rect 6843 8596 6860 8598
rect 6844 8591 6860 8596
rect 6834 8584 6840 8585
rect 6843 8584 6872 8591
rect 6761 8583 6872 8584
rect 6761 8582 6878 8583
rect 6437 8574 6488 8582
rect 6535 8574 6569 8582
rect 6437 8562 6462 8574
rect 6469 8562 6488 8574
rect 6542 8572 6569 8574
rect 6578 8572 6799 8582
rect 6834 8579 6840 8582
rect 6542 8568 6799 8572
rect 6437 8554 6488 8562
rect 6535 8554 6799 8568
rect 6843 8574 6878 8582
rect 6389 8506 6408 8540
rect 6453 8546 6482 8554
rect 6453 8540 6470 8546
rect 6453 8538 6487 8540
rect 6535 8538 6551 8554
rect 6552 8544 6760 8554
rect 6761 8544 6777 8554
rect 6825 8550 6840 8565
rect 6843 8562 6844 8574
rect 6851 8562 6878 8574
rect 6843 8554 6878 8562
rect 6843 8553 6872 8554
rect 6563 8540 6777 8544
rect 6578 8538 6777 8540
rect 6812 8540 6825 8550
rect 6843 8540 6860 8553
rect 6812 8538 6860 8540
rect 6454 8534 6487 8538
rect 6450 8532 6487 8534
rect 6450 8531 6517 8532
rect 6450 8526 6481 8531
rect 6487 8526 6517 8531
rect 6450 8522 6517 8526
rect 6423 8519 6517 8522
rect 6423 8512 6472 8519
rect 6423 8506 6453 8512
rect 6472 8507 6477 8512
rect 6389 8490 6469 8506
rect 6481 8498 6517 8519
rect 6578 8514 6767 8538
rect 6812 8537 6859 8538
rect 6825 8532 6859 8537
rect 6593 8511 6767 8514
rect 6586 8508 6767 8511
rect 6795 8531 6859 8532
rect 6389 8488 6408 8490
rect 6423 8488 6457 8490
rect 6389 8472 6469 8488
rect 6389 8466 6408 8472
rect 6105 8440 6208 8450
rect 6059 8438 6208 8440
rect 6229 8438 6264 8450
rect 5898 8436 6060 8438
rect 5910 8416 5929 8436
rect 5944 8434 5974 8436
rect 5793 8408 5834 8416
rect 5916 8412 5929 8416
rect 5981 8420 6060 8436
rect 6092 8436 6264 8438
rect 6092 8420 6171 8436
rect 6178 8434 6208 8436
rect 5756 8398 5785 8408
rect 5799 8398 5828 8408
rect 5843 8398 5873 8412
rect 5916 8398 5959 8412
rect 5981 8408 6171 8420
rect 6236 8416 6242 8436
rect 5966 8398 5996 8408
rect 5997 8398 6155 8408
rect 6159 8398 6189 8408
rect 6193 8398 6223 8412
rect 6251 8398 6264 8436
rect 6336 8450 6365 8466
rect 6379 8450 6408 8466
rect 6423 8456 6453 8472
rect 6481 8450 6487 8498
rect 6490 8492 6509 8498
rect 6524 8492 6554 8500
rect 6490 8484 6554 8492
rect 6490 8468 6570 8484
rect 6586 8477 6648 8508
rect 6664 8477 6726 8508
rect 6795 8506 6844 8531
rect 6859 8506 6889 8522
rect 6758 8492 6788 8500
rect 6795 8498 6905 8506
rect 6758 8484 6803 8492
rect 6490 8466 6509 8468
rect 6524 8466 6570 8468
rect 6490 8450 6570 8466
rect 6597 8464 6632 8477
rect 6673 8474 6710 8477
rect 6673 8472 6715 8474
rect 6602 8461 6632 8464
rect 6611 8457 6618 8461
rect 6618 8456 6619 8457
rect 6577 8450 6587 8456
rect 6336 8442 6371 8450
rect 6336 8416 6337 8442
rect 6344 8416 6371 8442
rect 6279 8398 6309 8412
rect 6336 8408 6371 8416
rect 6373 8442 6414 8450
rect 6373 8416 6388 8442
rect 6395 8416 6414 8442
rect 6478 8438 6509 8450
rect 6524 8438 6627 8450
rect 6639 8440 6665 8466
rect 6680 8461 6710 8472
rect 6742 8468 6804 8484
rect 6742 8466 6788 8468
rect 6742 8450 6804 8466
rect 6816 8450 6822 8498
rect 6825 8490 6905 8498
rect 6825 8488 6844 8490
rect 6859 8488 6893 8490
rect 6825 8472 6905 8488
rect 6825 8450 6844 8472
rect 6859 8456 6889 8472
rect 6917 8466 6923 8540
rect 6926 8466 6945 8610
rect 6960 8466 6966 8610
rect 6975 8540 6988 8610
rect 7033 8584 7062 8598
rect 7115 8584 7131 8598
rect 7169 8594 7175 8596
rect 7182 8594 7290 8610
rect 7297 8594 7303 8596
rect 7311 8594 7326 8610
rect 7392 8604 7411 8607
rect 7033 8582 7131 8584
rect 7158 8582 7326 8594
rect 7341 8584 7357 8598
rect 7392 8585 7414 8604
rect 7424 8598 7440 8599
rect 7423 8596 7440 8598
rect 7424 8591 7440 8596
rect 7414 8584 7420 8585
rect 7423 8584 7452 8591
rect 7341 8583 7452 8584
rect 7341 8582 7458 8583
rect 7017 8574 7068 8582
rect 7115 8574 7149 8582
rect 7017 8562 7042 8574
rect 7049 8562 7068 8574
rect 7122 8572 7149 8574
rect 7158 8572 7379 8582
rect 7414 8579 7420 8582
rect 7122 8568 7379 8572
rect 7017 8554 7068 8562
rect 7115 8554 7379 8568
rect 7423 8574 7458 8582
rect 6969 8506 6988 8540
rect 7033 8546 7062 8554
rect 7033 8540 7050 8546
rect 7033 8538 7067 8540
rect 7115 8538 7131 8554
rect 7132 8544 7340 8554
rect 7341 8544 7357 8554
rect 7405 8550 7420 8565
rect 7423 8562 7424 8574
rect 7431 8562 7458 8574
rect 7423 8554 7458 8562
rect 7423 8553 7452 8554
rect 7143 8540 7357 8544
rect 7158 8538 7357 8540
rect 7392 8540 7405 8550
rect 7423 8540 7440 8553
rect 7392 8538 7440 8540
rect 7034 8534 7067 8538
rect 7030 8532 7067 8534
rect 7030 8531 7097 8532
rect 7030 8526 7061 8531
rect 7067 8526 7097 8531
rect 7030 8522 7097 8526
rect 7003 8519 7097 8522
rect 7003 8512 7052 8519
rect 7003 8506 7033 8512
rect 7052 8507 7057 8512
rect 6969 8490 7049 8506
rect 7061 8498 7097 8519
rect 7158 8514 7347 8538
rect 7392 8537 7439 8538
rect 7405 8532 7439 8537
rect 7173 8511 7347 8514
rect 7166 8508 7347 8511
rect 7375 8531 7439 8532
rect 6969 8488 6988 8490
rect 7003 8488 7037 8490
rect 6969 8472 7049 8488
rect 6969 8466 6988 8472
rect 6685 8440 6788 8450
rect 6639 8438 6788 8440
rect 6809 8438 6844 8450
rect 6478 8436 6640 8438
rect 6490 8416 6509 8436
rect 6524 8434 6554 8436
rect 6373 8408 6414 8416
rect 6496 8412 6509 8416
rect 6561 8420 6640 8436
rect 6672 8436 6844 8438
rect 6672 8420 6751 8436
rect 6758 8434 6788 8436
rect 6336 8398 6365 8408
rect 6379 8398 6408 8408
rect 6423 8398 6453 8412
rect 6496 8398 6539 8412
rect 6561 8408 6751 8420
rect 6816 8416 6822 8436
rect 6546 8398 6576 8408
rect 6577 8398 6735 8408
rect 6739 8398 6769 8408
rect 6773 8398 6803 8412
rect 6831 8398 6844 8436
rect 6916 8450 6945 8466
rect 6959 8450 6988 8466
rect 7003 8456 7033 8472
rect 7061 8450 7067 8498
rect 7070 8492 7089 8498
rect 7104 8492 7134 8500
rect 7070 8484 7134 8492
rect 7070 8468 7150 8484
rect 7166 8477 7228 8508
rect 7244 8477 7306 8508
rect 7375 8506 7424 8531
rect 7439 8506 7469 8522
rect 7338 8492 7368 8500
rect 7375 8498 7485 8506
rect 7338 8484 7383 8492
rect 7070 8466 7089 8468
rect 7104 8466 7150 8468
rect 7070 8450 7150 8466
rect 7177 8464 7212 8477
rect 7253 8474 7290 8477
rect 7253 8472 7295 8474
rect 7182 8461 7212 8464
rect 7191 8457 7198 8461
rect 7198 8456 7199 8457
rect 7157 8450 7167 8456
rect 6916 8442 6951 8450
rect 6916 8416 6917 8442
rect 6924 8416 6951 8442
rect 6859 8398 6889 8412
rect 6916 8408 6951 8416
rect 6953 8442 6994 8450
rect 6953 8416 6968 8442
rect 6975 8416 6994 8442
rect 7058 8438 7089 8450
rect 7104 8438 7207 8450
rect 7219 8440 7245 8466
rect 7260 8461 7290 8472
rect 7322 8468 7384 8484
rect 7322 8466 7368 8468
rect 7322 8450 7384 8466
rect 7396 8450 7402 8498
rect 7405 8490 7485 8498
rect 7405 8488 7424 8490
rect 7439 8488 7473 8490
rect 7405 8472 7485 8488
rect 7405 8450 7424 8472
rect 7439 8456 7469 8472
rect 7497 8466 7503 8540
rect 7506 8466 7525 8610
rect 7540 8466 7546 8610
rect 7555 8540 7568 8610
rect 7613 8584 7642 8598
rect 7695 8584 7711 8598
rect 7749 8594 7755 8596
rect 7762 8594 7870 8610
rect 7877 8594 7883 8596
rect 7891 8594 7906 8610
rect 7972 8604 7991 8607
rect 7613 8582 7711 8584
rect 7738 8582 7906 8594
rect 7921 8584 7937 8598
rect 7972 8585 7994 8604
rect 8004 8598 8020 8599
rect 8003 8596 8020 8598
rect 8004 8591 8020 8596
rect 7994 8584 8000 8585
rect 8003 8584 8032 8591
rect 7921 8583 8032 8584
rect 7921 8582 8038 8583
rect 7597 8574 7648 8582
rect 7695 8574 7729 8582
rect 7597 8562 7622 8574
rect 7629 8562 7648 8574
rect 7702 8572 7729 8574
rect 7738 8572 7959 8582
rect 7994 8579 8000 8582
rect 7702 8568 7959 8572
rect 7597 8554 7648 8562
rect 7695 8554 7959 8568
rect 8003 8574 8038 8582
rect 7549 8506 7568 8540
rect 7613 8546 7642 8554
rect 7613 8540 7630 8546
rect 7613 8538 7647 8540
rect 7695 8538 7711 8554
rect 7712 8544 7920 8554
rect 7921 8544 7937 8554
rect 7985 8550 8000 8565
rect 8003 8562 8004 8574
rect 8011 8562 8038 8574
rect 8003 8554 8038 8562
rect 8003 8553 8032 8554
rect 7723 8540 7937 8544
rect 7738 8538 7937 8540
rect 7972 8540 7985 8550
rect 8003 8540 8020 8553
rect 7972 8538 8020 8540
rect 7614 8534 7647 8538
rect 7610 8532 7647 8534
rect 7610 8531 7677 8532
rect 7610 8526 7641 8531
rect 7647 8526 7677 8531
rect 7610 8522 7677 8526
rect 7583 8519 7677 8522
rect 7583 8512 7632 8519
rect 7583 8506 7613 8512
rect 7632 8507 7637 8512
rect 7549 8490 7629 8506
rect 7641 8498 7677 8519
rect 7738 8514 7927 8538
rect 7972 8537 8019 8538
rect 7985 8532 8019 8537
rect 7753 8511 7927 8514
rect 7746 8508 7927 8511
rect 7955 8531 8019 8532
rect 7549 8488 7568 8490
rect 7583 8488 7617 8490
rect 7549 8472 7629 8488
rect 7549 8466 7568 8472
rect 7265 8440 7368 8450
rect 7219 8438 7368 8440
rect 7389 8438 7424 8450
rect 7058 8436 7220 8438
rect 7070 8416 7089 8436
rect 7104 8434 7134 8436
rect 6953 8408 6994 8416
rect 7076 8412 7089 8416
rect 7141 8420 7220 8436
rect 7252 8436 7424 8438
rect 7252 8420 7331 8436
rect 7338 8434 7368 8436
rect 6916 8398 6945 8408
rect 6959 8398 6988 8408
rect 7003 8398 7033 8412
rect 7076 8398 7119 8412
rect 7141 8408 7331 8420
rect 7396 8416 7402 8436
rect 7126 8398 7156 8408
rect 7157 8398 7315 8408
rect 7319 8398 7349 8408
rect 7353 8398 7383 8412
rect 7411 8398 7424 8436
rect 7496 8450 7525 8466
rect 7539 8450 7568 8466
rect 7583 8456 7613 8472
rect 7641 8450 7647 8498
rect 7650 8492 7669 8498
rect 7684 8492 7714 8500
rect 7650 8484 7714 8492
rect 7650 8468 7730 8484
rect 7746 8477 7808 8508
rect 7824 8477 7886 8508
rect 7955 8506 8004 8531
rect 8019 8506 8049 8522
rect 7918 8492 7948 8500
rect 7955 8498 8065 8506
rect 7918 8484 7963 8492
rect 7650 8466 7669 8468
rect 7684 8466 7730 8468
rect 7650 8450 7730 8466
rect 7757 8464 7792 8477
rect 7833 8474 7870 8477
rect 7833 8472 7875 8474
rect 7762 8461 7792 8464
rect 7771 8457 7778 8461
rect 7778 8456 7779 8457
rect 7737 8450 7747 8456
rect 7496 8442 7531 8450
rect 7496 8416 7497 8442
rect 7504 8416 7531 8442
rect 7439 8398 7469 8412
rect 7496 8408 7531 8416
rect 7533 8442 7574 8450
rect 7533 8416 7548 8442
rect 7555 8416 7574 8442
rect 7638 8438 7669 8450
rect 7684 8438 7787 8450
rect 7799 8440 7825 8466
rect 7840 8461 7870 8472
rect 7902 8468 7964 8484
rect 7902 8466 7948 8468
rect 7902 8450 7964 8466
rect 7976 8450 7982 8498
rect 7985 8490 8065 8498
rect 7985 8488 8004 8490
rect 8019 8488 8053 8490
rect 7985 8472 8065 8488
rect 7985 8450 8004 8472
rect 8019 8456 8049 8472
rect 8077 8466 8083 8540
rect 8086 8466 8105 8610
rect 8120 8466 8126 8610
rect 8135 8540 8148 8610
rect 8193 8584 8222 8598
rect 8275 8584 8291 8598
rect 8329 8594 8335 8596
rect 8342 8594 8450 8610
rect 8457 8594 8463 8596
rect 8471 8594 8486 8610
rect 8552 8604 8571 8607
rect 8193 8582 8291 8584
rect 8318 8582 8486 8594
rect 8501 8584 8517 8598
rect 8552 8585 8574 8604
rect 8584 8598 8600 8599
rect 8583 8596 8600 8598
rect 8584 8591 8600 8596
rect 8574 8584 8580 8585
rect 8583 8584 8612 8591
rect 8501 8583 8612 8584
rect 8501 8582 8618 8583
rect 8177 8574 8228 8582
rect 8275 8574 8309 8582
rect 8177 8562 8202 8574
rect 8209 8562 8228 8574
rect 8282 8572 8309 8574
rect 8318 8572 8539 8582
rect 8574 8579 8580 8582
rect 8282 8568 8539 8572
rect 8177 8554 8228 8562
rect 8275 8554 8539 8568
rect 8583 8574 8618 8582
rect 8129 8506 8148 8540
rect 8193 8546 8222 8554
rect 8193 8540 8210 8546
rect 8193 8538 8227 8540
rect 8275 8538 8291 8554
rect 8292 8544 8500 8554
rect 8501 8544 8517 8554
rect 8565 8550 8580 8565
rect 8583 8562 8584 8574
rect 8591 8562 8618 8574
rect 8583 8554 8618 8562
rect 8583 8553 8612 8554
rect 8303 8540 8517 8544
rect 8318 8538 8517 8540
rect 8552 8540 8565 8550
rect 8583 8540 8600 8553
rect 8552 8538 8600 8540
rect 8194 8534 8227 8538
rect 8190 8532 8227 8534
rect 8190 8531 8257 8532
rect 8190 8526 8221 8531
rect 8227 8526 8257 8531
rect 8190 8522 8257 8526
rect 8163 8519 8257 8522
rect 8163 8512 8212 8519
rect 8163 8506 8193 8512
rect 8212 8507 8217 8512
rect 8129 8490 8209 8506
rect 8221 8498 8257 8519
rect 8318 8514 8507 8538
rect 8552 8537 8599 8538
rect 8565 8532 8599 8537
rect 8333 8511 8507 8514
rect 8326 8508 8507 8511
rect 8535 8531 8599 8532
rect 8129 8488 8148 8490
rect 8163 8488 8197 8490
rect 8129 8472 8209 8488
rect 8129 8466 8148 8472
rect 7845 8440 7948 8450
rect 7799 8438 7948 8440
rect 7969 8438 8004 8450
rect 7638 8436 7800 8438
rect 7650 8416 7669 8436
rect 7684 8434 7714 8436
rect 7533 8408 7574 8416
rect 7656 8412 7669 8416
rect 7721 8420 7800 8436
rect 7832 8436 8004 8438
rect 7832 8420 7911 8436
rect 7918 8434 7948 8436
rect 7496 8398 7525 8408
rect 7539 8398 7568 8408
rect 7583 8398 7613 8412
rect 7656 8398 7699 8412
rect 7721 8408 7911 8420
rect 7976 8416 7982 8436
rect 7706 8398 7736 8408
rect 7737 8398 7895 8408
rect 7899 8398 7929 8408
rect 7933 8398 7963 8412
rect 7991 8398 8004 8436
rect 8076 8450 8105 8466
rect 8119 8450 8148 8466
rect 8163 8456 8193 8472
rect 8221 8450 8227 8498
rect 8230 8492 8249 8498
rect 8264 8492 8294 8500
rect 8230 8484 8294 8492
rect 8230 8468 8310 8484
rect 8326 8477 8388 8508
rect 8404 8477 8466 8508
rect 8535 8506 8584 8531
rect 8599 8506 8629 8522
rect 8498 8492 8528 8500
rect 8535 8498 8645 8506
rect 8498 8484 8543 8492
rect 8230 8466 8249 8468
rect 8264 8466 8310 8468
rect 8230 8450 8310 8466
rect 8337 8464 8372 8477
rect 8413 8474 8450 8477
rect 8413 8472 8455 8474
rect 8342 8461 8372 8464
rect 8351 8457 8358 8461
rect 8358 8456 8359 8457
rect 8317 8450 8327 8456
rect 8076 8442 8111 8450
rect 8076 8416 8077 8442
rect 8084 8416 8111 8442
rect 8019 8398 8049 8412
rect 8076 8408 8111 8416
rect 8113 8442 8154 8450
rect 8113 8416 8128 8442
rect 8135 8416 8154 8442
rect 8218 8438 8249 8450
rect 8264 8438 8367 8450
rect 8379 8440 8405 8466
rect 8420 8461 8450 8472
rect 8482 8468 8544 8484
rect 8482 8466 8528 8468
rect 8482 8450 8544 8466
rect 8556 8450 8562 8498
rect 8565 8490 8645 8498
rect 8565 8488 8584 8490
rect 8599 8488 8633 8490
rect 8565 8472 8645 8488
rect 8565 8450 8584 8472
rect 8599 8456 8629 8472
rect 8657 8466 8663 8540
rect 8666 8466 8685 8610
rect 8700 8466 8706 8610
rect 8715 8540 8728 8610
rect 8773 8584 8802 8598
rect 8855 8584 8871 8598
rect 8909 8594 8915 8596
rect 8922 8594 9030 8610
rect 9037 8594 9043 8596
rect 9051 8594 9066 8610
rect 9132 8604 9151 8607
rect 8773 8582 8871 8584
rect 8898 8582 9066 8594
rect 9081 8584 9097 8598
rect 9132 8585 9154 8604
rect 9164 8598 9180 8599
rect 9163 8596 9180 8598
rect 9164 8591 9180 8596
rect 9154 8584 9160 8585
rect 9163 8584 9192 8591
rect 9081 8583 9192 8584
rect 9081 8582 9198 8583
rect 8757 8574 8808 8582
rect 8855 8574 8889 8582
rect 8757 8562 8782 8574
rect 8789 8562 8808 8574
rect 8862 8572 8889 8574
rect 8898 8572 9119 8582
rect 9154 8579 9160 8582
rect 8862 8568 9119 8572
rect 8757 8554 8808 8562
rect 8855 8554 9119 8568
rect 9163 8574 9198 8582
rect 8709 8506 8728 8540
rect 8773 8546 8802 8554
rect 8773 8540 8790 8546
rect 8773 8538 8807 8540
rect 8855 8538 8871 8554
rect 8872 8544 9080 8554
rect 9081 8544 9097 8554
rect 9145 8550 9160 8565
rect 9163 8562 9164 8574
rect 9171 8562 9198 8574
rect 9163 8554 9198 8562
rect 9163 8553 9192 8554
rect 8883 8540 9097 8544
rect 8898 8538 9097 8540
rect 9132 8540 9145 8550
rect 9163 8540 9180 8553
rect 9132 8538 9180 8540
rect 8774 8534 8807 8538
rect 8770 8532 8807 8534
rect 8770 8531 8837 8532
rect 8770 8526 8801 8531
rect 8807 8526 8837 8531
rect 8770 8522 8837 8526
rect 8743 8519 8837 8522
rect 8743 8512 8792 8519
rect 8743 8506 8773 8512
rect 8792 8507 8797 8512
rect 8709 8490 8789 8506
rect 8801 8498 8837 8519
rect 8898 8514 9087 8538
rect 9132 8537 9179 8538
rect 9145 8532 9179 8537
rect 8913 8511 9087 8514
rect 8906 8508 9087 8511
rect 9115 8531 9179 8532
rect 8709 8488 8728 8490
rect 8743 8488 8777 8490
rect 8709 8472 8789 8488
rect 8709 8466 8728 8472
rect 8425 8440 8528 8450
rect 8379 8438 8528 8440
rect 8549 8438 8584 8450
rect 8218 8436 8380 8438
rect 8230 8416 8249 8436
rect 8264 8434 8294 8436
rect 8113 8408 8154 8416
rect 8236 8412 8249 8416
rect 8301 8420 8380 8436
rect 8412 8436 8584 8438
rect 8412 8420 8491 8436
rect 8498 8434 8528 8436
rect 8076 8398 8105 8408
rect 8119 8398 8148 8408
rect 8163 8398 8193 8412
rect 8236 8398 8279 8412
rect 8301 8408 8491 8420
rect 8556 8416 8562 8436
rect 8286 8398 8316 8408
rect 8317 8398 8475 8408
rect 8479 8398 8509 8408
rect 8513 8398 8543 8412
rect 8571 8398 8584 8436
rect 8656 8450 8685 8466
rect 8699 8450 8728 8466
rect 8743 8456 8773 8472
rect 8801 8450 8807 8498
rect 8810 8492 8829 8498
rect 8844 8492 8874 8500
rect 8810 8484 8874 8492
rect 8810 8468 8890 8484
rect 8906 8477 8968 8508
rect 8984 8477 9046 8508
rect 9115 8506 9164 8531
rect 9179 8506 9209 8522
rect 9078 8492 9108 8500
rect 9115 8498 9225 8506
rect 9078 8484 9123 8492
rect 8810 8466 8829 8468
rect 8844 8466 8890 8468
rect 8810 8450 8890 8466
rect 8917 8464 8952 8477
rect 8993 8474 9030 8477
rect 8993 8472 9035 8474
rect 8922 8461 8952 8464
rect 8931 8457 8938 8461
rect 8938 8456 8939 8457
rect 8897 8450 8907 8456
rect 8656 8442 8691 8450
rect 8656 8416 8657 8442
rect 8664 8416 8691 8442
rect 8599 8398 8629 8412
rect 8656 8408 8691 8416
rect 8693 8442 8734 8450
rect 8693 8416 8708 8442
rect 8715 8416 8734 8442
rect 8798 8438 8829 8450
rect 8844 8438 8947 8450
rect 8959 8440 8985 8466
rect 9000 8461 9030 8472
rect 9062 8468 9124 8484
rect 9062 8466 9108 8468
rect 9062 8450 9124 8466
rect 9136 8450 9142 8498
rect 9145 8490 9225 8498
rect 9145 8488 9164 8490
rect 9179 8488 9213 8490
rect 9145 8472 9225 8488
rect 9145 8450 9164 8472
rect 9179 8456 9209 8472
rect 9237 8466 9243 8540
rect 9246 8466 9265 8610
rect 9280 8466 9286 8610
rect 9295 8540 9308 8610
rect 9353 8584 9382 8598
rect 9435 8584 9451 8598
rect 9489 8594 9495 8596
rect 9502 8594 9610 8610
rect 9617 8594 9623 8596
rect 9631 8594 9646 8610
rect 9712 8604 9731 8607
rect 9353 8582 9451 8584
rect 9478 8582 9646 8594
rect 9661 8584 9677 8598
rect 9712 8585 9734 8604
rect 9744 8598 9760 8599
rect 9743 8596 9760 8598
rect 9744 8591 9760 8596
rect 9734 8584 9740 8585
rect 9743 8584 9772 8591
rect 9661 8583 9772 8584
rect 9661 8582 9778 8583
rect 9337 8574 9388 8582
rect 9435 8574 9469 8582
rect 9337 8562 9362 8574
rect 9369 8562 9388 8574
rect 9442 8572 9469 8574
rect 9478 8572 9699 8582
rect 9734 8579 9740 8582
rect 9442 8568 9699 8572
rect 9337 8554 9388 8562
rect 9435 8554 9699 8568
rect 9743 8574 9778 8582
rect 9289 8506 9308 8540
rect 9353 8546 9382 8554
rect 9353 8540 9370 8546
rect 9353 8538 9387 8540
rect 9435 8538 9451 8554
rect 9452 8544 9660 8554
rect 9661 8544 9677 8554
rect 9725 8550 9740 8565
rect 9743 8562 9744 8574
rect 9751 8562 9778 8574
rect 9743 8554 9778 8562
rect 9743 8553 9772 8554
rect 9463 8540 9677 8544
rect 9478 8538 9677 8540
rect 9712 8540 9725 8550
rect 9743 8540 9760 8553
rect 9712 8538 9760 8540
rect 9354 8534 9387 8538
rect 9350 8532 9387 8534
rect 9350 8531 9417 8532
rect 9350 8526 9381 8531
rect 9387 8526 9417 8531
rect 9350 8522 9417 8526
rect 9323 8519 9417 8522
rect 9323 8512 9372 8519
rect 9323 8506 9353 8512
rect 9372 8507 9377 8512
rect 9289 8490 9369 8506
rect 9381 8498 9417 8519
rect 9478 8514 9667 8538
rect 9712 8537 9759 8538
rect 9725 8532 9759 8537
rect 9493 8511 9667 8514
rect 9486 8508 9667 8511
rect 9695 8531 9759 8532
rect 9289 8488 9308 8490
rect 9323 8488 9357 8490
rect 9289 8472 9369 8488
rect 9289 8466 9308 8472
rect 9005 8440 9108 8450
rect 8959 8438 9108 8440
rect 9129 8438 9164 8450
rect 8798 8436 8960 8438
rect 8810 8416 8829 8436
rect 8844 8434 8874 8436
rect 8693 8408 8734 8416
rect 8816 8412 8829 8416
rect 8881 8420 8960 8436
rect 8992 8436 9164 8438
rect 8992 8420 9071 8436
rect 9078 8434 9108 8436
rect 8656 8398 8685 8408
rect 8699 8398 8728 8408
rect 8743 8398 8773 8412
rect 8816 8398 8859 8412
rect 8881 8408 9071 8420
rect 9136 8416 9142 8436
rect 8866 8398 8896 8408
rect 8897 8398 9055 8408
rect 9059 8398 9089 8408
rect 9093 8398 9123 8412
rect 9151 8398 9164 8436
rect 9236 8450 9265 8466
rect 9279 8450 9308 8466
rect 9323 8456 9353 8472
rect 9381 8450 9387 8498
rect 9390 8492 9409 8498
rect 9424 8492 9454 8500
rect 9390 8484 9454 8492
rect 9390 8468 9470 8484
rect 9486 8477 9548 8508
rect 9564 8477 9626 8508
rect 9695 8506 9744 8531
rect 9759 8506 9789 8522
rect 9658 8492 9688 8500
rect 9695 8498 9805 8506
rect 9658 8484 9703 8492
rect 9390 8466 9409 8468
rect 9424 8466 9470 8468
rect 9390 8450 9470 8466
rect 9497 8464 9532 8477
rect 9573 8474 9610 8477
rect 9573 8472 9615 8474
rect 9502 8461 9532 8464
rect 9511 8457 9518 8461
rect 9518 8456 9519 8457
rect 9477 8450 9487 8456
rect 9236 8442 9271 8450
rect 9236 8416 9237 8442
rect 9244 8416 9271 8442
rect 9179 8398 9209 8412
rect 9236 8408 9271 8416
rect 9273 8442 9314 8450
rect 9273 8416 9288 8442
rect 9295 8416 9314 8442
rect 9378 8438 9409 8450
rect 9424 8438 9527 8450
rect 9539 8440 9565 8466
rect 9580 8461 9610 8472
rect 9642 8468 9704 8484
rect 9642 8466 9688 8468
rect 9642 8450 9704 8466
rect 9716 8450 9722 8498
rect 9725 8490 9805 8498
rect 9725 8488 9744 8490
rect 9759 8488 9793 8490
rect 9725 8472 9805 8488
rect 9725 8450 9744 8472
rect 9759 8456 9789 8472
rect 9817 8466 9823 8540
rect 9826 8466 9845 8610
rect 9860 8466 9866 8610
rect 9875 8540 9888 8610
rect 9933 8584 9962 8598
rect 10015 8584 10031 8598
rect 10069 8594 10075 8596
rect 10082 8594 10190 8610
rect 10197 8594 10203 8596
rect 10211 8594 10226 8610
rect 10292 8604 10311 8607
rect 9933 8582 10031 8584
rect 10058 8582 10226 8594
rect 10241 8584 10257 8598
rect 10292 8585 10314 8604
rect 10324 8598 10340 8599
rect 10323 8596 10340 8598
rect 10324 8591 10340 8596
rect 10314 8584 10320 8585
rect 10323 8584 10352 8591
rect 10241 8583 10352 8584
rect 10241 8582 10358 8583
rect 9917 8574 9968 8582
rect 10015 8574 10049 8582
rect 9917 8562 9942 8574
rect 9949 8562 9968 8574
rect 10022 8572 10049 8574
rect 10058 8572 10279 8582
rect 10314 8579 10320 8582
rect 10022 8568 10279 8572
rect 9917 8554 9968 8562
rect 10015 8554 10279 8568
rect 10323 8574 10358 8582
rect 9869 8506 9888 8540
rect 9933 8546 9962 8554
rect 9933 8540 9950 8546
rect 9933 8538 9967 8540
rect 10015 8538 10031 8554
rect 10032 8544 10240 8554
rect 10241 8544 10257 8554
rect 10305 8550 10320 8565
rect 10323 8562 10324 8574
rect 10331 8562 10358 8574
rect 10323 8554 10358 8562
rect 10323 8553 10352 8554
rect 10043 8540 10257 8544
rect 10058 8538 10257 8540
rect 10292 8540 10305 8550
rect 10323 8540 10340 8553
rect 10292 8538 10340 8540
rect 9934 8534 9967 8538
rect 9930 8532 9967 8534
rect 9930 8531 9997 8532
rect 9930 8526 9961 8531
rect 9967 8526 9997 8531
rect 9930 8522 9997 8526
rect 9903 8519 9997 8522
rect 9903 8512 9952 8519
rect 9903 8506 9933 8512
rect 9952 8507 9957 8512
rect 9869 8490 9949 8506
rect 9961 8498 9997 8519
rect 10058 8514 10247 8538
rect 10292 8537 10339 8538
rect 10305 8532 10339 8537
rect 10073 8511 10247 8514
rect 10066 8508 10247 8511
rect 10275 8531 10339 8532
rect 9869 8488 9888 8490
rect 9903 8488 9937 8490
rect 9869 8472 9949 8488
rect 9869 8466 9888 8472
rect 9585 8440 9688 8450
rect 9539 8438 9688 8440
rect 9709 8438 9744 8450
rect 9378 8436 9540 8438
rect 9390 8416 9409 8436
rect 9424 8434 9454 8436
rect 9273 8408 9314 8416
rect 9396 8412 9409 8416
rect 9461 8420 9540 8436
rect 9572 8436 9744 8438
rect 9572 8420 9651 8436
rect 9658 8434 9688 8436
rect 9236 8398 9265 8408
rect 9279 8398 9308 8408
rect 9323 8398 9353 8412
rect 9396 8398 9439 8412
rect 9461 8408 9651 8420
rect 9716 8416 9722 8436
rect 9446 8398 9476 8408
rect 9477 8398 9635 8408
rect 9639 8398 9669 8408
rect 9673 8398 9703 8412
rect 9731 8398 9744 8436
rect 9816 8450 9845 8466
rect 9859 8450 9888 8466
rect 9903 8456 9933 8472
rect 9961 8450 9967 8498
rect 9970 8492 9989 8498
rect 10004 8492 10034 8500
rect 9970 8484 10034 8492
rect 9970 8468 10050 8484
rect 10066 8477 10128 8508
rect 10144 8477 10206 8508
rect 10275 8506 10324 8531
rect 10339 8506 10369 8522
rect 10238 8492 10268 8500
rect 10275 8498 10385 8506
rect 10238 8484 10283 8492
rect 9970 8466 9989 8468
rect 10004 8466 10050 8468
rect 9970 8450 10050 8466
rect 10077 8464 10112 8477
rect 10153 8474 10190 8477
rect 10153 8472 10195 8474
rect 10082 8461 10112 8464
rect 10091 8457 10098 8461
rect 10098 8456 10099 8457
rect 10057 8450 10067 8456
rect 9816 8442 9851 8450
rect 9816 8416 9817 8442
rect 9824 8416 9851 8442
rect 9759 8398 9789 8412
rect 9816 8408 9851 8416
rect 9853 8442 9894 8450
rect 9853 8416 9868 8442
rect 9875 8416 9894 8442
rect 9958 8438 9989 8450
rect 10004 8438 10107 8450
rect 10119 8440 10145 8466
rect 10160 8461 10190 8472
rect 10222 8468 10284 8484
rect 10222 8466 10268 8468
rect 10222 8450 10284 8466
rect 10296 8450 10302 8498
rect 10305 8490 10385 8498
rect 10305 8488 10324 8490
rect 10339 8488 10373 8490
rect 10305 8472 10385 8488
rect 10305 8450 10324 8472
rect 10339 8456 10369 8472
rect 10397 8466 10403 8540
rect 10406 8466 10425 8610
rect 10440 8466 10446 8610
rect 10455 8540 10468 8610
rect 10513 8584 10542 8598
rect 10595 8584 10611 8598
rect 10649 8594 10655 8596
rect 10662 8594 10770 8610
rect 10777 8594 10783 8596
rect 10791 8594 10806 8610
rect 10872 8604 10891 8607
rect 10513 8582 10611 8584
rect 10638 8582 10806 8594
rect 10821 8584 10837 8598
rect 10872 8585 10894 8604
rect 10904 8598 10920 8599
rect 10903 8596 10920 8598
rect 10904 8591 10920 8596
rect 10894 8584 10900 8585
rect 10903 8584 10932 8591
rect 10821 8583 10932 8584
rect 10821 8582 10938 8583
rect 10497 8574 10548 8582
rect 10595 8574 10629 8582
rect 10497 8562 10522 8574
rect 10529 8562 10548 8574
rect 10602 8572 10629 8574
rect 10638 8572 10859 8582
rect 10894 8579 10900 8582
rect 10602 8568 10859 8572
rect 10497 8554 10548 8562
rect 10595 8554 10859 8568
rect 10903 8574 10938 8582
rect 10449 8506 10468 8540
rect 10513 8546 10542 8554
rect 10513 8540 10530 8546
rect 10513 8538 10547 8540
rect 10595 8538 10611 8554
rect 10612 8544 10820 8554
rect 10821 8544 10837 8554
rect 10885 8550 10900 8565
rect 10903 8562 10904 8574
rect 10911 8562 10938 8574
rect 10903 8554 10938 8562
rect 10903 8553 10932 8554
rect 10623 8540 10837 8544
rect 10638 8538 10837 8540
rect 10872 8540 10885 8550
rect 10903 8540 10920 8553
rect 10872 8538 10920 8540
rect 10514 8534 10547 8538
rect 10510 8532 10547 8534
rect 10510 8531 10577 8532
rect 10510 8526 10541 8531
rect 10547 8526 10577 8531
rect 10510 8522 10577 8526
rect 10483 8519 10577 8522
rect 10483 8512 10532 8519
rect 10483 8506 10513 8512
rect 10532 8507 10537 8512
rect 10449 8490 10529 8506
rect 10541 8498 10577 8519
rect 10638 8514 10827 8538
rect 10872 8537 10919 8538
rect 10885 8532 10919 8537
rect 10653 8511 10827 8514
rect 10646 8508 10827 8511
rect 10855 8531 10919 8532
rect 10449 8488 10468 8490
rect 10483 8488 10517 8490
rect 10449 8472 10529 8488
rect 10449 8466 10468 8472
rect 10165 8440 10268 8450
rect 10119 8438 10268 8440
rect 10289 8438 10324 8450
rect 9958 8436 10120 8438
rect 9970 8416 9989 8436
rect 10004 8434 10034 8436
rect 9853 8408 9894 8416
rect 9976 8412 9989 8416
rect 10041 8420 10120 8436
rect 10152 8436 10324 8438
rect 10152 8420 10231 8436
rect 10238 8434 10268 8436
rect 9816 8398 9845 8408
rect 9859 8398 9888 8408
rect 9903 8398 9933 8412
rect 9976 8398 10019 8412
rect 10041 8408 10231 8420
rect 10296 8416 10302 8436
rect 10026 8398 10056 8408
rect 10057 8398 10215 8408
rect 10219 8398 10249 8408
rect 10253 8398 10283 8412
rect 10311 8398 10324 8436
rect 10396 8450 10425 8466
rect 10439 8450 10468 8466
rect 10483 8456 10513 8472
rect 10541 8450 10547 8498
rect 10550 8492 10569 8498
rect 10584 8492 10614 8500
rect 10550 8484 10614 8492
rect 10550 8468 10630 8484
rect 10646 8477 10708 8508
rect 10724 8477 10786 8508
rect 10855 8506 10904 8531
rect 10919 8506 10949 8522
rect 10818 8492 10848 8500
rect 10855 8498 10965 8506
rect 10818 8484 10863 8492
rect 10550 8466 10569 8468
rect 10584 8466 10630 8468
rect 10550 8450 10630 8466
rect 10657 8464 10692 8477
rect 10733 8474 10770 8477
rect 10733 8472 10775 8474
rect 10662 8461 10692 8464
rect 10671 8457 10678 8461
rect 10678 8456 10679 8457
rect 10637 8450 10647 8456
rect 10396 8442 10431 8450
rect 10396 8416 10397 8442
rect 10404 8416 10431 8442
rect 10339 8398 10369 8412
rect 10396 8408 10431 8416
rect 10433 8442 10474 8450
rect 10433 8416 10448 8442
rect 10455 8416 10474 8442
rect 10538 8438 10569 8450
rect 10584 8438 10687 8450
rect 10699 8440 10725 8466
rect 10740 8461 10770 8472
rect 10802 8468 10864 8484
rect 10802 8466 10848 8468
rect 10802 8450 10864 8466
rect 10876 8450 10882 8498
rect 10885 8490 10965 8498
rect 10885 8488 10904 8490
rect 10919 8488 10953 8490
rect 10885 8472 10965 8488
rect 10885 8450 10904 8472
rect 10919 8456 10949 8472
rect 10977 8466 10983 8540
rect 10986 8466 11005 8610
rect 11020 8466 11026 8610
rect 11035 8540 11048 8610
rect 11093 8584 11122 8598
rect 11175 8584 11191 8598
rect 11229 8594 11235 8596
rect 11242 8594 11350 8610
rect 11357 8594 11363 8596
rect 11371 8594 11386 8610
rect 11452 8604 11471 8607
rect 11093 8582 11191 8584
rect 11218 8582 11386 8594
rect 11401 8584 11417 8598
rect 11452 8585 11474 8604
rect 11484 8598 11500 8599
rect 11483 8596 11500 8598
rect 11484 8591 11500 8596
rect 11474 8584 11480 8585
rect 11483 8584 11512 8591
rect 11401 8583 11512 8584
rect 11401 8582 11518 8583
rect 11077 8574 11128 8582
rect 11175 8574 11209 8582
rect 11077 8562 11102 8574
rect 11109 8562 11128 8574
rect 11182 8572 11209 8574
rect 11218 8572 11439 8582
rect 11474 8579 11480 8582
rect 11182 8568 11439 8572
rect 11077 8554 11128 8562
rect 11175 8554 11439 8568
rect 11483 8574 11518 8582
rect 11029 8506 11048 8540
rect 11093 8546 11122 8554
rect 11093 8540 11110 8546
rect 11093 8538 11127 8540
rect 11175 8538 11191 8554
rect 11192 8544 11400 8554
rect 11401 8544 11417 8554
rect 11465 8550 11480 8565
rect 11483 8562 11484 8574
rect 11491 8562 11518 8574
rect 11483 8554 11518 8562
rect 11483 8553 11512 8554
rect 11203 8540 11417 8544
rect 11218 8538 11417 8540
rect 11452 8540 11465 8550
rect 11483 8540 11500 8553
rect 11452 8538 11500 8540
rect 11094 8534 11127 8538
rect 11090 8532 11127 8534
rect 11090 8531 11157 8532
rect 11090 8526 11121 8531
rect 11127 8526 11157 8531
rect 11090 8522 11157 8526
rect 11063 8519 11157 8522
rect 11063 8512 11112 8519
rect 11063 8506 11093 8512
rect 11112 8507 11117 8512
rect 11029 8490 11109 8506
rect 11121 8498 11157 8519
rect 11218 8514 11407 8538
rect 11452 8537 11499 8538
rect 11465 8532 11499 8537
rect 11233 8511 11407 8514
rect 11226 8508 11407 8511
rect 11435 8531 11499 8532
rect 11029 8488 11048 8490
rect 11063 8488 11097 8490
rect 11029 8472 11109 8488
rect 11029 8466 11048 8472
rect 10745 8440 10848 8450
rect 10699 8438 10848 8440
rect 10869 8438 10904 8450
rect 10538 8436 10700 8438
rect 10550 8416 10569 8436
rect 10584 8434 10614 8436
rect 10433 8408 10474 8416
rect 10556 8412 10569 8416
rect 10621 8420 10700 8436
rect 10732 8436 10904 8438
rect 10732 8420 10811 8436
rect 10818 8434 10848 8436
rect 10396 8398 10425 8408
rect 10439 8398 10468 8408
rect 10483 8398 10513 8412
rect 10556 8398 10599 8412
rect 10621 8408 10811 8420
rect 10876 8416 10882 8436
rect 10606 8398 10636 8408
rect 10637 8398 10795 8408
rect 10799 8398 10829 8408
rect 10833 8398 10863 8412
rect 10891 8398 10904 8436
rect 10976 8450 11005 8466
rect 11019 8450 11048 8466
rect 11063 8456 11093 8472
rect 11121 8450 11127 8498
rect 11130 8492 11149 8498
rect 11164 8492 11194 8500
rect 11130 8484 11194 8492
rect 11130 8468 11210 8484
rect 11226 8477 11288 8508
rect 11304 8477 11366 8508
rect 11435 8506 11484 8531
rect 11499 8506 11529 8522
rect 11398 8492 11428 8500
rect 11435 8498 11545 8506
rect 11398 8484 11443 8492
rect 11130 8466 11149 8468
rect 11164 8466 11210 8468
rect 11130 8450 11210 8466
rect 11237 8464 11272 8477
rect 11313 8474 11350 8477
rect 11313 8472 11355 8474
rect 11242 8461 11272 8464
rect 11251 8457 11258 8461
rect 11258 8456 11259 8457
rect 11217 8450 11227 8456
rect 10976 8442 11011 8450
rect 10976 8416 10977 8442
rect 10984 8416 11011 8442
rect 10919 8398 10949 8412
rect 10976 8408 11011 8416
rect 11013 8442 11054 8450
rect 11013 8416 11028 8442
rect 11035 8416 11054 8442
rect 11118 8438 11149 8450
rect 11164 8438 11267 8450
rect 11279 8440 11305 8466
rect 11320 8461 11350 8472
rect 11382 8468 11444 8484
rect 11382 8466 11428 8468
rect 11382 8450 11444 8466
rect 11456 8450 11462 8498
rect 11465 8490 11545 8498
rect 11465 8488 11484 8490
rect 11499 8488 11533 8490
rect 11465 8472 11545 8488
rect 11465 8450 11484 8472
rect 11499 8456 11529 8472
rect 11557 8466 11563 8540
rect 11566 8466 11585 8610
rect 11600 8466 11606 8610
rect 11615 8540 11628 8610
rect 11673 8584 11702 8598
rect 11755 8584 11771 8598
rect 11809 8594 11815 8596
rect 11822 8594 11930 8610
rect 11937 8594 11943 8596
rect 11951 8594 11966 8610
rect 12032 8604 12051 8607
rect 11673 8582 11771 8584
rect 11798 8582 11966 8594
rect 11981 8584 11997 8598
rect 12032 8585 12054 8604
rect 12064 8598 12080 8599
rect 12063 8596 12080 8598
rect 12064 8591 12080 8596
rect 12054 8584 12060 8585
rect 12063 8584 12092 8591
rect 11981 8583 12092 8584
rect 11981 8582 12098 8583
rect 11657 8574 11708 8582
rect 11755 8574 11789 8582
rect 11657 8562 11682 8574
rect 11689 8562 11708 8574
rect 11762 8572 11789 8574
rect 11798 8572 12019 8582
rect 12054 8579 12060 8582
rect 11762 8568 12019 8572
rect 11657 8554 11708 8562
rect 11755 8554 12019 8568
rect 12063 8574 12098 8582
rect 11609 8506 11628 8540
rect 11673 8546 11702 8554
rect 11673 8540 11690 8546
rect 11673 8538 11707 8540
rect 11755 8538 11771 8554
rect 11772 8544 11980 8554
rect 11981 8544 11997 8554
rect 12045 8550 12060 8565
rect 12063 8562 12064 8574
rect 12071 8562 12098 8574
rect 12063 8554 12098 8562
rect 12063 8553 12092 8554
rect 11783 8540 11997 8544
rect 11798 8538 11997 8540
rect 12032 8540 12045 8550
rect 12063 8540 12080 8553
rect 12032 8538 12080 8540
rect 11674 8534 11707 8538
rect 11670 8532 11707 8534
rect 11670 8531 11737 8532
rect 11670 8526 11701 8531
rect 11707 8526 11737 8531
rect 11670 8522 11737 8526
rect 11643 8519 11737 8522
rect 11643 8512 11692 8519
rect 11643 8506 11673 8512
rect 11692 8507 11697 8512
rect 11609 8490 11689 8506
rect 11701 8498 11737 8519
rect 11798 8514 11987 8538
rect 12032 8537 12079 8538
rect 12045 8532 12079 8537
rect 11813 8511 11987 8514
rect 11806 8508 11987 8511
rect 12015 8531 12079 8532
rect 11609 8488 11628 8490
rect 11643 8488 11677 8490
rect 11609 8472 11689 8488
rect 11609 8466 11628 8472
rect 11325 8440 11428 8450
rect 11279 8438 11428 8440
rect 11449 8438 11484 8450
rect 11118 8436 11280 8438
rect 11130 8416 11149 8436
rect 11164 8434 11194 8436
rect 11013 8408 11054 8416
rect 11136 8412 11149 8416
rect 11201 8420 11280 8436
rect 11312 8436 11484 8438
rect 11312 8420 11391 8436
rect 11398 8434 11428 8436
rect 10976 8398 11005 8408
rect 11019 8398 11048 8408
rect 11063 8398 11093 8412
rect 11136 8398 11179 8412
rect 11201 8408 11391 8420
rect 11456 8416 11462 8436
rect 11186 8398 11216 8408
rect 11217 8398 11375 8408
rect 11379 8398 11409 8408
rect 11413 8398 11443 8412
rect 11471 8398 11484 8436
rect 11556 8450 11585 8466
rect 11599 8450 11628 8466
rect 11643 8456 11673 8472
rect 11701 8450 11707 8498
rect 11710 8492 11729 8498
rect 11744 8492 11774 8500
rect 11710 8484 11774 8492
rect 11710 8468 11790 8484
rect 11806 8477 11868 8508
rect 11884 8477 11946 8508
rect 12015 8506 12064 8531
rect 12079 8506 12109 8522
rect 11978 8492 12008 8500
rect 12015 8498 12125 8506
rect 11978 8484 12023 8492
rect 11710 8466 11729 8468
rect 11744 8466 11790 8468
rect 11710 8450 11790 8466
rect 11817 8464 11852 8477
rect 11893 8474 11930 8477
rect 11893 8472 11935 8474
rect 11822 8461 11852 8464
rect 11831 8457 11838 8461
rect 11838 8456 11839 8457
rect 11797 8450 11807 8456
rect 11556 8442 11591 8450
rect 11556 8416 11557 8442
rect 11564 8416 11591 8442
rect 11499 8398 11529 8412
rect 11556 8408 11591 8416
rect 11593 8442 11634 8450
rect 11593 8416 11608 8442
rect 11615 8416 11634 8442
rect 11698 8438 11729 8450
rect 11744 8438 11847 8450
rect 11859 8440 11885 8466
rect 11900 8461 11930 8472
rect 11962 8468 12024 8484
rect 11962 8466 12008 8468
rect 11962 8450 12024 8466
rect 12036 8450 12042 8498
rect 12045 8490 12125 8498
rect 12045 8488 12064 8490
rect 12079 8488 12113 8490
rect 12045 8472 12125 8488
rect 12045 8450 12064 8472
rect 12079 8456 12109 8472
rect 12137 8466 12143 8540
rect 12146 8466 12165 8610
rect 12180 8466 12186 8610
rect 12195 8540 12208 8610
rect 12253 8584 12282 8598
rect 12335 8584 12351 8598
rect 12389 8594 12395 8596
rect 12402 8594 12510 8610
rect 12517 8594 12523 8596
rect 12531 8594 12546 8610
rect 12612 8604 12631 8607
rect 12253 8582 12351 8584
rect 12378 8582 12546 8594
rect 12561 8584 12577 8598
rect 12612 8585 12634 8604
rect 12644 8598 12660 8599
rect 12643 8596 12660 8598
rect 12644 8591 12660 8596
rect 12634 8584 12640 8585
rect 12643 8584 12672 8591
rect 12561 8583 12672 8584
rect 12561 8582 12678 8583
rect 12237 8574 12288 8582
rect 12335 8574 12369 8582
rect 12237 8562 12262 8574
rect 12269 8562 12288 8574
rect 12342 8572 12369 8574
rect 12378 8572 12599 8582
rect 12634 8579 12640 8582
rect 12342 8568 12599 8572
rect 12237 8554 12288 8562
rect 12335 8554 12599 8568
rect 12643 8574 12678 8582
rect 12189 8506 12208 8540
rect 12253 8546 12282 8554
rect 12253 8540 12270 8546
rect 12253 8538 12287 8540
rect 12335 8538 12351 8554
rect 12352 8544 12560 8554
rect 12561 8544 12577 8554
rect 12625 8550 12640 8565
rect 12643 8562 12644 8574
rect 12651 8562 12678 8574
rect 12643 8554 12678 8562
rect 12643 8553 12672 8554
rect 12363 8540 12577 8544
rect 12378 8538 12577 8540
rect 12612 8540 12625 8550
rect 12643 8540 12660 8553
rect 12612 8538 12660 8540
rect 12254 8534 12287 8538
rect 12250 8532 12287 8534
rect 12250 8531 12317 8532
rect 12250 8526 12281 8531
rect 12287 8526 12317 8531
rect 12250 8522 12317 8526
rect 12223 8519 12317 8522
rect 12223 8512 12272 8519
rect 12223 8506 12253 8512
rect 12272 8507 12277 8512
rect 12189 8490 12269 8506
rect 12281 8498 12317 8519
rect 12378 8514 12567 8538
rect 12612 8537 12659 8538
rect 12625 8532 12659 8537
rect 12393 8511 12567 8514
rect 12386 8508 12567 8511
rect 12595 8531 12659 8532
rect 12189 8488 12208 8490
rect 12223 8488 12257 8490
rect 12189 8472 12269 8488
rect 12189 8466 12208 8472
rect 11905 8440 12008 8450
rect 11859 8438 12008 8440
rect 12029 8438 12064 8450
rect 11698 8436 11860 8438
rect 11710 8416 11729 8436
rect 11744 8434 11774 8436
rect 11593 8408 11634 8416
rect 11716 8412 11729 8416
rect 11781 8420 11860 8436
rect 11892 8436 12064 8438
rect 11892 8420 11971 8436
rect 11978 8434 12008 8436
rect 11556 8398 11585 8408
rect 11599 8398 11628 8408
rect 11643 8398 11673 8412
rect 11716 8398 11759 8412
rect 11781 8408 11971 8420
rect 12036 8416 12042 8436
rect 11766 8398 11796 8408
rect 11797 8398 11955 8408
rect 11959 8398 11989 8408
rect 11993 8398 12023 8412
rect 12051 8398 12064 8436
rect 12136 8450 12165 8466
rect 12179 8450 12208 8466
rect 12223 8456 12253 8472
rect 12281 8450 12287 8498
rect 12290 8492 12309 8498
rect 12324 8492 12354 8500
rect 12290 8484 12354 8492
rect 12290 8468 12370 8484
rect 12386 8477 12448 8508
rect 12464 8477 12526 8508
rect 12595 8506 12644 8531
rect 12659 8506 12689 8522
rect 12558 8492 12588 8500
rect 12595 8498 12705 8506
rect 12558 8484 12603 8492
rect 12290 8466 12309 8468
rect 12324 8466 12370 8468
rect 12290 8450 12370 8466
rect 12397 8464 12432 8477
rect 12473 8474 12510 8477
rect 12473 8472 12515 8474
rect 12402 8461 12432 8464
rect 12411 8457 12418 8461
rect 12418 8456 12419 8457
rect 12377 8450 12387 8456
rect 12136 8442 12171 8450
rect 12136 8416 12137 8442
rect 12144 8416 12171 8442
rect 12079 8398 12109 8412
rect 12136 8408 12171 8416
rect 12173 8442 12214 8450
rect 12173 8416 12188 8442
rect 12195 8416 12214 8442
rect 12278 8438 12309 8450
rect 12324 8438 12427 8450
rect 12439 8440 12465 8466
rect 12480 8461 12510 8472
rect 12542 8468 12604 8484
rect 12542 8466 12588 8468
rect 12542 8450 12604 8466
rect 12616 8450 12622 8498
rect 12625 8490 12705 8498
rect 12625 8488 12644 8490
rect 12659 8488 12693 8490
rect 12625 8472 12705 8488
rect 12625 8450 12644 8472
rect 12659 8456 12689 8472
rect 12717 8466 12723 8540
rect 12726 8466 12745 8610
rect 12760 8466 12766 8610
rect 12775 8540 12788 8610
rect 12833 8584 12862 8598
rect 12915 8584 12931 8598
rect 12969 8594 12975 8596
rect 12982 8594 13090 8610
rect 13097 8594 13103 8596
rect 13111 8594 13126 8610
rect 13192 8604 13211 8607
rect 12833 8582 12931 8584
rect 12958 8582 13126 8594
rect 13141 8584 13157 8598
rect 13192 8585 13214 8604
rect 13224 8598 13240 8599
rect 13223 8596 13240 8598
rect 13224 8591 13240 8596
rect 13214 8584 13220 8585
rect 13223 8584 13252 8591
rect 13141 8583 13252 8584
rect 13141 8582 13258 8583
rect 12817 8574 12868 8582
rect 12915 8574 12949 8582
rect 12817 8562 12842 8574
rect 12849 8562 12868 8574
rect 12922 8572 12949 8574
rect 12958 8572 13179 8582
rect 13214 8579 13220 8582
rect 12922 8568 13179 8572
rect 12817 8554 12868 8562
rect 12915 8554 13179 8568
rect 13223 8574 13258 8582
rect 12769 8506 12788 8540
rect 12833 8546 12862 8554
rect 12833 8540 12850 8546
rect 12833 8538 12867 8540
rect 12915 8538 12931 8554
rect 12932 8544 13140 8554
rect 13141 8544 13157 8554
rect 13205 8550 13220 8565
rect 13223 8562 13224 8574
rect 13231 8562 13258 8574
rect 13223 8554 13258 8562
rect 13223 8553 13252 8554
rect 12943 8540 13157 8544
rect 12958 8538 13157 8540
rect 13192 8540 13205 8550
rect 13223 8540 13240 8553
rect 13192 8538 13240 8540
rect 12834 8534 12867 8538
rect 12830 8532 12867 8534
rect 12830 8531 12897 8532
rect 12830 8526 12861 8531
rect 12867 8526 12897 8531
rect 12830 8522 12897 8526
rect 12803 8519 12897 8522
rect 12803 8512 12852 8519
rect 12803 8506 12833 8512
rect 12852 8507 12857 8512
rect 12769 8490 12849 8506
rect 12861 8498 12897 8519
rect 12958 8514 13147 8538
rect 13192 8537 13239 8538
rect 13205 8532 13239 8537
rect 12973 8511 13147 8514
rect 12966 8508 13147 8511
rect 13175 8531 13239 8532
rect 12769 8488 12788 8490
rect 12803 8488 12837 8490
rect 12769 8472 12849 8488
rect 12769 8466 12788 8472
rect 12485 8440 12588 8450
rect 12439 8438 12588 8440
rect 12609 8438 12644 8450
rect 12278 8436 12440 8438
rect 12290 8416 12309 8436
rect 12324 8434 12354 8436
rect 12173 8408 12214 8416
rect 12296 8412 12309 8416
rect 12361 8420 12440 8436
rect 12472 8436 12644 8438
rect 12472 8420 12551 8436
rect 12558 8434 12588 8436
rect 12136 8398 12165 8408
rect 12179 8398 12208 8408
rect 12223 8398 12253 8412
rect 12296 8398 12339 8412
rect 12361 8408 12551 8420
rect 12616 8416 12622 8436
rect 12346 8398 12376 8408
rect 12377 8398 12535 8408
rect 12539 8398 12569 8408
rect 12573 8398 12603 8412
rect 12631 8398 12644 8436
rect 12716 8450 12745 8466
rect 12759 8450 12788 8466
rect 12803 8456 12833 8472
rect 12861 8450 12867 8498
rect 12870 8492 12889 8498
rect 12904 8492 12934 8500
rect 12870 8484 12934 8492
rect 12870 8468 12950 8484
rect 12966 8477 13028 8508
rect 13044 8477 13106 8508
rect 13175 8506 13224 8531
rect 13239 8506 13269 8522
rect 13138 8492 13168 8500
rect 13175 8498 13285 8506
rect 13138 8484 13183 8492
rect 12870 8466 12889 8468
rect 12904 8466 12950 8468
rect 12870 8450 12950 8466
rect 12977 8464 13012 8477
rect 13053 8474 13090 8477
rect 13053 8472 13095 8474
rect 12982 8461 13012 8464
rect 12991 8457 12998 8461
rect 12998 8456 12999 8457
rect 12957 8450 12967 8456
rect 12716 8442 12751 8450
rect 12716 8416 12717 8442
rect 12724 8416 12751 8442
rect 12659 8398 12689 8412
rect 12716 8408 12751 8416
rect 12753 8442 12794 8450
rect 12753 8416 12768 8442
rect 12775 8416 12794 8442
rect 12858 8438 12889 8450
rect 12904 8438 13007 8450
rect 13019 8440 13045 8466
rect 13060 8461 13090 8472
rect 13122 8468 13184 8484
rect 13122 8466 13168 8468
rect 13122 8450 13184 8466
rect 13196 8450 13202 8498
rect 13205 8490 13285 8498
rect 13205 8488 13224 8490
rect 13239 8488 13273 8490
rect 13205 8472 13285 8488
rect 13205 8450 13224 8472
rect 13239 8456 13269 8472
rect 13297 8466 13303 8540
rect 13306 8466 13325 8610
rect 13340 8466 13346 8610
rect 13355 8540 13368 8610
rect 13413 8584 13442 8598
rect 13495 8584 13511 8598
rect 13549 8594 13555 8596
rect 13562 8594 13670 8610
rect 13677 8594 13683 8596
rect 13691 8594 13706 8610
rect 13772 8604 13791 8607
rect 13413 8582 13511 8584
rect 13538 8582 13706 8594
rect 13721 8584 13737 8598
rect 13772 8585 13794 8604
rect 13804 8598 13820 8599
rect 13803 8596 13820 8598
rect 13804 8591 13820 8596
rect 13794 8584 13800 8585
rect 13803 8584 13832 8591
rect 13721 8583 13832 8584
rect 13721 8582 13838 8583
rect 13397 8574 13448 8582
rect 13495 8574 13529 8582
rect 13397 8562 13422 8574
rect 13429 8562 13448 8574
rect 13502 8572 13529 8574
rect 13538 8572 13759 8582
rect 13794 8579 13800 8582
rect 13502 8568 13759 8572
rect 13397 8554 13448 8562
rect 13495 8554 13759 8568
rect 13803 8574 13838 8582
rect 13349 8506 13368 8540
rect 13413 8546 13442 8554
rect 13413 8540 13430 8546
rect 13413 8538 13447 8540
rect 13495 8538 13511 8554
rect 13512 8544 13720 8554
rect 13721 8544 13737 8554
rect 13785 8550 13800 8565
rect 13803 8562 13804 8574
rect 13811 8562 13838 8574
rect 13803 8554 13838 8562
rect 13803 8553 13832 8554
rect 13523 8540 13737 8544
rect 13538 8538 13737 8540
rect 13772 8540 13785 8550
rect 13803 8540 13820 8553
rect 13772 8538 13820 8540
rect 13414 8534 13447 8538
rect 13410 8532 13447 8534
rect 13410 8531 13477 8532
rect 13410 8526 13441 8531
rect 13447 8526 13477 8531
rect 13410 8522 13477 8526
rect 13383 8519 13477 8522
rect 13383 8512 13432 8519
rect 13383 8506 13413 8512
rect 13432 8507 13437 8512
rect 13349 8490 13429 8506
rect 13441 8498 13477 8519
rect 13538 8514 13727 8538
rect 13772 8537 13819 8538
rect 13785 8532 13819 8537
rect 13553 8511 13727 8514
rect 13546 8508 13727 8511
rect 13755 8531 13819 8532
rect 13349 8488 13368 8490
rect 13383 8488 13417 8490
rect 13349 8472 13429 8488
rect 13349 8466 13368 8472
rect 13065 8440 13168 8450
rect 13019 8438 13168 8440
rect 13189 8438 13224 8450
rect 12858 8436 13020 8438
rect 12870 8416 12889 8436
rect 12904 8434 12934 8436
rect 12753 8408 12794 8416
rect 12876 8412 12889 8416
rect 12941 8420 13020 8436
rect 13052 8436 13224 8438
rect 13052 8420 13131 8436
rect 13138 8434 13168 8436
rect 12716 8398 12745 8408
rect 12759 8398 12788 8408
rect 12803 8398 12833 8412
rect 12876 8398 12919 8412
rect 12941 8408 13131 8420
rect 13196 8416 13202 8436
rect 12926 8398 12956 8408
rect 12957 8398 13115 8408
rect 13119 8398 13149 8408
rect 13153 8398 13183 8412
rect 13211 8398 13224 8436
rect 13296 8450 13325 8466
rect 13339 8450 13368 8466
rect 13383 8456 13413 8472
rect 13441 8450 13447 8498
rect 13450 8492 13469 8498
rect 13484 8492 13514 8500
rect 13450 8484 13514 8492
rect 13450 8468 13530 8484
rect 13546 8477 13608 8508
rect 13624 8477 13686 8508
rect 13755 8506 13804 8531
rect 13819 8506 13849 8522
rect 13718 8492 13748 8500
rect 13755 8498 13865 8506
rect 13718 8484 13763 8492
rect 13450 8466 13469 8468
rect 13484 8466 13530 8468
rect 13450 8450 13530 8466
rect 13557 8464 13592 8477
rect 13633 8474 13670 8477
rect 13633 8472 13675 8474
rect 13562 8461 13592 8464
rect 13571 8457 13578 8461
rect 13578 8456 13579 8457
rect 13537 8450 13547 8456
rect 13296 8442 13331 8450
rect 13296 8416 13297 8442
rect 13304 8416 13331 8442
rect 13239 8398 13269 8412
rect 13296 8408 13331 8416
rect 13333 8442 13374 8450
rect 13333 8416 13348 8442
rect 13355 8416 13374 8442
rect 13438 8438 13469 8450
rect 13484 8438 13587 8450
rect 13599 8440 13625 8466
rect 13640 8461 13670 8472
rect 13702 8468 13764 8484
rect 13702 8466 13748 8468
rect 13702 8450 13764 8466
rect 13776 8450 13782 8498
rect 13785 8490 13865 8498
rect 13785 8488 13804 8490
rect 13819 8488 13853 8490
rect 13785 8472 13865 8488
rect 13785 8450 13804 8472
rect 13819 8456 13849 8472
rect 13877 8466 13883 8540
rect 13886 8466 13905 8610
rect 13920 8466 13926 8610
rect 13935 8540 13948 8610
rect 13993 8584 14022 8598
rect 14075 8584 14091 8598
rect 14129 8594 14135 8596
rect 14142 8594 14250 8610
rect 14257 8594 14263 8596
rect 14271 8594 14286 8610
rect 14352 8604 14371 8607
rect 13993 8582 14091 8584
rect 14118 8582 14286 8594
rect 14301 8584 14317 8598
rect 14352 8585 14374 8604
rect 14384 8598 14400 8599
rect 14383 8596 14400 8598
rect 14384 8591 14400 8596
rect 14374 8584 14380 8585
rect 14383 8584 14412 8591
rect 14301 8583 14412 8584
rect 14301 8582 14418 8583
rect 13977 8574 14028 8582
rect 14075 8574 14109 8582
rect 13977 8562 14002 8574
rect 14009 8562 14028 8574
rect 14082 8572 14109 8574
rect 14118 8572 14339 8582
rect 14374 8579 14380 8582
rect 14082 8568 14339 8572
rect 13977 8554 14028 8562
rect 14075 8554 14339 8568
rect 14383 8574 14418 8582
rect 13929 8506 13948 8540
rect 13993 8546 14022 8554
rect 13993 8540 14010 8546
rect 13993 8538 14027 8540
rect 14075 8538 14091 8554
rect 14092 8544 14300 8554
rect 14301 8544 14317 8554
rect 14365 8550 14380 8565
rect 14383 8562 14384 8574
rect 14391 8562 14418 8574
rect 14383 8554 14418 8562
rect 14383 8553 14412 8554
rect 14103 8540 14317 8544
rect 14118 8538 14317 8540
rect 14352 8540 14365 8550
rect 14383 8540 14400 8553
rect 14352 8538 14400 8540
rect 13994 8534 14027 8538
rect 13990 8532 14027 8534
rect 13990 8531 14057 8532
rect 13990 8526 14021 8531
rect 14027 8526 14057 8531
rect 13990 8522 14057 8526
rect 13963 8519 14057 8522
rect 13963 8512 14012 8519
rect 13963 8506 13993 8512
rect 14012 8507 14017 8512
rect 13929 8490 14009 8506
rect 14021 8498 14057 8519
rect 14118 8514 14307 8538
rect 14352 8537 14399 8538
rect 14365 8532 14399 8537
rect 14133 8511 14307 8514
rect 14126 8508 14307 8511
rect 14335 8531 14399 8532
rect 13929 8488 13948 8490
rect 13963 8488 13997 8490
rect 13929 8472 14009 8488
rect 13929 8466 13948 8472
rect 13645 8440 13748 8450
rect 13599 8438 13748 8440
rect 13769 8438 13804 8450
rect 13438 8436 13600 8438
rect 13450 8416 13469 8436
rect 13484 8434 13514 8436
rect 13333 8408 13374 8416
rect 13456 8412 13469 8416
rect 13521 8420 13600 8436
rect 13632 8436 13804 8438
rect 13632 8420 13711 8436
rect 13718 8434 13748 8436
rect 13296 8398 13325 8408
rect 13339 8398 13368 8408
rect 13383 8398 13413 8412
rect 13456 8398 13499 8412
rect 13521 8408 13711 8420
rect 13776 8416 13782 8436
rect 13506 8398 13536 8408
rect 13537 8398 13695 8408
rect 13699 8398 13729 8408
rect 13733 8398 13763 8412
rect 13791 8398 13804 8436
rect 13876 8450 13905 8466
rect 13919 8450 13948 8466
rect 13963 8456 13993 8472
rect 14021 8450 14027 8498
rect 14030 8492 14049 8498
rect 14064 8492 14094 8500
rect 14030 8484 14094 8492
rect 14030 8468 14110 8484
rect 14126 8477 14188 8508
rect 14204 8477 14266 8508
rect 14335 8506 14384 8531
rect 14399 8506 14429 8522
rect 14298 8492 14328 8500
rect 14335 8498 14445 8506
rect 14298 8484 14343 8492
rect 14030 8466 14049 8468
rect 14064 8466 14110 8468
rect 14030 8450 14110 8466
rect 14137 8464 14172 8477
rect 14213 8474 14250 8477
rect 14213 8472 14255 8474
rect 14142 8461 14172 8464
rect 14151 8457 14158 8461
rect 14158 8456 14159 8457
rect 14117 8450 14127 8456
rect 13876 8442 13911 8450
rect 13876 8416 13877 8442
rect 13884 8416 13911 8442
rect 13819 8398 13849 8412
rect 13876 8408 13911 8416
rect 13913 8442 13954 8450
rect 13913 8416 13928 8442
rect 13935 8416 13954 8442
rect 14018 8438 14049 8450
rect 14064 8438 14167 8450
rect 14179 8440 14205 8466
rect 14220 8461 14250 8472
rect 14282 8468 14344 8484
rect 14282 8466 14328 8468
rect 14282 8450 14344 8466
rect 14356 8450 14362 8498
rect 14365 8490 14445 8498
rect 14365 8488 14384 8490
rect 14399 8488 14433 8490
rect 14365 8472 14445 8488
rect 14365 8450 14384 8472
rect 14399 8456 14429 8472
rect 14457 8466 14463 8540
rect 14466 8466 14485 8610
rect 14500 8466 14506 8610
rect 14515 8540 14528 8610
rect 14573 8584 14602 8598
rect 14655 8584 14671 8598
rect 14709 8594 14715 8596
rect 14722 8594 14830 8610
rect 14837 8594 14843 8596
rect 14851 8594 14866 8610
rect 14932 8604 14951 8607
rect 14573 8582 14671 8584
rect 14698 8582 14866 8594
rect 14881 8584 14897 8598
rect 14932 8585 14954 8604
rect 14964 8598 14980 8599
rect 14963 8596 14980 8598
rect 14964 8591 14980 8596
rect 14954 8584 14960 8585
rect 14963 8584 14992 8591
rect 14881 8583 14992 8584
rect 14881 8582 14998 8583
rect 14557 8574 14608 8582
rect 14655 8574 14689 8582
rect 14557 8562 14582 8574
rect 14589 8562 14608 8574
rect 14662 8572 14689 8574
rect 14698 8572 14919 8582
rect 14954 8579 14960 8582
rect 14662 8568 14919 8572
rect 14557 8554 14608 8562
rect 14655 8554 14919 8568
rect 14963 8574 14998 8582
rect 14509 8506 14528 8540
rect 14573 8546 14602 8554
rect 14573 8540 14590 8546
rect 14573 8538 14607 8540
rect 14655 8538 14671 8554
rect 14672 8544 14880 8554
rect 14881 8544 14897 8554
rect 14945 8550 14960 8565
rect 14963 8562 14964 8574
rect 14971 8562 14998 8574
rect 14963 8554 14998 8562
rect 14963 8553 14992 8554
rect 14683 8540 14897 8544
rect 14698 8538 14897 8540
rect 14932 8540 14945 8550
rect 14963 8540 14980 8553
rect 14932 8538 14980 8540
rect 14574 8534 14607 8538
rect 14570 8532 14607 8534
rect 14570 8531 14637 8532
rect 14570 8526 14601 8531
rect 14607 8526 14637 8531
rect 14570 8522 14637 8526
rect 14543 8519 14637 8522
rect 14543 8512 14592 8519
rect 14543 8506 14573 8512
rect 14592 8507 14597 8512
rect 14509 8490 14589 8506
rect 14601 8498 14637 8519
rect 14698 8514 14887 8538
rect 14932 8537 14979 8538
rect 14945 8532 14979 8537
rect 14713 8511 14887 8514
rect 14706 8508 14887 8511
rect 14915 8531 14979 8532
rect 14509 8488 14528 8490
rect 14543 8488 14577 8490
rect 14509 8472 14589 8488
rect 14509 8466 14528 8472
rect 14225 8440 14328 8450
rect 14179 8438 14328 8440
rect 14349 8438 14384 8450
rect 14018 8436 14180 8438
rect 14030 8416 14049 8436
rect 14064 8434 14094 8436
rect 13913 8408 13954 8416
rect 14036 8412 14049 8416
rect 14101 8420 14180 8436
rect 14212 8436 14384 8438
rect 14212 8420 14291 8436
rect 14298 8434 14328 8436
rect 13876 8398 13905 8408
rect 13919 8398 13948 8408
rect 13963 8398 13993 8412
rect 14036 8398 14079 8412
rect 14101 8408 14291 8420
rect 14356 8416 14362 8436
rect 14086 8398 14116 8408
rect 14117 8398 14275 8408
rect 14279 8398 14309 8408
rect 14313 8398 14343 8412
rect 14371 8398 14384 8436
rect 14456 8450 14485 8466
rect 14499 8450 14528 8466
rect 14543 8456 14573 8472
rect 14601 8450 14607 8498
rect 14610 8492 14629 8498
rect 14644 8492 14674 8500
rect 14610 8484 14674 8492
rect 14610 8468 14690 8484
rect 14706 8477 14768 8508
rect 14784 8477 14846 8508
rect 14915 8506 14964 8531
rect 14979 8506 15009 8522
rect 14878 8492 14908 8500
rect 14915 8498 15025 8506
rect 14878 8484 14923 8492
rect 14610 8466 14629 8468
rect 14644 8466 14690 8468
rect 14610 8450 14690 8466
rect 14717 8464 14752 8477
rect 14793 8474 14830 8477
rect 14793 8472 14835 8474
rect 14722 8461 14752 8464
rect 14731 8457 14738 8461
rect 14738 8456 14739 8457
rect 14697 8450 14707 8456
rect 14456 8442 14491 8450
rect 14456 8416 14457 8442
rect 14464 8416 14491 8442
rect 14399 8398 14429 8412
rect 14456 8408 14491 8416
rect 14493 8442 14534 8450
rect 14493 8416 14508 8442
rect 14515 8416 14534 8442
rect 14598 8438 14629 8450
rect 14644 8438 14747 8450
rect 14759 8440 14785 8466
rect 14800 8461 14830 8472
rect 14862 8468 14924 8484
rect 14862 8466 14908 8468
rect 14862 8450 14924 8466
rect 14936 8450 14942 8498
rect 14945 8490 15025 8498
rect 14945 8488 14964 8490
rect 14979 8488 15013 8490
rect 14945 8472 15025 8488
rect 14945 8450 14964 8472
rect 14979 8456 15009 8472
rect 15037 8466 15043 8540
rect 15046 8466 15065 8610
rect 15080 8466 15086 8610
rect 15095 8540 15108 8610
rect 15153 8584 15182 8598
rect 15235 8584 15251 8598
rect 15289 8594 15295 8596
rect 15302 8594 15410 8610
rect 15417 8594 15423 8596
rect 15431 8594 15446 8610
rect 15512 8604 15531 8607
rect 15153 8582 15251 8584
rect 15278 8582 15446 8594
rect 15461 8584 15477 8598
rect 15512 8585 15534 8604
rect 15544 8598 15560 8599
rect 15543 8596 15560 8598
rect 15544 8591 15560 8596
rect 15534 8584 15540 8585
rect 15543 8584 15572 8591
rect 15461 8583 15572 8584
rect 15461 8582 15578 8583
rect 15137 8574 15188 8582
rect 15235 8574 15269 8582
rect 15137 8562 15162 8574
rect 15169 8562 15188 8574
rect 15242 8572 15269 8574
rect 15278 8572 15499 8582
rect 15534 8579 15540 8582
rect 15242 8568 15499 8572
rect 15137 8554 15188 8562
rect 15235 8554 15499 8568
rect 15543 8574 15578 8582
rect 15089 8506 15108 8540
rect 15153 8546 15182 8554
rect 15153 8540 15170 8546
rect 15153 8538 15187 8540
rect 15235 8538 15251 8554
rect 15252 8544 15460 8554
rect 15461 8544 15477 8554
rect 15525 8550 15540 8565
rect 15543 8562 15544 8574
rect 15551 8562 15578 8574
rect 15543 8554 15578 8562
rect 15543 8553 15572 8554
rect 15263 8540 15477 8544
rect 15278 8538 15477 8540
rect 15512 8540 15525 8550
rect 15543 8540 15560 8553
rect 15512 8538 15560 8540
rect 15154 8534 15187 8538
rect 15150 8532 15187 8534
rect 15150 8531 15217 8532
rect 15150 8526 15181 8531
rect 15187 8526 15217 8531
rect 15150 8522 15217 8526
rect 15123 8519 15217 8522
rect 15123 8512 15172 8519
rect 15123 8506 15153 8512
rect 15172 8507 15177 8512
rect 15089 8490 15169 8506
rect 15181 8498 15217 8519
rect 15278 8514 15467 8538
rect 15512 8537 15559 8538
rect 15525 8532 15559 8537
rect 15293 8511 15467 8514
rect 15286 8508 15467 8511
rect 15495 8531 15559 8532
rect 15089 8488 15108 8490
rect 15123 8488 15157 8490
rect 15089 8472 15169 8488
rect 15089 8466 15108 8472
rect 14805 8440 14908 8450
rect 14759 8438 14908 8440
rect 14929 8438 14964 8450
rect 14598 8436 14760 8438
rect 14610 8416 14629 8436
rect 14644 8434 14674 8436
rect 14493 8408 14534 8416
rect 14616 8412 14629 8416
rect 14681 8420 14760 8436
rect 14792 8436 14964 8438
rect 14792 8420 14871 8436
rect 14878 8434 14908 8436
rect 14456 8398 14485 8408
rect 14499 8398 14528 8408
rect 14543 8398 14573 8412
rect 14616 8398 14659 8412
rect 14681 8408 14871 8420
rect 14936 8416 14942 8436
rect 14666 8398 14696 8408
rect 14697 8398 14855 8408
rect 14859 8398 14889 8408
rect 14893 8398 14923 8412
rect 14951 8398 14964 8436
rect 15036 8450 15065 8466
rect 15079 8450 15108 8466
rect 15123 8456 15153 8472
rect 15181 8450 15187 8498
rect 15190 8492 15209 8498
rect 15224 8492 15254 8500
rect 15190 8484 15254 8492
rect 15190 8468 15270 8484
rect 15286 8477 15348 8508
rect 15364 8477 15426 8508
rect 15495 8506 15544 8531
rect 15559 8506 15589 8522
rect 15458 8492 15488 8500
rect 15495 8498 15605 8506
rect 15458 8484 15503 8492
rect 15190 8466 15209 8468
rect 15224 8466 15270 8468
rect 15190 8450 15270 8466
rect 15297 8464 15332 8477
rect 15373 8474 15410 8477
rect 15373 8472 15415 8474
rect 15302 8461 15332 8464
rect 15311 8457 15318 8461
rect 15318 8456 15319 8457
rect 15277 8450 15287 8456
rect 15036 8442 15071 8450
rect 15036 8416 15037 8442
rect 15044 8416 15071 8442
rect 14979 8398 15009 8412
rect 15036 8408 15071 8416
rect 15073 8442 15114 8450
rect 15073 8416 15088 8442
rect 15095 8416 15114 8442
rect 15178 8438 15209 8450
rect 15224 8438 15327 8450
rect 15339 8440 15365 8466
rect 15380 8461 15410 8472
rect 15442 8468 15504 8484
rect 15442 8466 15488 8468
rect 15442 8450 15504 8466
rect 15516 8450 15522 8498
rect 15525 8490 15605 8498
rect 15525 8488 15544 8490
rect 15559 8488 15593 8490
rect 15525 8472 15605 8488
rect 15525 8450 15544 8472
rect 15559 8456 15589 8472
rect 15617 8466 15623 8540
rect 15626 8466 15645 8610
rect 15660 8466 15666 8610
rect 15675 8540 15688 8610
rect 15733 8584 15762 8598
rect 15815 8584 15831 8598
rect 15869 8594 15875 8596
rect 15882 8594 15990 8610
rect 15997 8594 16003 8596
rect 16011 8594 16026 8610
rect 16092 8604 16111 8607
rect 15733 8582 15831 8584
rect 15858 8582 16026 8594
rect 16041 8584 16057 8598
rect 16092 8585 16114 8604
rect 16124 8598 16140 8599
rect 16123 8596 16140 8598
rect 16124 8591 16140 8596
rect 16114 8584 16120 8585
rect 16123 8584 16152 8591
rect 16041 8583 16152 8584
rect 16041 8582 16158 8583
rect 15717 8574 15768 8582
rect 15815 8574 15849 8582
rect 15717 8562 15742 8574
rect 15749 8562 15768 8574
rect 15822 8572 15849 8574
rect 15858 8572 16079 8582
rect 16114 8579 16120 8582
rect 15822 8568 16079 8572
rect 15717 8554 15768 8562
rect 15815 8554 16079 8568
rect 16123 8574 16158 8582
rect 15669 8506 15688 8540
rect 15733 8546 15762 8554
rect 15733 8540 15750 8546
rect 15733 8538 15767 8540
rect 15815 8538 15831 8554
rect 15832 8544 16040 8554
rect 16041 8544 16057 8554
rect 16105 8550 16120 8565
rect 16123 8562 16124 8574
rect 16131 8562 16158 8574
rect 16123 8554 16158 8562
rect 16123 8553 16152 8554
rect 15843 8540 16057 8544
rect 15858 8538 16057 8540
rect 16092 8540 16105 8550
rect 16123 8540 16140 8553
rect 16092 8538 16140 8540
rect 15734 8534 15767 8538
rect 15730 8532 15767 8534
rect 15730 8531 15797 8532
rect 15730 8526 15761 8531
rect 15767 8526 15797 8531
rect 15730 8522 15797 8526
rect 15703 8519 15797 8522
rect 15703 8512 15752 8519
rect 15703 8506 15733 8512
rect 15752 8507 15757 8512
rect 15669 8490 15749 8506
rect 15761 8498 15797 8519
rect 15858 8514 16047 8538
rect 16092 8537 16139 8538
rect 16105 8532 16139 8537
rect 15873 8511 16047 8514
rect 15866 8508 16047 8511
rect 16075 8531 16139 8532
rect 15669 8488 15688 8490
rect 15703 8488 15737 8490
rect 15669 8472 15749 8488
rect 15669 8466 15688 8472
rect 15385 8440 15488 8450
rect 15339 8438 15488 8440
rect 15509 8438 15544 8450
rect 15178 8436 15340 8438
rect 15190 8416 15209 8436
rect 15224 8434 15254 8436
rect 15073 8408 15114 8416
rect 15196 8412 15209 8416
rect 15261 8420 15340 8436
rect 15372 8436 15544 8438
rect 15372 8420 15451 8436
rect 15458 8434 15488 8436
rect 15036 8398 15065 8408
rect 15079 8398 15108 8408
rect 15123 8398 15153 8412
rect 15196 8398 15239 8412
rect 15261 8408 15451 8420
rect 15516 8416 15522 8436
rect 15246 8398 15276 8408
rect 15277 8398 15435 8408
rect 15439 8398 15469 8408
rect 15473 8398 15503 8412
rect 15531 8398 15544 8436
rect 15616 8450 15645 8466
rect 15659 8450 15688 8466
rect 15703 8456 15733 8472
rect 15761 8450 15767 8498
rect 15770 8492 15789 8498
rect 15804 8492 15834 8500
rect 15770 8484 15834 8492
rect 15770 8468 15850 8484
rect 15866 8477 15928 8508
rect 15944 8477 16006 8508
rect 16075 8506 16124 8531
rect 16139 8506 16169 8522
rect 16038 8492 16068 8500
rect 16075 8498 16185 8506
rect 16038 8484 16083 8492
rect 15770 8466 15789 8468
rect 15804 8466 15850 8468
rect 15770 8450 15850 8466
rect 15877 8464 15912 8477
rect 15953 8474 15990 8477
rect 15953 8472 15995 8474
rect 15882 8461 15912 8464
rect 15891 8457 15898 8461
rect 15898 8456 15899 8457
rect 15857 8450 15867 8456
rect 15616 8442 15651 8450
rect 15616 8416 15617 8442
rect 15624 8416 15651 8442
rect 15559 8398 15589 8412
rect 15616 8408 15651 8416
rect 15653 8442 15694 8450
rect 15653 8416 15668 8442
rect 15675 8416 15694 8442
rect 15758 8438 15789 8450
rect 15804 8438 15907 8450
rect 15919 8440 15945 8466
rect 15960 8461 15990 8472
rect 16022 8468 16084 8484
rect 16022 8466 16068 8468
rect 16022 8450 16084 8466
rect 16096 8450 16102 8498
rect 16105 8490 16185 8498
rect 16105 8488 16124 8490
rect 16139 8488 16173 8490
rect 16105 8472 16185 8488
rect 16105 8450 16124 8472
rect 16139 8456 16169 8472
rect 16197 8466 16203 8540
rect 16206 8466 16225 8610
rect 16240 8466 16246 8610
rect 16255 8540 16268 8610
rect 16313 8584 16342 8598
rect 16395 8584 16411 8598
rect 16449 8594 16455 8596
rect 16462 8594 16570 8610
rect 16577 8594 16583 8596
rect 16591 8594 16606 8610
rect 16672 8604 16691 8607
rect 16313 8582 16411 8584
rect 16438 8582 16606 8594
rect 16621 8584 16637 8598
rect 16672 8585 16694 8604
rect 16704 8598 16720 8599
rect 16703 8596 16720 8598
rect 16704 8591 16720 8596
rect 16694 8584 16700 8585
rect 16703 8584 16732 8591
rect 16621 8583 16732 8584
rect 16621 8582 16738 8583
rect 16297 8574 16348 8582
rect 16395 8574 16429 8582
rect 16297 8562 16322 8574
rect 16329 8562 16348 8574
rect 16402 8572 16429 8574
rect 16438 8572 16659 8582
rect 16694 8579 16700 8582
rect 16402 8568 16659 8572
rect 16297 8554 16348 8562
rect 16395 8554 16659 8568
rect 16703 8574 16738 8582
rect 16249 8506 16268 8540
rect 16313 8546 16342 8554
rect 16313 8540 16330 8546
rect 16313 8538 16347 8540
rect 16395 8538 16411 8554
rect 16412 8544 16620 8554
rect 16621 8544 16637 8554
rect 16685 8550 16700 8565
rect 16703 8562 16704 8574
rect 16711 8562 16738 8574
rect 16703 8554 16738 8562
rect 16703 8553 16732 8554
rect 16423 8540 16637 8544
rect 16438 8538 16637 8540
rect 16672 8540 16685 8550
rect 16703 8540 16720 8553
rect 16672 8538 16720 8540
rect 16314 8534 16347 8538
rect 16310 8532 16347 8534
rect 16310 8531 16377 8532
rect 16310 8526 16341 8531
rect 16347 8526 16377 8531
rect 16310 8522 16377 8526
rect 16283 8519 16377 8522
rect 16283 8512 16332 8519
rect 16283 8506 16313 8512
rect 16332 8507 16337 8512
rect 16249 8490 16329 8506
rect 16341 8498 16377 8519
rect 16438 8514 16627 8538
rect 16672 8537 16719 8538
rect 16685 8532 16719 8537
rect 16453 8511 16627 8514
rect 16446 8508 16627 8511
rect 16655 8531 16719 8532
rect 16249 8488 16268 8490
rect 16283 8488 16317 8490
rect 16249 8472 16329 8488
rect 16249 8466 16268 8472
rect 15965 8440 16068 8450
rect 15919 8438 16068 8440
rect 16089 8438 16124 8450
rect 15758 8436 15920 8438
rect 15770 8416 15789 8436
rect 15804 8434 15834 8436
rect 15653 8408 15694 8416
rect 15776 8412 15789 8416
rect 15841 8420 15920 8436
rect 15952 8436 16124 8438
rect 15952 8420 16031 8436
rect 16038 8434 16068 8436
rect 15616 8398 15645 8408
rect 15659 8398 15688 8408
rect 15703 8398 15733 8412
rect 15776 8398 15819 8412
rect 15841 8408 16031 8420
rect 16096 8416 16102 8436
rect 15826 8398 15856 8408
rect 15857 8398 16015 8408
rect 16019 8398 16049 8408
rect 16053 8398 16083 8412
rect 16111 8398 16124 8436
rect 16196 8450 16225 8466
rect 16239 8450 16268 8466
rect 16283 8456 16313 8472
rect 16341 8450 16347 8498
rect 16350 8492 16369 8498
rect 16384 8492 16414 8500
rect 16350 8484 16414 8492
rect 16350 8468 16430 8484
rect 16446 8477 16508 8508
rect 16524 8477 16586 8508
rect 16655 8506 16704 8531
rect 16719 8506 16749 8522
rect 16618 8492 16648 8500
rect 16655 8498 16765 8506
rect 16618 8484 16663 8492
rect 16350 8466 16369 8468
rect 16384 8466 16430 8468
rect 16350 8450 16430 8466
rect 16457 8464 16492 8477
rect 16533 8474 16570 8477
rect 16533 8472 16575 8474
rect 16462 8461 16492 8464
rect 16471 8457 16478 8461
rect 16478 8456 16479 8457
rect 16437 8450 16447 8456
rect 16196 8442 16231 8450
rect 16196 8416 16197 8442
rect 16204 8416 16231 8442
rect 16139 8398 16169 8412
rect 16196 8408 16231 8416
rect 16233 8442 16274 8450
rect 16233 8416 16248 8442
rect 16255 8416 16274 8442
rect 16338 8438 16369 8450
rect 16384 8438 16487 8450
rect 16499 8440 16525 8466
rect 16540 8461 16570 8472
rect 16602 8468 16664 8484
rect 16602 8466 16648 8468
rect 16602 8450 16664 8466
rect 16676 8450 16682 8498
rect 16685 8490 16765 8498
rect 16685 8488 16704 8490
rect 16719 8488 16753 8490
rect 16685 8472 16765 8488
rect 16685 8450 16704 8472
rect 16719 8456 16749 8472
rect 16777 8466 16783 8540
rect 16786 8466 16805 8610
rect 16820 8466 16826 8610
rect 16835 8540 16848 8610
rect 16893 8584 16922 8598
rect 16975 8584 16991 8598
rect 17029 8594 17035 8596
rect 17042 8594 17150 8610
rect 17157 8594 17163 8596
rect 17171 8594 17186 8610
rect 17252 8604 17271 8607
rect 16893 8582 16991 8584
rect 17018 8582 17186 8594
rect 17201 8584 17217 8598
rect 17252 8585 17274 8604
rect 17284 8598 17300 8599
rect 17283 8596 17300 8598
rect 17284 8591 17300 8596
rect 17274 8584 17280 8585
rect 17283 8584 17312 8591
rect 17201 8583 17312 8584
rect 17201 8582 17318 8583
rect 16877 8574 16928 8582
rect 16975 8574 17009 8582
rect 16877 8562 16902 8574
rect 16909 8562 16928 8574
rect 16982 8572 17009 8574
rect 17018 8572 17239 8582
rect 17274 8579 17280 8582
rect 16982 8568 17239 8572
rect 16877 8554 16928 8562
rect 16975 8554 17239 8568
rect 17283 8574 17318 8582
rect 16829 8506 16848 8540
rect 16893 8546 16922 8554
rect 16893 8540 16910 8546
rect 16893 8538 16927 8540
rect 16975 8538 16991 8554
rect 16992 8544 17200 8554
rect 17201 8544 17217 8554
rect 17265 8550 17280 8565
rect 17283 8562 17284 8574
rect 17291 8562 17318 8574
rect 17283 8554 17318 8562
rect 17283 8553 17312 8554
rect 17003 8540 17217 8544
rect 17018 8538 17217 8540
rect 17252 8540 17265 8550
rect 17283 8540 17300 8553
rect 17252 8538 17300 8540
rect 16894 8534 16927 8538
rect 16890 8532 16927 8534
rect 16890 8531 16957 8532
rect 16890 8526 16921 8531
rect 16927 8526 16957 8531
rect 16890 8522 16957 8526
rect 16863 8519 16957 8522
rect 16863 8512 16912 8519
rect 16863 8506 16893 8512
rect 16912 8507 16917 8512
rect 16829 8490 16909 8506
rect 16921 8498 16957 8519
rect 17018 8514 17207 8538
rect 17252 8537 17299 8538
rect 17265 8532 17299 8537
rect 17033 8511 17207 8514
rect 17026 8508 17207 8511
rect 17235 8531 17299 8532
rect 16829 8488 16848 8490
rect 16863 8488 16897 8490
rect 16829 8472 16909 8488
rect 16829 8466 16848 8472
rect 16545 8440 16648 8450
rect 16499 8438 16648 8440
rect 16669 8438 16704 8450
rect 16338 8436 16500 8438
rect 16350 8416 16369 8436
rect 16384 8434 16414 8436
rect 16233 8408 16274 8416
rect 16356 8412 16369 8416
rect 16421 8420 16500 8436
rect 16532 8436 16704 8438
rect 16532 8420 16611 8436
rect 16618 8434 16648 8436
rect 16196 8398 16225 8408
rect 16239 8398 16268 8408
rect 16283 8398 16313 8412
rect 16356 8398 16399 8412
rect 16421 8408 16611 8420
rect 16676 8416 16682 8436
rect 16406 8398 16436 8408
rect 16437 8398 16595 8408
rect 16599 8398 16629 8408
rect 16633 8398 16663 8412
rect 16691 8398 16704 8436
rect 16776 8450 16805 8466
rect 16819 8450 16848 8466
rect 16863 8456 16893 8472
rect 16921 8450 16927 8498
rect 16930 8492 16949 8498
rect 16964 8492 16994 8500
rect 16930 8484 16994 8492
rect 16930 8468 17010 8484
rect 17026 8477 17088 8508
rect 17104 8477 17166 8508
rect 17235 8506 17284 8531
rect 17299 8506 17329 8522
rect 17198 8492 17228 8500
rect 17235 8498 17345 8506
rect 17198 8484 17243 8492
rect 16930 8466 16949 8468
rect 16964 8466 17010 8468
rect 16930 8450 17010 8466
rect 17037 8464 17072 8477
rect 17113 8474 17150 8477
rect 17113 8472 17155 8474
rect 17042 8461 17072 8464
rect 17051 8457 17058 8461
rect 17058 8456 17059 8457
rect 17017 8450 17027 8456
rect 16776 8442 16811 8450
rect 16776 8416 16777 8442
rect 16784 8416 16811 8442
rect 16719 8398 16749 8412
rect 16776 8408 16811 8416
rect 16813 8442 16854 8450
rect 16813 8416 16828 8442
rect 16835 8416 16854 8442
rect 16918 8438 16949 8450
rect 16964 8438 17067 8450
rect 17079 8440 17105 8466
rect 17120 8461 17150 8472
rect 17182 8468 17244 8484
rect 17182 8466 17228 8468
rect 17182 8450 17244 8466
rect 17256 8450 17262 8498
rect 17265 8490 17345 8498
rect 17265 8488 17284 8490
rect 17299 8488 17333 8490
rect 17265 8472 17345 8488
rect 17265 8450 17284 8472
rect 17299 8456 17329 8472
rect 17357 8466 17363 8540
rect 17366 8466 17385 8610
rect 17400 8466 17406 8610
rect 17415 8540 17428 8610
rect 17473 8584 17502 8598
rect 17555 8584 17571 8598
rect 17609 8594 17615 8596
rect 17622 8594 17730 8610
rect 17737 8594 17743 8596
rect 17751 8594 17766 8610
rect 17832 8604 17851 8607
rect 17473 8582 17571 8584
rect 17598 8582 17766 8594
rect 17781 8584 17797 8598
rect 17832 8585 17854 8604
rect 17864 8598 17880 8599
rect 17863 8596 17880 8598
rect 17864 8591 17880 8596
rect 17854 8584 17860 8585
rect 17863 8584 17892 8591
rect 17781 8583 17892 8584
rect 17781 8582 17898 8583
rect 17457 8574 17508 8582
rect 17555 8574 17589 8582
rect 17457 8562 17482 8574
rect 17489 8562 17508 8574
rect 17562 8572 17589 8574
rect 17598 8572 17819 8582
rect 17854 8579 17860 8582
rect 17562 8568 17819 8572
rect 17457 8554 17508 8562
rect 17555 8554 17819 8568
rect 17863 8574 17898 8582
rect 17409 8506 17428 8540
rect 17473 8546 17502 8554
rect 17473 8540 17490 8546
rect 17473 8538 17507 8540
rect 17555 8538 17571 8554
rect 17572 8544 17780 8554
rect 17781 8544 17797 8554
rect 17845 8550 17860 8565
rect 17863 8562 17864 8574
rect 17871 8562 17898 8574
rect 17863 8554 17898 8562
rect 17863 8553 17892 8554
rect 17583 8540 17797 8544
rect 17598 8538 17797 8540
rect 17832 8540 17845 8550
rect 17863 8540 17880 8553
rect 17832 8538 17880 8540
rect 17474 8534 17507 8538
rect 17470 8532 17507 8534
rect 17470 8531 17537 8532
rect 17470 8526 17501 8531
rect 17507 8526 17537 8531
rect 17470 8522 17537 8526
rect 17443 8519 17537 8522
rect 17443 8512 17492 8519
rect 17443 8506 17473 8512
rect 17492 8507 17497 8512
rect 17409 8490 17489 8506
rect 17501 8498 17537 8519
rect 17598 8514 17787 8538
rect 17832 8537 17879 8538
rect 17845 8532 17879 8537
rect 17613 8511 17787 8514
rect 17606 8508 17787 8511
rect 17815 8531 17879 8532
rect 17409 8488 17428 8490
rect 17443 8488 17477 8490
rect 17409 8472 17489 8488
rect 17409 8466 17428 8472
rect 17125 8440 17228 8450
rect 17079 8438 17228 8440
rect 17249 8438 17284 8450
rect 16918 8436 17080 8438
rect 16930 8416 16949 8436
rect 16964 8434 16994 8436
rect 16813 8408 16854 8416
rect 16936 8412 16949 8416
rect 17001 8420 17080 8436
rect 17112 8436 17284 8438
rect 17112 8420 17191 8436
rect 17198 8434 17228 8436
rect 16776 8398 16805 8408
rect 16819 8398 16848 8408
rect 16863 8398 16893 8412
rect 16936 8398 16979 8412
rect 17001 8408 17191 8420
rect 17256 8416 17262 8436
rect 16986 8398 17016 8408
rect 17017 8398 17175 8408
rect 17179 8398 17209 8408
rect 17213 8398 17243 8412
rect 17271 8398 17284 8436
rect 17356 8450 17385 8466
rect 17399 8450 17428 8466
rect 17443 8456 17473 8472
rect 17501 8450 17507 8498
rect 17510 8492 17529 8498
rect 17544 8492 17574 8500
rect 17510 8484 17574 8492
rect 17510 8468 17590 8484
rect 17606 8477 17668 8508
rect 17684 8477 17746 8508
rect 17815 8506 17864 8531
rect 17879 8506 17909 8522
rect 17778 8492 17808 8500
rect 17815 8498 17925 8506
rect 17778 8484 17823 8492
rect 17510 8466 17529 8468
rect 17544 8466 17590 8468
rect 17510 8450 17590 8466
rect 17617 8464 17652 8477
rect 17693 8474 17730 8477
rect 17693 8472 17735 8474
rect 17622 8461 17652 8464
rect 17631 8457 17638 8461
rect 17638 8456 17639 8457
rect 17597 8450 17607 8456
rect 17356 8442 17391 8450
rect 17356 8416 17357 8442
rect 17364 8416 17391 8442
rect 17299 8398 17329 8412
rect 17356 8408 17391 8416
rect 17393 8442 17434 8450
rect 17393 8416 17408 8442
rect 17415 8416 17434 8442
rect 17498 8438 17529 8450
rect 17544 8438 17647 8450
rect 17659 8440 17685 8466
rect 17700 8461 17730 8472
rect 17762 8468 17824 8484
rect 17762 8466 17808 8468
rect 17762 8450 17824 8466
rect 17836 8450 17842 8498
rect 17845 8490 17925 8498
rect 17845 8488 17864 8490
rect 17879 8488 17913 8490
rect 17845 8472 17925 8488
rect 17845 8450 17864 8472
rect 17879 8456 17909 8472
rect 17937 8466 17943 8540
rect 17946 8466 17965 8610
rect 17980 8466 17986 8610
rect 17995 8540 18008 8610
rect 18053 8584 18082 8598
rect 18135 8584 18151 8598
rect 18189 8594 18195 8596
rect 18202 8594 18310 8610
rect 18317 8594 18323 8596
rect 18331 8594 18346 8610
rect 18412 8604 18431 8607
rect 18053 8582 18151 8584
rect 18178 8582 18346 8594
rect 18361 8584 18377 8598
rect 18412 8585 18434 8604
rect 18444 8598 18460 8599
rect 18443 8596 18460 8598
rect 18444 8591 18460 8596
rect 18434 8584 18440 8585
rect 18443 8584 18472 8591
rect 18361 8583 18472 8584
rect 18361 8582 18478 8583
rect 18037 8574 18088 8582
rect 18135 8574 18169 8582
rect 18037 8562 18062 8574
rect 18069 8562 18088 8574
rect 18142 8572 18169 8574
rect 18178 8572 18399 8582
rect 18434 8579 18440 8582
rect 18142 8568 18399 8572
rect 18037 8554 18088 8562
rect 18135 8554 18399 8568
rect 18443 8574 18478 8582
rect 17989 8506 18008 8540
rect 18053 8546 18082 8554
rect 18053 8540 18070 8546
rect 18053 8538 18087 8540
rect 18135 8538 18151 8554
rect 18152 8544 18360 8554
rect 18361 8544 18377 8554
rect 18425 8550 18440 8565
rect 18443 8562 18444 8574
rect 18451 8562 18478 8574
rect 18443 8554 18478 8562
rect 18443 8553 18472 8554
rect 18163 8540 18377 8544
rect 18178 8538 18377 8540
rect 18412 8540 18425 8550
rect 18443 8540 18460 8553
rect 18412 8538 18460 8540
rect 18054 8534 18087 8538
rect 18050 8532 18087 8534
rect 18050 8531 18117 8532
rect 18050 8526 18081 8531
rect 18087 8526 18117 8531
rect 18050 8522 18117 8526
rect 18023 8519 18117 8522
rect 18023 8512 18072 8519
rect 18023 8506 18053 8512
rect 18072 8507 18077 8512
rect 17989 8490 18069 8506
rect 18081 8498 18117 8519
rect 18178 8514 18367 8538
rect 18412 8537 18459 8538
rect 18425 8532 18459 8537
rect 18193 8511 18367 8514
rect 18186 8508 18367 8511
rect 18395 8531 18459 8532
rect 17989 8488 18008 8490
rect 18023 8488 18057 8490
rect 17989 8472 18069 8488
rect 17989 8466 18008 8472
rect 17705 8440 17808 8450
rect 17659 8438 17808 8440
rect 17829 8438 17864 8450
rect 17498 8436 17660 8438
rect 17510 8416 17529 8436
rect 17544 8434 17574 8436
rect 17393 8408 17434 8416
rect 17516 8412 17529 8416
rect 17581 8420 17660 8436
rect 17692 8436 17864 8438
rect 17692 8420 17771 8436
rect 17778 8434 17808 8436
rect 17356 8398 17385 8408
rect 17399 8398 17428 8408
rect 17443 8398 17473 8412
rect 17516 8398 17559 8412
rect 17581 8408 17771 8420
rect 17836 8416 17842 8436
rect 17566 8398 17596 8408
rect 17597 8398 17755 8408
rect 17759 8398 17789 8408
rect 17793 8398 17823 8412
rect 17851 8398 17864 8436
rect 17936 8450 17965 8466
rect 17979 8450 18008 8466
rect 18023 8456 18053 8472
rect 18081 8450 18087 8498
rect 18090 8492 18109 8498
rect 18124 8492 18154 8500
rect 18090 8484 18154 8492
rect 18090 8468 18170 8484
rect 18186 8477 18248 8508
rect 18264 8477 18326 8508
rect 18395 8506 18444 8531
rect 18459 8506 18489 8522
rect 18358 8492 18388 8500
rect 18395 8498 18505 8506
rect 18358 8484 18403 8492
rect 18090 8466 18109 8468
rect 18124 8466 18170 8468
rect 18090 8450 18170 8466
rect 18197 8464 18232 8477
rect 18273 8474 18310 8477
rect 18273 8472 18315 8474
rect 18202 8461 18232 8464
rect 18211 8457 18218 8461
rect 18218 8456 18219 8457
rect 18177 8450 18187 8456
rect 17936 8442 17971 8450
rect 17936 8416 17937 8442
rect 17944 8416 17971 8442
rect 17879 8398 17909 8412
rect 17936 8408 17971 8416
rect 17973 8442 18014 8450
rect 17973 8416 17988 8442
rect 17995 8416 18014 8442
rect 18078 8438 18109 8450
rect 18124 8438 18227 8450
rect 18239 8440 18265 8466
rect 18280 8461 18310 8472
rect 18342 8468 18404 8484
rect 18342 8466 18388 8468
rect 18342 8450 18404 8466
rect 18416 8450 18422 8498
rect 18425 8490 18505 8498
rect 18425 8488 18444 8490
rect 18459 8488 18493 8490
rect 18425 8472 18505 8488
rect 18425 8450 18444 8472
rect 18459 8456 18489 8472
rect 18517 8466 18523 8540
rect 18532 8466 18545 8610
rect 18285 8440 18388 8450
rect 18239 8438 18388 8440
rect 18409 8438 18444 8450
rect 18078 8436 18240 8438
rect 18090 8416 18109 8436
rect 18124 8434 18154 8436
rect 17973 8408 18014 8416
rect 18096 8412 18109 8416
rect 18161 8420 18240 8436
rect 18272 8436 18444 8438
rect 18272 8420 18351 8436
rect 18358 8434 18388 8436
rect 17936 8398 17965 8408
rect 17979 8398 18008 8408
rect 18023 8398 18053 8412
rect 18096 8398 18139 8412
rect 18161 8408 18351 8420
rect 18416 8416 18422 8436
rect 18146 8398 18176 8408
rect 18177 8398 18335 8408
rect 18339 8398 18369 8408
rect 18373 8398 18403 8412
rect 18431 8398 18444 8436
rect 18516 8450 18545 8466
rect 18516 8442 18551 8450
rect 18516 8416 18517 8442
rect 18524 8416 18551 8442
rect 18459 8398 18489 8412
rect 18516 8408 18551 8416
rect 18516 8398 18545 8408
rect -1 8392 18545 8398
rect 0 8384 18545 8392
rect 15 8354 28 8384
rect 43 8370 73 8384
rect 116 8370 159 8384
rect 166 8370 386 8384
rect 393 8370 423 8384
rect 83 8356 98 8368
rect 117 8356 130 8370
rect 198 8366 351 8370
rect 80 8354 102 8356
rect 180 8354 372 8366
rect 451 8354 464 8384
rect 479 8370 509 8384
rect 546 8354 565 8384
rect 580 8354 586 8384
rect 595 8354 608 8384
rect 623 8370 653 8384
rect 696 8370 739 8384
rect 746 8370 966 8384
rect 973 8370 1003 8384
rect 663 8356 678 8368
rect 697 8356 710 8370
rect 778 8366 931 8370
rect 660 8354 682 8356
rect 760 8354 952 8366
rect 1031 8354 1044 8384
rect 1059 8370 1089 8384
rect 1126 8354 1145 8384
rect 1160 8354 1166 8384
rect 1175 8354 1188 8384
rect 1203 8370 1233 8384
rect 1276 8370 1319 8384
rect 1326 8370 1546 8384
rect 1553 8370 1583 8384
rect 1243 8356 1258 8368
rect 1277 8356 1290 8370
rect 1358 8366 1511 8370
rect 1240 8354 1262 8356
rect 1340 8354 1532 8366
rect 1611 8354 1624 8384
rect 1639 8370 1669 8384
rect 1706 8354 1725 8384
rect 1740 8354 1746 8384
rect 1755 8354 1768 8384
rect 1783 8370 1813 8384
rect 1856 8370 1899 8384
rect 1906 8370 2126 8384
rect 2133 8370 2163 8384
rect 1823 8356 1838 8368
rect 1857 8356 1870 8370
rect 1938 8366 2091 8370
rect 1820 8354 1842 8356
rect 1920 8354 2112 8366
rect 2191 8354 2204 8384
rect 2219 8370 2249 8384
rect 2286 8354 2305 8384
rect 2320 8354 2326 8384
rect 2335 8354 2348 8384
rect 2363 8370 2393 8384
rect 2436 8370 2479 8384
rect 2486 8370 2706 8384
rect 2713 8370 2743 8384
rect 2403 8356 2418 8368
rect 2437 8356 2450 8370
rect 2518 8366 2671 8370
rect 2400 8354 2422 8356
rect 2500 8354 2692 8366
rect 2771 8354 2784 8384
rect 2799 8370 2829 8384
rect 2866 8354 2885 8384
rect 2900 8354 2906 8384
rect 2915 8354 2928 8384
rect 2943 8370 2973 8384
rect 3016 8370 3059 8384
rect 3066 8370 3286 8384
rect 3293 8370 3323 8384
rect 2983 8356 2998 8368
rect 3017 8356 3030 8370
rect 3098 8366 3251 8370
rect 2980 8354 3002 8356
rect 3080 8354 3272 8366
rect 3351 8354 3364 8384
rect 3379 8370 3409 8384
rect 3446 8354 3465 8384
rect 3480 8354 3486 8384
rect 3495 8354 3508 8384
rect 3523 8370 3553 8384
rect 3596 8370 3639 8384
rect 3646 8370 3866 8384
rect 3873 8370 3903 8384
rect 3563 8356 3578 8368
rect 3597 8356 3610 8370
rect 3678 8366 3831 8370
rect 3560 8354 3582 8356
rect 3660 8354 3852 8366
rect 3931 8354 3944 8384
rect 3959 8370 3989 8384
rect 4026 8354 4045 8384
rect 4060 8354 4066 8384
rect 4075 8354 4088 8384
rect 4103 8370 4133 8384
rect 4176 8370 4219 8384
rect 4226 8370 4446 8384
rect 4453 8370 4483 8384
rect 4143 8356 4158 8368
rect 4177 8356 4190 8370
rect 4258 8366 4411 8370
rect 4140 8354 4162 8356
rect 4240 8354 4432 8366
rect 4511 8354 4524 8384
rect 4539 8370 4569 8384
rect 4606 8354 4625 8384
rect 4640 8354 4646 8384
rect 4655 8354 4668 8384
rect 4683 8370 4713 8384
rect 4756 8370 4799 8384
rect 4806 8370 5026 8384
rect 5033 8370 5063 8384
rect 4723 8356 4738 8368
rect 4757 8356 4770 8370
rect 4838 8366 4991 8370
rect 4720 8354 4742 8356
rect 4820 8354 5012 8366
rect 5091 8354 5104 8384
rect 5119 8370 5149 8384
rect 5186 8354 5205 8384
rect 5220 8354 5226 8384
rect 5235 8354 5248 8384
rect 5263 8370 5293 8384
rect 5336 8370 5379 8384
rect 5386 8370 5606 8384
rect 5613 8370 5643 8384
rect 5303 8356 5318 8368
rect 5337 8356 5350 8370
rect 5418 8366 5571 8370
rect 5300 8354 5322 8356
rect 5400 8354 5592 8366
rect 5671 8354 5684 8384
rect 5699 8370 5729 8384
rect 5766 8354 5785 8384
rect 5800 8354 5806 8384
rect 5815 8354 5828 8384
rect 5843 8370 5873 8384
rect 5916 8370 5959 8384
rect 5966 8370 6186 8384
rect 6193 8370 6223 8384
rect 5883 8356 5898 8368
rect 5917 8356 5930 8370
rect 5998 8366 6151 8370
rect 5880 8354 5902 8356
rect 5980 8354 6172 8366
rect 6251 8354 6264 8384
rect 6279 8370 6309 8384
rect 6346 8354 6365 8384
rect 6380 8354 6386 8384
rect 6395 8354 6408 8384
rect 6423 8370 6453 8384
rect 6496 8370 6539 8384
rect 6546 8370 6766 8384
rect 6773 8370 6803 8384
rect 6463 8356 6478 8368
rect 6497 8356 6510 8370
rect 6578 8366 6731 8370
rect 6460 8354 6482 8356
rect 6560 8354 6752 8366
rect 6831 8354 6844 8384
rect 6859 8370 6889 8384
rect 6926 8354 6945 8384
rect 6960 8354 6966 8384
rect 6975 8354 6988 8384
rect 7003 8370 7033 8384
rect 7076 8370 7119 8384
rect 7126 8370 7346 8384
rect 7353 8370 7383 8384
rect 7043 8356 7058 8368
rect 7077 8356 7090 8370
rect 7158 8366 7311 8370
rect 7040 8354 7062 8356
rect 7140 8354 7332 8366
rect 7411 8354 7424 8384
rect 7439 8370 7469 8384
rect 7506 8354 7525 8384
rect 7540 8354 7546 8384
rect 7555 8354 7568 8384
rect 7583 8370 7613 8384
rect 7656 8370 7699 8384
rect 7706 8370 7926 8384
rect 7933 8370 7963 8384
rect 7623 8356 7638 8368
rect 7657 8356 7670 8370
rect 7738 8366 7891 8370
rect 7620 8354 7642 8356
rect 7720 8354 7912 8366
rect 7991 8354 8004 8384
rect 8019 8370 8049 8384
rect 8086 8354 8105 8384
rect 8120 8354 8126 8384
rect 8135 8354 8148 8384
rect 8163 8370 8193 8384
rect 8236 8370 8279 8384
rect 8286 8370 8506 8384
rect 8513 8370 8543 8384
rect 8203 8356 8218 8368
rect 8237 8356 8250 8370
rect 8318 8366 8471 8370
rect 8200 8354 8222 8356
rect 8300 8354 8492 8366
rect 8571 8354 8584 8384
rect 8599 8370 8629 8384
rect 8666 8354 8685 8384
rect 8700 8354 8706 8384
rect 8715 8354 8728 8384
rect 8743 8370 8773 8384
rect 8816 8370 8859 8384
rect 8866 8370 9086 8384
rect 9093 8370 9123 8384
rect 8783 8356 8798 8368
rect 8817 8356 8830 8370
rect 8898 8366 9051 8370
rect 8780 8354 8802 8356
rect 8880 8354 9072 8366
rect 9151 8354 9164 8384
rect 9179 8370 9209 8384
rect 9246 8354 9265 8384
rect 9280 8354 9286 8384
rect 9295 8354 9308 8384
rect 9323 8370 9353 8384
rect 9396 8370 9439 8384
rect 9446 8370 9666 8384
rect 9673 8370 9703 8384
rect 9363 8356 9378 8368
rect 9397 8356 9410 8370
rect 9478 8366 9631 8370
rect 9360 8354 9382 8356
rect 9460 8354 9652 8366
rect 9731 8354 9744 8384
rect 9759 8370 9789 8384
rect 9826 8354 9845 8384
rect 9860 8354 9866 8384
rect 9875 8354 9888 8384
rect 9903 8370 9933 8384
rect 9976 8370 10019 8384
rect 10026 8370 10246 8384
rect 10253 8370 10283 8384
rect 9943 8356 9958 8368
rect 9977 8356 9990 8370
rect 10058 8366 10211 8370
rect 9940 8354 9962 8356
rect 10040 8354 10232 8366
rect 10311 8354 10324 8384
rect 10339 8370 10369 8384
rect 10406 8354 10425 8384
rect 10440 8354 10446 8384
rect 10455 8354 10468 8384
rect 10483 8370 10513 8384
rect 10556 8370 10599 8384
rect 10606 8370 10826 8384
rect 10833 8370 10863 8384
rect 10523 8356 10538 8368
rect 10557 8356 10570 8370
rect 10638 8366 10791 8370
rect 10520 8354 10542 8356
rect 10620 8354 10812 8366
rect 10891 8354 10904 8384
rect 10919 8370 10949 8384
rect 10986 8354 11005 8384
rect 11020 8354 11026 8384
rect 11035 8354 11048 8384
rect 11063 8370 11093 8384
rect 11136 8370 11179 8384
rect 11186 8370 11406 8384
rect 11413 8370 11443 8384
rect 11103 8356 11118 8368
rect 11137 8356 11150 8370
rect 11218 8366 11371 8370
rect 11100 8354 11122 8356
rect 11200 8354 11392 8366
rect 11471 8354 11484 8384
rect 11499 8370 11529 8384
rect 11566 8354 11585 8384
rect 11600 8354 11606 8384
rect 11615 8354 11628 8384
rect 11643 8370 11673 8384
rect 11716 8370 11759 8384
rect 11766 8370 11986 8384
rect 11993 8370 12023 8384
rect 11683 8356 11698 8368
rect 11717 8356 11730 8370
rect 11798 8366 11951 8370
rect 11680 8354 11702 8356
rect 11780 8354 11972 8366
rect 12051 8354 12064 8384
rect 12079 8370 12109 8384
rect 12146 8354 12165 8384
rect 12180 8354 12186 8384
rect 12195 8354 12208 8384
rect 12223 8370 12253 8384
rect 12296 8370 12339 8384
rect 12346 8370 12566 8384
rect 12573 8370 12603 8384
rect 12263 8356 12278 8368
rect 12297 8356 12310 8370
rect 12378 8366 12531 8370
rect 12260 8354 12282 8356
rect 12360 8354 12552 8366
rect 12631 8354 12644 8384
rect 12659 8370 12689 8384
rect 12726 8354 12745 8384
rect 12760 8354 12766 8384
rect 12775 8354 12788 8384
rect 12803 8370 12833 8384
rect 12876 8370 12919 8384
rect 12926 8370 13146 8384
rect 13153 8370 13183 8384
rect 12843 8356 12858 8368
rect 12877 8356 12890 8370
rect 12958 8366 13111 8370
rect 12840 8354 12862 8356
rect 12940 8354 13132 8366
rect 13211 8354 13224 8384
rect 13239 8370 13269 8384
rect 13306 8354 13325 8384
rect 13340 8354 13346 8384
rect 13355 8354 13368 8384
rect 13383 8370 13413 8384
rect 13456 8370 13499 8384
rect 13506 8370 13726 8384
rect 13733 8370 13763 8384
rect 13423 8356 13438 8368
rect 13457 8356 13470 8370
rect 13538 8366 13691 8370
rect 13420 8354 13442 8356
rect 13520 8354 13712 8366
rect 13791 8354 13804 8384
rect 13819 8370 13849 8384
rect 13886 8354 13905 8384
rect 13920 8354 13926 8384
rect 13935 8354 13948 8384
rect 13963 8370 13993 8384
rect 14036 8370 14079 8384
rect 14086 8370 14306 8384
rect 14313 8370 14343 8384
rect 14003 8356 14018 8368
rect 14037 8356 14050 8370
rect 14118 8366 14271 8370
rect 14000 8354 14022 8356
rect 14100 8354 14292 8366
rect 14371 8354 14384 8384
rect 14399 8370 14429 8384
rect 14466 8354 14485 8384
rect 14500 8354 14506 8384
rect 14515 8354 14528 8384
rect 14543 8370 14573 8384
rect 14616 8370 14659 8384
rect 14666 8370 14886 8384
rect 14893 8370 14923 8384
rect 14583 8356 14598 8368
rect 14617 8356 14630 8370
rect 14698 8366 14851 8370
rect 14580 8354 14602 8356
rect 14680 8354 14872 8366
rect 14951 8354 14964 8384
rect 14979 8370 15009 8384
rect 15046 8354 15065 8384
rect 15080 8354 15086 8384
rect 15095 8354 15108 8384
rect 15123 8370 15153 8384
rect 15196 8370 15239 8384
rect 15246 8370 15466 8384
rect 15473 8370 15503 8384
rect 15163 8356 15178 8368
rect 15197 8356 15210 8370
rect 15278 8366 15431 8370
rect 15160 8354 15182 8356
rect 15260 8354 15452 8366
rect 15531 8354 15544 8384
rect 15559 8370 15589 8384
rect 15626 8354 15645 8384
rect 15660 8354 15666 8384
rect 15675 8354 15688 8384
rect 15703 8370 15733 8384
rect 15776 8370 15819 8384
rect 15826 8370 16046 8384
rect 16053 8370 16083 8384
rect 15743 8356 15758 8368
rect 15777 8356 15790 8370
rect 15858 8366 16011 8370
rect 15740 8354 15762 8356
rect 15840 8354 16032 8366
rect 16111 8354 16124 8384
rect 16139 8370 16169 8384
rect 16206 8354 16225 8384
rect 16240 8354 16246 8384
rect 16255 8354 16268 8384
rect 16283 8370 16313 8384
rect 16356 8370 16399 8384
rect 16406 8370 16626 8384
rect 16633 8370 16663 8384
rect 16323 8356 16338 8368
rect 16357 8356 16370 8370
rect 16438 8366 16591 8370
rect 16320 8354 16342 8356
rect 16420 8354 16612 8366
rect 16691 8354 16704 8384
rect 16719 8370 16749 8384
rect 16786 8354 16805 8384
rect 16820 8354 16826 8384
rect 16835 8354 16848 8384
rect 16863 8370 16893 8384
rect 16936 8370 16979 8384
rect 16986 8370 17206 8384
rect 17213 8370 17243 8384
rect 16903 8356 16918 8368
rect 16937 8356 16950 8370
rect 17018 8366 17171 8370
rect 16900 8354 16922 8356
rect 17000 8354 17192 8366
rect 17271 8354 17284 8384
rect 17299 8370 17329 8384
rect 17366 8354 17385 8384
rect 17400 8354 17406 8384
rect 17415 8354 17428 8384
rect 17443 8370 17473 8384
rect 17516 8370 17559 8384
rect 17566 8370 17786 8384
rect 17793 8370 17823 8384
rect 17483 8356 17498 8368
rect 17517 8356 17530 8370
rect 17598 8366 17751 8370
rect 17480 8354 17502 8356
rect 17580 8354 17772 8366
rect 17851 8354 17864 8384
rect 17879 8370 17909 8384
rect 17946 8354 17965 8384
rect 17980 8354 17986 8384
rect 17995 8354 18008 8384
rect 18023 8370 18053 8384
rect 18096 8370 18139 8384
rect 18146 8370 18366 8384
rect 18373 8370 18403 8384
rect 18063 8356 18078 8368
rect 18097 8356 18110 8370
rect 18178 8366 18331 8370
rect 18060 8354 18082 8356
rect 18160 8354 18352 8366
rect 18431 8354 18444 8384
rect 18459 8370 18489 8384
rect 18532 8354 18545 8384
rect 0 8340 18545 8354
rect 15 8270 28 8340
rect 80 8336 102 8340
rect 73 8314 102 8328
rect 155 8314 171 8328
rect 209 8324 215 8326
rect 222 8324 330 8340
rect 337 8324 343 8326
rect 351 8324 366 8340
rect 432 8334 451 8337
rect 73 8312 171 8314
rect 198 8312 366 8324
rect 381 8314 397 8328
rect 432 8315 454 8334
rect 464 8328 480 8329
rect 463 8326 480 8328
rect 464 8321 480 8326
rect 454 8314 460 8315
rect 463 8314 492 8321
rect 381 8313 492 8314
rect 381 8312 498 8313
rect 57 8304 108 8312
rect 155 8304 189 8312
rect 57 8292 82 8304
rect 89 8292 108 8304
rect 162 8302 189 8304
rect 198 8302 419 8312
rect 454 8309 460 8312
rect 162 8298 419 8302
rect 57 8284 108 8292
rect 155 8284 419 8298
rect 463 8304 498 8312
rect 9 8236 28 8270
rect 73 8276 102 8284
rect 73 8270 90 8276
rect 73 8268 107 8270
rect 155 8268 171 8284
rect 172 8274 380 8284
rect 381 8274 397 8284
rect 445 8280 460 8295
rect 463 8292 464 8304
rect 471 8292 498 8304
rect 463 8284 498 8292
rect 463 8283 492 8284
rect 183 8270 397 8274
rect 198 8268 397 8270
rect 432 8270 445 8280
rect 463 8270 480 8283
rect 432 8268 480 8270
rect 74 8264 107 8268
rect 70 8262 107 8264
rect 70 8261 137 8262
rect 70 8256 101 8261
rect 107 8256 137 8261
rect 70 8252 137 8256
rect 43 8249 137 8252
rect 43 8242 92 8249
rect 43 8236 73 8242
rect 92 8237 97 8242
rect 9 8220 89 8236
rect 101 8228 137 8249
rect 198 8244 387 8268
rect 432 8267 479 8268
rect 445 8262 479 8267
rect 213 8241 387 8244
rect 206 8238 387 8241
rect 415 8261 479 8262
rect 9 8218 28 8220
rect 43 8218 77 8220
rect 9 8202 89 8218
rect 9 8196 28 8202
rect -1 8180 28 8196
rect 43 8186 73 8202
rect 101 8180 107 8228
rect 110 8222 129 8228
rect 144 8222 174 8230
rect 110 8214 174 8222
rect 110 8198 190 8214
rect 206 8207 268 8238
rect 284 8207 346 8238
rect 415 8236 464 8261
rect 479 8236 509 8252
rect 378 8222 408 8230
rect 415 8228 525 8236
rect 378 8214 423 8222
rect 110 8196 129 8198
rect 144 8196 190 8198
rect 110 8180 190 8196
rect 217 8194 252 8207
rect 293 8204 330 8207
rect 293 8202 335 8204
rect 222 8191 252 8194
rect 231 8187 238 8191
rect 238 8186 239 8187
rect 197 8180 207 8186
rect -7 8172 34 8180
rect -7 8146 8 8172
rect 15 8146 34 8172
rect 98 8168 129 8180
rect 144 8168 247 8180
rect 259 8170 285 8196
rect 300 8191 330 8202
rect 362 8198 424 8214
rect 362 8196 408 8198
rect 362 8180 424 8196
rect 436 8180 442 8228
rect 445 8220 525 8228
rect 445 8218 464 8220
rect 479 8218 513 8220
rect 445 8202 525 8218
rect 445 8180 464 8202
rect 479 8186 509 8202
rect 537 8196 543 8270
rect 546 8196 565 8340
rect 580 8196 586 8340
rect 595 8270 608 8340
rect 660 8336 682 8340
rect 653 8314 682 8328
rect 735 8314 751 8328
rect 789 8324 795 8326
rect 802 8324 910 8340
rect 917 8324 923 8326
rect 931 8324 946 8340
rect 1012 8334 1031 8337
rect 653 8312 751 8314
rect 778 8312 946 8324
rect 961 8314 977 8328
rect 1012 8315 1034 8334
rect 1044 8328 1060 8329
rect 1043 8326 1060 8328
rect 1044 8321 1060 8326
rect 1034 8314 1040 8315
rect 1043 8314 1072 8321
rect 961 8313 1072 8314
rect 961 8312 1078 8313
rect 637 8304 688 8312
rect 735 8304 769 8312
rect 637 8292 662 8304
rect 669 8292 688 8304
rect 742 8302 769 8304
rect 778 8302 999 8312
rect 1034 8309 1040 8312
rect 742 8298 999 8302
rect 637 8284 688 8292
rect 735 8284 999 8298
rect 1043 8304 1078 8312
rect 589 8236 608 8270
rect 653 8276 682 8284
rect 653 8270 670 8276
rect 653 8268 687 8270
rect 735 8268 751 8284
rect 752 8274 960 8284
rect 961 8274 977 8284
rect 1025 8280 1040 8295
rect 1043 8292 1044 8304
rect 1051 8292 1078 8304
rect 1043 8284 1078 8292
rect 1043 8283 1072 8284
rect 763 8270 977 8274
rect 778 8268 977 8270
rect 1012 8270 1025 8280
rect 1043 8270 1060 8283
rect 1012 8268 1060 8270
rect 654 8264 687 8268
rect 650 8262 687 8264
rect 650 8261 717 8262
rect 650 8256 681 8261
rect 687 8256 717 8261
rect 650 8252 717 8256
rect 623 8249 717 8252
rect 623 8242 672 8249
rect 623 8236 653 8242
rect 672 8237 677 8242
rect 589 8220 669 8236
rect 681 8228 717 8249
rect 778 8244 967 8268
rect 1012 8267 1059 8268
rect 1025 8262 1059 8267
rect 793 8241 967 8244
rect 786 8238 967 8241
rect 995 8261 1059 8262
rect 589 8218 608 8220
rect 623 8218 657 8220
rect 589 8202 669 8218
rect 589 8196 608 8202
rect 305 8170 408 8180
rect 259 8168 408 8170
rect 429 8168 464 8180
rect 98 8166 260 8168
rect 110 8146 129 8166
rect 144 8164 174 8166
rect -7 8138 34 8146
rect 116 8142 129 8146
rect 181 8150 260 8166
rect 292 8166 464 8168
rect 292 8150 371 8166
rect 378 8164 408 8166
rect -1 8128 28 8138
rect 43 8128 73 8142
rect 116 8128 159 8142
rect 181 8138 371 8150
rect 436 8146 442 8166
rect 166 8128 196 8138
rect 197 8128 355 8138
rect 359 8128 389 8138
rect 393 8128 423 8142
rect 451 8128 464 8166
rect 536 8180 565 8196
rect 579 8180 608 8196
rect 623 8186 653 8202
rect 681 8180 687 8228
rect 690 8222 709 8228
rect 724 8222 754 8230
rect 690 8214 754 8222
rect 690 8198 770 8214
rect 786 8207 848 8238
rect 864 8207 926 8238
rect 995 8236 1044 8261
rect 1059 8236 1089 8252
rect 958 8222 988 8230
rect 995 8228 1105 8236
rect 958 8214 1003 8222
rect 690 8196 709 8198
rect 724 8196 770 8198
rect 690 8180 770 8196
rect 797 8194 832 8207
rect 873 8204 910 8207
rect 873 8202 915 8204
rect 802 8191 832 8194
rect 811 8187 818 8191
rect 818 8186 819 8187
rect 777 8180 787 8186
rect 536 8172 571 8180
rect 536 8146 537 8172
rect 544 8146 571 8172
rect 479 8128 509 8142
rect 536 8138 571 8146
rect 573 8172 614 8180
rect 573 8146 588 8172
rect 595 8146 614 8172
rect 678 8168 709 8180
rect 724 8168 827 8180
rect 839 8170 865 8196
rect 880 8191 910 8202
rect 942 8198 1004 8214
rect 942 8196 988 8198
rect 942 8180 1004 8196
rect 1016 8180 1022 8228
rect 1025 8220 1105 8228
rect 1025 8218 1044 8220
rect 1059 8218 1093 8220
rect 1025 8202 1105 8218
rect 1025 8180 1044 8202
rect 1059 8186 1089 8202
rect 1117 8196 1123 8270
rect 1126 8196 1145 8340
rect 1160 8196 1166 8340
rect 1175 8270 1188 8340
rect 1240 8336 1262 8340
rect 1233 8314 1262 8328
rect 1315 8314 1331 8328
rect 1369 8324 1375 8326
rect 1382 8324 1490 8340
rect 1497 8324 1503 8326
rect 1511 8324 1526 8340
rect 1592 8334 1611 8337
rect 1233 8312 1331 8314
rect 1358 8312 1526 8324
rect 1541 8314 1557 8328
rect 1592 8315 1614 8334
rect 1624 8328 1640 8329
rect 1623 8326 1640 8328
rect 1624 8321 1640 8326
rect 1614 8314 1620 8315
rect 1623 8314 1652 8321
rect 1541 8313 1652 8314
rect 1541 8312 1658 8313
rect 1217 8304 1268 8312
rect 1315 8304 1349 8312
rect 1217 8292 1242 8304
rect 1249 8292 1268 8304
rect 1322 8302 1349 8304
rect 1358 8302 1579 8312
rect 1614 8309 1620 8312
rect 1322 8298 1579 8302
rect 1217 8284 1268 8292
rect 1315 8284 1579 8298
rect 1623 8304 1658 8312
rect 1169 8236 1188 8270
rect 1233 8276 1262 8284
rect 1233 8270 1250 8276
rect 1233 8268 1267 8270
rect 1315 8268 1331 8284
rect 1332 8274 1540 8284
rect 1541 8274 1557 8284
rect 1605 8280 1620 8295
rect 1623 8292 1624 8304
rect 1631 8292 1658 8304
rect 1623 8284 1658 8292
rect 1623 8283 1652 8284
rect 1343 8270 1557 8274
rect 1358 8268 1557 8270
rect 1592 8270 1605 8280
rect 1623 8270 1640 8283
rect 1592 8268 1640 8270
rect 1234 8264 1267 8268
rect 1230 8262 1267 8264
rect 1230 8261 1297 8262
rect 1230 8256 1261 8261
rect 1267 8256 1297 8261
rect 1230 8252 1297 8256
rect 1203 8249 1297 8252
rect 1203 8242 1252 8249
rect 1203 8236 1233 8242
rect 1252 8237 1257 8242
rect 1169 8220 1249 8236
rect 1261 8228 1297 8249
rect 1358 8244 1547 8268
rect 1592 8267 1639 8268
rect 1605 8262 1639 8267
rect 1373 8241 1547 8244
rect 1366 8238 1547 8241
rect 1575 8261 1639 8262
rect 1169 8218 1188 8220
rect 1203 8218 1237 8220
rect 1169 8202 1249 8218
rect 1169 8196 1188 8202
rect 885 8170 988 8180
rect 839 8168 988 8170
rect 1009 8168 1044 8180
rect 678 8166 840 8168
rect 690 8146 709 8166
rect 724 8164 754 8166
rect 573 8138 614 8146
rect 696 8142 709 8146
rect 761 8150 840 8166
rect 872 8166 1044 8168
rect 872 8150 951 8166
rect 958 8164 988 8166
rect 536 8128 565 8138
rect 579 8128 608 8138
rect 623 8128 653 8142
rect 696 8128 739 8142
rect 761 8138 951 8150
rect 1016 8146 1022 8166
rect 746 8128 776 8138
rect 777 8128 935 8138
rect 939 8128 969 8138
rect 973 8128 1003 8142
rect 1031 8128 1044 8166
rect 1116 8180 1145 8196
rect 1159 8180 1188 8196
rect 1203 8186 1233 8202
rect 1261 8180 1267 8228
rect 1270 8222 1289 8228
rect 1304 8222 1334 8230
rect 1270 8214 1334 8222
rect 1270 8198 1350 8214
rect 1366 8207 1428 8238
rect 1444 8207 1506 8238
rect 1575 8236 1624 8261
rect 1639 8236 1669 8252
rect 1538 8222 1568 8230
rect 1575 8228 1685 8236
rect 1538 8214 1583 8222
rect 1270 8196 1289 8198
rect 1304 8196 1350 8198
rect 1270 8180 1350 8196
rect 1377 8194 1412 8207
rect 1453 8204 1490 8207
rect 1453 8202 1495 8204
rect 1382 8191 1412 8194
rect 1391 8187 1398 8191
rect 1398 8186 1399 8187
rect 1357 8180 1367 8186
rect 1116 8172 1151 8180
rect 1116 8146 1117 8172
rect 1124 8146 1151 8172
rect 1059 8128 1089 8142
rect 1116 8138 1151 8146
rect 1153 8172 1194 8180
rect 1153 8146 1168 8172
rect 1175 8146 1194 8172
rect 1258 8168 1289 8180
rect 1304 8168 1407 8180
rect 1419 8170 1445 8196
rect 1460 8191 1490 8202
rect 1522 8198 1584 8214
rect 1522 8196 1568 8198
rect 1522 8180 1584 8196
rect 1596 8180 1602 8228
rect 1605 8220 1685 8228
rect 1605 8218 1624 8220
rect 1639 8218 1673 8220
rect 1605 8202 1685 8218
rect 1605 8180 1624 8202
rect 1639 8186 1669 8202
rect 1697 8196 1703 8270
rect 1706 8196 1725 8340
rect 1740 8196 1746 8340
rect 1755 8270 1768 8340
rect 1820 8336 1842 8340
rect 1813 8314 1842 8328
rect 1895 8314 1911 8328
rect 1949 8324 1955 8326
rect 1962 8324 2070 8340
rect 2077 8324 2083 8326
rect 2091 8324 2106 8340
rect 2172 8334 2191 8337
rect 1813 8312 1911 8314
rect 1938 8312 2106 8324
rect 2121 8314 2137 8328
rect 2172 8315 2194 8334
rect 2204 8328 2220 8329
rect 2203 8326 2220 8328
rect 2204 8321 2220 8326
rect 2194 8314 2200 8315
rect 2203 8314 2232 8321
rect 2121 8313 2232 8314
rect 2121 8312 2238 8313
rect 1797 8304 1848 8312
rect 1895 8304 1929 8312
rect 1797 8292 1822 8304
rect 1829 8292 1848 8304
rect 1902 8302 1929 8304
rect 1938 8302 2159 8312
rect 2194 8309 2200 8312
rect 1902 8298 2159 8302
rect 1797 8284 1848 8292
rect 1895 8284 2159 8298
rect 2203 8304 2238 8312
rect 1749 8236 1768 8270
rect 1813 8276 1842 8284
rect 1813 8270 1830 8276
rect 1813 8268 1847 8270
rect 1895 8268 1911 8284
rect 1912 8274 2120 8284
rect 2121 8274 2137 8284
rect 2185 8280 2200 8295
rect 2203 8292 2204 8304
rect 2211 8292 2238 8304
rect 2203 8284 2238 8292
rect 2203 8283 2232 8284
rect 1923 8270 2137 8274
rect 1938 8268 2137 8270
rect 2172 8270 2185 8280
rect 2203 8270 2220 8283
rect 2172 8268 2220 8270
rect 1814 8264 1847 8268
rect 1810 8262 1847 8264
rect 1810 8261 1877 8262
rect 1810 8256 1841 8261
rect 1847 8256 1877 8261
rect 1810 8252 1877 8256
rect 1783 8249 1877 8252
rect 1783 8242 1832 8249
rect 1783 8236 1813 8242
rect 1832 8237 1837 8242
rect 1749 8220 1829 8236
rect 1841 8228 1877 8249
rect 1938 8244 2127 8268
rect 2172 8267 2219 8268
rect 2185 8262 2219 8267
rect 1953 8241 2127 8244
rect 1946 8238 2127 8241
rect 2155 8261 2219 8262
rect 1749 8218 1768 8220
rect 1783 8218 1817 8220
rect 1749 8202 1829 8218
rect 1749 8196 1768 8202
rect 1465 8170 1568 8180
rect 1419 8168 1568 8170
rect 1589 8168 1624 8180
rect 1258 8166 1420 8168
rect 1270 8146 1289 8166
rect 1304 8164 1334 8166
rect 1153 8138 1194 8146
rect 1276 8142 1289 8146
rect 1341 8150 1420 8166
rect 1452 8166 1624 8168
rect 1452 8150 1531 8166
rect 1538 8164 1568 8166
rect 1116 8128 1145 8138
rect 1159 8128 1188 8138
rect 1203 8128 1233 8142
rect 1276 8128 1319 8142
rect 1341 8138 1531 8150
rect 1596 8146 1602 8166
rect 1326 8128 1356 8138
rect 1357 8128 1515 8138
rect 1519 8128 1549 8138
rect 1553 8128 1583 8142
rect 1611 8128 1624 8166
rect 1696 8180 1725 8196
rect 1739 8180 1768 8196
rect 1783 8186 1813 8202
rect 1841 8180 1847 8228
rect 1850 8222 1869 8228
rect 1884 8222 1914 8230
rect 1850 8214 1914 8222
rect 1850 8198 1930 8214
rect 1946 8207 2008 8238
rect 2024 8207 2086 8238
rect 2155 8236 2204 8261
rect 2219 8236 2249 8252
rect 2118 8222 2148 8230
rect 2155 8228 2265 8236
rect 2118 8214 2163 8222
rect 1850 8196 1869 8198
rect 1884 8196 1930 8198
rect 1850 8180 1930 8196
rect 1957 8194 1992 8207
rect 2033 8204 2070 8207
rect 2033 8202 2075 8204
rect 1962 8191 1992 8194
rect 1971 8187 1978 8191
rect 1978 8186 1979 8187
rect 1937 8180 1947 8186
rect 1696 8172 1731 8180
rect 1696 8146 1697 8172
rect 1704 8146 1731 8172
rect 1639 8128 1669 8142
rect 1696 8138 1731 8146
rect 1733 8172 1774 8180
rect 1733 8146 1748 8172
rect 1755 8146 1774 8172
rect 1838 8168 1869 8180
rect 1884 8168 1987 8180
rect 1999 8170 2025 8196
rect 2040 8191 2070 8202
rect 2102 8198 2164 8214
rect 2102 8196 2148 8198
rect 2102 8180 2164 8196
rect 2176 8180 2182 8228
rect 2185 8220 2265 8228
rect 2185 8218 2204 8220
rect 2219 8218 2253 8220
rect 2185 8202 2265 8218
rect 2185 8180 2204 8202
rect 2219 8186 2249 8202
rect 2277 8196 2283 8270
rect 2286 8196 2305 8340
rect 2320 8196 2326 8340
rect 2335 8270 2348 8340
rect 2400 8336 2422 8340
rect 2393 8314 2422 8328
rect 2475 8314 2491 8328
rect 2529 8324 2535 8326
rect 2542 8324 2650 8340
rect 2657 8324 2663 8326
rect 2671 8324 2686 8340
rect 2752 8334 2771 8337
rect 2393 8312 2491 8314
rect 2518 8312 2686 8324
rect 2701 8314 2717 8328
rect 2752 8315 2774 8334
rect 2784 8328 2800 8329
rect 2783 8326 2800 8328
rect 2784 8321 2800 8326
rect 2774 8314 2780 8315
rect 2783 8314 2812 8321
rect 2701 8313 2812 8314
rect 2701 8312 2818 8313
rect 2377 8304 2428 8312
rect 2475 8304 2509 8312
rect 2377 8292 2402 8304
rect 2409 8292 2428 8304
rect 2482 8302 2509 8304
rect 2518 8302 2739 8312
rect 2774 8309 2780 8312
rect 2482 8298 2739 8302
rect 2377 8284 2428 8292
rect 2475 8284 2739 8298
rect 2783 8304 2818 8312
rect 2329 8236 2348 8270
rect 2393 8276 2422 8284
rect 2393 8270 2410 8276
rect 2393 8268 2427 8270
rect 2475 8268 2491 8284
rect 2492 8274 2700 8284
rect 2701 8274 2717 8284
rect 2765 8280 2780 8295
rect 2783 8292 2784 8304
rect 2791 8292 2818 8304
rect 2783 8284 2818 8292
rect 2783 8283 2812 8284
rect 2503 8270 2717 8274
rect 2518 8268 2717 8270
rect 2752 8270 2765 8280
rect 2783 8270 2800 8283
rect 2752 8268 2800 8270
rect 2394 8264 2427 8268
rect 2390 8262 2427 8264
rect 2390 8261 2457 8262
rect 2390 8256 2421 8261
rect 2427 8256 2457 8261
rect 2390 8252 2457 8256
rect 2363 8249 2457 8252
rect 2363 8242 2412 8249
rect 2363 8236 2393 8242
rect 2412 8237 2417 8242
rect 2329 8220 2409 8236
rect 2421 8228 2457 8249
rect 2518 8244 2707 8268
rect 2752 8267 2799 8268
rect 2765 8262 2799 8267
rect 2533 8241 2707 8244
rect 2526 8238 2707 8241
rect 2735 8261 2799 8262
rect 2329 8218 2348 8220
rect 2363 8218 2397 8220
rect 2329 8202 2409 8218
rect 2329 8196 2348 8202
rect 2045 8170 2148 8180
rect 1999 8168 2148 8170
rect 2169 8168 2204 8180
rect 1838 8166 2000 8168
rect 1850 8146 1869 8166
rect 1884 8164 1914 8166
rect 1733 8138 1774 8146
rect 1856 8142 1869 8146
rect 1921 8150 2000 8166
rect 2032 8166 2204 8168
rect 2032 8150 2111 8166
rect 2118 8164 2148 8166
rect 1696 8128 1725 8138
rect 1739 8128 1768 8138
rect 1783 8128 1813 8142
rect 1856 8128 1899 8142
rect 1921 8138 2111 8150
rect 2176 8146 2182 8166
rect 1906 8128 1936 8138
rect 1937 8128 2095 8138
rect 2099 8128 2129 8138
rect 2133 8128 2163 8142
rect 2191 8128 2204 8166
rect 2276 8180 2305 8196
rect 2319 8180 2348 8196
rect 2363 8186 2393 8202
rect 2421 8180 2427 8228
rect 2430 8222 2449 8228
rect 2464 8222 2494 8230
rect 2430 8214 2494 8222
rect 2430 8198 2510 8214
rect 2526 8207 2588 8238
rect 2604 8207 2666 8238
rect 2735 8236 2784 8261
rect 2799 8236 2829 8252
rect 2698 8222 2728 8230
rect 2735 8228 2845 8236
rect 2698 8214 2743 8222
rect 2430 8196 2449 8198
rect 2464 8196 2510 8198
rect 2430 8180 2510 8196
rect 2537 8194 2572 8207
rect 2613 8204 2650 8207
rect 2613 8202 2655 8204
rect 2542 8191 2572 8194
rect 2551 8187 2558 8191
rect 2558 8186 2559 8187
rect 2517 8180 2527 8186
rect 2276 8172 2311 8180
rect 2276 8146 2277 8172
rect 2284 8146 2311 8172
rect 2219 8128 2249 8142
rect 2276 8138 2311 8146
rect 2313 8172 2354 8180
rect 2313 8146 2328 8172
rect 2335 8146 2354 8172
rect 2418 8168 2449 8180
rect 2464 8168 2567 8180
rect 2579 8170 2605 8196
rect 2620 8191 2650 8202
rect 2682 8198 2744 8214
rect 2682 8196 2728 8198
rect 2682 8180 2744 8196
rect 2756 8180 2762 8228
rect 2765 8220 2845 8228
rect 2765 8218 2784 8220
rect 2799 8218 2833 8220
rect 2765 8202 2845 8218
rect 2765 8180 2784 8202
rect 2799 8186 2829 8202
rect 2857 8196 2863 8270
rect 2866 8196 2885 8340
rect 2900 8196 2906 8340
rect 2915 8270 2928 8340
rect 2980 8336 3002 8340
rect 2973 8314 3002 8328
rect 3055 8314 3071 8328
rect 3109 8324 3115 8326
rect 3122 8324 3230 8340
rect 3237 8324 3243 8326
rect 3251 8324 3266 8340
rect 3332 8334 3351 8337
rect 2973 8312 3071 8314
rect 3098 8312 3266 8324
rect 3281 8314 3297 8328
rect 3332 8315 3354 8334
rect 3364 8328 3380 8329
rect 3363 8326 3380 8328
rect 3364 8321 3380 8326
rect 3354 8314 3360 8315
rect 3363 8314 3392 8321
rect 3281 8313 3392 8314
rect 3281 8312 3398 8313
rect 2957 8304 3008 8312
rect 3055 8304 3089 8312
rect 2957 8292 2982 8304
rect 2989 8292 3008 8304
rect 3062 8302 3089 8304
rect 3098 8302 3319 8312
rect 3354 8309 3360 8312
rect 3062 8298 3319 8302
rect 2957 8284 3008 8292
rect 3055 8284 3319 8298
rect 3363 8304 3398 8312
rect 2909 8236 2928 8270
rect 2973 8276 3002 8284
rect 2973 8270 2990 8276
rect 2973 8268 3007 8270
rect 3055 8268 3071 8284
rect 3072 8274 3280 8284
rect 3281 8274 3297 8284
rect 3345 8280 3360 8295
rect 3363 8292 3364 8304
rect 3371 8292 3398 8304
rect 3363 8284 3398 8292
rect 3363 8283 3392 8284
rect 3083 8270 3297 8274
rect 3098 8268 3297 8270
rect 3332 8270 3345 8280
rect 3363 8270 3380 8283
rect 3332 8268 3380 8270
rect 2974 8264 3007 8268
rect 2970 8262 3007 8264
rect 2970 8261 3037 8262
rect 2970 8256 3001 8261
rect 3007 8256 3037 8261
rect 2970 8252 3037 8256
rect 2943 8249 3037 8252
rect 2943 8242 2992 8249
rect 2943 8236 2973 8242
rect 2992 8237 2997 8242
rect 2909 8220 2989 8236
rect 3001 8228 3037 8249
rect 3098 8244 3287 8268
rect 3332 8267 3379 8268
rect 3345 8262 3379 8267
rect 3113 8241 3287 8244
rect 3106 8238 3287 8241
rect 3315 8261 3379 8262
rect 2909 8218 2928 8220
rect 2943 8218 2977 8220
rect 2909 8202 2989 8218
rect 2909 8196 2928 8202
rect 2625 8170 2728 8180
rect 2579 8168 2728 8170
rect 2749 8168 2784 8180
rect 2418 8166 2580 8168
rect 2430 8146 2449 8166
rect 2464 8164 2494 8166
rect 2313 8138 2354 8146
rect 2436 8142 2449 8146
rect 2501 8150 2580 8166
rect 2612 8166 2784 8168
rect 2612 8150 2691 8166
rect 2698 8164 2728 8166
rect 2276 8128 2305 8138
rect 2319 8128 2348 8138
rect 2363 8128 2393 8142
rect 2436 8128 2479 8142
rect 2501 8138 2691 8150
rect 2756 8146 2762 8166
rect 2486 8128 2516 8138
rect 2517 8128 2675 8138
rect 2679 8128 2709 8138
rect 2713 8128 2743 8142
rect 2771 8128 2784 8166
rect 2856 8180 2885 8196
rect 2899 8180 2928 8196
rect 2943 8186 2973 8202
rect 3001 8180 3007 8228
rect 3010 8222 3029 8228
rect 3044 8222 3074 8230
rect 3010 8214 3074 8222
rect 3010 8198 3090 8214
rect 3106 8207 3168 8238
rect 3184 8207 3246 8238
rect 3315 8236 3364 8261
rect 3379 8236 3409 8252
rect 3278 8222 3308 8230
rect 3315 8228 3425 8236
rect 3278 8214 3323 8222
rect 3010 8196 3029 8198
rect 3044 8196 3090 8198
rect 3010 8180 3090 8196
rect 3117 8194 3152 8207
rect 3193 8204 3230 8207
rect 3193 8202 3235 8204
rect 3122 8191 3152 8194
rect 3131 8187 3138 8191
rect 3138 8186 3139 8187
rect 3097 8180 3107 8186
rect 2856 8172 2891 8180
rect 2856 8146 2857 8172
rect 2864 8146 2891 8172
rect 2799 8128 2829 8142
rect 2856 8138 2891 8146
rect 2893 8172 2934 8180
rect 2893 8146 2908 8172
rect 2915 8146 2934 8172
rect 2998 8168 3029 8180
rect 3044 8168 3147 8180
rect 3159 8170 3185 8196
rect 3200 8191 3230 8202
rect 3262 8198 3324 8214
rect 3262 8196 3308 8198
rect 3262 8180 3324 8196
rect 3336 8180 3342 8228
rect 3345 8220 3425 8228
rect 3345 8218 3364 8220
rect 3379 8218 3413 8220
rect 3345 8202 3425 8218
rect 3345 8180 3364 8202
rect 3379 8186 3409 8202
rect 3437 8196 3443 8270
rect 3446 8196 3465 8340
rect 3480 8196 3486 8340
rect 3495 8270 3508 8340
rect 3560 8336 3582 8340
rect 3553 8314 3582 8328
rect 3635 8314 3651 8328
rect 3689 8324 3695 8326
rect 3702 8324 3810 8340
rect 3817 8324 3823 8326
rect 3831 8324 3846 8340
rect 3912 8334 3931 8337
rect 3553 8312 3651 8314
rect 3678 8312 3846 8324
rect 3861 8314 3877 8328
rect 3912 8315 3934 8334
rect 3944 8328 3960 8329
rect 3943 8326 3960 8328
rect 3944 8321 3960 8326
rect 3934 8314 3940 8315
rect 3943 8314 3972 8321
rect 3861 8313 3972 8314
rect 3861 8312 3978 8313
rect 3537 8304 3588 8312
rect 3635 8304 3669 8312
rect 3537 8292 3562 8304
rect 3569 8292 3588 8304
rect 3642 8302 3669 8304
rect 3678 8302 3899 8312
rect 3934 8309 3940 8312
rect 3642 8298 3899 8302
rect 3537 8284 3588 8292
rect 3635 8284 3899 8298
rect 3943 8304 3978 8312
rect 3489 8236 3508 8270
rect 3553 8276 3582 8284
rect 3553 8270 3570 8276
rect 3553 8268 3587 8270
rect 3635 8268 3651 8284
rect 3652 8274 3860 8284
rect 3861 8274 3877 8284
rect 3925 8280 3940 8295
rect 3943 8292 3944 8304
rect 3951 8292 3978 8304
rect 3943 8284 3978 8292
rect 3943 8283 3972 8284
rect 3663 8270 3877 8274
rect 3678 8268 3877 8270
rect 3912 8270 3925 8280
rect 3943 8270 3960 8283
rect 3912 8268 3960 8270
rect 3554 8264 3587 8268
rect 3550 8262 3587 8264
rect 3550 8261 3617 8262
rect 3550 8256 3581 8261
rect 3587 8256 3617 8261
rect 3550 8252 3617 8256
rect 3523 8249 3617 8252
rect 3523 8242 3572 8249
rect 3523 8236 3553 8242
rect 3572 8237 3577 8242
rect 3489 8220 3569 8236
rect 3581 8228 3617 8249
rect 3678 8244 3867 8268
rect 3912 8267 3959 8268
rect 3925 8262 3959 8267
rect 3693 8241 3867 8244
rect 3686 8238 3867 8241
rect 3895 8261 3959 8262
rect 3489 8218 3508 8220
rect 3523 8218 3557 8220
rect 3489 8202 3569 8218
rect 3489 8196 3508 8202
rect 3205 8170 3308 8180
rect 3159 8168 3308 8170
rect 3329 8168 3364 8180
rect 2998 8166 3160 8168
rect 3010 8146 3029 8166
rect 3044 8164 3074 8166
rect 2893 8138 2934 8146
rect 3016 8142 3029 8146
rect 3081 8150 3160 8166
rect 3192 8166 3364 8168
rect 3192 8150 3271 8166
rect 3278 8164 3308 8166
rect 2856 8128 2885 8138
rect 2899 8128 2928 8138
rect 2943 8128 2973 8142
rect 3016 8128 3059 8142
rect 3081 8138 3271 8150
rect 3336 8146 3342 8166
rect 3066 8128 3096 8138
rect 3097 8128 3255 8138
rect 3259 8128 3289 8138
rect 3293 8128 3323 8142
rect 3351 8128 3364 8166
rect 3436 8180 3465 8196
rect 3479 8180 3508 8196
rect 3523 8186 3553 8202
rect 3581 8180 3587 8228
rect 3590 8222 3609 8228
rect 3624 8222 3654 8230
rect 3590 8214 3654 8222
rect 3590 8198 3670 8214
rect 3686 8207 3748 8238
rect 3764 8207 3826 8238
rect 3895 8236 3944 8261
rect 3959 8236 3989 8252
rect 3858 8222 3888 8230
rect 3895 8228 4005 8236
rect 3858 8214 3903 8222
rect 3590 8196 3609 8198
rect 3624 8196 3670 8198
rect 3590 8180 3670 8196
rect 3697 8194 3732 8207
rect 3773 8204 3810 8207
rect 3773 8202 3815 8204
rect 3702 8191 3732 8194
rect 3711 8187 3718 8191
rect 3718 8186 3719 8187
rect 3677 8180 3687 8186
rect 3436 8172 3471 8180
rect 3436 8146 3437 8172
rect 3444 8146 3471 8172
rect 3379 8128 3409 8142
rect 3436 8138 3471 8146
rect 3473 8172 3514 8180
rect 3473 8146 3488 8172
rect 3495 8146 3514 8172
rect 3578 8168 3609 8180
rect 3624 8168 3727 8180
rect 3739 8170 3765 8196
rect 3780 8191 3810 8202
rect 3842 8198 3904 8214
rect 3842 8196 3888 8198
rect 3842 8180 3904 8196
rect 3916 8180 3922 8228
rect 3925 8220 4005 8228
rect 3925 8218 3944 8220
rect 3959 8218 3993 8220
rect 3925 8202 4005 8218
rect 3925 8180 3944 8202
rect 3959 8186 3989 8202
rect 4017 8196 4023 8270
rect 4026 8196 4045 8340
rect 4060 8196 4066 8340
rect 4075 8270 4088 8340
rect 4140 8336 4162 8340
rect 4133 8314 4162 8328
rect 4215 8314 4231 8328
rect 4269 8324 4275 8326
rect 4282 8324 4390 8340
rect 4397 8324 4403 8326
rect 4411 8324 4426 8340
rect 4492 8334 4511 8337
rect 4133 8312 4231 8314
rect 4258 8312 4426 8324
rect 4441 8314 4457 8328
rect 4492 8315 4514 8334
rect 4524 8328 4540 8329
rect 4523 8326 4540 8328
rect 4524 8321 4540 8326
rect 4514 8314 4520 8315
rect 4523 8314 4552 8321
rect 4441 8313 4552 8314
rect 4441 8312 4558 8313
rect 4117 8304 4168 8312
rect 4215 8304 4249 8312
rect 4117 8292 4142 8304
rect 4149 8292 4168 8304
rect 4222 8302 4249 8304
rect 4258 8302 4479 8312
rect 4514 8309 4520 8312
rect 4222 8298 4479 8302
rect 4117 8284 4168 8292
rect 4215 8284 4479 8298
rect 4523 8304 4558 8312
rect 4069 8236 4088 8270
rect 4133 8276 4162 8284
rect 4133 8270 4150 8276
rect 4133 8268 4167 8270
rect 4215 8268 4231 8284
rect 4232 8274 4440 8284
rect 4441 8274 4457 8284
rect 4505 8280 4520 8295
rect 4523 8292 4524 8304
rect 4531 8292 4558 8304
rect 4523 8284 4558 8292
rect 4523 8283 4552 8284
rect 4243 8270 4457 8274
rect 4258 8268 4457 8270
rect 4492 8270 4505 8280
rect 4523 8270 4540 8283
rect 4492 8268 4540 8270
rect 4134 8264 4167 8268
rect 4130 8262 4167 8264
rect 4130 8261 4197 8262
rect 4130 8256 4161 8261
rect 4167 8256 4197 8261
rect 4130 8252 4197 8256
rect 4103 8249 4197 8252
rect 4103 8242 4152 8249
rect 4103 8236 4133 8242
rect 4152 8237 4157 8242
rect 4069 8220 4149 8236
rect 4161 8228 4197 8249
rect 4258 8244 4447 8268
rect 4492 8267 4539 8268
rect 4505 8262 4539 8267
rect 4273 8241 4447 8244
rect 4266 8238 4447 8241
rect 4475 8261 4539 8262
rect 4069 8218 4088 8220
rect 4103 8218 4137 8220
rect 4069 8202 4149 8218
rect 4069 8196 4088 8202
rect 3785 8170 3888 8180
rect 3739 8168 3888 8170
rect 3909 8168 3944 8180
rect 3578 8166 3740 8168
rect 3590 8146 3609 8166
rect 3624 8164 3654 8166
rect 3473 8138 3514 8146
rect 3596 8142 3609 8146
rect 3661 8150 3740 8166
rect 3772 8166 3944 8168
rect 3772 8150 3851 8166
rect 3858 8164 3888 8166
rect 3436 8128 3465 8138
rect 3479 8128 3508 8138
rect 3523 8128 3553 8142
rect 3596 8128 3639 8142
rect 3661 8138 3851 8150
rect 3916 8146 3922 8166
rect 3646 8128 3676 8138
rect 3677 8128 3835 8138
rect 3839 8128 3869 8138
rect 3873 8128 3903 8142
rect 3931 8128 3944 8166
rect 4016 8180 4045 8196
rect 4059 8180 4088 8196
rect 4103 8186 4133 8202
rect 4161 8180 4167 8228
rect 4170 8222 4189 8228
rect 4204 8222 4234 8230
rect 4170 8214 4234 8222
rect 4170 8198 4250 8214
rect 4266 8207 4328 8238
rect 4344 8207 4406 8238
rect 4475 8236 4524 8261
rect 4539 8236 4569 8252
rect 4438 8222 4468 8230
rect 4475 8228 4585 8236
rect 4438 8214 4483 8222
rect 4170 8196 4189 8198
rect 4204 8196 4250 8198
rect 4170 8180 4250 8196
rect 4277 8194 4312 8207
rect 4353 8204 4390 8207
rect 4353 8202 4395 8204
rect 4282 8191 4312 8194
rect 4291 8187 4298 8191
rect 4298 8186 4299 8187
rect 4257 8180 4267 8186
rect 4016 8172 4051 8180
rect 4016 8146 4017 8172
rect 4024 8146 4051 8172
rect 3959 8128 3989 8142
rect 4016 8138 4051 8146
rect 4053 8172 4094 8180
rect 4053 8146 4068 8172
rect 4075 8146 4094 8172
rect 4158 8168 4189 8180
rect 4204 8168 4307 8180
rect 4319 8170 4345 8196
rect 4360 8191 4390 8202
rect 4422 8198 4484 8214
rect 4422 8196 4468 8198
rect 4422 8180 4484 8196
rect 4496 8180 4502 8228
rect 4505 8220 4585 8228
rect 4505 8218 4524 8220
rect 4539 8218 4573 8220
rect 4505 8202 4585 8218
rect 4505 8180 4524 8202
rect 4539 8186 4569 8202
rect 4597 8196 4603 8270
rect 4606 8196 4625 8340
rect 4640 8196 4646 8340
rect 4655 8270 4668 8340
rect 4720 8336 4742 8340
rect 4713 8314 4742 8328
rect 4795 8314 4811 8328
rect 4849 8324 4855 8326
rect 4862 8324 4970 8340
rect 4977 8324 4983 8326
rect 4991 8324 5006 8340
rect 5072 8334 5091 8337
rect 4713 8312 4811 8314
rect 4838 8312 5006 8324
rect 5021 8314 5037 8328
rect 5072 8315 5094 8334
rect 5104 8328 5120 8329
rect 5103 8326 5120 8328
rect 5104 8321 5120 8326
rect 5094 8314 5100 8315
rect 5103 8314 5132 8321
rect 5021 8313 5132 8314
rect 5021 8312 5138 8313
rect 4697 8304 4748 8312
rect 4795 8304 4829 8312
rect 4697 8292 4722 8304
rect 4729 8292 4748 8304
rect 4802 8302 4829 8304
rect 4838 8302 5059 8312
rect 5094 8309 5100 8312
rect 4802 8298 5059 8302
rect 4697 8284 4748 8292
rect 4795 8284 5059 8298
rect 5103 8304 5138 8312
rect 4649 8236 4668 8270
rect 4713 8276 4742 8284
rect 4713 8270 4730 8276
rect 4713 8268 4747 8270
rect 4795 8268 4811 8284
rect 4812 8274 5020 8284
rect 5021 8274 5037 8284
rect 5085 8280 5100 8295
rect 5103 8292 5104 8304
rect 5111 8292 5138 8304
rect 5103 8284 5138 8292
rect 5103 8283 5132 8284
rect 4823 8270 5037 8274
rect 4838 8268 5037 8270
rect 5072 8270 5085 8280
rect 5103 8270 5120 8283
rect 5072 8268 5120 8270
rect 4714 8264 4747 8268
rect 4710 8262 4747 8264
rect 4710 8261 4777 8262
rect 4710 8256 4741 8261
rect 4747 8256 4777 8261
rect 4710 8252 4777 8256
rect 4683 8249 4777 8252
rect 4683 8242 4732 8249
rect 4683 8236 4713 8242
rect 4732 8237 4737 8242
rect 4649 8220 4729 8236
rect 4741 8228 4777 8249
rect 4838 8244 5027 8268
rect 5072 8267 5119 8268
rect 5085 8262 5119 8267
rect 4853 8241 5027 8244
rect 4846 8238 5027 8241
rect 5055 8261 5119 8262
rect 4649 8218 4668 8220
rect 4683 8218 4717 8220
rect 4649 8202 4729 8218
rect 4649 8196 4668 8202
rect 4365 8170 4468 8180
rect 4319 8168 4468 8170
rect 4489 8168 4524 8180
rect 4158 8166 4320 8168
rect 4170 8146 4189 8166
rect 4204 8164 4234 8166
rect 4053 8138 4094 8146
rect 4176 8142 4189 8146
rect 4241 8150 4320 8166
rect 4352 8166 4524 8168
rect 4352 8150 4431 8166
rect 4438 8164 4468 8166
rect 4016 8128 4045 8138
rect 4059 8128 4088 8138
rect 4103 8128 4133 8142
rect 4176 8128 4219 8142
rect 4241 8138 4431 8150
rect 4496 8146 4502 8166
rect 4226 8128 4256 8138
rect 4257 8128 4415 8138
rect 4419 8128 4449 8138
rect 4453 8128 4483 8142
rect 4511 8128 4524 8166
rect 4596 8180 4625 8196
rect 4639 8180 4668 8196
rect 4683 8186 4713 8202
rect 4741 8180 4747 8228
rect 4750 8222 4769 8228
rect 4784 8222 4814 8230
rect 4750 8214 4814 8222
rect 4750 8198 4830 8214
rect 4846 8207 4908 8238
rect 4924 8207 4986 8238
rect 5055 8236 5104 8261
rect 5119 8236 5149 8252
rect 5018 8222 5048 8230
rect 5055 8228 5165 8236
rect 5018 8214 5063 8222
rect 4750 8196 4769 8198
rect 4784 8196 4830 8198
rect 4750 8180 4830 8196
rect 4857 8194 4892 8207
rect 4933 8204 4970 8207
rect 4933 8202 4975 8204
rect 4862 8191 4892 8194
rect 4871 8187 4878 8191
rect 4878 8186 4879 8187
rect 4837 8180 4847 8186
rect 4596 8172 4631 8180
rect 4596 8146 4597 8172
rect 4604 8146 4631 8172
rect 4539 8128 4569 8142
rect 4596 8138 4631 8146
rect 4633 8172 4674 8180
rect 4633 8146 4648 8172
rect 4655 8146 4674 8172
rect 4738 8168 4769 8180
rect 4784 8168 4887 8180
rect 4899 8170 4925 8196
rect 4940 8191 4970 8202
rect 5002 8198 5064 8214
rect 5002 8196 5048 8198
rect 5002 8180 5064 8196
rect 5076 8180 5082 8228
rect 5085 8220 5165 8228
rect 5085 8218 5104 8220
rect 5119 8218 5153 8220
rect 5085 8202 5165 8218
rect 5085 8180 5104 8202
rect 5119 8186 5149 8202
rect 5177 8196 5183 8270
rect 5186 8196 5205 8340
rect 5220 8196 5226 8340
rect 5235 8270 5248 8340
rect 5300 8336 5322 8340
rect 5293 8314 5322 8328
rect 5375 8314 5391 8328
rect 5429 8324 5435 8326
rect 5442 8324 5550 8340
rect 5557 8324 5563 8326
rect 5571 8324 5586 8340
rect 5652 8334 5671 8337
rect 5293 8312 5391 8314
rect 5418 8312 5586 8324
rect 5601 8314 5617 8328
rect 5652 8315 5674 8334
rect 5684 8328 5700 8329
rect 5683 8326 5700 8328
rect 5684 8321 5700 8326
rect 5674 8314 5680 8315
rect 5683 8314 5712 8321
rect 5601 8313 5712 8314
rect 5601 8312 5718 8313
rect 5277 8304 5328 8312
rect 5375 8304 5409 8312
rect 5277 8292 5302 8304
rect 5309 8292 5328 8304
rect 5382 8302 5409 8304
rect 5418 8302 5639 8312
rect 5674 8309 5680 8312
rect 5382 8298 5639 8302
rect 5277 8284 5328 8292
rect 5375 8284 5639 8298
rect 5683 8304 5718 8312
rect 5229 8236 5248 8270
rect 5293 8276 5322 8284
rect 5293 8270 5310 8276
rect 5293 8268 5327 8270
rect 5375 8268 5391 8284
rect 5392 8274 5600 8284
rect 5601 8274 5617 8284
rect 5665 8280 5680 8295
rect 5683 8292 5684 8304
rect 5691 8292 5718 8304
rect 5683 8284 5718 8292
rect 5683 8283 5712 8284
rect 5403 8270 5617 8274
rect 5418 8268 5617 8270
rect 5652 8270 5665 8280
rect 5683 8270 5700 8283
rect 5652 8268 5700 8270
rect 5294 8264 5327 8268
rect 5290 8262 5327 8264
rect 5290 8261 5357 8262
rect 5290 8256 5321 8261
rect 5327 8256 5357 8261
rect 5290 8252 5357 8256
rect 5263 8249 5357 8252
rect 5263 8242 5312 8249
rect 5263 8236 5293 8242
rect 5312 8237 5317 8242
rect 5229 8220 5309 8236
rect 5321 8228 5357 8249
rect 5418 8244 5607 8268
rect 5652 8267 5699 8268
rect 5665 8262 5699 8267
rect 5433 8241 5607 8244
rect 5426 8238 5607 8241
rect 5635 8261 5699 8262
rect 5229 8218 5248 8220
rect 5263 8218 5297 8220
rect 5229 8202 5309 8218
rect 5229 8196 5248 8202
rect 4945 8170 5048 8180
rect 4899 8168 5048 8170
rect 5069 8168 5104 8180
rect 4738 8166 4900 8168
rect 4750 8146 4769 8166
rect 4784 8164 4814 8166
rect 4633 8138 4674 8146
rect 4756 8142 4769 8146
rect 4821 8150 4900 8166
rect 4932 8166 5104 8168
rect 4932 8150 5011 8166
rect 5018 8164 5048 8166
rect 4596 8128 4625 8138
rect 4639 8128 4668 8138
rect 4683 8128 4713 8142
rect 4756 8128 4799 8142
rect 4821 8138 5011 8150
rect 5076 8146 5082 8166
rect 4806 8128 4836 8138
rect 4837 8128 4995 8138
rect 4999 8128 5029 8138
rect 5033 8128 5063 8142
rect 5091 8128 5104 8166
rect 5176 8180 5205 8196
rect 5219 8180 5248 8196
rect 5263 8186 5293 8202
rect 5321 8180 5327 8228
rect 5330 8222 5349 8228
rect 5364 8222 5394 8230
rect 5330 8214 5394 8222
rect 5330 8198 5410 8214
rect 5426 8207 5488 8238
rect 5504 8207 5566 8238
rect 5635 8236 5684 8261
rect 5699 8236 5729 8252
rect 5598 8222 5628 8230
rect 5635 8228 5745 8236
rect 5598 8214 5643 8222
rect 5330 8196 5349 8198
rect 5364 8196 5410 8198
rect 5330 8180 5410 8196
rect 5437 8194 5472 8207
rect 5513 8204 5550 8207
rect 5513 8202 5555 8204
rect 5442 8191 5472 8194
rect 5451 8187 5458 8191
rect 5458 8186 5459 8187
rect 5417 8180 5427 8186
rect 5176 8172 5211 8180
rect 5176 8146 5177 8172
rect 5184 8146 5211 8172
rect 5119 8128 5149 8142
rect 5176 8138 5211 8146
rect 5213 8172 5254 8180
rect 5213 8146 5228 8172
rect 5235 8146 5254 8172
rect 5318 8168 5349 8180
rect 5364 8168 5467 8180
rect 5479 8170 5505 8196
rect 5520 8191 5550 8202
rect 5582 8198 5644 8214
rect 5582 8196 5628 8198
rect 5582 8180 5644 8196
rect 5656 8180 5662 8228
rect 5665 8220 5745 8228
rect 5665 8218 5684 8220
rect 5699 8218 5733 8220
rect 5665 8202 5745 8218
rect 5665 8180 5684 8202
rect 5699 8186 5729 8202
rect 5757 8196 5763 8270
rect 5766 8196 5785 8340
rect 5800 8196 5806 8340
rect 5815 8270 5828 8340
rect 5880 8336 5902 8340
rect 5873 8314 5902 8328
rect 5955 8314 5971 8328
rect 6009 8324 6015 8326
rect 6022 8324 6130 8340
rect 6137 8324 6143 8326
rect 6151 8324 6166 8340
rect 6232 8334 6251 8337
rect 5873 8312 5971 8314
rect 5998 8312 6166 8324
rect 6181 8314 6197 8328
rect 6232 8315 6254 8334
rect 6264 8328 6280 8329
rect 6263 8326 6280 8328
rect 6264 8321 6280 8326
rect 6254 8314 6260 8315
rect 6263 8314 6292 8321
rect 6181 8313 6292 8314
rect 6181 8312 6298 8313
rect 5857 8304 5908 8312
rect 5955 8304 5989 8312
rect 5857 8292 5882 8304
rect 5889 8292 5908 8304
rect 5962 8302 5989 8304
rect 5998 8302 6219 8312
rect 6254 8309 6260 8312
rect 5962 8298 6219 8302
rect 5857 8284 5908 8292
rect 5955 8284 6219 8298
rect 6263 8304 6298 8312
rect 5809 8236 5828 8270
rect 5873 8276 5902 8284
rect 5873 8270 5890 8276
rect 5873 8268 5907 8270
rect 5955 8268 5971 8284
rect 5972 8274 6180 8284
rect 6181 8274 6197 8284
rect 6245 8280 6260 8295
rect 6263 8292 6264 8304
rect 6271 8292 6298 8304
rect 6263 8284 6298 8292
rect 6263 8283 6292 8284
rect 5983 8270 6197 8274
rect 5998 8268 6197 8270
rect 6232 8270 6245 8280
rect 6263 8270 6280 8283
rect 6232 8268 6280 8270
rect 5874 8264 5907 8268
rect 5870 8262 5907 8264
rect 5870 8261 5937 8262
rect 5870 8256 5901 8261
rect 5907 8256 5937 8261
rect 5870 8252 5937 8256
rect 5843 8249 5937 8252
rect 5843 8242 5892 8249
rect 5843 8236 5873 8242
rect 5892 8237 5897 8242
rect 5809 8220 5889 8236
rect 5901 8228 5937 8249
rect 5998 8244 6187 8268
rect 6232 8267 6279 8268
rect 6245 8262 6279 8267
rect 6013 8241 6187 8244
rect 6006 8238 6187 8241
rect 6215 8261 6279 8262
rect 5809 8218 5828 8220
rect 5843 8218 5877 8220
rect 5809 8202 5889 8218
rect 5809 8196 5828 8202
rect 5525 8170 5628 8180
rect 5479 8168 5628 8170
rect 5649 8168 5684 8180
rect 5318 8166 5480 8168
rect 5330 8146 5349 8166
rect 5364 8164 5394 8166
rect 5213 8138 5254 8146
rect 5336 8142 5349 8146
rect 5401 8150 5480 8166
rect 5512 8166 5684 8168
rect 5512 8150 5591 8166
rect 5598 8164 5628 8166
rect 5176 8128 5205 8138
rect 5219 8128 5248 8138
rect 5263 8128 5293 8142
rect 5336 8128 5379 8142
rect 5401 8138 5591 8150
rect 5656 8146 5662 8166
rect 5386 8128 5416 8138
rect 5417 8128 5575 8138
rect 5579 8128 5609 8138
rect 5613 8128 5643 8142
rect 5671 8128 5684 8166
rect 5756 8180 5785 8196
rect 5799 8180 5828 8196
rect 5843 8186 5873 8202
rect 5901 8180 5907 8228
rect 5910 8222 5929 8228
rect 5944 8222 5974 8230
rect 5910 8214 5974 8222
rect 5910 8198 5990 8214
rect 6006 8207 6068 8238
rect 6084 8207 6146 8238
rect 6215 8236 6264 8261
rect 6279 8236 6309 8252
rect 6178 8222 6208 8230
rect 6215 8228 6325 8236
rect 6178 8214 6223 8222
rect 5910 8196 5929 8198
rect 5944 8196 5990 8198
rect 5910 8180 5990 8196
rect 6017 8194 6052 8207
rect 6093 8204 6130 8207
rect 6093 8202 6135 8204
rect 6022 8191 6052 8194
rect 6031 8187 6038 8191
rect 6038 8186 6039 8187
rect 5997 8180 6007 8186
rect 5756 8172 5791 8180
rect 5756 8146 5757 8172
rect 5764 8146 5791 8172
rect 5699 8128 5729 8142
rect 5756 8138 5791 8146
rect 5793 8172 5834 8180
rect 5793 8146 5808 8172
rect 5815 8146 5834 8172
rect 5898 8168 5929 8180
rect 5944 8168 6047 8180
rect 6059 8170 6085 8196
rect 6100 8191 6130 8202
rect 6162 8198 6224 8214
rect 6162 8196 6208 8198
rect 6162 8180 6224 8196
rect 6236 8180 6242 8228
rect 6245 8220 6325 8228
rect 6245 8218 6264 8220
rect 6279 8218 6313 8220
rect 6245 8202 6325 8218
rect 6245 8180 6264 8202
rect 6279 8186 6309 8202
rect 6337 8196 6343 8270
rect 6346 8196 6365 8340
rect 6380 8196 6386 8340
rect 6395 8270 6408 8340
rect 6460 8336 6482 8340
rect 6453 8314 6482 8328
rect 6535 8314 6551 8328
rect 6589 8324 6595 8326
rect 6602 8324 6710 8340
rect 6717 8324 6723 8326
rect 6731 8324 6746 8340
rect 6812 8334 6831 8337
rect 6453 8312 6551 8314
rect 6578 8312 6746 8324
rect 6761 8314 6777 8328
rect 6812 8315 6834 8334
rect 6844 8328 6860 8329
rect 6843 8326 6860 8328
rect 6844 8321 6860 8326
rect 6834 8314 6840 8315
rect 6843 8314 6872 8321
rect 6761 8313 6872 8314
rect 6761 8312 6878 8313
rect 6437 8304 6488 8312
rect 6535 8304 6569 8312
rect 6437 8292 6462 8304
rect 6469 8292 6488 8304
rect 6542 8302 6569 8304
rect 6578 8302 6799 8312
rect 6834 8309 6840 8312
rect 6542 8298 6799 8302
rect 6437 8284 6488 8292
rect 6535 8284 6799 8298
rect 6843 8304 6878 8312
rect 6389 8236 6408 8270
rect 6453 8276 6482 8284
rect 6453 8270 6470 8276
rect 6453 8268 6487 8270
rect 6535 8268 6551 8284
rect 6552 8274 6760 8284
rect 6761 8274 6777 8284
rect 6825 8280 6840 8295
rect 6843 8292 6844 8304
rect 6851 8292 6878 8304
rect 6843 8284 6878 8292
rect 6843 8283 6872 8284
rect 6563 8270 6777 8274
rect 6578 8268 6777 8270
rect 6812 8270 6825 8280
rect 6843 8270 6860 8283
rect 6812 8268 6860 8270
rect 6454 8264 6487 8268
rect 6450 8262 6487 8264
rect 6450 8261 6517 8262
rect 6450 8256 6481 8261
rect 6487 8256 6517 8261
rect 6450 8252 6517 8256
rect 6423 8249 6517 8252
rect 6423 8242 6472 8249
rect 6423 8236 6453 8242
rect 6472 8237 6477 8242
rect 6389 8220 6469 8236
rect 6481 8228 6517 8249
rect 6578 8244 6767 8268
rect 6812 8267 6859 8268
rect 6825 8262 6859 8267
rect 6593 8241 6767 8244
rect 6586 8238 6767 8241
rect 6795 8261 6859 8262
rect 6389 8218 6408 8220
rect 6423 8218 6457 8220
rect 6389 8202 6469 8218
rect 6389 8196 6408 8202
rect 6105 8170 6208 8180
rect 6059 8168 6208 8170
rect 6229 8168 6264 8180
rect 5898 8166 6060 8168
rect 5910 8146 5929 8166
rect 5944 8164 5974 8166
rect 5793 8138 5834 8146
rect 5916 8142 5929 8146
rect 5981 8150 6060 8166
rect 6092 8166 6264 8168
rect 6092 8150 6171 8166
rect 6178 8164 6208 8166
rect 5756 8128 5785 8138
rect 5799 8128 5828 8138
rect 5843 8128 5873 8142
rect 5916 8128 5959 8142
rect 5981 8138 6171 8150
rect 6236 8146 6242 8166
rect 5966 8128 5996 8138
rect 5997 8128 6155 8138
rect 6159 8128 6189 8138
rect 6193 8128 6223 8142
rect 6251 8128 6264 8166
rect 6336 8180 6365 8196
rect 6379 8180 6408 8196
rect 6423 8186 6453 8202
rect 6481 8180 6487 8228
rect 6490 8222 6509 8228
rect 6524 8222 6554 8230
rect 6490 8214 6554 8222
rect 6490 8198 6570 8214
rect 6586 8207 6648 8238
rect 6664 8207 6726 8238
rect 6795 8236 6844 8261
rect 6859 8236 6889 8252
rect 6758 8222 6788 8230
rect 6795 8228 6905 8236
rect 6758 8214 6803 8222
rect 6490 8196 6509 8198
rect 6524 8196 6570 8198
rect 6490 8180 6570 8196
rect 6597 8194 6632 8207
rect 6673 8204 6710 8207
rect 6673 8202 6715 8204
rect 6602 8191 6632 8194
rect 6611 8187 6618 8191
rect 6618 8186 6619 8187
rect 6577 8180 6587 8186
rect 6336 8172 6371 8180
rect 6336 8146 6337 8172
rect 6344 8146 6371 8172
rect 6279 8128 6309 8142
rect 6336 8138 6371 8146
rect 6373 8172 6414 8180
rect 6373 8146 6388 8172
rect 6395 8146 6414 8172
rect 6478 8168 6509 8180
rect 6524 8168 6627 8180
rect 6639 8170 6665 8196
rect 6680 8191 6710 8202
rect 6742 8198 6804 8214
rect 6742 8196 6788 8198
rect 6742 8180 6804 8196
rect 6816 8180 6822 8228
rect 6825 8220 6905 8228
rect 6825 8218 6844 8220
rect 6859 8218 6893 8220
rect 6825 8202 6905 8218
rect 6825 8180 6844 8202
rect 6859 8186 6889 8202
rect 6917 8196 6923 8270
rect 6926 8196 6945 8340
rect 6960 8196 6966 8340
rect 6975 8270 6988 8340
rect 7040 8336 7062 8340
rect 7033 8314 7062 8328
rect 7115 8314 7131 8328
rect 7169 8324 7175 8326
rect 7182 8324 7290 8340
rect 7297 8324 7303 8326
rect 7311 8324 7326 8340
rect 7392 8334 7411 8337
rect 7033 8312 7131 8314
rect 7158 8312 7326 8324
rect 7341 8314 7357 8328
rect 7392 8315 7414 8334
rect 7424 8328 7440 8329
rect 7423 8326 7440 8328
rect 7424 8321 7440 8326
rect 7414 8314 7420 8315
rect 7423 8314 7452 8321
rect 7341 8313 7452 8314
rect 7341 8312 7458 8313
rect 7017 8304 7068 8312
rect 7115 8304 7149 8312
rect 7017 8292 7042 8304
rect 7049 8292 7068 8304
rect 7122 8302 7149 8304
rect 7158 8302 7379 8312
rect 7414 8309 7420 8312
rect 7122 8298 7379 8302
rect 7017 8284 7068 8292
rect 7115 8284 7379 8298
rect 7423 8304 7458 8312
rect 6969 8236 6988 8270
rect 7033 8276 7062 8284
rect 7033 8270 7050 8276
rect 7033 8268 7067 8270
rect 7115 8268 7131 8284
rect 7132 8274 7340 8284
rect 7341 8274 7357 8284
rect 7405 8280 7420 8295
rect 7423 8292 7424 8304
rect 7431 8292 7458 8304
rect 7423 8284 7458 8292
rect 7423 8283 7452 8284
rect 7143 8270 7357 8274
rect 7158 8268 7357 8270
rect 7392 8270 7405 8280
rect 7423 8270 7440 8283
rect 7392 8268 7440 8270
rect 7034 8264 7067 8268
rect 7030 8262 7067 8264
rect 7030 8261 7097 8262
rect 7030 8256 7061 8261
rect 7067 8256 7097 8261
rect 7030 8252 7097 8256
rect 7003 8249 7097 8252
rect 7003 8242 7052 8249
rect 7003 8236 7033 8242
rect 7052 8237 7057 8242
rect 6969 8220 7049 8236
rect 7061 8228 7097 8249
rect 7158 8244 7347 8268
rect 7392 8267 7439 8268
rect 7405 8262 7439 8267
rect 7173 8241 7347 8244
rect 7166 8238 7347 8241
rect 7375 8261 7439 8262
rect 6969 8218 6988 8220
rect 7003 8218 7037 8220
rect 6969 8202 7049 8218
rect 6969 8196 6988 8202
rect 6685 8170 6788 8180
rect 6639 8168 6788 8170
rect 6809 8168 6844 8180
rect 6478 8166 6640 8168
rect 6490 8146 6509 8166
rect 6524 8164 6554 8166
rect 6373 8138 6414 8146
rect 6496 8142 6509 8146
rect 6561 8150 6640 8166
rect 6672 8166 6844 8168
rect 6672 8150 6751 8166
rect 6758 8164 6788 8166
rect 6336 8128 6365 8138
rect 6379 8128 6408 8138
rect 6423 8128 6453 8142
rect 6496 8128 6539 8142
rect 6561 8138 6751 8150
rect 6816 8146 6822 8166
rect 6546 8128 6576 8138
rect 6577 8128 6735 8138
rect 6739 8128 6769 8138
rect 6773 8128 6803 8142
rect 6831 8128 6844 8166
rect 6916 8180 6945 8196
rect 6959 8180 6988 8196
rect 7003 8186 7033 8202
rect 7061 8180 7067 8228
rect 7070 8222 7089 8228
rect 7104 8222 7134 8230
rect 7070 8214 7134 8222
rect 7070 8198 7150 8214
rect 7166 8207 7228 8238
rect 7244 8207 7306 8238
rect 7375 8236 7424 8261
rect 7439 8236 7469 8252
rect 7338 8222 7368 8230
rect 7375 8228 7485 8236
rect 7338 8214 7383 8222
rect 7070 8196 7089 8198
rect 7104 8196 7150 8198
rect 7070 8180 7150 8196
rect 7177 8194 7212 8207
rect 7253 8204 7290 8207
rect 7253 8202 7295 8204
rect 7182 8191 7212 8194
rect 7191 8187 7198 8191
rect 7198 8186 7199 8187
rect 7157 8180 7167 8186
rect 6916 8172 6951 8180
rect 6916 8146 6917 8172
rect 6924 8146 6951 8172
rect 6859 8128 6889 8142
rect 6916 8138 6951 8146
rect 6953 8172 6994 8180
rect 6953 8146 6968 8172
rect 6975 8146 6994 8172
rect 7058 8168 7089 8180
rect 7104 8168 7207 8180
rect 7219 8170 7245 8196
rect 7260 8191 7290 8202
rect 7322 8198 7384 8214
rect 7322 8196 7368 8198
rect 7322 8180 7384 8196
rect 7396 8180 7402 8228
rect 7405 8220 7485 8228
rect 7405 8218 7424 8220
rect 7439 8218 7473 8220
rect 7405 8202 7485 8218
rect 7405 8180 7424 8202
rect 7439 8186 7469 8202
rect 7497 8196 7503 8270
rect 7506 8196 7525 8340
rect 7540 8196 7546 8340
rect 7555 8270 7568 8340
rect 7620 8336 7642 8340
rect 7613 8314 7642 8328
rect 7695 8314 7711 8328
rect 7749 8324 7755 8326
rect 7762 8324 7870 8340
rect 7877 8324 7883 8326
rect 7891 8324 7906 8340
rect 7972 8334 7991 8337
rect 7613 8312 7711 8314
rect 7738 8312 7906 8324
rect 7921 8314 7937 8328
rect 7972 8315 7994 8334
rect 8004 8328 8020 8329
rect 8003 8326 8020 8328
rect 8004 8321 8020 8326
rect 7994 8314 8000 8315
rect 8003 8314 8032 8321
rect 7921 8313 8032 8314
rect 7921 8312 8038 8313
rect 7597 8304 7648 8312
rect 7695 8304 7729 8312
rect 7597 8292 7622 8304
rect 7629 8292 7648 8304
rect 7702 8302 7729 8304
rect 7738 8302 7959 8312
rect 7994 8309 8000 8312
rect 7702 8298 7959 8302
rect 7597 8284 7648 8292
rect 7695 8284 7959 8298
rect 8003 8304 8038 8312
rect 7549 8236 7568 8270
rect 7613 8276 7642 8284
rect 7613 8270 7630 8276
rect 7613 8268 7647 8270
rect 7695 8268 7711 8284
rect 7712 8274 7920 8284
rect 7921 8274 7937 8284
rect 7985 8280 8000 8295
rect 8003 8292 8004 8304
rect 8011 8292 8038 8304
rect 8003 8284 8038 8292
rect 8003 8283 8032 8284
rect 7723 8270 7937 8274
rect 7738 8268 7937 8270
rect 7972 8270 7985 8280
rect 8003 8270 8020 8283
rect 7972 8268 8020 8270
rect 7614 8264 7647 8268
rect 7610 8262 7647 8264
rect 7610 8261 7677 8262
rect 7610 8256 7641 8261
rect 7647 8256 7677 8261
rect 7610 8252 7677 8256
rect 7583 8249 7677 8252
rect 7583 8242 7632 8249
rect 7583 8236 7613 8242
rect 7632 8237 7637 8242
rect 7549 8220 7629 8236
rect 7641 8228 7677 8249
rect 7738 8244 7927 8268
rect 7972 8267 8019 8268
rect 7985 8262 8019 8267
rect 7753 8241 7927 8244
rect 7746 8238 7927 8241
rect 7955 8261 8019 8262
rect 7549 8218 7568 8220
rect 7583 8218 7617 8220
rect 7549 8202 7629 8218
rect 7549 8196 7568 8202
rect 7265 8170 7368 8180
rect 7219 8168 7368 8170
rect 7389 8168 7424 8180
rect 7058 8166 7220 8168
rect 7070 8146 7089 8166
rect 7104 8164 7134 8166
rect 6953 8138 6994 8146
rect 7076 8142 7089 8146
rect 7141 8150 7220 8166
rect 7252 8166 7424 8168
rect 7252 8150 7331 8166
rect 7338 8164 7368 8166
rect 6916 8128 6945 8138
rect 6959 8128 6988 8138
rect 7003 8128 7033 8142
rect 7076 8128 7119 8142
rect 7141 8138 7331 8150
rect 7396 8146 7402 8166
rect 7126 8128 7156 8138
rect 7157 8128 7315 8138
rect 7319 8128 7349 8138
rect 7353 8128 7383 8142
rect 7411 8128 7424 8166
rect 7496 8180 7525 8196
rect 7539 8180 7568 8196
rect 7583 8186 7613 8202
rect 7641 8180 7647 8228
rect 7650 8222 7669 8228
rect 7684 8222 7714 8230
rect 7650 8214 7714 8222
rect 7650 8198 7730 8214
rect 7746 8207 7808 8238
rect 7824 8207 7886 8238
rect 7955 8236 8004 8261
rect 8019 8236 8049 8252
rect 7918 8222 7948 8230
rect 7955 8228 8065 8236
rect 7918 8214 7963 8222
rect 7650 8196 7669 8198
rect 7684 8196 7730 8198
rect 7650 8180 7730 8196
rect 7757 8194 7792 8207
rect 7833 8204 7870 8207
rect 7833 8202 7875 8204
rect 7762 8191 7792 8194
rect 7771 8187 7778 8191
rect 7778 8186 7779 8187
rect 7737 8180 7747 8186
rect 7496 8172 7531 8180
rect 7496 8146 7497 8172
rect 7504 8146 7531 8172
rect 7439 8128 7469 8142
rect 7496 8138 7531 8146
rect 7533 8172 7574 8180
rect 7533 8146 7548 8172
rect 7555 8146 7574 8172
rect 7638 8168 7669 8180
rect 7684 8168 7787 8180
rect 7799 8170 7825 8196
rect 7840 8191 7870 8202
rect 7902 8198 7964 8214
rect 7902 8196 7948 8198
rect 7902 8180 7964 8196
rect 7976 8180 7982 8228
rect 7985 8220 8065 8228
rect 7985 8218 8004 8220
rect 8019 8218 8053 8220
rect 7985 8202 8065 8218
rect 7985 8180 8004 8202
rect 8019 8186 8049 8202
rect 8077 8196 8083 8270
rect 8086 8196 8105 8340
rect 8120 8196 8126 8340
rect 8135 8270 8148 8340
rect 8200 8336 8222 8340
rect 8193 8314 8222 8328
rect 8275 8314 8291 8328
rect 8329 8324 8335 8326
rect 8342 8324 8450 8340
rect 8457 8324 8463 8326
rect 8471 8324 8486 8340
rect 8552 8334 8571 8337
rect 8193 8312 8291 8314
rect 8318 8312 8486 8324
rect 8501 8314 8517 8328
rect 8552 8315 8574 8334
rect 8584 8328 8600 8329
rect 8583 8326 8600 8328
rect 8584 8321 8600 8326
rect 8574 8314 8580 8315
rect 8583 8314 8612 8321
rect 8501 8313 8612 8314
rect 8501 8312 8618 8313
rect 8177 8304 8228 8312
rect 8275 8304 8309 8312
rect 8177 8292 8202 8304
rect 8209 8292 8228 8304
rect 8282 8302 8309 8304
rect 8318 8302 8539 8312
rect 8574 8309 8580 8312
rect 8282 8298 8539 8302
rect 8177 8284 8228 8292
rect 8275 8284 8539 8298
rect 8583 8304 8618 8312
rect 8129 8236 8148 8270
rect 8193 8276 8222 8284
rect 8193 8270 8210 8276
rect 8193 8268 8227 8270
rect 8275 8268 8291 8284
rect 8292 8274 8500 8284
rect 8501 8274 8517 8284
rect 8565 8280 8580 8295
rect 8583 8292 8584 8304
rect 8591 8292 8618 8304
rect 8583 8284 8618 8292
rect 8583 8283 8612 8284
rect 8303 8270 8517 8274
rect 8318 8268 8517 8270
rect 8552 8270 8565 8280
rect 8583 8270 8600 8283
rect 8552 8268 8600 8270
rect 8194 8264 8227 8268
rect 8190 8262 8227 8264
rect 8190 8261 8257 8262
rect 8190 8256 8221 8261
rect 8227 8256 8257 8261
rect 8190 8252 8257 8256
rect 8163 8249 8257 8252
rect 8163 8242 8212 8249
rect 8163 8236 8193 8242
rect 8212 8237 8217 8242
rect 8129 8220 8209 8236
rect 8221 8228 8257 8249
rect 8318 8244 8507 8268
rect 8552 8267 8599 8268
rect 8565 8262 8599 8267
rect 8333 8241 8507 8244
rect 8326 8238 8507 8241
rect 8535 8261 8599 8262
rect 8129 8218 8148 8220
rect 8163 8218 8197 8220
rect 8129 8202 8209 8218
rect 8129 8196 8148 8202
rect 7845 8170 7948 8180
rect 7799 8168 7948 8170
rect 7969 8168 8004 8180
rect 7638 8166 7800 8168
rect 7650 8146 7669 8166
rect 7684 8164 7714 8166
rect 7533 8138 7574 8146
rect 7656 8142 7669 8146
rect 7721 8150 7800 8166
rect 7832 8166 8004 8168
rect 7832 8150 7911 8166
rect 7918 8164 7948 8166
rect 7496 8128 7525 8138
rect 7539 8128 7568 8138
rect 7583 8128 7613 8142
rect 7656 8128 7699 8142
rect 7721 8138 7911 8150
rect 7976 8146 7982 8166
rect 7706 8128 7736 8138
rect 7737 8128 7895 8138
rect 7899 8128 7929 8138
rect 7933 8128 7963 8142
rect 7991 8128 8004 8166
rect 8076 8180 8105 8196
rect 8119 8180 8148 8196
rect 8163 8186 8193 8202
rect 8221 8180 8227 8228
rect 8230 8222 8249 8228
rect 8264 8222 8294 8230
rect 8230 8214 8294 8222
rect 8230 8198 8310 8214
rect 8326 8207 8388 8238
rect 8404 8207 8466 8238
rect 8535 8236 8584 8261
rect 8599 8236 8629 8252
rect 8498 8222 8528 8230
rect 8535 8228 8645 8236
rect 8498 8214 8543 8222
rect 8230 8196 8249 8198
rect 8264 8196 8310 8198
rect 8230 8180 8310 8196
rect 8337 8194 8372 8207
rect 8413 8204 8450 8207
rect 8413 8202 8455 8204
rect 8342 8191 8372 8194
rect 8351 8187 8358 8191
rect 8358 8186 8359 8187
rect 8317 8180 8327 8186
rect 8076 8172 8111 8180
rect 8076 8146 8077 8172
rect 8084 8146 8111 8172
rect 8019 8128 8049 8142
rect 8076 8138 8111 8146
rect 8113 8172 8154 8180
rect 8113 8146 8128 8172
rect 8135 8146 8154 8172
rect 8218 8168 8249 8180
rect 8264 8168 8367 8180
rect 8379 8170 8405 8196
rect 8420 8191 8450 8202
rect 8482 8198 8544 8214
rect 8482 8196 8528 8198
rect 8482 8180 8544 8196
rect 8556 8180 8562 8228
rect 8565 8220 8645 8228
rect 8565 8218 8584 8220
rect 8599 8218 8633 8220
rect 8565 8202 8645 8218
rect 8565 8180 8584 8202
rect 8599 8186 8629 8202
rect 8657 8196 8663 8270
rect 8666 8196 8685 8340
rect 8700 8196 8706 8340
rect 8715 8270 8728 8340
rect 8780 8336 8802 8340
rect 8773 8314 8802 8328
rect 8855 8314 8871 8328
rect 8909 8324 8915 8326
rect 8922 8324 9030 8340
rect 9037 8324 9043 8326
rect 9051 8324 9066 8340
rect 9132 8334 9151 8337
rect 8773 8312 8871 8314
rect 8898 8312 9066 8324
rect 9081 8314 9097 8328
rect 9132 8315 9154 8334
rect 9164 8328 9180 8329
rect 9163 8326 9180 8328
rect 9164 8321 9180 8326
rect 9154 8314 9160 8315
rect 9163 8314 9192 8321
rect 9081 8313 9192 8314
rect 9081 8312 9198 8313
rect 8757 8304 8808 8312
rect 8855 8304 8889 8312
rect 8757 8292 8782 8304
rect 8789 8292 8808 8304
rect 8862 8302 8889 8304
rect 8898 8302 9119 8312
rect 9154 8309 9160 8312
rect 8862 8298 9119 8302
rect 8757 8284 8808 8292
rect 8855 8284 9119 8298
rect 9163 8304 9198 8312
rect 8709 8236 8728 8270
rect 8773 8276 8802 8284
rect 8773 8270 8790 8276
rect 8773 8268 8807 8270
rect 8855 8268 8871 8284
rect 8872 8274 9080 8284
rect 9081 8274 9097 8284
rect 9145 8280 9160 8295
rect 9163 8292 9164 8304
rect 9171 8292 9198 8304
rect 9163 8284 9198 8292
rect 9163 8283 9192 8284
rect 8883 8270 9097 8274
rect 8898 8268 9097 8270
rect 9132 8270 9145 8280
rect 9163 8270 9180 8283
rect 9132 8268 9180 8270
rect 8774 8264 8807 8268
rect 8770 8262 8807 8264
rect 8770 8261 8837 8262
rect 8770 8256 8801 8261
rect 8807 8256 8837 8261
rect 8770 8252 8837 8256
rect 8743 8249 8837 8252
rect 8743 8242 8792 8249
rect 8743 8236 8773 8242
rect 8792 8237 8797 8242
rect 8709 8220 8789 8236
rect 8801 8228 8837 8249
rect 8898 8244 9087 8268
rect 9132 8267 9179 8268
rect 9145 8262 9179 8267
rect 8913 8241 9087 8244
rect 8906 8238 9087 8241
rect 9115 8261 9179 8262
rect 8709 8218 8728 8220
rect 8743 8218 8777 8220
rect 8709 8202 8789 8218
rect 8709 8196 8728 8202
rect 8425 8170 8528 8180
rect 8379 8168 8528 8170
rect 8549 8168 8584 8180
rect 8218 8166 8380 8168
rect 8230 8146 8249 8166
rect 8264 8164 8294 8166
rect 8113 8138 8154 8146
rect 8236 8142 8249 8146
rect 8301 8150 8380 8166
rect 8412 8166 8584 8168
rect 8412 8150 8491 8166
rect 8498 8164 8528 8166
rect 8076 8128 8105 8138
rect 8119 8128 8148 8138
rect 8163 8128 8193 8142
rect 8236 8128 8279 8142
rect 8301 8138 8491 8150
rect 8556 8146 8562 8166
rect 8286 8128 8316 8138
rect 8317 8128 8475 8138
rect 8479 8128 8509 8138
rect 8513 8128 8543 8142
rect 8571 8128 8584 8166
rect 8656 8180 8685 8196
rect 8699 8180 8728 8196
rect 8743 8186 8773 8202
rect 8801 8180 8807 8228
rect 8810 8222 8829 8228
rect 8844 8222 8874 8230
rect 8810 8214 8874 8222
rect 8810 8198 8890 8214
rect 8906 8207 8968 8238
rect 8984 8207 9046 8238
rect 9115 8236 9164 8261
rect 9179 8236 9209 8252
rect 9078 8222 9108 8230
rect 9115 8228 9225 8236
rect 9078 8214 9123 8222
rect 8810 8196 8829 8198
rect 8844 8196 8890 8198
rect 8810 8180 8890 8196
rect 8917 8194 8952 8207
rect 8993 8204 9030 8207
rect 8993 8202 9035 8204
rect 8922 8191 8952 8194
rect 8931 8187 8938 8191
rect 8938 8186 8939 8187
rect 8897 8180 8907 8186
rect 8656 8172 8691 8180
rect 8656 8146 8657 8172
rect 8664 8146 8691 8172
rect 8599 8128 8629 8142
rect 8656 8138 8691 8146
rect 8693 8172 8734 8180
rect 8693 8146 8708 8172
rect 8715 8146 8734 8172
rect 8798 8168 8829 8180
rect 8844 8168 8947 8180
rect 8959 8170 8985 8196
rect 9000 8191 9030 8202
rect 9062 8198 9124 8214
rect 9062 8196 9108 8198
rect 9062 8180 9124 8196
rect 9136 8180 9142 8228
rect 9145 8220 9225 8228
rect 9145 8218 9164 8220
rect 9179 8218 9213 8220
rect 9145 8202 9225 8218
rect 9145 8180 9164 8202
rect 9179 8186 9209 8202
rect 9237 8196 9243 8270
rect 9246 8196 9265 8340
rect 9280 8196 9286 8340
rect 9295 8270 9308 8340
rect 9360 8336 9382 8340
rect 9353 8314 9382 8328
rect 9435 8314 9451 8328
rect 9489 8324 9495 8326
rect 9502 8324 9610 8340
rect 9617 8324 9623 8326
rect 9631 8324 9646 8340
rect 9712 8334 9731 8337
rect 9353 8312 9451 8314
rect 9478 8312 9646 8324
rect 9661 8314 9677 8328
rect 9712 8315 9734 8334
rect 9744 8328 9760 8329
rect 9743 8326 9760 8328
rect 9744 8321 9760 8326
rect 9734 8314 9740 8315
rect 9743 8314 9772 8321
rect 9661 8313 9772 8314
rect 9661 8312 9778 8313
rect 9337 8304 9388 8312
rect 9435 8304 9469 8312
rect 9337 8292 9362 8304
rect 9369 8292 9388 8304
rect 9442 8302 9469 8304
rect 9478 8302 9699 8312
rect 9734 8309 9740 8312
rect 9442 8298 9699 8302
rect 9337 8284 9388 8292
rect 9435 8284 9699 8298
rect 9743 8304 9778 8312
rect 9289 8236 9308 8270
rect 9353 8276 9382 8284
rect 9353 8270 9370 8276
rect 9353 8268 9387 8270
rect 9435 8268 9451 8284
rect 9452 8274 9660 8284
rect 9661 8274 9677 8284
rect 9725 8280 9740 8295
rect 9743 8292 9744 8304
rect 9751 8292 9778 8304
rect 9743 8284 9778 8292
rect 9743 8283 9772 8284
rect 9463 8270 9677 8274
rect 9478 8268 9677 8270
rect 9712 8270 9725 8280
rect 9743 8270 9760 8283
rect 9712 8268 9760 8270
rect 9354 8264 9387 8268
rect 9350 8262 9387 8264
rect 9350 8261 9417 8262
rect 9350 8256 9381 8261
rect 9387 8256 9417 8261
rect 9350 8252 9417 8256
rect 9323 8249 9417 8252
rect 9323 8242 9372 8249
rect 9323 8236 9353 8242
rect 9372 8237 9377 8242
rect 9289 8220 9369 8236
rect 9381 8228 9417 8249
rect 9478 8244 9667 8268
rect 9712 8267 9759 8268
rect 9725 8262 9759 8267
rect 9493 8241 9667 8244
rect 9486 8238 9667 8241
rect 9695 8261 9759 8262
rect 9289 8218 9308 8220
rect 9323 8218 9357 8220
rect 9289 8202 9369 8218
rect 9289 8196 9308 8202
rect 9005 8170 9108 8180
rect 8959 8168 9108 8170
rect 9129 8168 9164 8180
rect 8798 8166 8960 8168
rect 8810 8146 8829 8166
rect 8844 8164 8874 8166
rect 8693 8138 8734 8146
rect 8816 8142 8829 8146
rect 8881 8150 8960 8166
rect 8992 8166 9164 8168
rect 8992 8150 9071 8166
rect 9078 8164 9108 8166
rect 8656 8128 8685 8138
rect 8699 8128 8728 8138
rect 8743 8128 8773 8142
rect 8816 8128 8859 8142
rect 8881 8138 9071 8150
rect 9136 8146 9142 8166
rect 8866 8128 8896 8138
rect 8897 8128 9055 8138
rect 9059 8128 9089 8138
rect 9093 8128 9123 8142
rect 9151 8128 9164 8166
rect 9236 8180 9265 8196
rect 9279 8180 9308 8196
rect 9323 8186 9353 8202
rect 9381 8180 9387 8228
rect 9390 8222 9409 8228
rect 9424 8222 9454 8230
rect 9390 8214 9454 8222
rect 9390 8198 9470 8214
rect 9486 8207 9548 8238
rect 9564 8207 9626 8238
rect 9695 8236 9744 8261
rect 9759 8236 9789 8252
rect 9658 8222 9688 8230
rect 9695 8228 9805 8236
rect 9658 8214 9703 8222
rect 9390 8196 9409 8198
rect 9424 8196 9470 8198
rect 9390 8180 9470 8196
rect 9497 8194 9532 8207
rect 9573 8204 9610 8207
rect 9573 8202 9615 8204
rect 9502 8191 9532 8194
rect 9511 8187 9518 8191
rect 9518 8186 9519 8187
rect 9477 8180 9487 8186
rect 9236 8172 9271 8180
rect 9236 8146 9237 8172
rect 9244 8146 9271 8172
rect 9179 8128 9209 8142
rect 9236 8138 9271 8146
rect 9273 8172 9314 8180
rect 9273 8146 9288 8172
rect 9295 8146 9314 8172
rect 9378 8168 9409 8180
rect 9424 8168 9527 8180
rect 9539 8170 9565 8196
rect 9580 8191 9610 8202
rect 9642 8198 9704 8214
rect 9642 8196 9688 8198
rect 9642 8180 9704 8196
rect 9716 8180 9722 8228
rect 9725 8220 9805 8228
rect 9725 8218 9744 8220
rect 9759 8218 9793 8220
rect 9725 8202 9805 8218
rect 9725 8180 9744 8202
rect 9759 8186 9789 8202
rect 9817 8196 9823 8270
rect 9826 8196 9845 8340
rect 9860 8196 9866 8340
rect 9875 8270 9888 8340
rect 9940 8336 9962 8340
rect 9933 8314 9962 8328
rect 10015 8314 10031 8328
rect 10069 8324 10075 8326
rect 10082 8324 10190 8340
rect 10197 8324 10203 8326
rect 10211 8324 10226 8340
rect 10292 8334 10311 8337
rect 9933 8312 10031 8314
rect 10058 8312 10226 8324
rect 10241 8314 10257 8328
rect 10292 8315 10314 8334
rect 10324 8328 10340 8329
rect 10323 8326 10340 8328
rect 10324 8321 10340 8326
rect 10314 8314 10320 8315
rect 10323 8314 10352 8321
rect 10241 8313 10352 8314
rect 10241 8312 10358 8313
rect 9917 8304 9968 8312
rect 10015 8304 10049 8312
rect 9917 8292 9942 8304
rect 9949 8292 9968 8304
rect 10022 8302 10049 8304
rect 10058 8302 10279 8312
rect 10314 8309 10320 8312
rect 10022 8298 10279 8302
rect 9917 8284 9968 8292
rect 10015 8284 10279 8298
rect 10323 8304 10358 8312
rect 9869 8236 9888 8270
rect 9933 8276 9962 8284
rect 9933 8270 9950 8276
rect 9933 8268 9967 8270
rect 10015 8268 10031 8284
rect 10032 8274 10240 8284
rect 10241 8274 10257 8284
rect 10305 8280 10320 8295
rect 10323 8292 10324 8304
rect 10331 8292 10358 8304
rect 10323 8284 10358 8292
rect 10323 8283 10352 8284
rect 10043 8270 10257 8274
rect 10058 8268 10257 8270
rect 10292 8270 10305 8280
rect 10323 8270 10340 8283
rect 10292 8268 10340 8270
rect 9934 8264 9967 8268
rect 9930 8262 9967 8264
rect 9930 8261 9997 8262
rect 9930 8256 9961 8261
rect 9967 8256 9997 8261
rect 9930 8252 9997 8256
rect 9903 8249 9997 8252
rect 9903 8242 9952 8249
rect 9903 8236 9933 8242
rect 9952 8237 9957 8242
rect 9869 8220 9949 8236
rect 9961 8228 9997 8249
rect 10058 8244 10247 8268
rect 10292 8267 10339 8268
rect 10305 8262 10339 8267
rect 10073 8241 10247 8244
rect 10066 8238 10247 8241
rect 10275 8261 10339 8262
rect 9869 8218 9888 8220
rect 9903 8218 9937 8220
rect 9869 8202 9949 8218
rect 9869 8196 9888 8202
rect 9585 8170 9688 8180
rect 9539 8168 9688 8170
rect 9709 8168 9744 8180
rect 9378 8166 9540 8168
rect 9390 8146 9409 8166
rect 9424 8164 9454 8166
rect 9273 8138 9314 8146
rect 9396 8142 9409 8146
rect 9461 8150 9540 8166
rect 9572 8166 9744 8168
rect 9572 8150 9651 8166
rect 9658 8164 9688 8166
rect 9236 8128 9265 8138
rect 9279 8128 9308 8138
rect 9323 8128 9353 8142
rect 9396 8128 9439 8142
rect 9461 8138 9651 8150
rect 9716 8146 9722 8166
rect 9446 8128 9476 8138
rect 9477 8128 9635 8138
rect 9639 8128 9669 8138
rect 9673 8128 9703 8142
rect 9731 8128 9744 8166
rect 9816 8180 9845 8196
rect 9859 8180 9888 8196
rect 9903 8186 9933 8202
rect 9961 8180 9967 8228
rect 9970 8222 9989 8228
rect 10004 8222 10034 8230
rect 9970 8214 10034 8222
rect 9970 8198 10050 8214
rect 10066 8207 10128 8238
rect 10144 8207 10206 8238
rect 10275 8236 10324 8261
rect 10339 8236 10369 8252
rect 10238 8222 10268 8230
rect 10275 8228 10385 8236
rect 10238 8214 10283 8222
rect 9970 8196 9989 8198
rect 10004 8196 10050 8198
rect 9970 8180 10050 8196
rect 10077 8194 10112 8207
rect 10153 8204 10190 8207
rect 10153 8202 10195 8204
rect 10082 8191 10112 8194
rect 10091 8187 10098 8191
rect 10098 8186 10099 8187
rect 10057 8180 10067 8186
rect 9816 8172 9851 8180
rect 9816 8146 9817 8172
rect 9824 8146 9851 8172
rect 9759 8128 9789 8142
rect 9816 8138 9851 8146
rect 9853 8172 9894 8180
rect 9853 8146 9868 8172
rect 9875 8146 9894 8172
rect 9958 8168 9989 8180
rect 10004 8168 10107 8180
rect 10119 8170 10145 8196
rect 10160 8191 10190 8202
rect 10222 8198 10284 8214
rect 10222 8196 10268 8198
rect 10222 8180 10284 8196
rect 10296 8180 10302 8228
rect 10305 8220 10385 8228
rect 10305 8218 10324 8220
rect 10339 8218 10373 8220
rect 10305 8202 10385 8218
rect 10305 8180 10324 8202
rect 10339 8186 10369 8202
rect 10397 8196 10403 8270
rect 10406 8196 10425 8340
rect 10440 8196 10446 8340
rect 10455 8270 10468 8340
rect 10520 8336 10542 8340
rect 10513 8314 10542 8328
rect 10595 8314 10611 8328
rect 10649 8324 10655 8326
rect 10662 8324 10770 8340
rect 10777 8324 10783 8326
rect 10791 8324 10806 8340
rect 10872 8334 10891 8337
rect 10513 8312 10611 8314
rect 10638 8312 10806 8324
rect 10821 8314 10837 8328
rect 10872 8315 10894 8334
rect 10904 8328 10920 8329
rect 10903 8326 10920 8328
rect 10904 8321 10920 8326
rect 10894 8314 10900 8315
rect 10903 8314 10932 8321
rect 10821 8313 10932 8314
rect 10821 8312 10938 8313
rect 10497 8304 10548 8312
rect 10595 8304 10629 8312
rect 10497 8292 10522 8304
rect 10529 8292 10548 8304
rect 10602 8302 10629 8304
rect 10638 8302 10859 8312
rect 10894 8309 10900 8312
rect 10602 8298 10859 8302
rect 10497 8284 10548 8292
rect 10595 8284 10859 8298
rect 10903 8304 10938 8312
rect 10449 8236 10468 8270
rect 10513 8276 10542 8284
rect 10513 8270 10530 8276
rect 10513 8268 10547 8270
rect 10595 8268 10611 8284
rect 10612 8274 10820 8284
rect 10821 8274 10837 8284
rect 10885 8280 10900 8295
rect 10903 8292 10904 8304
rect 10911 8292 10938 8304
rect 10903 8284 10938 8292
rect 10903 8283 10932 8284
rect 10623 8270 10837 8274
rect 10638 8268 10837 8270
rect 10872 8270 10885 8280
rect 10903 8270 10920 8283
rect 10872 8268 10920 8270
rect 10514 8264 10547 8268
rect 10510 8262 10547 8264
rect 10510 8261 10577 8262
rect 10510 8256 10541 8261
rect 10547 8256 10577 8261
rect 10510 8252 10577 8256
rect 10483 8249 10577 8252
rect 10483 8242 10532 8249
rect 10483 8236 10513 8242
rect 10532 8237 10537 8242
rect 10449 8220 10529 8236
rect 10541 8228 10577 8249
rect 10638 8244 10827 8268
rect 10872 8267 10919 8268
rect 10885 8262 10919 8267
rect 10653 8241 10827 8244
rect 10646 8238 10827 8241
rect 10855 8261 10919 8262
rect 10449 8218 10468 8220
rect 10483 8218 10517 8220
rect 10449 8202 10529 8218
rect 10449 8196 10468 8202
rect 10165 8170 10268 8180
rect 10119 8168 10268 8170
rect 10289 8168 10324 8180
rect 9958 8166 10120 8168
rect 9970 8146 9989 8166
rect 10004 8164 10034 8166
rect 9853 8138 9894 8146
rect 9976 8142 9989 8146
rect 10041 8150 10120 8166
rect 10152 8166 10324 8168
rect 10152 8150 10231 8166
rect 10238 8164 10268 8166
rect 9816 8128 9845 8138
rect 9859 8128 9888 8138
rect 9903 8128 9933 8142
rect 9976 8128 10019 8142
rect 10041 8138 10231 8150
rect 10296 8146 10302 8166
rect 10026 8128 10056 8138
rect 10057 8128 10215 8138
rect 10219 8128 10249 8138
rect 10253 8128 10283 8142
rect 10311 8128 10324 8166
rect 10396 8180 10425 8196
rect 10439 8180 10468 8196
rect 10483 8186 10513 8202
rect 10541 8180 10547 8228
rect 10550 8222 10569 8228
rect 10584 8222 10614 8230
rect 10550 8214 10614 8222
rect 10550 8198 10630 8214
rect 10646 8207 10708 8238
rect 10724 8207 10786 8238
rect 10855 8236 10904 8261
rect 10919 8236 10949 8252
rect 10818 8222 10848 8230
rect 10855 8228 10965 8236
rect 10818 8214 10863 8222
rect 10550 8196 10569 8198
rect 10584 8196 10630 8198
rect 10550 8180 10630 8196
rect 10657 8194 10692 8207
rect 10733 8204 10770 8207
rect 10733 8202 10775 8204
rect 10662 8191 10692 8194
rect 10671 8187 10678 8191
rect 10678 8186 10679 8187
rect 10637 8180 10647 8186
rect 10396 8172 10431 8180
rect 10396 8146 10397 8172
rect 10404 8146 10431 8172
rect 10339 8128 10369 8142
rect 10396 8138 10431 8146
rect 10433 8172 10474 8180
rect 10433 8146 10448 8172
rect 10455 8146 10474 8172
rect 10538 8168 10569 8180
rect 10584 8168 10687 8180
rect 10699 8170 10725 8196
rect 10740 8191 10770 8202
rect 10802 8198 10864 8214
rect 10802 8196 10848 8198
rect 10802 8180 10864 8196
rect 10876 8180 10882 8228
rect 10885 8220 10965 8228
rect 10885 8218 10904 8220
rect 10919 8218 10953 8220
rect 10885 8202 10965 8218
rect 10885 8180 10904 8202
rect 10919 8186 10949 8202
rect 10977 8196 10983 8270
rect 10986 8196 11005 8340
rect 11020 8196 11026 8340
rect 11035 8270 11048 8340
rect 11100 8336 11122 8340
rect 11093 8314 11122 8328
rect 11175 8314 11191 8328
rect 11229 8324 11235 8326
rect 11242 8324 11350 8340
rect 11357 8324 11363 8326
rect 11371 8324 11386 8340
rect 11452 8334 11471 8337
rect 11093 8312 11191 8314
rect 11218 8312 11386 8324
rect 11401 8314 11417 8328
rect 11452 8315 11474 8334
rect 11484 8328 11500 8329
rect 11483 8326 11500 8328
rect 11484 8321 11500 8326
rect 11474 8314 11480 8315
rect 11483 8314 11512 8321
rect 11401 8313 11512 8314
rect 11401 8312 11518 8313
rect 11077 8304 11128 8312
rect 11175 8304 11209 8312
rect 11077 8292 11102 8304
rect 11109 8292 11128 8304
rect 11182 8302 11209 8304
rect 11218 8302 11439 8312
rect 11474 8309 11480 8312
rect 11182 8298 11439 8302
rect 11077 8284 11128 8292
rect 11175 8284 11439 8298
rect 11483 8304 11518 8312
rect 11029 8236 11048 8270
rect 11093 8276 11122 8284
rect 11093 8270 11110 8276
rect 11093 8268 11127 8270
rect 11175 8268 11191 8284
rect 11192 8274 11400 8284
rect 11401 8274 11417 8284
rect 11465 8280 11480 8295
rect 11483 8292 11484 8304
rect 11491 8292 11518 8304
rect 11483 8284 11518 8292
rect 11483 8283 11512 8284
rect 11203 8270 11417 8274
rect 11218 8268 11417 8270
rect 11452 8270 11465 8280
rect 11483 8270 11500 8283
rect 11452 8268 11500 8270
rect 11094 8264 11127 8268
rect 11090 8262 11127 8264
rect 11090 8261 11157 8262
rect 11090 8256 11121 8261
rect 11127 8256 11157 8261
rect 11090 8252 11157 8256
rect 11063 8249 11157 8252
rect 11063 8242 11112 8249
rect 11063 8236 11093 8242
rect 11112 8237 11117 8242
rect 11029 8220 11109 8236
rect 11121 8228 11157 8249
rect 11218 8244 11407 8268
rect 11452 8267 11499 8268
rect 11465 8262 11499 8267
rect 11233 8241 11407 8244
rect 11226 8238 11407 8241
rect 11435 8261 11499 8262
rect 11029 8218 11048 8220
rect 11063 8218 11097 8220
rect 11029 8202 11109 8218
rect 11029 8196 11048 8202
rect 10745 8170 10848 8180
rect 10699 8168 10848 8170
rect 10869 8168 10904 8180
rect 10538 8166 10700 8168
rect 10550 8146 10569 8166
rect 10584 8164 10614 8166
rect 10433 8138 10474 8146
rect 10556 8142 10569 8146
rect 10621 8150 10700 8166
rect 10732 8166 10904 8168
rect 10732 8150 10811 8166
rect 10818 8164 10848 8166
rect 10396 8128 10425 8138
rect 10439 8128 10468 8138
rect 10483 8128 10513 8142
rect 10556 8128 10599 8142
rect 10621 8138 10811 8150
rect 10876 8146 10882 8166
rect 10606 8128 10636 8138
rect 10637 8128 10795 8138
rect 10799 8128 10829 8138
rect 10833 8128 10863 8142
rect 10891 8128 10904 8166
rect 10976 8180 11005 8196
rect 11019 8180 11048 8196
rect 11063 8186 11093 8202
rect 11121 8180 11127 8228
rect 11130 8222 11149 8228
rect 11164 8222 11194 8230
rect 11130 8214 11194 8222
rect 11130 8198 11210 8214
rect 11226 8207 11288 8238
rect 11304 8207 11366 8238
rect 11435 8236 11484 8261
rect 11499 8236 11529 8252
rect 11398 8222 11428 8230
rect 11435 8228 11545 8236
rect 11398 8214 11443 8222
rect 11130 8196 11149 8198
rect 11164 8196 11210 8198
rect 11130 8180 11210 8196
rect 11237 8194 11272 8207
rect 11313 8204 11350 8207
rect 11313 8202 11355 8204
rect 11242 8191 11272 8194
rect 11251 8187 11258 8191
rect 11258 8186 11259 8187
rect 11217 8180 11227 8186
rect 10976 8172 11011 8180
rect 10976 8146 10977 8172
rect 10984 8146 11011 8172
rect 10919 8128 10949 8142
rect 10976 8138 11011 8146
rect 11013 8172 11054 8180
rect 11013 8146 11028 8172
rect 11035 8146 11054 8172
rect 11118 8168 11149 8180
rect 11164 8168 11267 8180
rect 11279 8170 11305 8196
rect 11320 8191 11350 8202
rect 11382 8198 11444 8214
rect 11382 8196 11428 8198
rect 11382 8180 11444 8196
rect 11456 8180 11462 8228
rect 11465 8220 11545 8228
rect 11465 8218 11484 8220
rect 11499 8218 11533 8220
rect 11465 8202 11545 8218
rect 11465 8180 11484 8202
rect 11499 8186 11529 8202
rect 11557 8196 11563 8270
rect 11566 8196 11585 8340
rect 11600 8196 11606 8340
rect 11615 8270 11628 8340
rect 11680 8336 11702 8340
rect 11673 8314 11702 8328
rect 11755 8314 11771 8328
rect 11809 8324 11815 8326
rect 11822 8324 11930 8340
rect 11937 8324 11943 8326
rect 11951 8324 11966 8340
rect 12032 8334 12051 8337
rect 11673 8312 11771 8314
rect 11798 8312 11966 8324
rect 11981 8314 11997 8328
rect 12032 8315 12054 8334
rect 12064 8328 12080 8329
rect 12063 8326 12080 8328
rect 12064 8321 12080 8326
rect 12054 8314 12060 8315
rect 12063 8314 12092 8321
rect 11981 8313 12092 8314
rect 11981 8312 12098 8313
rect 11657 8304 11708 8312
rect 11755 8304 11789 8312
rect 11657 8292 11682 8304
rect 11689 8292 11708 8304
rect 11762 8302 11789 8304
rect 11798 8302 12019 8312
rect 12054 8309 12060 8312
rect 11762 8298 12019 8302
rect 11657 8284 11708 8292
rect 11755 8284 12019 8298
rect 12063 8304 12098 8312
rect 11609 8236 11628 8270
rect 11673 8276 11702 8284
rect 11673 8270 11690 8276
rect 11673 8268 11707 8270
rect 11755 8268 11771 8284
rect 11772 8274 11980 8284
rect 11981 8274 11997 8284
rect 12045 8280 12060 8295
rect 12063 8292 12064 8304
rect 12071 8292 12098 8304
rect 12063 8284 12098 8292
rect 12063 8283 12092 8284
rect 11783 8270 11997 8274
rect 11798 8268 11997 8270
rect 12032 8270 12045 8280
rect 12063 8270 12080 8283
rect 12032 8268 12080 8270
rect 11674 8264 11707 8268
rect 11670 8262 11707 8264
rect 11670 8261 11737 8262
rect 11670 8256 11701 8261
rect 11707 8256 11737 8261
rect 11670 8252 11737 8256
rect 11643 8249 11737 8252
rect 11643 8242 11692 8249
rect 11643 8236 11673 8242
rect 11692 8237 11697 8242
rect 11609 8220 11689 8236
rect 11701 8228 11737 8249
rect 11798 8244 11987 8268
rect 12032 8267 12079 8268
rect 12045 8262 12079 8267
rect 11813 8241 11987 8244
rect 11806 8238 11987 8241
rect 12015 8261 12079 8262
rect 11609 8218 11628 8220
rect 11643 8218 11677 8220
rect 11609 8202 11689 8218
rect 11609 8196 11628 8202
rect 11325 8170 11428 8180
rect 11279 8168 11428 8170
rect 11449 8168 11484 8180
rect 11118 8166 11280 8168
rect 11130 8146 11149 8166
rect 11164 8164 11194 8166
rect 11013 8138 11054 8146
rect 11136 8142 11149 8146
rect 11201 8150 11280 8166
rect 11312 8166 11484 8168
rect 11312 8150 11391 8166
rect 11398 8164 11428 8166
rect 10976 8128 11005 8138
rect 11019 8128 11048 8138
rect 11063 8128 11093 8142
rect 11136 8128 11179 8142
rect 11201 8138 11391 8150
rect 11456 8146 11462 8166
rect 11186 8128 11216 8138
rect 11217 8128 11375 8138
rect 11379 8128 11409 8138
rect 11413 8128 11443 8142
rect 11471 8128 11484 8166
rect 11556 8180 11585 8196
rect 11599 8180 11628 8196
rect 11643 8186 11673 8202
rect 11701 8180 11707 8228
rect 11710 8222 11729 8228
rect 11744 8222 11774 8230
rect 11710 8214 11774 8222
rect 11710 8198 11790 8214
rect 11806 8207 11868 8238
rect 11884 8207 11946 8238
rect 12015 8236 12064 8261
rect 12079 8236 12109 8252
rect 11978 8222 12008 8230
rect 12015 8228 12125 8236
rect 11978 8214 12023 8222
rect 11710 8196 11729 8198
rect 11744 8196 11790 8198
rect 11710 8180 11790 8196
rect 11817 8194 11852 8207
rect 11893 8204 11930 8207
rect 11893 8202 11935 8204
rect 11822 8191 11852 8194
rect 11831 8187 11838 8191
rect 11838 8186 11839 8187
rect 11797 8180 11807 8186
rect 11556 8172 11591 8180
rect 11556 8146 11557 8172
rect 11564 8146 11591 8172
rect 11499 8128 11529 8142
rect 11556 8138 11591 8146
rect 11593 8172 11634 8180
rect 11593 8146 11608 8172
rect 11615 8146 11634 8172
rect 11698 8168 11729 8180
rect 11744 8168 11847 8180
rect 11859 8170 11885 8196
rect 11900 8191 11930 8202
rect 11962 8198 12024 8214
rect 11962 8196 12008 8198
rect 11962 8180 12024 8196
rect 12036 8180 12042 8228
rect 12045 8220 12125 8228
rect 12045 8218 12064 8220
rect 12079 8218 12113 8220
rect 12045 8202 12125 8218
rect 12045 8180 12064 8202
rect 12079 8186 12109 8202
rect 12137 8196 12143 8270
rect 12146 8196 12165 8340
rect 12180 8196 12186 8340
rect 12195 8270 12208 8340
rect 12260 8336 12282 8340
rect 12253 8314 12282 8328
rect 12335 8314 12351 8328
rect 12389 8324 12395 8326
rect 12402 8324 12510 8340
rect 12517 8324 12523 8326
rect 12531 8324 12546 8340
rect 12612 8334 12631 8337
rect 12253 8312 12351 8314
rect 12378 8312 12546 8324
rect 12561 8314 12577 8328
rect 12612 8315 12634 8334
rect 12644 8328 12660 8329
rect 12643 8326 12660 8328
rect 12644 8321 12660 8326
rect 12634 8314 12640 8315
rect 12643 8314 12672 8321
rect 12561 8313 12672 8314
rect 12561 8312 12678 8313
rect 12237 8304 12288 8312
rect 12335 8304 12369 8312
rect 12237 8292 12262 8304
rect 12269 8292 12288 8304
rect 12342 8302 12369 8304
rect 12378 8302 12599 8312
rect 12634 8309 12640 8312
rect 12342 8298 12599 8302
rect 12237 8284 12288 8292
rect 12335 8284 12599 8298
rect 12643 8304 12678 8312
rect 12189 8236 12208 8270
rect 12253 8276 12282 8284
rect 12253 8270 12270 8276
rect 12253 8268 12287 8270
rect 12335 8268 12351 8284
rect 12352 8274 12560 8284
rect 12561 8274 12577 8284
rect 12625 8280 12640 8295
rect 12643 8292 12644 8304
rect 12651 8292 12678 8304
rect 12643 8284 12678 8292
rect 12643 8283 12672 8284
rect 12363 8270 12577 8274
rect 12378 8268 12577 8270
rect 12612 8270 12625 8280
rect 12643 8270 12660 8283
rect 12612 8268 12660 8270
rect 12254 8264 12287 8268
rect 12250 8262 12287 8264
rect 12250 8261 12317 8262
rect 12250 8256 12281 8261
rect 12287 8256 12317 8261
rect 12250 8252 12317 8256
rect 12223 8249 12317 8252
rect 12223 8242 12272 8249
rect 12223 8236 12253 8242
rect 12272 8237 12277 8242
rect 12189 8220 12269 8236
rect 12281 8228 12317 8249
rect 12378 8244 12567 8268
rect 12612 8267 12659 8268
rect 12625 8262 12659 8267
rect 12393 8241 12567 8244
rect 12386 8238 12567 8241
rect 12595 8261 12659 8262
rect 12189 8218 12208 8220
rect 12223 8218 12257 8220
rect 12189 8202 12269 8218
rect 12189 8196 12208 8202
rect 11905 8170 12008 8180
rect 11859 8168 12008 8170
rect 12029 8168 12064 8180
rect 11698 8166 11860 8168
rect 11710 8146 11729 8166
rect 11744 8164 11774 8166
rect 11593 8138 11634 8146
rect 11716 8142 11729 8146
rect 11781 8150 11860 8166
rect 11892 8166 12064 8168
rect 11892 8150 11971 8166
rect 11978 8164 12008 8166
rect 11556 8128 11585 8138
rect 11599 8128 11628 8138
rect 11643 8128 11673 8142
rect 11716 8128 11759 8142
rect 11781 8138 11971 8150
rect 12036 8146 12042 8166
rect 11766 8128 11796 8138
rect 11797 8128 11955 8138
rect 11959 8128 11989 8138
rect 11993 8128 12023 8142
rect 12051 8128 12064 8166
rect 12136 8180 12165 8196
rect 12179 8180 12208 8196
rect 12223 8186 12253 8202
rect 12281 8180 12287 8228
rect 12290 8222 12309 8228
rect 12324 8222 12354 8230
rect 12290 8214 12354 8222
rect 12290 8198 12370 8214
rect 12386 8207 12448 8238
rect 12464 8207 12526 8238
rect 12595 8236 12644 8261
rect 12659 8236 12689 8252
rect 12558 8222 12588 8230
rect 12595 8228 12705 8236
rect 12558 8214 12603 8222
rect 12290 8196 12309 8198
rect 12324 8196 12370 8198
rect 12290 8180 12370 8196
rect 12397 8194 12432 8207
rect 12473 8204 12510 8207
rect 12473 8202 12515 8204
rect 12402 8191 12432 8194
rect 12411 8187 12418 8191
rect 12418 8186 12419 8187
rect 12377 8180 12387 8186
rect 12136 8172 12171 8180
rect 12136 8146 12137 8172
rect 12144 8146 12171 8172
rect 12079 8128 12109 8142
rect 12136 8138 12171 8146
rect 12173 8172 12214 8180
rect 12173 8146 12188 8172
rect 12195 8146 12214 8172
rect 12278 8168 12309 8180
rect 12324 8168 12427 8180
rect 12439 8170 12465 8196
rect 12480 8191 12510 8202
rect 12542 8198 12604 8214
rect 12542 8196 12588 8198
rect 12542 8180 12604 8196
rect 12616 8180 12622 8228
rect 12625 8220 12705 8228
rect 12625 8218 12644 8220
rect 12659 8218 12693 8220
rect 12625 8202 12705 8218
rect 12625 8180 12644 8202
rect 12659 8186 12689 8202
rect 12717 8196 12723 8270
rect 12726 8196 12745 8340
rect 12760 8196 12766 8340
rect 12775 8270 12788 8340
rect 12840 8336 12862 8340
rect 12833 8314 12862 8328
rect 12915 8314 12931 8328
rect 12969 8324 12975 8326
rect 12982 8324 13090 8340
rect 13097 8324 13103 8326
rect 13111 8324 13126 8340
rect 13192 8334 13211 8337
rect 12833 8312 12931 8314
rect 12958 8312 13126 8324
rect 13141 8314 13157 8328
rect 13192 8315 13214 8334
rect 13224 8328 13240 8329
rect 13223 8326 13240 8328
rect 13224 8321 13240 8326
rect 13214 8314 13220 8315
rect 13223 8314 13252 8321
rect 13141 8313 13252 8314
rect 13141 8312 13258 8313
rect 12817 8304 12868 8312
rect 12915 8304 12949 8312
rect 12817 8292 12842 8304
rect 12849 8292 12868 8304
rect 12922 8302 12949 8304
rect 12958 8302 13179 8312
rect 13214 8309 13220 8312
rect 12922 8298 13179 8302
rect 12817 8284 12868 8292
rect 12915 8284 13179 8298
rect 13223 8304 13258 8312
rect 12769 8236 12788 8270
rect 12833 8276 12862 8284
rect 12833 8270 12850 8276
rect 12833 8268 12867 8270
rect 12915 8268 12931 8284
rect 12932 8274 13140 8284
rect 13141 8274 13157 8284
rect 13205 8280 13220 8295
rect 13223 8292 13224 8304
rect 13231 8292 13258 8304
rect 13223 8284 13258 8292
rect 13223 8283 13252 8284
rect 12943 8270 13157 8274
rect 12958 8268 13157 8270
rect 13192 8270 13205 8280
rect 13223 8270 13240 8283
rect 13192 8268 13240 8270
rect 12834 8264 12867 8268
rect 12830 8262 12867 8264
rect 12830 8261 12897 8262
rect 12830 8256 12861 8261
rect 12867 8256 12897 8261
rect 12830 8252 12897 8256
rect 12803 8249 12897 8252
rect 12803 8242 12852 8249
rect 12803 8236 12833 8242
rect 12852 8237 12857 8242
rect 12769 8220 12849 8236
rect 12861 8228 12897 8249
rect 12958 8244 13147 8268
rect 13192 8267 13239 8268
rect 13205 8262 13239 8267
rect 12973 8241 13147 8244
rect 12966 8238 13147 8241
rect 13175 8261 13239 8262
rect 12769 8218 12788 8220
rect 12803 8218 12837 8220
rect 12769 8202 12849 8218
rect 12769 8196 12788 8202
rect 12485 8170 12588 8180
rect 12439 8168 12588 8170
rect 12609 8168 12644 8180
rect 12278 8166 12440 8168
rect 12290 8146 12309 8166
rect 12324 8164 12354 8166
rect 12173 8138 12214 8146
rect 12296 8142 12309 8146
rect 12361 8150 12440 8166
rect 12472 8166 12644 8168
rect 12472 8150 12551 8166
rect 12558 8164 12588 8166
rect 12136 8128 12165 8138
rect 12179 8128 12208 8138
rect 12223 8128 12253 8142
rect 12296 8128 12339 8142
rect 12361 8138 12551 8150
rect 12616 8146 12622 8166
rect 12346 8128 12376 8138
rect 12377 8128 12535 8138
rect 12539 8128 12569 8138
rect 12573 8128 12603 8142
rect 12631 8128 12644 8166
rect 12716 8180 12745 8196
rect 12759 8180 12788 8196
rect 12803 8186 12833 8202
rect 12861 8180 12867 8228
rect 12870 8222 12889 8228
rect 12904 8222 12934 8230
rect 12870 8214 12934 8222
rect 12870 8198 12950 8214
rect 12966 8207 13028 8238
rect 13044 8207 13106 8238
rect 13175 8236 13224 8261
rect 13239 8236 13269 8252
rect 13138 8222 13168 8230
rect 13175 8228 13285 8236
rect 13138 8214 13183 8222
rect 12870 8196 12889 8198
rect 12904 8196 12950 8198
rect 12870 8180 12950 8196
rect 12977 8194 13012 8207
rect 13053 8204 13090 8207
rect 13053 8202 13095 8204
rect 12982 8191 13012 8194
rect 12991 8187 12998 8191
rect 12998 8186 12999 8187
rect 12957 8180 12967 8186
rect 12716 8172 12751 8180
rect 12716 8146 12717 8172
rect 12724 8146 12751 8172
rect 12659 8128 12689 8142
rect 12716 8138 12751 8146
rect 12753 8172 12794 8180
rect 12753 8146 12768 8172
rect 12775 8146 12794 8172
rect 12858 8168 12889 8180
rect 12904 8168 13007 8180
rect 13019 8170 13045 8196
rect 13060 8191 13090 8202
rect 13122 8198 13184 8214
rect 13122 8196 13168 8198
rect 13122 8180 13184 8196
rect 13196 8180 13202 8228
rect 13205 8220 13285 8228
rect 13205 8218 13224 8220
rect 13239 8218 13273 8220
rect 13205 8202 13285 8218
rect 13205 8180 13224 8202
rect 13239 8186 13269 8202
rect 13297 8196 13303 8270
rect 13306 8196 13325 8340
rect 13340 8196 13346 8340
rect 13355 8270 13368 8340
rect 13420 8336 13442 8340
rect 13413 8314 13442 8328
rect 13495 8314 13511 8328
rect 13549 8324 13555 8326
rect 13562 8324 13670 8340
rect 13677 8324 13683 8326
rect 13691 8324 13706 8340
rect 13772 8334 13791 8337
rect 13413 8312 13511 8314
rect 13538 8312 13706 8324
rect 13721 8314 13737 8328
rect 13772 8315 13794 8334
rect 13804 8328 13820 8329
rect 13803 8326 13820 8328
rect 13804 8321 13820 8326
rect 13794 8314 13800 8315
rect 13803 8314 13832 8321
rect 13721 8313 13832 8314
rect 13721 8312 13838 8313
rect 13397 8304 13448 8312
rect 13495 8304 13529 8312
rect 13397 8292 13422 8304
rect 13429 8292 13448 8304
rect 13502 8302 13529 8304
rect 13538 8302 13759 8312
rect 13794 8309 13800 8312
rect 13502 8298 13759 8302
rect 13397 8284 13448 8292
rect 13495 8284 13759 8298
rect 13803 8304 13838 8312
rect 13349 8236 13368 8270
rect 13413 8276 13442 8284
rect 13413 8270 13430 8276
rect 13413 8268 13447 8270
rect 13495 8268 13511 8284
rect 13512 8274 13720 8284
rect 13721 8274 13737 8284
rect 13785 8280 13800 8295
rect 13803 8292 13804 8304
rect 13811 8292 13838 8304
rect 13803 8284 13838 8292
rect 13803 8283 13832 8284
rect 13523 8270 13737 8274
rect 13538 8268 13737 8270
rect 13772 8270 13785 8280
rect 13803 8270 13820 8283
rect 13772 8268 13820 8270
rect 13414 8264 13447 8268
rect 13410 8262 13447 8264
rect 13410 8261 13477 8262
rect 13410 8256 13441 8261
rect 13447 8256 13477 8261
rect 13410 8252 13477 8256
rect 13383 8249 13477 8252
rect 13383 8242 13432 8249
rect 13383 8236 13413 8242
rect 13432 8237 13437 8242
rect 13349 8220 13429 8236
rect 13441 8228 13477 8249
rect 13538 8244 13727 8268
rect 13772 8267 13819 8268
rect 13785 8262 13819 8267
rect 13553 8241 13727 8244
rect 13546 8238 13727 8241
rect 13755 8261 13819 8262
rect 13349 8218 13368 8220
rect 13383 8218 13417 8220
rect 13349 8202 13429 8218
rect 13349 8196 13368 8202
rect 13065 8170 13168 8180
rect 13019 8168 13168 8170
rect 13189 8168 13224 8180
rect 12858 8166 13020 8168
rect 12870 8146 12889 8166
rect 12904 8164 12934 8166
rect 12753 8138 12794 8146
rect 12876 8142 12889 8146
rect 12941 8150 13020 8166
rect 13052 8166 13224 8168
rect 13052 8150 13131 8166
rect 13138 8164 13168 8166
rect 12716 8128 12745 8138
rect 12759 8128 12788 8138
rect 12803 8128 12833 8142
rect 12876 8128 12919 8142
rect 12941 8138 13131 8150
rect 13196 8146 13202 8166
rect 12926 8128 12956 8138
rect 12957 8128 13115 8138
rect 13119 8128 13149 8138
rect 13153 8128 13183 8142
rect 13211 8128 13224 8166
rect 13296 8180 13325 8196
rect 13339 8180 13368 8196
rect 13383 8186 13413 8202
rect 13441 8180 13447 8228
rect 13450 8222 13469 8228
rect 13484 8222 13514 8230
rect 13450 8214 13514 8222
rect 13450 8198 13530 8214
rect 13546 8207 13608 8238
rect 13624 8207 13686 8238
rect 13755 8236 13804 8261
rect 13819 8236 13849 8252
rect 13718 8222 13748 8230
rect 13755 8228 13865 8236
rect 13718 8214 13763 8222
rect 13450 8196 13469 8198
rect 13484 8196 13530 8198
rect 13450 8180 13530 8196
rect 13557 8194 13592 8207
rect 13633 8204 13670 8207
rect 13633 8202 13675 8204
rect 13562 8191 13592 8194
rect 13571 8187 13578 8191
rect 13578 8186 13579 8187
rect 13537 8180 13547 8186
rect 13296 8172 13331 8180
rect 13296 8146 13297 8172
rect 13304 8146 13331 8172
rect 13239 8128 13269 8142
rect 13296 8138 13331 8146
rect 13333 8172 13374 8180
rect 13333 8146 13348 8172
rect 13355 8146 13374 8172
rect 13438 8168 13469 8180
rect 13484 8168 13587 8180
rect 13599 8170 13625 8196
rect 13640 8191 13670 8202
rect 13702 8198 13764 8214
rect 13702 8196 13748 8198
rect 13702 8180 13764 8196
rect 13776 8180 13782 8228
rect 13785 8220 13865 8228
rect 13785 8218 13804 8220
rect 13819 8218 13853 8220
rect 13785 8202 13865 8218
rect 13785 8180 13804 8202
rect 13819 8186 13849 8202
rect 13877 8196 13883 8270
rect 13886 8196 13905 8340
rect 13920 8196 13926 8340
rect 13935 8270 13948 8340
rect 14000 8336 14022 8340
rect 13993 8314 14022 8328
rect 14075 8314 14091 8328
rect 14129 8324 14135 8326
rect 14142 8324 14250 8340
rect 14257 8324 14263 8326
rect 14271 8324 14286 8340
rect 14352 8334 14371 8337
rect 13993 8312 14091 8314
rect 14118 8312 14286 8324
rect 14301 8314 14317 8328
rect 14352 8315 14374 8334
rect 14384 8328 14400 8329
rect 14383 8326 14400 8328
rect 14384 8321 14400 8326
rect 14374 8314 14380 8315
rect 14383 8314 14412 8321
rect 14301 8313 14412 8314
rect 14301 8312 14418 8313
rect 13977 8304 14028 8312
rect 14075 8304 14109 8312
rect 13977 8292 14002 8304
rect 14009 8292 14028 8304
rect 14082 8302 14109 8304
rect 14118 8302 14339 8312
rect 14374 8309 14380 8312
rect 14082 8298 14339 8302
rect 13977 8284 14028 8292
rect 14075 8284 14339 8298
rect 14383 8304 14418 8312
rect 13929 8236 13948 8270
rect 13993 8276 14022 8284
rect 13993 8270 14010 8276
rect 13993 8268 14027 8270
rect 14075 8268 14091 8284
rect 14092 8274 14300 8284
rect 14301 8274 14317 8284
rect 14365 8280 14380 8295
rect 14383 8292 14384 8304
rect 14391 8292 14418 8304
rect 14383 8284 14418 8292
rect 14383 8283 14412 8284
rect 14103 8270 14317 8274
rect 14118 8268 14317 8270
rect 14352 8270 14365 8280
rect 14383 8270 14400 8283
rect 14352 8268 14400 8270
rect 13994 8264 14027 8268
rect 13990 8262 14027 8264
rect 13990 8261 14057 8262
rect 13990 8256 14021 8261
rect 14027 8256 14057 8261
rect 13990 8252 14057 8256
rect 13963 8249 14057 8252
rect 13963 8242 14012 8249
rect 13963 8236 13993 8242
rect 14012 8237 14017 8242
rect 13929 8220 14009 8236
rect 14021 8228 14057 8249
rect 14118 8244 14307 8268
rect 14352 8267 14399 8268
rect 14365 8262 14399 8267
rect 14133 8241 14307 8244
rect 14126 8238 14307 8241
rect 14335 8261 14399 8262
rect 13929 8218 13948 8220
rect 13963 8218 13997 8220
rect 13929 8202 14009 8218
rect 13929 8196 13948 8202
rect 13645 8170 13748 8180
rect 13599 8168 13748 8170
rect 13769 8168 13804 8180
rect 13438 8166 13600 8168
rect 13450 8146 13469 8166
rect 13484 8164 13514 8166
rect 13333 8138 13374 8146
rect 13456 8142 13469 8146
rect 13521 8150 13600 8166
rect 13632 8166 13804 8168
rect 13632 8150 13711 8166
rect 13718 8164 13748 8166
rect 13296 8128 13325 8138
rect 13339 8128 13368 8138
rect 13383 8128 13413 8142
rect 13456 8128 13499 8142
rect 13521 8138 13711 8150
rect 13776 8146 13782 8166
rect 13506 8128 13536 8138
rect 13537 8128 13695 8138
rect 13699 8128 13729 8138
rect 13733 8128 13763 8142
rect 13791 8128 13804 8166
rect 13876 8180 13905 8196
rect 13919 8180 13948 8196
rect 13963 8186 13993 8202
rect 14021 8180 14027 8228
rect 14030 8222 14049 8228
rect 14064 8222 14094 8230
rect 14030 8214 14094 8222
rect 14030 8198 14110 8214
rect 14126 8207 14188 8238
rect 14204 8207 14266 8238
rect 14335 8236 14384 8261
rect 14399 8236 14429 8252
rect 14298 8222 14328 8230
rect 14335 8228 14445 8236
rect 14298 8214 14343 8222
rect 14030 8196 14049 8198
rect 14064 8196 14110 8198
rect 14030 8180 14110 8196
rect 14137 8194 14172 8207
rect 14213 8204 14250 8207
rect 14213 8202 14255 8204
rect 14142 8191 14172 8194
rect 14151 8187 14158 8191
rect 14158 8186 14159 8187
rect 14117 8180 14127 8186
rect 13876 8172 13911 8180
rect 13876 8146 13877 8172
rect 13884 8146 13911 8172
rect 13819 8128 13849 8142
rect 13876 8138 13911 8146
rect 13913 8172 13954 8180
rect 13913 8146 13928 8172
rect 13935 8146 13954 8172
rect 14018 8168 14049 8180
rect 14064 8168 14167 8180
rect 14179 8170 14205 8196
rect 14220 8191 14250 8202
rect 14282 8198 14344 8214
rect 14282 8196 14328 8198
rect 14282 8180 14344 8196
rect 14356 8180 14362 8228
rect 14365 8220 14445 8228
rect 14365 8218 14384 8220
rect 14399 8218 14433 8220
rect 14365 8202 14445 8218
rect 14365 8180 14384 8202
rect 14399 8186 14429 8202
rect 14457 8196 14463 8270
rect 14466 8196 14485 8340
rect 14500 8196 14506 8340
rect 14515 8270 14528 8340
rect 14580 8336 14602 8340
rect 14573 8314 14602 8328
rect 14655 8314 14671 8328
rect 14709 8324 14715 8326
rect 14722 8324 14830 8340
rect 14837 8324 14843 8326
rect 14851 8324 14866 8340
rect 14932 8334 14951 8337
rect 14573 8312 14671 8314
rect 14698 8312 14866 8324
rect 14881 8314 14897 8328
rect 14932 8315 14954 8334
rect 14964 8328 14980 8329
rect 14963 8326 14980 8328
rect 14964 8321 14980 8326
rect 14954 8314 14960 8315
rect 14963 8314 14992 8321
rect 14881 8313 14992 8314
rect 14881 8312 14998 8313
rect 14557 8304 14608 8312
rect 14655 8304 14689 8312
rect 14557 8292 14582 8304
rect 14589 8292 14608 8304
rect 14662 8302 14689 8304
rect 14698 8302 14919 8312
rect 14954 8309 14960 8312
rect 14662 8298 14919 8302
rect 14557 8284 14608 8292
rect 14655 8284 14919 8298
rect 14963 8304 14998 8312
rect 14509 8236 14528 8270
rect 14573 8276 14602 8284
rect 14573 8270 14590 8276
rect 14573 8268 14607 8270
rect 14655 8268 14671 8284
rect 14672 8274 14880 8284
rect 14881 8274 14897 8284
rect 14945 8280 14960 8295
rect 14963 8292 14964 8304
rect 14971 8292 14998 8304
rect 14963 8284 14998 8292
rect 14963 8283 14992 8284
rect 14683 8270 14897 8274
rect 14698 8268 14897 8270
rect 14932 8270 14945 8280
rect 14963 8270 14980 8283
rect 14932 8268 14980 8270
rect 14574 8264 14607 8268
rect 14570 8262 14607 8264
rect 14570 8261 14637 8262
rect 14570 8256 14601 8261
rect 14607 8256 14637 8261
rect 14570 8252 14637 8256
rect 14543 8249 14637 8252
rect 14543 8242 14592 8249
rect 14543 8236 14573 8242
rect 14592 8237 14597 8242
rect 14509 8220 14589 8236
rect 14601 8228 14637 8249
rect 14698 8244 14887 8268
rect 14932 8267 14979 8268
rect 14945 8262 14979 8267
rect 14713 8241 14887 8244
rect 14706 8238 14887 8241
rect 14915 8261 14979 8262
rect 14509 8218 14528 8220
rect 14543 8218 14577 8220
rect 14509 8202 14589 8218
rect 14509 8196 14528 8202
rect 14225 8170 14328 8180
rect 14179 8168 14328 8170
rect 14349 8168 14384 8180
rect 14018 8166 14180 8168
rect 14030 8146 14049 8166
rect 14064 8164 14094 8166
rect 13913 8138 13954 8146
rect 14036 8142 14049 8146
rect 14101 8150 14180 8166
rect 14212 8166 14384 8168
rect 14212 8150 14291 8166
rect 14298 8164 14328 8166
rect 13876 8128 13905 8138
rect 13919 8128 13948 8138
rect 13963 8128 13993 8142
rect 14036 8128 14079 8142
rect 14101 8138 14291 8150
rect 14356 8146 14362 8166
rect 14086 8128 14116 8138
rect 14117 8128 14275 8138
rect 14279 8128 14309 8138
rect 14313 8128 14343 8142
rect 14371 8128 14384 8166
rect 14456 8180 14485 8196
rect 14499 8180 14528 8196
rect 14543 8186 14573 8202
rect 14601 8180 14607 8228
rect 14610 8222 14629 8228
rect 14644 8222 14674 8230
rect 14610 8214 14674 8222
rect 14610 8198 14690 8214
rect 14706 8207 14768 8238
rect 14784 8207 14846 8238
rect 14915 8236 14964 8261
rect 14979 8236 15009 8252
rect 14878 8222 14908 8230
rect 14915 8228 15025 8236
rect 14878 8214 14923 8222
rect 14610 8196 14629 8198
rect 14644 8196 14690 8198
rect 14610 8180 14690 8196
rect 14717 8194 14752 8207
rect 14793 8204 14830 8207
rect 14793 8202 14835 8204
rect 14722 8191 14752 8194
rect 14731 8187 14738 8191
rect 14738 8186 14739 8187
rect 14697 8180 14707 8186
rect 14456 8172 14491 8180
rect 14456 8146 14457 8172
rect 14464 8146 14491 8172
rect 14399 8128 14429 8142
rect 14456 8138 14491 8146
rect 14493 8172 14534 8180
rect 14493 8146 14508 8172
rect 14515 8146 14534 8172
rect 14598 8168 14629 8180
rect 14644 8168 14747 8180
rect 14759 8170 14785 8196
rect 14800 8191 14830 8202
rect 14862 8198 14924 8214
rect 14862 8196 14908 8198
rect 14862 8180 14924 8196
rect 14936 8180 14942 8228
rect 14945 8220 15025 8228
rect 14945 8218 14964 8220
rect 14979 8218 15013 8220
rect 14945 8202 15025 8218
rect 14945 8180 14964 8202
rect 14979 8186 15009 8202
rect 15037 8196 15043 8270
rect 15046 8196 15065 8340
rect 15080 8196 15086 8340
rect 15095 8270 15108 8340
rect 15160 8336 15182 8340
rect 15153 8314 15182 8328
rect 15235 8314 15251 8328
rect 15289 8324 15295 8326
rect 15302 8324 15410 8340
rect 15417 8324 15423 8326
rect 15431 8324 15446 8340
rect 15512 8334 15531 8337
rect 15153 8312 15251 8314
rect 15278 8312 15446 8324
rect 15461 8314 15477 8328
rect 15512 8315 15534 8334
rect 15544 8328 15560 8329
rect 15543 8326 15560 8328
rect 15544 8321 15560 8326
rect 15534 8314 15540 8315
rect 15543 8314 15572 8321
rect 15461 8313 15572 8314
rect 15461 8312 15578 8313
rect 15137 8304 15188 8312
rect 15235 8304 15269 8312
rect 15137 8292 15162 8304
rect 15169 8292 15188 8304
rect 15242 8302 15269 8304
rect 15278 8302 15499 8312
rect 15534 8309 15540 8312
rect 15242 8298 15499 8302
rect 15137 8284 15188 8292
rect 15235 8284 15499 8298
rect 15543 8304 15578 8312
rect 15089 8236 15108 8270
rect 15153 8276 15182 8284
rect 15153 8270 15170 8276
rect 15153 8268 15187 8270
rect 15235 8268 15251 8284
rect 15252 8274 15460 8284
rect 15461 8274 15477 8284
rect 15525 8280 15540 8295
rect 15543 8292 15544 8304
rect 15551 8292 15578 8304
rect 15543 8284 15578 8292
rect 15543 8283 15572 8284
rect 15263 8270 15477 8274
rect 15278 8268 15477 8270
rect 15512 8270 15525 8280
rect 15543 8270 15560 8283
rect 15512 8268 15560 8270
rect 15154 8264 15187 8268
rect 15150 8262 15187 8264
rect 15150 8261 15217 8262
rect 15150 8256 15181 8261
rect 15187 8256 15217 8261
rect 15150 8252 15217 8256
rect 15123 8249 15217 8252
rect 15123 8242 15172 8249
rect 15123 8236 15153 8242
rect 15172 8237 15177 8242
rect 15089 8220 15169 8236
rect 15181 8228 15217 8249
rect 15278 8244 15467 8268
rect 15512 8267 15559 8268
rect 15525 8262 15559 8267
rect 15293 8241 15467 8244
rect 15286 8238 15467 8241
rect 15495 8261 15559 8262
rect 15089 8218 15108 8220
rect 15123 8218 15157 8220
rect 15089 8202 15169 8218
rect 15089 8196 15108 8202
rect 14805 8170 14908 8180
rect 14759 8168 14908 8170
rect 14929 8168 14964 8180
rect 14598 8166 14760 8168
rect 14610 8146 14629 8166
rect 14644 8164 14674 8166
rect 14493 8138 14534 8146
rect 14616 8142 14629 8146
rect 14681 8150 14760 8166
rect 14792 8166 14964 8168
rect 14792 8150 14871 8166
rect 14878 8164 14908 8166
rect 14456 8128 14485 8138
rect 14499 8128 14528 8138
rect 14543 8128 14573 8142
rect 14616 8128 14659 8142
rect 14681 8138 14871 8150
rect 14936 8146 14942 8166
rect 14666 8128 14696 8138
rect 14697 8128 14855 8138
rect 14859 8128 14889 8138
rect 14893 8128 14923 8142
rect 14951 8128 14964 8166
rect 15036 8180 15065 8196
rect 15079 8180 15108 8196
rect 15123 8186 15153 8202
rect 15181 8180 15187 8228
rect 15190 8222 15209 8228
rect 15224 8222 15254 8230
rect 15190 8214 15254 8222
rect 15190 8198 15270 8214
rect 15286 8207 15348 8238
rect 15364 8207 15426 8238
rect 15495 8236 15544 8261
rect 15559 8236 15589 8252
rect 15458 8222 15488 8230
rect 15495 8228 15605 8236
rect 15458 8214 15503 8222
rect 15190 8196 15209 8198
rect 15224 8196 15270 8198
rect 15190 8180 15270 8196
rect 15297 8194 15332 8207
rect 15373 8204 15410 8207
rect 15373 8202 15415 8204
rect 15302 8191 15332 8194
rect 15311 8187 15318 8191
rect 15318 8186 15319 8187
rect 15277 8180 15287 8186
rect 15036 8172 15071 8180
rect 15036 8146 15037 8172
rect 15044 8146 15071 8172
rect 14979 8128 15009 8142
rect 15036 8138 15071 8146
rect 15073 8172 15114 8180
rect 15073 8146 15088 8172
rect 15095 8146 15114 8172
rect 15178 8168 15209 8180
rect 15224 8168 15327 8180
rect 15339 8170 15365 8196
rect 15380 8191 15410 8202
rect 15442 8198 15504 8214
rect 15442 8196 15488 8198
rect 15442 8180 15504 8196
rect 15516 8180 15522 8228
rect 15525 8220 15605 8228
rect 15525 8218 15544 8220
rect 15559 8218 15593 8220
rect 15525 8202 15605 8218
rect 15525 8180 15544 8202
rect 15559 8186 15589 8202
rect 15617 8196 15623 8270
rect 15626 8196 15645 8340
rect 15660 8196 15666 8340
rect 15675 8270 15688 8340
rect 15740 8336 15762 8340
rect 15733 8314 15762 8328
rect 15815 8314 15831 8328
rect 15869 8324 15875 8326
rect 15882 8324 15990 8340
rect 15997 8324 16003 8326
rect 16011 8324 16026 8340
rect 16092 8334 16111 8337
rect 15733 8312 15831 8314
rect 15858 8312 16026 8324
rect 16041 8314 16057 8328
rect 16092 8315 16114 8334
rect 16124 8328 16140 8329
rect 16123 8326 16140 8328
rect 16124 8321 16140 8326
rect 16114 8314 16120 8315
rect 16123 8314 16152 8321
rect 16041 8313 16152 8314
rect 16041 8312 16158 8313
rect 15717 8304 15768 8312
rect 15815 8304 15849 8312
rect 15717 8292 15742 8304
rect 15749 8292 15768 8304
rect 15822 8302 15849 8304
rect 15858 8302 16079 8312
rect 16114 8309 16120 8312
rect 15822 8298 16079 8302
rect 15717 8284 15768 8292
rect 15815 8284 16079 8298
rect 16123 8304 16158 8312
rect 15669 8236 15688 8270
rect 15733 8276 15762 8284
rect 15733 8270 15750 8276
rect 15733 8268 15767 8270
rect 15815 8268 15831 8284
rect 15832 8274 16040 8284
rect 16041 8274 16057 8284
rect 16105 8280 16120 8295
rect 16123 8292 16124 8304
rect 16131 8292 16158 8304
rect 16123 8284 16158 8292
rect 16123 8283 16152 8284
rect 15843 8270 16057 8274
rect 15858 8268 16057 8270
rect 16092 8270 16105 8280
rect 16123 8270 16140 8283
rect 16092 8268 16140 8270
rect 15734 8264 15767 8268
rect 15730 8262 15767 8264
rect 15730 8261 15797 8262
rect 15730 8256 15761 8261
rect 15767 8256 15797 8261
rect 15730 8252 15797 8256
rect 15703 8249 15797 8252
rect 15703 8242 15752 8249
rect 15703 8236 15733 8242
rect 15752 8237 15757 8242
rect 15669 8220 15749 8236
rect 15761 8228 15797 8249
rect 15858 8244 16047 8268
rect 16092 8267 16139 8268
rect 16105 8262 16139 8267
rect 15873 8241 16047 8244
rect 15866 8238 16047 8241
rect 16075 8261 16139 8262
rect 15669 8218 15688 8220
rect 15703 8218 15737 8220
rect 15669 8202 15749 8218
rect 15669 8196 15688 8202
rect 15385 8170 15488 8180
rect 15339 8168 15488 8170
rect 15509 8168 15544 8180
rect 15178 8166 15340 8168
rect 15190 8146 15209 8166
rect 15224 8164 15254 8166
rect 15073 8138 15114 8146
rect 15196 8142 15209 8146
rect 15261 8150 15340 8166
rect 15372 8166 15544 8168
rect 15372 8150 15451 8166
rect 15458 8164 15488 8166
rect 15036 8128 15065 8138
rect 15079 8128 15108 8138
rect 15123 8128 15153 8142
rect 15196 8128 15239 8142
rect 15261 8138 15451 8150
rect 15516 8146 15522 8166
rect 15246 8128 15276 8138
rect 15277 8128 15435 8138
rect 15439 8128 15469 8138
rect 15473 8128 15503 8142
rect 15531 8128 15544 8166
rect 15616 8180 15645 8196
rect 15659 8180 15688 8196
rect 15703 8186 15733 8202
rect 15761 8180 15767 8228
rect 15770 8222 15789 8228
rect 15804 8222 15834 8230
rect 15770 8214 15834 8222
rect 15770 8198 15850 8214
rect 15866 8207 15928 8238
rect 15944 8207 16006 8238
rect 16075 8236 16124 8261
rect 16139 8236 16169 8252
rect 16038 8222 16068 8230
rect 16075 8228 16185 8236
rect 16038 8214 16083 8222
rect 15770 8196 15789 8198
rect 15804 8196 15850 8198
rect 15770 8180 15850 8196
rect 15877 8194 15912 8207
rect 15953 8204 15990 8207
rect 15953 8202 15995 8204
rect 15882 8191 15912 8194
rect 15891 8187 15898 8191
rect 15898 8186 15899 8187
rect 15857 8180 15867 8186
rect 15616 8172 15651 8180
rect 15616 8146 15617 8172
rect 15624 8146 15651 8172
rect 15559 8128 15589 8142
rect 15616 8138 15651 8146
rect 15653 8172 15694 8180
rect 15653 8146 15668 8172
rect 15675 8146 15694 8172
rect 15758 8168 15789 8180
rect 15804 8168 15907 8180
rect 15919 8170 15945 8196
rect 15960 8191 15990 8202
rect 16022 8198 16084 8214
rect 16022 8196 16068 8198
rect 16022 8180 16084 8196
rect 16096 8180 16102 8228
rect 16105 8220 16185 8228
rect 16105 8218 16124 8220
rect 16139 8218 16173 8220
rect 16105 8202 16185 8218
rect 16105 8180 16124 8202
rect 16139 8186 16169 8202
rect 16197 8196 16203 8270
rect 16206 8196 16225 8340
rect 16240 8196 16246 8340
rect 16255 8270 16268 8340
rect 16320 8336 16342 8340
rect 16313 8314 16342 8328
rect 16395 8314 16411 8328
rect 16449 8324 16455 8326
rect 16462 8324 16570 8340
rect 16577 8324 16583 8326
rect 16591 8324 16606 8340
rect 16672 8334 16691 8337
rect 16313 8312 16411 8314
rect 16438 8312 16606 8324
rect 16621 8314 16637 8328
rect 16672 8315 16694 8334
rect 16704 8328 16720 8329
rect 16703 8326 16720 8328
rect 16704 8321 16720 8326
rect 16694 8314 16700 8315
rect 16703 8314 16732 8321
rect 16621 8313 16732 8314
rect 16621 8312 16738 8313
rect 16297 8304 16348 8312
rect 16395 8304 16429 8312
rect 16297 8292 16322 8304
rect 16329 8292 16348 8304
rect 16402 8302 16429 8304
rect 16438 8302 16659 8312
rect 16694 8309 16700 8312
rect 16402 8298 16659 8302
rect 16297 8284 16348 8292
rect 16395 8284 16659 8298
rect 16703 8304 16738 8312
rect 16249 8236 16268 8270
rect 16313 8276 16342 8284
rect 16313 8270 16330 8276
rect 16313 8268 16347 8270
rect 16395 8268 16411 8284
rect 16412 8274 16620 8284
rect 16621 8274 16637 8284
rect 16685 8280 16700 8295
rect 16703 8292 16704 8304
rect 16711 8292 16738 8304
rect 16703 8284 16738 8292
rect 16703 8283 16732 8284
rect 16423 8270 16637 8274
rect 16438 8268 16637 8270
rect 16672 8270 16685 8280
rect 16703 8270 16720 8283
rect 16672 8268 16720 8270
rect 16314 8264 16347 8268
rect 16310 8262 16347 8264
rect 16310 8261 16377 8262
rect 16310 8256 16341 8261
rect 16347 8256 16377 8261
rect 16310 8252 16377 8256
rect 16283 8249 16377 8252
rect 16283 8242 16332 8249
rect 16283 8236 16313 8242
rect 16332 8237 16337 8242
rect 16249 8220 16329 8236
rect 16341 8228 16377 8249
rect 16438 8244 16627 8268
rect 16672 8267 16719 8268
rect 16685 8262 16719 8267
rect 16453 8241 16627 8244
rect 16446 8238 16627 8241
rect 16655 8261 16719 8262
rect 16249 8218 16268 8220
rect 16283 8218 16317 8220
rect 16249 8202 16329 8218
rect 16249 8196 16268 8202
rect 15965 8170 16068 8180
rect 15919 8168 16068 8170
rect 16089 8168 16124 8180
rect 15758 8166 15920 8168
rect 15770 8146 15789 8166
rect 15804 8164 15834 8166
rect 15653 8138 15694 8146
rect 15776 8142 15789 8146
rect 15841 8150 15920 8166
rect 15952 8166 16124 8168
rect 15952 8150 16031 8166
rect 16038 8164 16068 8166
rect 15616 8128 15645 8138
rect 15659 8128 15688 8138
rect 15703 8128 15733 8142
rect 15776 8128 15819 8142
rect 15841 8138 16031 8150
rect 16096 8146 16102 8166
rect 15826 8128 15856 8138
rect 15857 8128 16015 8138
rect 16019 8128 16049 8138
rect 16053 8128 16083 8142
rect 16111 8128 16124 8166
rect 16196 8180 16225 8196
rect 16239 8180 16268 8196
rect 16283 8186 16313 8202
rect 16341 8180 16347 8228
rect 16350 8222 16369 8228
rect 16384 8222 16414 8230
rect 16350 8214 16414 8222
rect 16350 8198 16430 8214
rect 16446 8207 16508 8238
rect 16524 8207 16586 8238
rect 16655 8236 16704 8261
rect 16719 8236 16749 8252
rect 16618 8222 16648 8230
rect 16655 8228 16765 8236
rect 16618 8214 16663 8222
rect 16350 8196 16369 8198
rect 16384 8196 16430 8198
rect 16350 8180 16430 8196
rect 16457 8194 16492 8207
rect 16533 8204 16570 8207
rect 16533 8202 16575 8204
rect 16462 8191 16492 8194
rect 16471 8187 16478 8191
rect 16478 8186 16479 8187
rect 16437 8180 16447 8186
rect 16196 8172 16231 8180
rect 16196 8146 16197 8172
rect 16204 8146 16231 8172
rect 16139 8128 16169 8142
rect 16196 8138 16231 8146
rect 16233 8172 16274 8180
rect 16233 8146 16248 8172
rect 16255 8146 16274 8172
rect 16338 8168 16369 8180
rect 16384 8168 16487 8180
rect 16499 8170 16525 8196
rect 16540 8191 16570 8202
rect 16602 8198 16664 8214
rect 16602 8196 16648 8198
rect 16602 8180 16664 8196
rect 16676 8180 16682 8228
rect 16685 8220 16765 8228
rect 16685 8218 16704 8220
rect 16719 8218 16753 8220
rect 16685 8202 16765 8218
rect 16685 8180 16704 8202
rect 16719 8186 16749 8202
rect 16777 8196 16783 8270
rect 16786 8196 16805 8340
rect 16820 8196 16826 8340
rect 16835 8270 16848 8340
rect 16900 8336 16922 8340
rect 16893 8314 16922 8328
rect 16975 8314 16991 8328
rect 17029 8324 17035 8326
rect 17042 8324 17150 8340
rect 17157 8324 17163 8326
rect 17171 8324 17186 8340
rect 17252 8334 17271 8337
rect 16893 8312 16991 8314
rect 17018 8312 17186 8324
rect 17201 8314 17217 8328
rect 17252 8315 17274 8334
rect 17284 8328 17300 8329
rect 17283 8326 17300 8328
rect 17284 8321 17300 8326
rect 17274 8314 17280 8315
rect 17283 8314 17312 8321
rect 17201 8313 17312 8314
rect 17201 8312 17318 8313
rect 16877 8304 16928 8312
rect 16975 8304 17009 8312
rect 16877 8292 16902 8304
rect 16909 8292 16928 8304
rect 16982 8302 17009 8304
rect 17018 8302 17239 8312
rect 17274 8309 17280 8312
rect 16982 8298 17239 8302
rect 16877 8284 16928 8292
rect 16975 8284 17239 8298
rect 17283 8304 17318 8312
rect 16829 8236 16848 8270
rect 16893 8276 16922 8284
rect 16893 8270 16910 8276
rect 16893 8268 16927 8270
rect 16975 8268 16991 8284
rect 16992 8274 17200 8284
rect 17201 8274 17217 8284
rect 17265 8280 17280 8295
rect 17283 8292 17284 8304
rect 17291 8292 17318 8304
rect 17283 8284 17318 8292
rect 17283 8283 17312 8284
rect 17003 8270 17217 8274
rect 17018 8268 17217 8270
rect 17252 8270 17265 8280
rect 17283 8270 17300 8283
rect 17252 8268 17300 8270
rect 16894 8264 16927 8268
rect 16890 8262 16927 8264
rect 16890 8261 16957 8262
rect 16890 8256 16921 8261
rect 16927 8256 16957 8261
rect 16890 8252 16957 8256
rect 16863 8249 16957 8252
rect 16863 8242 16912 8249
rect 16863 8236 16893 8242
rect 16912 8237 16917 8242
rect 16829 8220 16909 8236
rect 16921 8228 16957 8249
rect 17018 8244 17207 8268
rect 17252 8267 17299 8268
rect 17265 8262 17299 8267
rect 17033 8241 17207 8244
rect 17026 8238 17207 8241
rect 17235 8261 17299 8262
rect 16829 8218 16848 8220
rect 16863 8218 16897 8220
rect 16829 8202 16909 8218
rect 16829 8196 16848 8202
rect 16545 8170 16648 8180
rect 16499 8168 16648 8170
rect 16669 8168 16704 8180
rect 16338 8166 16500 8168
rect 16350 8146 16369 8166
rect 16384 8164 16414 8166
rect 16233 8138 16274 8146
rect 16356 8142 16369 8146
rect 16421 8150 16500 8166
rect 16532 8166 16704 8168
rect 16532 8150 16611 8166
rect 16618 8164 16648 8166
rect 16196 8128 16225 8138
rect 16239 8128 16268 8138
rect 16283 8128 16313 8142
rect 16356 8128 16399 8142
rect 16421 8138 16611 8150
rect 16676 8146 16682 8166
rect 16406 8128 16436 8138
rect 16437 8128 16595 8138
rect 16599 8128 16629 8138
rect 16633 8128 16663 8142
rect 16691 8128 16704 8166
rect 16776 8180 16805 8196
rect 16819 8180 16848 8196
rect 16863 8186 16893 8202
rect 16921 8180 16927 8228
rect 16930 8222 16949 8228
rect 16964 8222 16994 8230
rect 16930 8214 16994 8222
rect 16930 8198 17010 8214
rect 17026 8207 17088 8238
rect 17104 8207 17166 8238
rect 17235 8236 17284 8261
rect 17299 8236 17329 8252
rect 17198 8222 17228 8230
rect 17235 8228 17345 8236
rect 17198 8214 17243 8222
rect 16930 8196 16949 8198
rect 16964 8196 17010 8198
rect 16930 8180 17010 8196
rect 17037 8194 17072 8207
rect 17113 8204 17150 8207
rect 17113 8202 17155 8204
rect 17042 8191 17072 8194
rect 17051 8187 17058 8191
rect 17058 8186 17059 8187
rect 17017 8180 17027 8186
rect 16776 8172 16811 8180
rect 16776 8146 16777 8172
rect 16784 8146 16811 8172
rect 16719 8128 16749 8142
rect 16776 8138 16811 8146
rect 16813 8172 16854 8180
rect 16813 8146 16828 8172
rect 16835 8146 16854 8172
rect 16918 8168 16949 8180
rect 16964 8168 17067 8180
rect 17079 8170 17105 8196
rect 17120 8191 17150 8202
rect 17182 8198 17244 8214
rect 17182 8196 17228 8198
rect 17182 8180 17244 8196
rect 17256 8180 17262 8228
rect 17265 8220 17345 8228
rect 17265 8218 17284 8220
rect 17299 8218 17333 8220
rect 17265 8202 17345 8218
rect 17265 8180 17284 8202
rect 17299 8186 17329 8202
rect 17357 8196 17363 8270
rect 17366 8196 17385 8340
rect 17400 8196 17406 8340
rect 17415 8270 17428 8340
rect 17480 8336 17502 8340
rect 17473 8314 17502 8328
rect 17555 8314 17571 8328
rect 17609 8324 17615 8326
rect 17622 8324 17730 8340
rect 17737 8324 17743 8326
rect 17751 8324 17766 8340
rect 17832 8334 17851 8337
rect 17473 8312 17571 8314
rect 17598 8312 17766 8324
rect 17781 8314 17797 8328
rect 17832 8315 17854 8334
rect 17864 8328 17880 8329
rect 17863 8326 17880 8328
rect 17864 8321 17880 8326
rect 17854 8314 17860 8315
rect 17863 8314 17892 8321
rect 17781 8313 17892 8314
rect 17781 8312 17898 8313
rect 17457 8304 17508 8312
rect 17555 8304 17589 8312
rect 17457 8292 17482 8304
rect 17489 8292 17508 8304
rect 17562 8302 17589 8304
rect 17598 8302 17819 8312
rect 17854 8309 17860 8312
rect 17562 8298 17819 8302
rect 17457 8284 17508 8292
rect 17555 8284 17819 8298
rect 17863 8304 17898 8312
rect 17409 8236 17428 8270
rect 17473 8276 17502 8284
rect 17473 8270 17490 8276
rect 17473 8268 17507 8270
rect 17555 8268 17571 8284
rect 17572 8274 17780 8284
rect 17781 8274 17797 8284
rect 17845 8280 17860 8295
rect 17863 8292 17864 8304
rect 17871 8292 17898 8304
rect 17863 8284 17898 8292
rect 17863 8283 17892 8284
rect 17583 8270 17797 8274
rect 17598 8268 17797 8270
rect 17832 8270 17845 8280
rect 17863 8270 17880 8283
rect 17832 8268 17880 8270
rect 17474 8264 17507 8268
rect 17470 8262 17507 8264
rect 17470 8261 17537 8262
rect 17470 8256 17501 8261
rect 17507 8256 17537 8261
rect 17470 8252 17537 8256
rect 17443 8249 17537 8252
rect 17443 8242 17492 8249
rect 17443 8236 17473 8242
rect 17492 8237 17497 8242
rect 17409 8220 17489 8236
rect 17501 8228 17537 8249
rect 17598 8244 17787 8268
rect 17832 8267 17879 8268
rect 17845 8262 17879 8267
rect 17613 8241 17787 8244
rect 17606 8238 17787 8241
rect 17815 8261 17879 8262
rect 17409 8218 17428 8220
rect 17443 8218 17477 8220
rect 17409 8202 17489 8218
rect 17409 8196 17428 8202
rect 17125 8170 17228 8180
rect 17079 8168 17228 8170
rect 17249 8168 17284 8180
rect 16918 8166 17080 8168
rect 16930 8146 16949 8166
rect 16964 8164 16994 8166
rect 16813 8138 16854 8146
rect 16936 8142 16949 8146
rect 17001 8150 17080 8166
rect 17112 8166 17284 8168
rect 17112 8150 17191 8166
rect 17198 8164 17228 8166
rect 16776 8128 16805 8138
rect 16819 8128 16848 8138
rect 16863 8128 16893 8142
rect 16936 8128 16979 8142
rect 17001 8138 17191 8150
rect 17256 8146 17262 8166
rect 16986 8128 17016 8138
rect 17017 8128 17175 8138
rect 17179 8128 17209 8138
rect 17213 8128 17243 8142
rect 17271 8128 17284 8166
rect 17356 8180 17385 8196
rect 17399 8180 17428 8196
rect 17443 8186 17473 8202
rect 17501 8180 17507 8228
rect 17510 8222 17529 8228
rect 17544 8222 17574 8230
rect 17510 8214 17574 8222
rect 17510 8198 17590 8214
rect 17606 8207 17668 8238
rect 17684 8207 17746 8238
rect 17815 8236 17864 8261
rect 17879 8236 17909 8252
rect 17778 8222 17808 8230
rect 17815 8228 17925 8236
rect 17778 8214 17823 8222
rect 17510 8196 17529 8198
rect 17544 8196 17590 8198
rect 17510 8180 17590 8196
rect 17617 8194 17652 8207
rect 17693 8204 17730 8207
rect 17693 8202 17735 8204
rect 17622 8191 17652 8194
rect 17631 8187 17638 8191
rect 17638 8186 17639 8187
rect 17597 8180 17607 8186
rect 17356 8172 17391 8180
rect 17356 8146 17357 8172
rect 17364 8146 17391 8172
rect 17299 8128 17329 8142
rect 17356 8138 17391 8146
rect 17393 8172 17434 8180
rect 17393 8146 17408 8172
rect 17415 8146 17434 8172
rect 17498 8168 17529 8180
rect 17544 8168 17647 8180
rect 17659 8170 17685 8196
rect 17700 8191 17730 8202
rect 17762 8198 17824 8214
rect 17762 8196 17808 8198
rect 17762 8180 17824 8196
rect 17836 8180 17842 8228
rect 17845 8220 17925 8228
rect 17845 8218 17864 8220
rect 17879 8218 17913 8220
rect 17845 8202 17925 8218
rect 17845 8180 17864 8202
rect 17879 8186 17909 8202
rect 17937 8196 17943 8270
rect 17946 8196 17965 8340
rect 17980 8196 17986 8340
rect 17995 8270 18008 8340
rect 18060 8336 18082 8340
rect 18053 8314 18082 8328
rect 18135 8314 18151 8328
rect 18189 8324 18195 8326
rect 18202 8324 18310 8340
rect 18317 8324 18323 8326
rect 18331 8324 18346 8340
rect 18412 8334 18431 8337
rect 18053 8312 18151 8314
rect 18178 8312 18346 8324
rect 18361 8314 18377 8328
rect 18412 8315 18434 8334
rect 18444 8328 18460 8329
rect 18443 8326 18460 8328
rect 18444 8321 18460 8326
rect 18434 8314 18440 8315
rect 18443 8314 18472 8321
rect 18361 8313 18472 8314
rect 18361 8312 18478 8313
rect 18037 8304 18088 8312
rect 18135 8304 18169 8312
rect 18037 8292 18062 8304
rect 18069 8292 18088 8304
rect 18142 8302 18169 8304
rect 18178 8302 18399 8312
rect 18434 8309 18440 8312
rect 18142 8298 18399 8302
rect 18037 8284 18088 8292
rect 18135 8284 18399 8298
rect 18443 8304 18478 8312
rect 17989 8236 18008 8270
rect 18053 8276 18082 8284
rect 18053 8270 18070 8276
rect 18053 8268 18087 8270
rect 18135 8268 18151 8284
rect 18152 8274 18360 8284
rect 18361 8274 18377 8284
rect 18425 8280 18440 8295
rect 18443 8292 18444 8304
rect 18451 8292 18478 8304
rect 18443 8284 18478 8292
rect 18443 8283 18472 8284
rect 18163 8270 18377 8274
rect 18178 8268 18377 8270
rect 18412 8270 18425 8280
rect 18443 8270 18460 8283
rect 18412 8268 18460 8270
rect 18054 8264 18087 8268
rect 18050 8262 18087 8264
rect 18050 8261 18117 8262
rect 18050 8256 18081 8261
rect 18087 8256 18117 8261
rect 18050 8252 18117 8256
rect 18023 8249 18117 8252
rect 18023 8242 18072 8249
rect 18023 8236 18053 8242
rect 18072 8237 18077 8242
rect 17989 8220 18069 8236
rect 18081 8228 18117 8249
rect 18178 8244 18367 8268
rect 18412 8267 18459 8268
rect 18425 8262 18459 8267
rect 18193 8241 18367 8244
rect 18186 8238 18367 8241
rect 18395 8261 18459 8262
rect 17989 8218 18008 8220
rect 18023 8218 18057 8220
rect 17989 8202 18069 8218
rect 17989 8196 18008 8202
rect 17705 8170 17808 8180
rect 17659 8168 17808 8170
rect 17829 8168 17864 8180
rect 17498 8166 17660 8168
rect 17510 8146 17529 8166
rect 17544 8164 17574 8166
rect 17393 8138 17434 8146
rect 17516 8142 17529 8146
rect 17581 8150 17660 8166
rect 17692 8166 17864 8168
rect 17692 8150 17771 8166
rect 17778 8164 17808 8166
rect 17356 8128 17385 8138
rect 17399 8128 17428 8138
rect 17443 8128 17473 8142
rect 17516 8128 17559 8142
rect 17581 8138 17771 8150
rect 17836 8146 17842 8166
rect 17566 8128 17596 8138
rect 17597 8128 17755 8138
rect 17759 8128 17789 8138
rect 17793 8128 17823 8142
rect 17851 8128 17864 8166
rect 17936 8180 17965 8196
rect 17979 8180 18008 8196
rect 18023 8186 18053 8202
rect 18081 8180 18087 8228
rect 18090 8222 18109 8228
rect 18124 8222 18154 8230
rect 18090 8214 18154 8222
rect 18090 8198 18170 8214
rect 18186 8207 18248 8238
rect 18264 8207 18326 8238
rect 18395 8236 18444 8261
rect 18459 8236 18489 8252
rect 18358 8222 18388 8230
rect 18395 8228 18505 8236
rect 18358 8214 18403 8222
rect 18090 8196 18109 8198
rect 18124 8196 18170 8198
rect 18090 8180 18170 8196
rect 18197 8194 18232 8207
rect 18273 8204 18310 8207
rect 18273 8202 18315 8204
rect 18202 8191 18232 8194
rect 18211 8187 18218 8191
rect 18218 8186 18219 8187
rect 18177 8180 18187 8186
rect 17936 8172 17971 8180
rect 17936 8146 17937 8172
rect 17944 8146 17971 8172
rect 17879 8128 17909 8142
rect 17936 8138 17971 8146
rect 17973 8172 18014 8180
rect 17973 8146 17988 8172
rect 17995 8146 18014 8172
rect 18078 8168 18109 8180
rect 18124 8168 18227 8180
rect 18239 8170 18265 8196
rect 18280 8191 18310 8202
rect 18342 8198 18404 8214
rect 18342 8196 18388 8198
rect 18342 8180 18404 8196
rect 18416 8180 18422 8228
rect 18425 8220 18505 8228
rect 18425 8218 18444 8220
rect 18459 8218 18493 8220
rect 18425 8202 18505 8218
rect 18425 8180 18444 8202
rect 18459 8186 18489 8202
rect 18517 8196 18523 8270
rect 18532 8196 18545 8340
rect 18285 8170 18388 8180
rect 18239 8168 18388 8170
rect 18409 8168 18444 8180
rect 18078 8166 18240 8168
rect 18090 8146 18109 8166
rect 18124 8164 18154 8166
rect 17973 8138 18014 8146
rect 18096 8142 18109 8146
rect 18161 8150 18240 8166
rect 18272 8166 18444 8168
rect 18272 8150 18351 8166
rect 18358 8164 18388 8166
rect 17936 8128 17965 8138
rect 17979 8128 18008 8138
rect 18023 8128 18053 8142
rect 18096 8128 18139 8142
rect 18161 8138 18351 8150
rect 18416 8146 18422 8166
rect 18146 8128 18176 8138
rect 18177 8128 18335 8138
rect 18339 8128 18369 8138
rect 18373 8128 18403 8142
rect 18431 8128 18444 8166
rect 18516 8180 18545 8196
rect 18516 8172 18551 8180
rect 18516 8146 18517 8172
rect 18524 8146 18551 8172
rect 18459 8128 18489 8142
rect 18516 8138 18551 8146
rect 18516 8128 18545 8138
rect -1 8122 18545 8128
rect 0 8114 18545 8122
rect 15 8084 28 8114
rect 43 8100 73 8114
rect 116 8100 159 8114
rect 166 8100 386 8114
rect 393 8100 423 8114
rect 83 8086 98 8098
rect 117 8086 130 8100
rect 198 8096 351 8100
rect 80 8084 102 8086
rect 180 8084 372 8096
rect 451 8084 464 8114
rect 479 8100 509 8114
rect 546 8084 565 8114
rect 580 8084 586 8114
rect 595 8084 608 8114
rect 623 8100 653 8114
rect 696 8100 739 8114
rect 746 8100 966 8114
rect 973 8100 1003 8114
rect 663 8086 678 8098
rect 697 8086 710 8100
rect 778 8096 931 8100
rect 660 8084 682 8086
rect 760 8084 952 8096
rect 1031 8084 1044 8114
rect 1059 8100 1089 8114
rect 1126 8084 1145 8114
rect 1160 8084 1166 8114
rect 1175 8084 1188 8114
rect 1203 8100 1233 8114
rect 1276 8100 1319 8114
rect 1326 8100 1546 8114
rect 1553 8100 1583 8114
rect 1243 8086 1258 8098
rect 1277 8086 1290 8100
rect 1358 8096 1511 8100
rect 1240 8084 1262 8086
rect 1340 8084 1532 8096
rect 1611 8084 1624 8114
rect 1639 8100 1669 8114
rect 1706 8084 1725 8114
rect 1740 8084 1746 8114
rect 1755 8084 1768 8114
rect 1783 8100 1813 8114
rect 1856 8100 1899 8114
rect 1906 8100 2126 8114
rect 2133 8100 2163 8114
rect 1823 8086 1838 8098
rect 1857 8086 1870 8100
rect 1938 8096 2091 8100
rect 1820 8084 1842 8086
rect 1920 8084 2112 8096
rect 2191 8084 2204 8114
rect 2219 8100 2249 8114
rect 2286 8084 2305 8114
rect 2320 8084 2326 8114
rect 2335 8084 2348 8114
rect 2363 8100 2393 8114
rect 2436 8100 2479 8114
rect 2486 8100 2706 8114
rect 2713 8100 2743 8114
rect 2403 8086 2418 8098
rect 2437 8086 2450 8100
rect 2518 8096 2671 8100
rect 2400 8084 2422 8086
rect 2500 8084 2692 8096
rect 2771 8084 2784 8114
rect 2799 8100 2829 8114
rect 2866 8084 2885 8114
rect 2900 8084 2906 8114
rect 2915 8084 2928 8114
rect 2943 8100 2973 8114
rect 3016 8100 3059 8114
rect 3066 8100 3286 8114
rect 3293 8100 3323 8114
rect 2983 8086 2998 8098
rect 3017 8086 3030 8100
rect 3098 8096 3251 8100
rect 2980 8084 3002 8086
rect 3080 8084 3272 8096
rect 3351 8084 3364 8114
rect 3379 8100 3409 8114
rect 3446 8084 3465 8114
rect 3480 8084 3486 8114
rect 3495 8084 3508 8114
rect 3523 8100 3553 8114
rect 3596 8100 3639 8114
rect 3646 8100 3866 8114
rect 3873 8100 3903 8114
rect 3563 8086 3578 8098
rect 3597 8086 3610 8100
rect 3678 8096 3831 8100
rect 3560 8084 3582 8086
rect 3660 8084 3852 8096
rect 3931 8084 3944 8114
rect 3959 8100 3989 8114
rect 4026 8084 4045 8114
rect 4060 8084 4066 8114
rect 4075 8084 4088 8114
rect 4103 8100 4133 8114
rect 4176 8100 4219 8114
rect 4226 8100 4446 8114
rect 4453 8100 4483 8114
rect 4143 8086 4158 8098
rect 4177 8086 4190 8100
rect 4258 8096 4411 8100
rect 4140 8084 4162 8086
rect 4240 8084 4432 8096
rect 4511 8084 4524 8114
rect 4539 8100 4569 8114
rect 4606 8084 4625 8114
rect 4640 8084 4646 8114
rect 4655 8084 4668 8114
rect 4683 8100 4713 8114
rect 4756 8100 4799 8114
rect 4806 8100 5026 8114
rect 5033 8100 5063 8114
rect 4723 8086 4738 8098
rect 4757 8086 4770 8100
rect 4838 8096 4991 8100
rect 4720 8084 4742 8086
rect 4820 8084 5012 8096
rect 5091 8084 5104 8114
rect 5119 8100 5149 8114
rect 5186 8084 5205 8114
rect 5220 8084 5226 8114
rect 5235 8084 5248 8114
rect 5263 8100 5293 8114
rect 5336 8100 5379 8114
rect 5386 8100 5606 8114
rect 5613 8100 5643 8114
rect 5303 8086 5318 8098
rect 5337 8086 5350 8100
rect 5418 8096 5571 8100
rect 5300 8084 5322 8086
rect 5400 8084 5592 8096
rect 5671 8084 5684 8114
rect 5699 8100 5729 8114
rect 5766 8084 5785 8114
rect 5800 8084 5806 8114
rect 5815 8084 5828 8114
rect 5843 8100 5873 8114
rect 5916 8100 5959 8114
rect 5966 8100 6186 8114
rect 6193 8100 6223 8114
rect 5883 8086 5898 8098
rect 5917 8086 5930 8100
rect 5998 8096 6151 8100
rect 5880 8084 5902 8086
rect 5980 8084 6172 8096
rect 6251 8084 6264 8114
rect 6279 8100 6309 8114
rect 6346 8084 6365 8114
rect 6380 8084 6386 8114
rect 6395 8084 6408 8114
rect 6423 8100 6453 8114
rect 6496 8100 6539 8114
rect 6546 8100 6766 8114
rect 6773 8100 6803 8114
rect 6463 8086 6478 8098
rect 6497 8086 6510 8100
rect 6578 8096 6731 8100
rect 6460 8084 6482 8086
rect 6560 8084 6752 8096
rect 6831 8084 6844 8114
rect 6859 8100 6889 8114
rect 6926 8084 6945 8114
rect 6960 8084 6966 8114
rect 6975 8084 6988 8114
rect 7003 8100 7033 8114
rect 7076 8100 7119 8114
rect 7126 8100 7346 8114
rect 7353 8100 7383 8114
rect 7043 8086 7058 8098
rect 7077 8086 7090 8100
rect 7158 8096 7311 8100
rect 7040 8084 7062 8086
rect 7140 8084 7332 8096
rect 7411 8084 7424 8114
rect 7439 8100 7469 8114
rect 7506 8084 7525 8114
rect 7540 8084 7546 8114
rect 7555 8084 7568 8114
rect 7583 8100 7613 8114
rect 7656 8100 7699 8114
rect 7706 8100 7926 8114
rect 7933 8100 7963 8114
rect 7623 8086 7638 8098
rect 7657 8086 7670 8100
rect 7738 8096 7891 8100
rect 7620 8084 7642 8086
rect 7720 8084 7912 8096
rect 7991 8084 8004 8114
rect 8019 8100 8049 8114
rect 8086 8084 8105 8114
rect 8120 8084 8126 8114
rect 8135 8084 8148 8114
rect 8163 8100 8193 8114
rect 8236 8100 8279 8114
rect 8286 8100 8506 8114
rect 8513 8100 8543 8114
rect 8203 8086 8218 8098
rect 8237 8086 8250 8100
rect 8318 8096 8471 8100
rect 8200 8084 8222 8086
rect 8300 8084 8492 8096
rect 8571 8084 8584 8114
rect 8599 8100 8629 8114
rect 8666 8084 8685 8114
rect 8700 8084 8706 8114
rect 8715 8084 8728 8114
rect 8743 8100 8773 8114
rect 8816 8100 8859 8114
rect 8866 8100 9086 8114
rect 9093 8100 9123 8114
rect 8783 8086 8798 8098
rect 8817 8086 8830 8100
rect 8898 8096 9051 8100
rect 8780 8084 8802 8086
rect 8880 8084 9072 8096
rect 9151 8084 9164 8114
rect 9179 8100 9209 8114
rect 9246 8084 9265 8114
rect 9280 8084 9286 8114
rect 9295 8084 9308 8114
rect 9323 8100 9353 8114
rect 9396 8100 9439 8114
rect 9446 8100 9666 8114
rect 9673 8100 9703 8114
rect 9363 8086 9378 8098
rect 9397 8086 9410 8100
rect 9478 8096 9631 8100
rect 9360 8084 9382 8086
rect 9460 8084 9652 8096
rect 9731 8084 9744 8114
rect 9759 8100 9789 8114
rect 9826 8084 9845 8114
rect 9860 8084 9866 8114
rect 9875 8084 9888 8114
rect 9903 8100 9933 8114
rect 9976 8100 10019 8114
rect 10026 8100 10246 8114
rect 10253 8100 10283 8114
rect 9943 8086 9958 8098
rect 9977 8086 9990 8100
rect 10058 8096 10211 8100
rect 9940 8084 9962 8086
rect 10040 8084 10232 8096
rect 10311 8084 10324 8114
rect 10339 8100 10369 8114
rect 10406 8084 10425 8114
rect 10440 8084 10446 8114
rect 10455 8084 10468 8114
rect 10483 8100 10513 8114
rect 10556 8100 10599 8114
rect 10606 8100 10826 8114
rect 10833 8100 10863 8114
rect 10523 8086 10538 8098
rect 10557 8086 10570 8100
rect 10638 8096 10791 8100
rect 10520 8084 10542 8086
rect 10620 8084 10812 8096
rect 10891 8084 10904 8114
rect 10919 8100 10949 8114
rect 10986 8084 11005 8114
rect 11020 8084 11026 8114
rect 11035 8084 11048 8114
rect 11063 8100 11093 8114
rect 11136 8100 11179 8114
rect 11186 8100 11406 8114
rect 11413 8100 11443 8114
rect 11103 8086 11118 8098
rect 11137 8086 11150 8100
rect 11218 8096 11371 8100
rect 11100 8084 11122 8086
rect 11200 8084 11392 8096
rect 11471 8084 11484 8114
rect 11499 8100 11529 8114
rect 11566 8084 11585 8114
rect 11600 8084 11606 8114
rect 11615 8084 11628 8114
rect 11643 8100 11673 8114
rect 11716 8100 11759 8114
rect 11766 8100 11986 8114
rect 11993 8100 12023 8114
rect 11683 8086 11698 8098
rect 11717 8086 11730 8100
rect 11798 8096 11951 8100
rect 11680 8084 11702 8086
rect 11780 8084 11972 8096
rect 12051 8084 12064 8114
rect 12079 8100 12109 8114
rect 12146 8084 12165 8114
rect 12180 8084 12186 8114
rect 12195 8084 12208 8114
rect 12223 8100 12253 8114
rect 12296 8100 12339 8114
rect 12346 8100 12566 8114
rect 12573 8100 12603 8114
rect 12263 8086 12278 8098
rect 12297 8086 12310 8100
rect 12378 8096 12531 8100
rect 12260 8084 12282 8086
rect 12360 8084 12552 8096
rect 12631 8084 12644 8114
rect 12659 8100 12689 8114
rect 12726 8084 12745 8114
rect 12760 8084 12766 8114
rect 12775 8084 12788 8114
rect 12803 8100 12833 8114
rect 12876 8100 12919 8114
rect 12926 8100 13146 8114
rect 13153 8100 13183 8114
rect 12843 8086 12858 8098
rect 12877 8086 12890 8100
rect 12958 8096 13111 8100
rect 12840 8084 12862 8086
rect 12940 8084 13132 8096
rect 13211 8084 13224 8114
rect 13239 8100 13269 8114
rect 13306 8084 13325 8114
rect 13340 8084 13346 8114
rect 13355 8084 13368 8114
rect 13383 8100 13413 8114
rect 13456 8100 13499 8114
rect 13506 8100 13726 8114
rect 13733 8100 13763 8114
rect 13423 8086 13438 8098
rect 13457 8086 13470 8100
rect 13538 8096 13691 8100
rect 13420 8084 13442 8086
rect 13520 8084 13712 8096
rect 13791 8084 13804 8114
rect 13819 8100 13849 8114
rect 13886 8084 13905 8114
rect 13920 8084 13926 8114
rect 13935 8084 13948 8114
rect 13963 8100 13993 8114
rect 14036 8100 14079 8114
rect 14086 8100 14306 8114
rect 14313 8100 14343 8114
rect 14003 8086 14018 8098
rect 14037 8086 14050 8100
rect 14118 8096 14271 8100
rect 14000 8084 14022 8086
rect 14100 8084 14292 8096
rect 14371 8084 14384 8114
rect 14399 8100 14429 8114
rect 14466 8084 14485 8114
rect 14500 8084 14506 8114
rect 14515 8084 14528 8114
rect 14543 8100 14573 8114
rect 14616 8100 14659 8114
rect 14666 8100 14886 8114
rect 14893 8100 14923 8114
rect 14583 8086 14598 8098
rect 14617 8086 14630 8100
rect 14698 8096 14851 8100
rect 14580 8084 14602 8086
rect 14680 8084 14872 8096
rect 14951 8084 14964 8114
rect 14979 8100 15009 8114
rect 15046 8084 15065 8114
rect 15080 8084 15086 8114
rect 15095 8084 15108 8114
rect 15123 8100 15153 8114
rect 15196 8100 15239 8114
rect 15246 8100 15466 8114
rect 15473 8100 15503 8114
rect 15163 8086 15178 8098
rect 15197 8086 15210 8100
rect 15278 8096 15431 8100
rect 15160 8084 15182 8086
rect 15260 8084 15452 8096
rect 15531 8084 15544 8114
rect 15559 8100 15589 8114
rect 15626 8084 15645 8114
rect 15660 8084 15666 8114
rect 15675 8084 15688 8114
rect 15703 8100 15733 8114
rect 15776 8100 15819 8114
rect 15826 8100 16046 8114
rect 16053 8100 16083 8114
rect 15743 8086 15758 8098
rect 15777 8086 15790 8100
rect 15858 8096 16011 8100
rect 15740 8084 15762 8086
rect 15840 8084 16032 8096
rect 16111 8084 16124 8114
rect 16139 8100 16169 8114
rect 16206 8084 16225 8114
rect 16240 8084 16246 8114
rect 16255 8084 16268 8114
rect 16283 8100 16313 8114
rect 16356 8100 16399 8114
rect 16406 8100 16626 8114
rect 16633 8100 16663 8114
rect 16323 8086 16338 8098
rect 16357 8086 16370 8100
rect 16438 8096 16591 8100
rect 16320 8084 16342 8086
rect 16420 8084 16612 8096
rect 16691 8084 16704 8114
rect 16719 8100 16749 8114
rect 16786 8084 16805 8114
rect 16820 8084 16826 8114
rect 16835 8084 16848 8114
rect 16863 8100 16893 8114
rect 16936 8100 16979 8114
rect 16986 8100 17206 8114
rect 17213 8100 17243 8114
rect 16903 8086 16918 8098
rect 16937 8086 16950 8100
rect 17018 8096 17171 8100
rect 16900 8084 16922 8086
rect 17000 8084 17192 8096
rect 17271 8084 17284 8114
rect 17299 8100 17329 8114
rect 17366 8084 17385 8114
rect 17400 8084 17406 8114
rect 17415 8084 17428 8114
rect 17443 8100 17473 8114
rect 17516 8100 17559 8114
rect 17566 8100 17786 8114
rect 17793 8100 17823 8114
rect 17483 8086 17498 8098
rect 17517 8086 17530 8100
rect 17598 8096 17751 8100
rect 17480 8084 17502 8086
rect 17580 8084 17772 8096
rect 17851 8084 17864 8114
rect 17879 8100 17909 8114
rect 17946 8084 17965 8114
rect 17980 8084 17986 8114
rect 17995 8084 18008 8114
rect 18023 8100 18053 8114
rect 18096 8100 18139 8114
rect 18146 8100 18366 8114
rect 18373 8100 18403 8114
rect 18063 8086 18078 8098
rect 18097 8086 18110 8100
rect 18178 8096 18331 8100
rect 18060 8084 18082 8086
rect 18160 8084 18352 8096
rect 18431 8084 18444 8114
rect 18459 8100 18489 8114
rect 18532 8084 18545 8114
rect 0 8070 18545 8084
rect 15 8000 28 8070
rect 80 8066 102 8070
rect 73 8044 102 8058
rect 155 8044 171 8058
rect 209 8054 215 8056
rect 222 8054 330 8070
rect 337 8054 343 8056
rect 351 8054 366 8070
rect 432 8064 451 8067
rect 73 8042 171 8044
rect 198 8042 366 8054
rect 381 8044 397 8058
rect 432 8045 454 8064
rect 464 8058 480 8059
rect 463 8056 480 8058
rect 464 8051 480 8056
rect 454 8044 460 8045
rect 463 8044 492 8051
rect 381 8043 492 8044
rect 381 8042 498 8043
rect 57 8034 108 8042
rect 155 8034 189 8042
rect 57 8022 82 8034
rect 89 8022 108 8034
rect 162 8032 189 8034
rect 198 8032 419 8042
rect 454 8039 460 8042
rect 162 8028 419 8032
rect 57 8014 108 8022
rect 155 8014 419 8028
rect 463 8034 498 8042
rect 9 7966 28 8000
rect 73 8006 102 8014
rect 73 8000 90 8006
rect 73 7998 107 8000
rect 155 7998 171 8014
rect 172 8004 380 8014
rect 381 8004 397 8014
rect 445 8010 460 8025
rect 463 8022 464 8034
rect 471 8022 498 8034
rect 463 8014 498 8022
rect 463 8013 492 8014
rect 183 8000 397 8004
rect 198 7998 397 8000
rect 432 8000 445 8010
rect 463 8000 480 8013
rect 432 7998 480 8000
rect 74 7994 107 7998
rect 70 7992 107 7994
rect 70 7991 137 7992
rect 70 7986 101 7991
rect 107 7986 137 7991
rect 70 7982 137 7986
rect 43 7979 137 7982
rect 43 7972 92 7979
rect 43 7966 73 7972
rect 92 7967 97 7972
rect 9 7950 89 7966
rect 101 7958 137 7979
rect 198 7974 387 7998
rect 432 7997 479 7998
rect 445 7992 479 7997
rect 213 7971 387 7974
rect 206 7968 387 7971
rect 415 7991 479 7992
rect 9 7948 28 7950
rect 43 7948 77 7950
rect 9 7932 89 7948
rect 9 7926 28 7932
rect -1 7910 28 7926
rect 43 7916 73 7932
rect 101 7910 107 7958
rect 110 7952 129 7958
rect 144 7952 174 7960
rect 110 7944 174 7952
rect 110 7928 190 7944
rect 206 7937 268 7968
rect 284 7937 346 7968
rect 415 7966 464 7991
rect 479 7966 509 7982
rect 378 7952 408 7960
rect 415 7958 525 7966
rect 378 7944 423 7952
rect 110 7926 129 7928
rect 144 7926 190 7928
rect 110 7910 190 7926
rect 217 7924 252 7937
rect 293 7934 330 7937
rect 293 7932 335 7934
rect 222 7921 252 7924
rect 231 7917 238 7921
rect 238 7916 239 7917
rect 197 7910 207 7916
rect -7 7902 34 7910
rect -7 7876 8 7902
rect 15 7876 34 7902
rect 98 7898 129 7910
rect 144 7898 247 7910
rect 259 7900 285 7926
rect 300 7921 330 7932
rect 362 7928 424 7944
rect 362 7926 408 7928
rect 362 7910 424 7926
rect 436 7910 442 7958
rect 445 7950 525 7958
rect 445 7948 464 7950
rect 479 7948 513 7950
rect 445 7932 525 7948
rect 445 7910 464 7932
rect 479 7916 509 7932
rect 537 7926 543 8000
rect 546 7926 565 8070
rect 580 7926 586 8070
rect 595 8000 608 8070
rect 660 8066 682 8070
rect 653 8044 682 8058
rect 735 8044 751 8058
rect 789 8054 795 8056
rect 802 8054 910 8070
rect 917 8054 923 8056
rect 931 8054 946 8070
rect 1012 8064 1031 8067
rect 653 8042 751 8044
rect 778 8042 946 8054
rect 961 8044 977 8058
rect 1012 8045 1034 8064
rect 1044 8058 1060 8059
rect 1043 8056 1060 8058
rect 1044 8051 1060 8056
rect 1034 8044 1040 8045
rect 1043 8044 1072 8051
rect 961 8043 1072 8044
rect 961 8042 1078 8043
rect 637 8034 688 8042
rect 735 8034 769 8042
rect 637 8022 662 8034
rect 669 8022 688 8034
rect 742 8032 769 8034
rect 778 8032 999 8042
rect 1034 8039 1040 8042
rect 742 8028 999 8032
rect 637 8014 688 8022
rect 735 8014 999 8028
rect 1043 8034 1078 8042
rect 589 7966 608 8000
rect 653 8006 682 8014
rect 653 8000 670 8006
rect 653 7998 687 8000
rect 735 7998 751 8014
rect 752 8004 960 8014
rect 961 8004 977 8014
rect 1025 8010 1040 8025
rect 1043 8022 1044 8034
rect 1051 8022 1078 8034
rect 1043 8014 1078 8022
rect 1043 8013 1072 8014
rect 763 8000 977 8004
rect 778 7998 977 8000
rect 1012 8000 1025 8010
rect 1043 8000 1060 8013
rect 1012 7998 1060 8000
rect 654 7994 687 7998
rect 650 7992 687 7994
rect 650 7991 717 7992
rect 650 7986 681 7991
rect 687 7986 717 7991
rect 650 7982 717 7986
rect 623 7979 717 7982
rect 623 7972 672 7979
rect 623 7966 653 7972
rect 672 7967 677 7972
rect 589 7950 669 7966
rect 681 7958 717 7979
rect 778 7974 967 7998
rect 1012 7997 1059 7998
rect 1025 7992 1059 7997
rect 793 7971 967 7974
rect 786 7968 967 7971
rect 995 7991 1059 7992
rect 589 7948 608 7950
rect 623 7948 657 7950
rect 589 7932 669 7948
rect 589 7926 608 7932
rect 305 7900 408 7910
rect 259 7898 408 7900
rect 429 7898 464 7910
rect 98 7896 260 7898
rect 110 7876 129 7896
rect 144 7894 174 7896
rect -7 7868 34 7876
rect 116 7872 129 7876
rect 181 7880 260 7896
rect 292 7896 464 7898
rect 292 7880 371 7896
rect 378 7894 408 7896
rect -1 7858 28 7868
rect 43 7858 73 7872
rect 116 7858 159 7872
rect 181 7868 371 7880
rect 436 7876 442 7896
rect 166 7858 196 7868
rect 197 7858 355 7868
rect 359 7858 389 7868
rect 393 7858 423 7872
rect 451 7858 464 7896
rect 536 7910 565 7926
rect 579 7910 608 7926
rect 623 7916 653 7932
rect 681 7910 687 7958
rect 690 7952 709 7958
rect 724 7952 754 7960
rect 690 7944 754 7952
rect 690 7928 770 7944
rect 786 7937 848 7968
rect 864 7937 926 7968
rect 995 7966 1044 7991
rect 1059 7966 1089 7982
rect 958 7952 988 7960
rect 995 7958 1105 7966
rect 958 7944 1003 7952
rect 690 7926 709 7928
rect 724 7926 770 7928
rect 690 7910 770 7926
rect 797 7924 832 7937
rect 873 7934 910 7937
rect 873 7932 915 7934
rect 802 7921 832 7924
rect 811 7917 818 7921
rect 818 7916 819 7917
rect 777 7910 787 7916
rect 536 7902 571 7910
rect 536 7876 537 7902
rect 544 7876 571 7902
rect 479 7858 509 7872
rect 536 7868 571 7876
rect 573 7902 614 7910
rect 573 7876 588 7902
rect 595 7876 614 7902
rect 678 7898 709 7910
rect 724 7898 827 7910
rect 839 7900 865 7926
rect 880 7921 910 7932
rect 942 7928 1004 7944
rect 942 7926 988 7928
rect 942 7910 1004 7926
rect 1016 7910 1022 7958
rect 1025 7950 1105 7958
rect 1025 7948 1044 7950
rect 1059 7948 1093 7950
rect 1025 7932 1105 7948
rect 1025 7910 1044 7932
rect 1059 7916 1089 7932
rect 1117 7926 1123 8000
rect 1126 7926 1145 8070
rect 1160 7926 1166 8070
rect 1175 8000 1188 8070
rect 1240 8066 1262 8070
rect 1233 8044 1262 8058
rect 1315 8044 1331 8058
rect 1369 8054 1375 8056
rect 1382 8054 1490 8070
rect 1497 8054 1503 8056
rect 1511 8054 1526 8070
rect 1592 8064 1611 8067
rect 1233 8042 1331 8044
rect 1358 8042 1526 8054
rect 1541 8044 1557 8058
rect 1592 8045 1614 8064
rect 1624 8058 1640 8059
rect 1623 8056 1640 8058
rect 1624 8051 1640 8056
rect 1614 8044 1620 8045
rect 1623 8044 1652 8051
rect 1541 8043 1652 8044
rect 1541 8042 1658 8043
rect 1217 8034 1268 8042
rect 1315 8034 1349 8042
rect 1217 8022 1242 8034
rect 1249 8022 1268 8034
rect 1322 8032 1349 8034
rect 1358 8032 1579 8042
rect 1614 8039 1620 8042
rect 1322 8028 1579 8032
rect 1217 8014 1268 8022
rect 1315 8014 1579 8028
rect 1623 8034 1658 8042
rect 1169 7966 1188 8000
rect 1233 8006 1262 8014
rect 1233 8000 1250 8006
rect 1233 7998 1267 8000
rect 1315 7998 1331 8014
rect 1332 8004 1540 8014
rect 1541 8004 1557 8014
rect 1605 8010 1620 8025
rect 1623 8022 1624 8034
rect 1631 8022 1658 8034
rect 1623 8014 1658 8022
rect 1623 8013 1652 8014
rect 1343 8000 1557 8004
rect 1358 7998 1557 8000
rect 1592 8000 1605 8010
rect 1623 8000 1640 8013
rect 1592 7998 1640 8000
rect 1234 7994 1267 7998
rect 1230 7992 1267 7994
rect 1230 7991 1297 7992
rect 1230 7986 1261 7991
rect 1267 7986 1297 7991
rect 1230 7982 1297 7986
rect 1203 7979 1297 7982
rect 1203 7972 1252 7979
rect 1203 7966 1233 7972
rect 1252 7967 1257 7972
rect 1169 7950 1249 7966
rect 1261 7958 1297 7979
rect 1358 7974 1547 7998
rect 1592 7997 1639 7998
rect 1605 7992 1639 7997
rect 1373 7971 1547 7974
rect 1366 7968 1547 7971
rect 1575 7991 1639 7992
rect 1169 7948 1188 7950
rect 1203 7948 1237 7950
rect 1169 7932 1249 7948
rect 1169 7926 1188 7932
rect 885 7900 988 7910
rect 839 7898 988 7900
rect 1009 7898 1044 7910
rect 678 7896 840 7898
rect 690 7876 709 7896
rect 724 7894 754 7896
rect 573 7868 614 7876
rect 696 7872 709 7876
rect 761 7880 840 7896
rect 872 7896 1044 7898
rect 872 7880 951 7896
rect 958 7894 988 7896
rect 536 7858 565 7868
rect 579 7858 608 7868
rect 623 7858 653 7872
rect 696 7858 739 7872
rect 761 7868 951 7880
rect 1016 7876 1022 7896
rect 746 7858 776 7868
rect 777 7858 935 7868
rect 939 7858 969 7868
rect 973 7858 1003 7872
rect 1031 7858 1044 7896
rect 1116 7910 1145 7926
rect 1159 7910 1188 7926
rect 1203 7916 1233 7932
rect 1261 7910 1267 7958
rect 1270 7952 1289 7958
rect 1304 7952 1334 7960
rect 1270 7944 1334 7952
rect 1270 7928 1350 7944
rect 1366 7937 1428 7968
rect 1444 7937 1506 7968
rect 1575 7966 1624 7991
rect 1639 7966 1669 7982
rect 1538 7952 1568 7960
rect 1575 7958 1685 7966
rect 1538 7944 1583 7952
rect 1270 7926 1289 7928
rect 1304 7926 1350 7928
rect 1270 7910 1350 7926
rect 1377 7924 1412 7937
rect 1453 7934 1490 7937
rect 1453 7932 1495 7934
rect 1382 7921 1412 7924
rect 1391 7917 1398 7921
rect 1398 7916 1399 7917
rect 1357 7910 1367 7916
rect 1116 7902 1151 7910
rect 1116 7876 1117 7902
rect 1124 7876 1151 7902
rect 1059 7858 1089 7872
rect 1116 7868 1151 7876
rect 1153 7902 1194 7910
rect 1153 7876 1168 7902
rect 1175 7876 1194 7902
rect 1258 7898 1289 7910
rect 1304 7898 1407 7910
rect 1419 7900 1445 7926
rect 1460 7921 1490 7932
rect 1522 7928 1584 7944
rect 1522 7926 1568 7928
rect 1522 7910 1584 7926
rect 1596 7910 1602 7958
rect 1605 7950 1685 7958
rect 1605 7948 1624 7950
rect 1639 7948 1673 7950
rect 1605 7932 1685 7948
rect 1605 7910 1624 7932
rect 1639 7916 1669 7932
rect 1697 7926 1703 8000
rect 1706 7926 1725 8070
rect 1740 7926 1746 8070
rect 1755 8000 1768 8070
rect 1820 8066 1842 8070
rect 1813 8044 1842 8058
rect 1895 8044 1911 8058
rect 1949 8054 1955 8056
rect 1962 8054 2070 8070
rect 2077 8054 2083 8056
rect 2091 8054 2106 8070
rect 2172 8064 2191 8067
rect 1813 8042 1911 8044
rect 1938 8042 2106 8054
rect 2121 8044 2137 8058
rect 2172 8045 2194 8064
rect 2204 8058 2220 8059
rect 2203 8056 2220 8058
rect 2204 8051 2220 8056
rect 2194 8044 2200 8045
rect 2203 8044 2232 8051
rect 2121 8043 2232 8044
rect 2121 8042 2238 8043
rect 1797 8034 1848 8042
rect 1895 8034 1929 8042
rect 1797 8022 1822 8034
rect 1829 8022 1848 8034
rect 1902 8032 1929 8034
rect 1938 8032 2159 8042
rect 2194 8039 2200 8042
rect 1902 8028 2159 8032
rect 1797 8014 1848 8022
rect 1895 8014 2159 8028
rect 2203 8034 2238 8042
rect 1749 7966 1768 8000
rect 1813 8006 1842 8014
rect 1813 8000 1830 8006
rect 1813 7998 1847 8000
rect 1895 7998 1911 8014
rect 1912 8004 2120 8014
rect 2121 8004 2137 8014
rect 2185 8010 2200 8025
rect 2203 8022 2204 8034
rect 2211 8022 2238 8034
rect 2203 8014 2238 8022
rect 2203 8013 2232 8014
rect 1923 8000 2137 8004
rect 1938 7998 2137 8000
rect 2172 8000 2185 8010
rect 2203 8000 2220 8013
rect 2172 7998 2220 8000
rect 1814 7994 1847 7998
rect 1810 7992 1847 7994
rect 1810 7991 1877 7992
rect 1810 7986 1841 7991
rect 1847 7986 1877 7991
rect 1810 7982 1877 7986
rect 1783 7979 1877 7982
rect 1783 7972 1832 7979
rect 1783 7966 1813 7972
rect 1832 7967 1837 7972
rect 1749 7950 1829 7966
rect 1841 7958 1877 7979
rect 1938 7974 2127 7998
rect 2172 7997 2219 7998
rect 2185 7992 2219 7997
rect 1953 7971 2127 7974
rect 1946 7968 2127 7971
rect 2155 7991 2219 7992
rect 1749 7948 1768 7950
rect 1783 7948 1817 7950
rect 1749 7932 1829 7948
rect 1749 7926 1768 7932
rect 1465 7900 1568 7910
rect 1419 7898 1568 7900
rect 1589 7898 1624 7910
rect 1258 7896 1420 7898
rect 1270 7876 1289 7896
rect 1304 7894 1334 7896
rect 1153 7868 1194 7876
rect 1276 7872 1289 7876
rect 1341 7880 1420 7896
rect 1452 7896 1624 7898
rect 1452 7880 1531 7896
rect 1538 7894 1568 7896
rect 1116 7858 1145 7868
rect 1159 7858 1188 7868
rect 1203 7858 1233 7872
rect 1276 7858 1319 7872
rect 1341 7868 1531 7880
rect 1596 7876 1602 7896
rect 1326 7858 1356 7868
rect 1357 7858 1515 7868
rect 1519 7858 1549 7868
rect 1553 7858 1583 7872
rect 1611 7858 1624 7896
rect 1696 7910 1725 7926
rect 1739 7910 1768 7926
rect 1783 7916 1813 7932
rect 1841 7910 1847 7958
rect 1850 7952 1869 7958
rect 1884 7952 1914 7960
rect 1850 7944 1914 7952
rect 1850 7928 1930 7944
rect 1946 7937 2008 7968
rect 2024 7937 2086 7968
rect 2155 7966 2204 7991
rect 2219 7966 2249 7982
rect 2118 7952 2148 7960
rect 2155 7958 2265 7966
rect 2118 7944 2163 7952
rect 1850 7926 1869 7928
rect 1884 7926 1930 7928
rect 1850 7910 1930 7926
rect 1957 7924 1992 7937
rect 2033 7934 2070 7937
rect 2033 7932 2075 7934
rect 1962 7921 1992 7924
rect 1971 7917 1978 7921
rect 1978 7916 1979 7917
rect 1937 7910 1947 7916
rect 1696 7902 1731 7910
rect 1696 7876 1697 7902
rect 1704 7876 1731 7902
rect 1639 7858 1669 7872
rect 1696 7868 1731 7876
rect 1733 7902 1774 7910
rect 1733 7876 1748 7902
rect 1755 7876 1774 7902
rect 1838 7898 1869 7910
rect 1884 7898 1987 7910
rect 1999 7900 2025 7926
rect 2040 7921 2070 7932
rect 2102 7928 2164 7944
rect 2102 7926 2148 7928
rect 2102 7910 2164 7926
rect 2176 7910 2182 7958
rect 2185 7950 2265 7958
rect 2185 7948 2204 7950
rect 2219 7948 2253 7950
rect 2185 7932 2265 7948
rect 2185 7910 2204 7932
rect 2219 7916 2249 7932
rect 2277 7926 2283 8000
rect 2286 7926 2305 8070
rect 2320 7926 2326 8070
rect 2335 8000 2348 8070
rect 2400 8066 2422 8070
rect 2393 8044 2422 8058
rect 2475 8044 2491 8058
rect 2529 8054 2535 8056
rect 2542 8054 2650 8070
rect 2657 8054 2663 8056
rect 2671 8054 2686 8070
rect 2752 8064 2771 8067
rect 2393 8042 2491 8044
rect 2518 8042 2686 8054
rect 2701 8044 2717 8058
rect 2752 8045 2774 8064
rect 2784 8058 2800 8059
rect 2783 8056 2800 8058
rect 2784 8051 2800 8056
rect 2774 8044 2780 8045
rect 2783 8044 2812 8051
rect 2701 8043 2812 8044
rect 2701 8042 2818 8043
rect 2377 8034 2428 8042
rect 2475 8034 2509 8042
rect 2377 8022 2402 8034
rect 2409 8022 2428 8034
rect 2482 8032 2509 8034
rect 2518 8032 2739 8042
rect 2774 8039 2780 8042
rect 2482 8028 2739 8032
rect 2377 8014 2428 8022
rect 2475 8014 2739 8028
rect 2783 8034 2818 8042
rect 2329 7966 2348 8000
rect 2393 8006 2422 8014
rect 2393 8000 2410 8006
rect 2393 7998 2427 8000
rect 2475 7998 2491 8014
rect 2492 8004 2700 8014
rect 2701 8004 2717 8014
rect 2765 8010 2780 8025
rect 2783 8022 2784 8034
rect 2791 8022 2818 8034
rect 2783 8014 2818 8022
rect 2783 8013 2812 8014
rect 2503 8000 2717 8004
rect 2518 7998 2717 8000
rect 2752 8000 2765 8010
rect 2783 8000 2800 8013
rect 2752 7998 2800 8000
rect 2394 7994 2427 7998
rect 2390 7992 2427 7994
rect 2390 7991 2457 7992
rect 2390 7986 2421 7991
rect 2427 7986 2457 7991
rect 2390 7982 2457 7986
rect 2363 7979 2457 7982
rect 2363 7972 2412 7979
rect 2363 7966 2393 7972
rect 2412 7967 2417 7972
rect 2329 7950 2409 7966
rect 2421 7958 2457 7979
rect 2518 7974 2707 7998
rect 2752 7997 2799 7998
rect 2765 7992 2799 7997
rect 2533 7971 2707 7974
rect 2526 7968 2707 7971
rect 2735 7991 2799 7992
rect 2329 7948 2348 7950
rect 2363 7948 2397 7950
rect 2329 7932 2409 7948
rect 2329 7926 2348 7932
rect 2045 7900 2148 7910
rect 1999 7898 2148 7900
rect 2169 7898 2204 7910
rect 1838 7896 2000 7898
rect 1850 7876 1869 7896
rect 1884 7894 1914 7896
rect 1733 7868 1774 7876
rect 1856 7872 1869 7876
rect 1921 7880 2000 7896
rect 2032 7896 2204 7898
rect 2032 7880 2111 7896
rect 2118 7894 2148 7896
rect 1696 7858 1725 7868
rect 1739 7858 1768 7868
rect 1783 7858 1813 7872
rect 1856 7858 1899 7872
rect 1921 7868 2111 7880
rect 2176 7876 2182 7896
rect 1906 7858 1936 7868
rect 1937 7858 2095 7868
rect 2099 7858 2129 7868
rect 2133 7858 2163 7872
rect 2191 7858 2204 7896
rect 2276 7910 2305 7926
rect 2319 7910 2348 7926
rect 2363 7916 2393 7932
rect 2421 7910 2427 7958
rect 2430 7952 2449 7958
rect 2464 7952 2494 7960
rect 2430 7944 2494 7952
rect 2430 7928 2510 7944
rect 2526 7937 2588 7968
rect 2604 7937 2666 7968
rect 2735 7966 2784 7991
rect 2799 7966 2829 7982
rect 2698 7952 2728 7960
rect 2735 7958 2845 7966
rect 2698 7944 2743 7952
rect 2430 7926 2449 7928
rect 2464 7926 2510 7928
rect 2430 7910 2510 7926
rect 2537 7924 2572 7937
rect 2613 7934 2650 7937
rect 2613 7932 2655 7934
rect 2542 7921 2572 7924
rect 2551 7917 2558 7921
rect 2558 7916 2559 7917
rect 2517 7910 2527 7916
rect 2276 7902 2311 7910
rect 2276 7876 2277 7902
rect 2284 7876 2311 7902
rect 2219 7858 2249 7872
rect 2276 7868 2311 7876
rect 2313 7902 2354 7910
rect 2313 7876 2328 7902
rect 2335 7876 2354 7902
rect 2418 7898 2449 7910
rect 2464 7898 2567 7910
rect 2579 7900 2605 7926
rect 2620 7921 2650 7932
rect 2682 7928 2744 7944
rect 2682 7926 2728 7928
rect 2682 7910 2744 7926
rect 2756 7910 2762 7958
rect 2765 7950 2845 7958
rect 2765 7948 2784 7950
rect 2799 7948 2833 7950
rect 2765 7932 2845 7948
rect 2765 7910 2784 7932
rect 2799 7916 2829 7932
rect 2857 7926 2863 8000
rect 2866 7926 2885 8070
rect 2900 7926 2906 8070
rect 2915 8000 2928 8070
rect 2980 8066 3002 8070
rect 2973 8044 3002 8058
rect 3055 8044 3071 8058
rect 3109 8054 3115 8056
rect 3122 8054 3230 8070
rect 3237 8054 3243 8056
rect 3251 8054 3266 8070
rect 3332 8064 3351 8067
rect 2973 8042 3071 8044
rect 3098 8042 3266 8054
rect 3281 8044 3297 8058
rect 3332 8045 3354 8064
rect 3364 8058 3380 8059
rect 3363 8056 3380 8058
rect 3364 8051 3380 8056
rect 3354 8044 3360 8045
rect 3363 8044 3392 8051
rect 3281 8043 3392 8044
rect 3281 8042 3398 8043
rect 2957 8034 3008 8042
rect 3055 8034 3089 8042
rect 2957 8022 2982 8034
rect 2989 8022 3008 8034
rect 3062 8032 3089 8034
rect 3098 8032 3319 8042
rect 3354 8039 3360 8042
rect 3062 8028 3319 8032
rect 2957 8014 3008 8022
rect 3055 8014 3319 8028
rect 3363 8034 3398 8042
rect 2909 7966 2928 8000
rect 2973 8006 3002 8014
rect 2973 8000 2990 8006
rect 2973 7998 3007 8000
rect 3055 7998 3071 8014
rect 3072 8004 3280 8014
rect 3281 8004 3297 8014
rect 3345 8010 3360 8025
rect 3363 8022 3364 8034
rect 3371 8022 3398 8034
rect 3363 8014 3398 8022
rect 3363 8013 3392 8014
rect 3083 8000 3297 8004
rect 3098 7998 3297 8000
rect 3332 8000 3345 8010
rect 3363 8000 3380 8013
rect 3332 7998 3380 8000
rect 2974 7994 3007 7998
rect 2970 7992 3007 7994
rect 2970 7991 3037 7992
rect 2970 7986 3001 7991
rect 3007 7986 3037 7991
rect 2970 7982 3037 7986
rect 2943 7979 3037 7982
rect 2943 7972 2992 7979
rect 2943 7966 2973 7972
rect 2992 7967 2997 7972
rect 2909 7950 2989 7966
rect 3001 7958 3037 7979
rect 3098 7974 3287 7998
rect 3332 7997 3379 7998
rect 3345 7992 3379 7997
rect 3113 7971 3287 7974
rect 3106 7968 3287 7971
rect 3315 7991 3379 7992
rect 2909 7948 2928 7950
rect 2943 7948 2977 7950
rect 2909 7932 2989 7948
rect 2909 7926 2928 7932
rect 2625 7900 2728 7910
rect 2579 7898 2728 7900
rect 2749 7898 2784 7910
rect 2418 7896 2580 7898
rect 2430 7876 2449 7896
rect 2464 7894 2494 7896
rect 2313 7868 2354 7876
rect 2436 7872 2449 7876
rect 2501 7880 2580 7896
rect 2612 7896 2784 7898
rect 2612 7880 2691 7896
rect 2698 7894 2728 7896
rect 2276 7858 2305 7868
rect 2319 7858 2348 7868
rect 2363 7858 2393 7872
rect 2436 7858 2479 7872
rect 2501 7868 2691 7880
rect 2756 7876 2762 7896
rect 2486 7858 2516 7868
rect 2517 7858 2675 7868
rect 2679 7858 2709 7868
rect 2713 7858 2743 7872
rect 2771 7858 2784 7896
rect 2856 7910 2885 7926
rect 2899 7910 2928 7926
rect 2943 7916 2973 7932
rect 3001 7910 3007 7958
rect 3010 7952 3029 7958
rect 3044 7952 3074 7960
rect 3010 7944 3074 7952
rect 3010 7928 3090 7944
rect 3106 7937 3168 7968
rect 3184 7937 3246 7968
rect 3315 7966 3364 7991
rect 3379 7966 3409 7982
rect 3278 7952 3308 7960
rect 3315 7958 3425 7966
rect 3278 7944 3323 7952
rect 3010 7926 3029 7928
rect 3044 7926 3090 7928
rect 3010 7910 3090 7926
rect 3117 7924 3152 7937
rect 3193 7934 3230 7937
rect 3193 7932 3235 7934
rect 3122 7921 3152 7924
rect 3131 7917 3138 7921
rect 3138 7916 3139 7917
rect 3097 7910 3107 7916
rect 2856 7902 2891 7910
rect 2856 7876 2857 7902
rect 2864 7876 2891 7902
rect 2799 7858 2829 7872
rect 2856 7868 2891 7876
rect 2893 7902 2934 7910
rect 2893 7876 2908 7902
rect 2915 7876 2934 7902
rect 2998 7898 3029 7910
rect 3044 7898 3147 7910
rect 3159 7900 3185 7926
rect 3200 7921 3230 7932
rect 3262 7928 3324 7944
rect 3262 7926 3308 7928
rect 3262 7910 3324 7926
rect 3336 7910 3342 7958
rect 3345 7950 3425 7958
rect 3345 7948 3364 7950
rect 3379 7948 3413 7950
rect 3345 7932 3425 7948
rect 3345 7910 3364 7932
rect 3379 7916 3409 7932
rect 3437 7926 3443 8000
rect 3446 7926 3465 8070
rect 3480 7926 3486 8070
rect 3495 8000 3508 8070
rect 3560 8066 3582 8070
rect 3553 8044 3582 8058
rect 3635 8044 3651 8058
rect 3689 8054 3695 8056
rect 3702 8054 3810 8070
rect 3817 8054 3823 8056
rect 3831 8054 3846 8070
rect 3912 8064 3931 8067
rect 3553 8042 3651 8044
rect 3678 8042 3846 8054
rect 3861 8044 3877 8058
rect 3912 8045 3934 8064
rect 3944 8058 3960 8059
rect 3943 8056 3960 8058
rect 3944 8051 3960 8056
rect 3934 8044 3940 8045
rect 3943 8044 3972 8051
rect 3861 8043 3972 8044
rect 3861 8042 3978 8043
rect 3537 8034 3588 8042
rect 3635 8034 3669 8042
rect 3537 8022 3562 8034
rect 3569 8022 3588 8034
rect 3642 8032 3669 8034
rect 3678 8032 3899 8042
rect 3934 8039 3940 8042
rect 3642 8028 3899 8032
rect 3537 8014 3588 8022
rect 3635 8014 3899 8028
rect 3943 8034 3978 8042
rect 3489 7966 3508 8000
rect 3553 8006 3582 8014
rect 3553 8000 3570 8006
rect 3553 7998 3587 8000
rect 3635 7998 3651 8014
rect 3652 8004 3860 8014
rect 3861 8004 3877 8014
rect 3925 8010 3940 8025
rect 3943 8022 3944 8034
rect 3951 8022 3978 8034
rect 3943 8014 3978 8022
rect 3943 8013 3972 8014
rect 3663 8000 3877 8004
rect 3678 7998 3877 8000
rect 3912 8000 3925 8010
rect 3943 8000 3960 8013
rect 3912 7998 3960 8000
rect 3554 7994 3587 7998
rect 3550 7992 3587 7994
rect 3550 7991 3617 7992
rect 3550 7986 3581 7991
rect 3587 7986 3617 7991
rect 3550 7982 3617 7986
rect 3523 7979 3617 7982
rect 3523 7972 3572 7979
rect 3523 7966 3553 7972
rect 3572 7967 3577 7972
rect 3489 7950 3569 7966
rect 3581 7958 3617 7979
rect 3678 7974 3867 7998
rect 3912 7997 3959 7998
rect 3925 7992 3959 7997
rect 3693 7971 3867 7974
rect 3686 7968 3867 7971
rect 3895 7991 3959 7992
rect 3489 7948 3508 7950
rect 3523 7948 3557 7950
rect 3489 7932 3569 7948
rect 3489 7926 3508 7932
rect 3205 7900 3308 7910
rect 3159 7898 3308 7900
rect 3329 7898 3364 7910
rect 2998 7896 3160 7898
rect 3010 7876 3029 7896
rect 3044 7894 3074 7896
rect 2893 7868 2934 7876
rect 3016 7872 3029 7876
rect 3081 7880 3160 7896
rect 3192 7896 3364 7898
rect 3192 7880 3271 7896
rect 3278 7894 3308 7896
rect 2856 7858 2885 7868
rect 2899 7858 2928 7868
rect 2943 7858 2973 7872
rect 3016 7858 3059 7872
rect 3081 7868 3271 7880
rect 3336 7876 3342 7896
rect 3066 7858 3096 7868
rect 3097 7858 3255 7868
rect 3259 7858 3289 7868
rect 3293 7858 3323 7872
rect 3351 7858 3364 7896
rect 3436 7910 3465 7926
rect 3479 7910 3508 7926
rect 3523 7916 3553 7932
rect 3581 7910 3587 7958
rect 3590 7952 3609 7958
rect 3624 7952 3654 7960
rect 3590 7944 3654 7952
rect 3590 7928 3670 7944
rect 3686 7937 3748 7968
rect 3764 7937 3826 7968
rect 3895 7966 3944 7991
rect 3959 7966 3989 7982
rect 3858 7952 3888 7960
rect 3895 7958 4005 7966
rect 3858 7944 3903 7952
rect 3590 7926 3609 7928
rect 3624 7926 3670 7928
rect 3590 7910 3670 7926
rect 3697 7924 3732 7937
rect 3773 7934 3810 7937
rect 3773 7932 3815 7934
rect 3702 7921 3732 7924
rect 3711 7917 3718 7921
rect 3718 7916 3719 7917
rect 3677 7910 3687 7916
rect 3436 7902 3471 7910
rect 3436 7876 3437 7902
rect 3444 7876 3471 7902
rect 3379 7858 3409 7872
rect 3436 7868 3471 7876
rect 3473 7902 3514 7910
rect 3473 7876 3488 7902
rect 3495 7876 3514 7902
rect 3578 7898 3609 7910
rect 3624 7898 3727 7910
rect 3739 7900 3765 7926
rect 3780 7921 3810 7932
rect 3842 7928 3904 7944
rect 3842 7926 3888 7928
rect 3842 7910 3904 7926
rect 3916 7910 3922 7958
rect 3925 7950 4005 7958
rect 3925 7948 3944 7950
rect 3959 7948 3993 7950
rect 3925 7932 4005 7948
rect 3925 7910 3944 7932
rect 3959 7916 3989 7932
rect 4017 7926 4023 8000
rect 4026 7926 4045 8070
rect 4060 7926 4066 8070
rect 4075 8000 4088 8070
rect 4140 8066 4162 8070
rect 4133 8044 4162 8058
rect 4215 8044 4231 8058
rect 4269 8054 4275 8056
rect 4282 8054 4390 8070
rect 4397 8054 4403 8056
rect 4411 8054 4426 8070
rect 4492 8064 4511 8067
rect 4133 8042 4231 8044
rect 4258 8042 4426 8054
rect 4441 8044 4457 8058
rect 4492 8045 4514 8064
rect 4524 8058 4540 8059
rect 4523 8056 4540 8058
rect 4524 8051 4540 8056
rect 4514 8044 4520 8045
rect 4523 8044 4552 8051
rect 4441 8043 4552 8044
rect 4441 8042 4558 8043
rect 4117 8034 4168 8042
rect 4215 8034 4249 8042
rect 4117 8022 4142 8034
rect 4149 8022 4168 8034
rect 4222 8032 4249 8034
rect 4258 8032 4479 8042
rect 4514 8039 4520 8042
rect 4222 8028 4479 8032
rect 4117 8014 4168 8022
rect 4215 8014 4479 8028
rect 4523 8034 4558 8042
rect 4069 7966 4088 8000
rect 4133 8006 4162 8014
rect 4133 8000 4150 8006
rect 4133 7998 4167 8000
rect 4215 7998 4231 8014
rect 4232 8004 4440 8014
rect 4441 8004 4457 8014
rect 4505 8010 4520 8025
rect 4523 8022 4524 8034
rect 4531 8022 4558 8034
rect 4523 8014 4558 8022
rect 4523 8013 4552 8014
rect 4243 8000 4457 8004
rect 4258 7998 4457 8000
rect 4492 8000 4505 8010
rect 4523 8000 4540 8013
rect 4492 7998 4540 8000
rect 4134 7994 4167 7998
rect 4130 7992 4167 7994
rect 4130 7991 4197 7992
rect 4130 7986 4161 7991
rect 4167 7986 4197 7991
rect 4130 7982 4197 7986
rect 4103 7979 4197 7982
rect 4103 7972 4152 7979
rect 4103 7966 4133 7972
rect 4152 7967 4157 7972
rect 4069 7950 4149 7966
rect 4161 7958 4197 7979
rect 4258 7974 4447 7998
rect 4492 7997 4539 7998
rect 4505 7992 4539 7997
rect 4273 7971 4447 7974
rect 4266 7968 4447 7971
rect 4475 7991 4539 7992
rect 4069 7948 4088 7950
rect 4103 7948 4137 7950
rect 4069 7932 4149 7948
rect 4069 7926 4088 7932
rect 3785 7900 3888 7910
rect 3739 7898 3888 7900
rect 3909 7898 3944 7910
rect 3578 7896 3740 7898
rect 3590 7876 3609 7896
rect 3624 7894 3654 7896
rect 3473 7868 3514 7876
rect 3596 7872 3609 7876
rect 3661 7880 3740 7896
rect 3772 7896 3944 7898
rect 3772 7880 3851 7896
rect 3858 7894 3888 7896
rect 3436 7858 3465 7868
rect 3479 7858 3508 7868
rect 3523 7858 3553 7872
rect 3596 7858 3639 7872
rect 3661 7868 3851 7880
rect 3916 7876 3922 7896
rect 3646 7858 3676 7868
rect 3677 7858 3835 7868
rect 3839 7858 3869 7868
rect 3873 7858 3903 7872
rect 3931 7858 3944 7896
rect 4016 7910 4045 7926
rect 4059 7910 4088 7926
rect 4103 7916 4133 7932
rect 4161 7910 4167 7958
rect 4170 7952 4189 7958
rect 4204 7952 4234 7960
rect 4170 7944 4234 7952
rect 4170 7928 4250 7944
rect 4266 7937 4328 7968
rect 4344 7937 4406 7968
rect 4475 7966 4524 7991
rect 4539 7966 4569 7982
rect 4438 7952 4468 7960
rect 4475 7958 4585 7966
rect 4438 7944 4483 7952
rect 4170 7926 4189 7928
rect 4204 7926 4250 7928
rect 4170 7910 4250 7926
rect 4277 7924 4312 7937
rect 4353 7934 4390 7937
rect 4353 7932 4395 7934
rect 4282 7921 4312 7924
rect 4291 7917 4298 7921
rect 4298 7916 4299 7917
rect 4257 7910 4267 7916
rect 4016 7902 4051 7910
rect 4016 7876 4017 7902
rect 4024 7876 4051 7902
rect 3959 7858 3989 7872
rect 4016 7868 4051 7876
rect 4053 7902 4094 7910
rect 4053 7876 4068 7902
rect 4075 7876 4094 7902
rect 4158 7898 4189 7910
rect 4204 7898 4307 7910
rect 4319 7900 4345 7926
rect 4360 7921 4390 7932
rect 4422 7928 4484 7944
rect 4422 7926 4468 7928
rect 4422 7910 4484 7926
rect 4496 7910 4502 7958
rect 4505 7950 4585 7958
rect 4505 7948 4524 7950
rect 4539 7948 4573 7950
rect 4505 7932 4585 7948
rect 4505 7910 4524 7932
rect 4539 7916 4569 7932
rect 4597 7926 4603 8000
rect 4606 7926 4625 8070
rect 4640 7926 4646 8070
rect 4655 8000 4668 8070
rect 4720 8066 4742 8070
rect 4713 8044 4742 8058
rect 4795 8044 4811 8058
rect 4849 8054 4855 8056
rect 4862 8054 4970 8070
rect 4977 8054 4983 8056
rect 4991 8054 5006 8070
rect 5072 8064 5091 8067
rect 4713 8042 4811 8044
rect 4838 8042 5006 8054
rect 5021 8044 5037 8058
rect 5072 8045 5094 8064
rect 5104 8058 5120 8059
rect 5103 8056 5120 8058
rect 5104 8051 5120 8056
rect 5094 8044 5100 8045
rect 5103 8044 5132 8051
rect 5021 8043 5132 8044
rect 5021 8042 5138 8043
rect 4697 8034 4748 8042
rect 4795 8034 4829 8042
rect 4697 8022 4722 8034
rect 4729 8022 4748 8034
rect 4802 8032 4829 8034
rect 4838 8032 5059 8042
rect 5094 8039 5100 8042
rect 4802 8028 5059 8032
rect 4697 8014 4748 8022
rect 4795 8014 5059 8028
rect 5103 8034 5138 8042
rect 4649 7966 4668 8000
rect 4713 8006 4742 8014
rect 4713 8000 4730 8006
rect 4713 7998 4747 8000
rect 4795 7998 4811 8014
rect 4812 8004 5020 8014
rect 5021 8004 5037 8014
rect 5085 8010 5100 8025
rect 5103 8022 5104 8034
rect 5111 8022 5138 8034
rect 5103 8014 5138 8022
rect 5103 8013 5132 8014
rect 4823 8000 5037 8004
rect 4838 7998 5037 8000
rect 5072 8000 5085 8010
rect 5103 8000 5120 8013
rect 5072 7998 5120 8000
rect 4714 7994 4747 7998
rect 4710 7992 4747 7994
rect 4710 7991 4777 7992
rect 4710 7986 4741 7991
rect 4747 7986 4777 7991
rect 4710 7982 4777 7986
rect 4683 7979 4777 7982
rect 4683 7972 4732 7979
rect 4683 7966 4713 7972
rect 4732 7967 4737 7972
rect 4649 7950 4729 7966
rect 4741 7958 4777 7979
rect 4838 7974 5027 7998
rect 5072 7997 5119 7998
rect 5085 7992 5119 7997
rect 4853 7971 5027 7974
rect 4846 7968 5027 7971
rect 5055 7991 5119 7992
rect 4649 7948 4668 7950
rect 4683 7948 4717 7950
rect 4649 7932 4729 7948
rect 4649 7926 4668 7932
rect 4365 7900 4468 7910
rect 4319 7898 4468 7900
rect 4489 7898 4524 7910
rect 4158 7896 4320 7898
rect 4170 7876 4189 7896
rect 4204 7894 4234 7896
rect 4053 7868 4094 7876
rect 4176 7872 4189 7876
rect 4241 7880 4320 7896
rect 4352 7896 4524 7898
rect 4352 7880 4431 7896
rect 4438 7894 4468 7896
rect 4016 7858 4045 7868
rect 4059 7858 4088 7868
rect 4103 7858 4133 7872
rect 4176 7858 4219 7872
rect 4241 7868 4431 7880
rect 4496 7876 4502 7896
rect 4226 7858 4256 7868
rect 4257 7858 4415 7868
rect 4419 7858 4449 7868
rect 4453 7858 4483 7872
rect 4511 7858 4524 7896
rect 4596 7910 4625 7926
rect 4639 7910 4668 7926
rect 4683 7916 4713 7932
rect 4741 7910 4747 7958
rect 4750 7952 4769 7958
rect 4784 7952 4814 7960
rect 4750 7944 4814 7952
rect 4750 7928 4830 7944
rect 4846 7937 4908 7968
rect 4924 7937 4986 7968
rect 5055 7966 5104 7991
rect 5119 7966 5149 7982
rect 5018 7952 5048 7960
rect 5055 7958 5165 7966
rect 5018 7944 5063 7952
rect 4750 7926 4769 7928
rect 4784 7926 4830 7928
rect 4750 7910 4830 7926
rect 4857 7924 4892 7937
rect 4933 7934 4970 7937
rect 4933 7932 4975 7934
rect 4862 7921 4892 7924
rect 4871 7917 4878 7921
rect 4878 7916 4879 7917
rect 4837 7910 4847 7916
rect 4596 7902 4631 7910
rect 4596 7876 4597 7902
rect 4604 7876 4631 7902
rect 4539 7858 4569 7872
rect 4596 7868 4631 7876
rect 4633 7902 4674 7910
rect 4633 7876 4648 7902
rect 4655 7876 4674 7902
rect 4738 7898 4769 7910
rect 4784 7898 4887 7910
rect 4899 7900 4925 7926
rect 4940 7921 4970 7932
rect 5002 7928 5064 7944
rect 5002 7926 5048 7928
rect 5002 7910 5064 7926
rect 5076 7910 5082 7958
rect 5085 7950 5165 7958
rect 5085 7948 5104 7950
rect 5119 7948 5153 7950
rect 5085 7932 5165 7948
rect 5085 7910 5104 7932
rect 5119 7916 5149 7932
rect 5177 7926 5183 8000
rect 5186 7926 5205 8070
rect 5220 7926 5226 8070
rect 5235 8000 5248 8070
rect 5300 8066 5322 8070
rect 5293 8044 5322 8058
rect 5375 8044 5391 8058
rect 5429 8054 5435 8056
rect 5442 8054 5550 8070
rect 5557 8054 5563 8056
rect 5571 8054 5586 8070
rect 5652 8064 5671 8067
rect 5293 8042 5391 8044
rect 5418 8042 5586 8054
rect 5601 8044 5617 8058
rect 5652 8045 5674 8064
rect 5684 8058 5700 8059
rect 5683 8056 5700 8058
rect 5684 8051 5700 8056
rect 5674 8044 5680 8045
rect 5683 8044 5712 8051
rect 5601 8043 5712 8044
rect 5601 8042 5718 8043
rect 5277 8034 5328 8042
rect 5375 8034 5409 8042
rect 5277 8022 5302 8034
rect 5309 8022 5328 8034
rect 5382 8032 5409 8034
rect 5418 8032 5639 8042
rect 5674 8039 5680 8042
rect 5382 8028 5639 8032
rect 5277 8014 5328 8022
rect 5375 8014 5639 8028
rect 5683 8034 5718 8042
rect 5229 7966 5248 8000
rect 5293 8006 5322 8014
rect 5293 8000 5310 8006
rect 5293 7998 5327 8000
rect 5375 7998 5391 8014
rect 5392 8004 5600 8014
rect 5601 8004 5617 8014
rect 5665 8010 5680 8025
rect 5683 8022 5684 8034
rect 5691 8022 5718 8034
rect 5683 8014 5718 8022
rect 5683 8013 5712 8014
rect 5403 8000 5617 8004
rect 5418 7998 5617 8000
rect 5652 8000 5665 8010
rect 5683 8000 5700 8013
rect 5652 7998 5700 8000
rect 5294 7994 5327 7998
rect 5290 7992 5327 7994
rect 5290 7991 5357 7992
rect 5290 7986 5321 7991
rect 5327 7986 5357 7991
rect 5290 7982 5357 7986
rect 5263 7979 5357 7982
rect 5263 7972 5312 7979
rect 5263 7966 5293 7972
rect 5312 7967 5317 7972
rect 5229 7950 5309 7966
rect 5321 7958 5357 7979
rect 5418 7974 5607 7998
rect 5652 7997 5699 7998
rect 5665 7992 5699 7997
rect 5433 7971 5607 7974
rect 5426 7968 5607 7971
rect 5635 7991 5699 7992
rect 5229 7948 5248 7950
rect 5263 7948 5297 7950
rect 5229 7932 5309 7948
rect 5229 7926 5248 7932
rect 4945 7900 5048 7910
rect 4899 7898 5048 7900
rect 5069 7898 5104 7910
rect 4738 7896 4900 7898
rect 4750 7876 4769 7896
rect 4784 7894 4814 7896
rect 4633 7868 4674 7876
rect 4756 7872 4769 7876
rect 4821 7880 4900 7896
rect 4932 7896 5104 7898
rect 4932 7880 5011 7896
rect 5018 7894 5048 7896
rect 4596 7858 4625 7868
rect 4639 7858 4668 7868
rect 4683 7858 4713 7872
rect 4756 7858 4799 7872
rect 4821 7868 5011 7880
rect 5076 7876 5082 7896
rect 4806 7858 4836 7868
rect 4837 7858 4995 7868
rect 4999 7858 5029 7868
rect 5033 7858 5063 7872
rect 5091 7858 5104 7896
rect 5176 7910 5205 7926
rect 5219 7910 5248 7926
rect 5263 7916 5293 7932
rect 5321 7910 5327 7958
rect 5330 7952 5349 7958
rect 5364 7952 5394 7960
rect 5330 7944 5394 7952
rect 5330 7928 5410 7944
rect 5426 7937 5488 7968
rect 5504 7937 5566 7968
rect 5635 7966 5684 7991
rect 5699 7966 5729 7982
rect 5598 7952 5628 7960
rect 5635 7958 5745 7966
rect 5598 7944 5643 7952
rect 5330 7926 5349 7928
rect 5364 7926 5410 7928
rect 5330 7910 5410 7926
rect 5437 7924 5472 7937
rect 5513 7934 5550 7937
rect 5513 7932 5555 7934
rect 5442 7921 5472 7924
rect 5451 7917 5458 7921
rect 5458 7916 5459 7917
rect 5417 7910 5427 7916
rect 5176 7902 5211 7910
rect 5176 7876 5177 7902
rect 5184 7876 5211 7902
rect 5119 7858 5149 7872
rect 5176 7868 5211 7876
rect 5213 7902 5254 7910
rect 5213 7876 5228 7902
rect 5235 7876 5254 7902
rect 5318 7898 5349 7910
rect 5364 7898 5467 7910
rect 5479 7900 5505 7926
rect 5520 7921 5550 7932
rect 5582 7928 5644 7944
rect 5582 7926 5628 7928
rect 5582 7910 5644 7926
rect 5656 7910 5662 7958
rect 5665 7950 5745 7958
rect 5665 7948 5684 7950
rect 5699 7948 5733 7950
rect 5665 7932 5745 7948
rect 5665 7910 5684 7932
rect 5699 7916 5729 7932
rect 5757 7926 5763 8000
rect 5766 7926 5785 8070
rect 5800 7926 5806 8070
rect 5815 8000 5828 8070
rect 5880 8066 5902 8070
rect 5873 8044 5902 8058
rect 5955 8044 5971 8058
rect 6009 8054 6015 8056
rect 6022 8054 6130 8070
rect 6137 8054 6143 8056
rect 6151 8054 6166 8070
rect 6232 8064 6251 8067
rect 5873 8042 5971 8044
rect 5998 8042 6166 8054
rect 6181 8044 6197 8058
rect 6232 8045 6254 8064
rect 6264 8058 6280 8059
rect 6263 8056 6280 8058
rect 6264 8051 6280 8056
rect 6254 8044 6260 8045
rect 6263 8044 6292 8051
rect 6181 8043 6292 8044
rect 6181 8042 6298 8043
rect 5857 8034 5908 8042
rect 5955 8034 5989 8042
rect 5857 8022 5882 8034
rect 5889 8022 5908 8034
rect 5962 8032 5989 8034
rect 5998 8032 6219 8042
rect 6254 8039 6260 8042
rect 5962 8028 6219 8032
rect 5857 8014 5908 8022
rect 5955 8014 6219 8028
rect 6263 8034 6298 8042
rect 5809 7966 5828 8000
rect 5873 8006 5902 8014
rect 5873 8000 5890 8006
rect 5873 7998 5907 8000
rect 5955 7998 5971 8014
rect 5972 8004 6180 8014
rect 6181 8004 6197 8014
rect 6245 8010 6260 8025
rect 6263 8022 6264 8034
rect 6271 8022 6298 8034
rect 6263 8014 6298 8022
rect 6263 8013 6292 8014
rect 5983 8000 6197 8004
rect 5998 7998 6197 8000
rect 6232 8000 6245 8010
rect 6263 8000 6280 8013
rect 6232 7998 6280 8000
rect 5874 7994 5907 7998
rect 5870 7992 5907 7994
rect 5870 7991 5937 7992
rect 5870 7986 5901 7991
rect 5907 7986 5937 7991
rect 5870 7982 5937 7986
rect 5843 7979 5937 7982
rect 5843 7972 5892 7979
rect 5843 7966 5873 7972
rect 5892 7967 5897 7972
rect 5809 7950 5889 7966
rect 5901 7958 5937 7979
rect 5998 7974 6187 7998
rect 6232 7997 6279 7998
rect 6245 7992 6279 7997
rect 6013 7971 6187 7974
rect 6006 7968 6187 7971
rect 6215 7991 6279 7992
rect 5809 7948 5828 7950
rect 5843 7948 5877 7950
rect 5809 7932 5889 7948
rect 5809 7926 5828 7932
rect 5525 7900 5628 7910
rect 5479 7898 5628 7900
rect 5649 7898 5684 7910
rect 5318 7896 5480 7898
rect 5330 7876 5349 7896
rect 5364 7894 5394 7896
rect 5213 7868 5254 7876
rect 5336 7872 5349 7876
rect 5401 7880 5480 7896
rect 5512 7896 5684 7898
rect 5512 7880 5591 7896
rect 5598 7894 5628 7896
rect 5176 7858 5205 7868
rect 5219 7858 5248 7868
rect 5263 7858 5293 7872
rect 5336 7858 5379 7872
rect 5401 7868 5591 7880
rect 5656 7876 5662 7896
rect 5386 7858 5416 7868
rect 5417 7858 5575 7868
rect 5579 7858 5609 7868
rect 5613 7858 5643 7872
rect 5671 7858 5684 7896
rect 5756 7910 5785 7926
rect 5799 7910 5828 7926
rect 5843 7916 5873 7932
rect 5901 7910 5907 7958
rect 5910 7952 5929 7958
rect 5944 7952 5974 7960
rect 5910 7944 5974 7952
rect 5910 7928 5990 7944
rect 6006 7937 6068 7968
rect 6084 7937 6146 7968
rect 6215 7966 6264 7991
rect 6279 7966 6309 7982
rect 6178 7952 6208 7960
rect 6215 7958 6325 7966
rect 6178 7944 6223 7952
rect 5910 7926 5929 7928
rect 5944 7926 5990 7928
rect 5910 7910 5990 7926
rect 6017 7924 6052 7937
rect 6093 7934 6130 7937
rect 6093 7932 6135 7934
rect 6022 7921 6052 7924
rect 6031 7917 6038 7921
rect 6038 7916 6039 7917
rect 5997 7910 6007 7916
rect 5756 7902 5791 7910
rect 5756 7876 5757 7902
rect 5764 7876 5791 7902
rect 5699 7858 5729 7872
rect 5756 7868 5791 7876
rect 5793 7902 5834 7910
rect 5793 7876 5808 7902
rect 5815 7876 5834 7902
rect 5898 7898 5929 7910
rect 5944 7898 6047 7910
rect 6059 7900 6085 7926
rect 6100 7921 6130 7932
rect 6162 7928 6224 7944
rect 6162 7926 6208 7928
rect 6162 7910 6224 7926
rect 6236 7910 6242 7958
rect 6245 7950 6325 7958
rect 6245 7948 6264 7950
rect 6279 7948 6313 7950
rect 6245 7932 6325 7948
rect 6245 7910 6264 7932
rect 6279 7916 6309 7932
rect 6337 7926 6343 8000
rect 6346 7926 6365 8070
rect 6380 7926 6386 8070
rect 6395 8000 6408 8070
rect 6460 8066 6482 8070
rect 6453 8044 6482 8058
rect 6535 8044 6551 8058
rect 6589 8054 6595 8056
rect 6602 8054 6710 8070
rect 6717 8054 6723 8056
rect 6731 8054 6746 8070
rect 6812 8064 6831 8067
rect 6453 8042 6551 8044
rect 6578 8042 6746 8054
rect 6761 8044 6777 8058
rect 6812 8045 6834 8064
rect 6844 8058 6860 8059
rect 6843 8056 6860 8058
rect 6844 8051 6860 8056
rect 6834 8044 6840 8045
rect 6843 8044 6872 8051
rect 6761 8043 6872 8044
rect 6761 8042 6878 8043
rect 6437 8034 6488 8042
rect 6535 8034 6569 8042
rect 6437 8022 6462 8034
rect 6469 8022 6488 8034
rect 6542 8032 6569 8034
rect 6578 8032 6799 8042
rect 6834 8039 6840 8042
rect 6542 8028 6799 8032
rect 6437 8014 6488 8022
rect 6535 8014 6799 8028
rect 6843 8034 6878 8042
rect 6389 7966 6408 8000
rect 6453 8006 6482 8014
rect 6453 8000 6470 8006
rect 6453 7998 6487 8000
rect 6535 7998 6551 8014
rect 6552 8004 6760 8014
rect 6761 8004 6777 8014
rect 6825 8010 6840 8025
rect 6843 8022 6844 8034
rect 6851 8022 6878 8034
rect 6843 8014 6878 8022
rect 6843 8013 6872 8014
rect 6563 8000 6777 8004
rect 6578 7998 6777 8000
rect 6812 8000 6825 8010
rect 6843 8000 6860 8013
rect 6812 7998 6860 8000
rect 6454 7994 6487 7998
rect 6450 7992 6487 7994
rect 6450 7991 6517 7992
rect 6450 7986 6481 7991
rect 6487 7986 6517 7991
rect 6450 7982 6517 7986
rect 6423 7979 6517 7982
rect 6423 7972 6472 7979
rect 6423 7966 6453 7972
rect 6472 7967 6477 7972
rect 6389 7950 6469 7966
rect 6481 7958 6517 7979
rect 6578 7974 6767 7998
rect 6812 7997 6859 7998
rect 6825 7992 6859 7997
rect 6593 7971 6767 7974
rect 6586 7968 6767 7971
rect 6795 7991 6859 7992
rect 6389 7948 6408 7950
rect 6423 7948 6457 7950
rect 6389 7932 6469 7948
rect 6389 7926 6408 7932
rect 6105 7900 6208 7910
rect 6059 7898 6208 7900
rect 6229 7898 6264 7910
rect 5898 7896 6060 7898
rect 5910 7876 5929 7896
rect 5944 7894 5974 7896
rect 5793 7868 5834 7876
rect 5916 7872 5929 7876
rect 5981 7880 6060 7896
rect 6092 7896 6264 7898
rect 6092 7880 6171 7896
rect 6178 7894 6208 7896
rect 5756 7858 5785 7868
rect 5799 7858 5828 7868
rect 5843 7858 5873 7872
rect 5916 7858 5959 7872
rect 5981 7868 6171 7880
rect 6236 7876 6242 7896
rect 5966 7858 5996 7868
rect 5997 7858 6155 7868
rect 6159 7858 6189 7868
rect 6193 7858 6223 7872
rect 6251 7858 6264 7896
rect 6336 7910 6365 7926
rect 6379 7910 6408 7926
rect 6423 7916 6453 7932
rect 6481 7910 6487 7958
rect 6490 7952 6509 7958
rect 6524 7952 6554 7960
rect 6490 7944 6554 7952
rect 6490 7928 6570 7944
rect 6586 7937 6648 7968
rect 6664 7937 6726 7968
rect 6795 7966 6844 7991
rect 6859 7966 6889 7982
rect 6758 7952 6788 7960
rect 6795 7958 6905 7966
rect 6758 7944 6803 7952
rect 6490 7926 6509 7928
rect 6524 7926 6570 7928
rect 6490 7910 6570 7926
rect 6597 7924 6632 7937
rect 6673 7934 6710 7937
rect 6673 7932 6715 7934
rect 6602 7921 6632 7924
rect 6611 7917 6618 7921
rect 6618 7916 6619 7917
rect 6577 7910 6587 7916
rect 6336 7902 6371 7910
rect 6336 7876 6337 7902
rect 6344 7876 6371 7902
rect 6279 7858 6309 7872
rect 6336 7868 6371 7876
rect 6373 7902 6414 7910
rect 6373 7876 6388 7902
rect 6395 7876 6414 7902
rect 6478 7898 6509 7910
rect 6524 7898 6627 7910
rect 6639 7900 6665 7926
rect 6680 7921 6710 7932
rect 6742 7928 6804 7944
rect 6742 7926 6788 7928
rect 6742 7910 6804 7926
rect 6816 7910 6822 7958
rect 6825 7950 6905 7958
rect 6825 7948 6844 7950
rect 6859 7948 6893 7950
rect 6825 7932 6905 7948
rect 6825 7910 6844 7932
rect 6859 7916 6889 7932
rect 6917 7926 6923 8000
rect 6926 7926 6945 8070
rect 6960 7926 6966 8070
rect 6975 8000 6988 8070
rect 7040 8066 7062 8070
rect 7033 8044 7062 8058
rect 7115 8044 7131 8058
rect 7169 8054 7175 8056
rect 7182 8054 7290 8070
rect 7297 8054 7303 8056
rect 7311 8054 7326 8070
rect 7392 8064 7411 8067
rect 7033 8042 7131 8044
rect 7158 8042 7326 8054
rect 7341 8044 7357 8058
rect 7392 8045 7414 8064
rect 7424 8058 7440 8059
rect 7423 8056 7440 8058
rect 7424 8051 7440 8056
rect 7414 8044 7420 8045
rect 7423 8044 7452 8051
rect 7341 8043 7452 8044
rect 7341 8042 7458 8043
rect 7017 8034 7068 8042
rect 7115 8034 7149 8042
rect 7017 8022 7042 8034
rect 7049 8022 7068 8034
rect 7122 8032 7149 8034
rect 7158 8032 7379 8042
rect 7414 8039 7420 8042
rect 7122 8028 7379 8032
rect 7017 8014 7068 8022
rect 7115 8014 7379 8028
rect 7423 8034 7458 8042
rect 6969 7966 6988 8000
rect 7033 8006 7062 8014
rect 7033 8000 7050 8006
rect 7033 7998 7067 8000
rect 7115 7998 7131 8014
rect 7132 8004 7340 8014
rect 7341 8004 7357 8014
rect 7405 8010 7420 8025
rect 7423 8022 7424 8034
rect 7431 8022 7458 8034
rect 7423 8014 7458 8022
rect 7423 8013 7452 8014
rect 7143 8000 7357 8004
rect 7158 7998 7357 8000
rect 7392 8000 7405 8010
rect 7423 8000 7440 8013
rect 7392 7998 7440 8000
rect 7034 7994 7067 7998
rect 7030 7992 7067 7994
rect 7030 7991 7097 7992
rect 7030 7986 7061 7991
rect 7067 7986 7097 7991
rect 7030 7982 7097 7986
rect 7003 7979 7097 7982
rect 7003 7972 7052 7979
rect 7003 7966 7033 7972
rect 7052 7967 7057 7972
rect 6969 7950 7049 7966
rect 7061 7958 7097 7979
rect 7158 7974 7347 7998
rect 7392 7997 7439 7998
rect 7405 7992 7439 7997
rect 7173 7971 7347 7974
rect 7166 7968 7347 7971
rect 7375 7991 7439 7992
rect 6969 7948 6988 7950
rect 7003 7948 7037 7950
rect 6969 7932 7049 7948
rect 6969 7926 6988 7932
rect 6685 7900 6788 7910
rect 6639 7898 6788 7900
rect 6809 7898 6844 7910
rect 6478 7896 6640 7898
rect 6490 7876 6509 7896
rect 6524 7894 6554 7896
rect 6373 7868 6414 7876
rect 6496 7872 6509 7876
rect 6561 7880 6640 7896
rect 6672 7896 6844 7898
rect 6672 7880 6751 7896
rect 6758 7894 6788 7896
rect 6336 7858 6365 7868
rect 6379 7858 6408 7868
rect 6423 7858 6453 7872
rect 6496 7858 6539 7872
rect 6561 7868 6751 7880
rect 6816 7876 6822 7896
rect 6546 7858 6576 7868
rect 6577 7858 6735 7868
rect 6739 7858 6769 7868
rect 6773 7858 6803 7872
rect 6831 7858 6844 7896
rect 6916 7910 6945 7926
rect 6959 7910 6988 7926
rect 7003 7916 7033 7932
rect 7061 7910 7067 7958
rect 7070 7952 7089 7958
rect 7104 7952 7134 7960
rect 7070 7944 7134 7952
rect 7070 7928 7150 7944
rect 7166 7937 7228 7968
rect 7244 7937 7306 7968
rect 7375 7966 7424 7991
rect 7439 7966 7469 7982
rect 7338 7952 7368 7960
rect 7375 7958 7485 7966
rect 7338 7944 7383 7952
rect 7070 7926 7089 7928
rect 7104 7926 7150 7928
rect 7070 7910 7150 7926
rect 7177 7924 7212 7937
rect 7253 7934 7290 7937
rect 7253 7932 7295 7934
rect 7182 7921 7212 7924
rect 7191 7917 7198 7921
rect 7198 7916 7199 7917
rect 7157 7910 7167 7916
rect 6916 7902 6951 7910
rect 6916 7876 6917 7902
rect 6924 7876 6951 7902
rect 6859 7858 6889 7872
rect 6916 7868 6951 7876
rect 6953 7902 6994 7910
rect 6953 7876 6968 7902
rect 6975 7876 6994 7902
rect 7058 7898 7089 7910
rect 7104 7898 7207 7910
rect 7219 7900 7245 7926
rect 7260 7921 7290 7932
rect 7322 7928 7384 7944
rect 7322 7926 7368 7928
rect 7322 7910 7384 7926
rect 7396 7910 7402 7958
rect 7405 7950 7485 7958
rect 7405 7948 7424 7950
rect 7439 7948 7473 7950
rect 7405 7932 7485 7948
rect 7405 7910 7424 7932
rect 7439 7916 7469 7932
rect 7497 7926 7503 8000
rect 7506 7926 7525 8070
rect 7540 7926 7546 8070
rect 7555 8000 7568 8070
rect 7620 8066 7642 8070
rect 7613 8044 7642 8058
rect 7695 8044 7711 8058
rect 7749 8054 7755 8056
rect 7762 8054 7870 8070
rect 7877 8054 7883 8056
rect 7891 8054 7906 8070
rect 7972 8064 7991 8067
rect 7613 8042 7711 8044
rect 7738 8042 7906 8054
rect 7921 8044 7937 8058
rect 7972 8045 7994 8064
rect 8004 8058 8020 8059
rect 8003 8056 8020 8058
rect 8004 8051 8020 8056
rect 7994 8044 8000 8045
rect 8003 8044 8032 8051
rect 7921 8043 8032 8044
rect 7921 8042 8038 8043
rect 7597 8034 7648 8042
rect 7695 8034 7729 8042
rect 7597 8022 7622 8034
rect 7629 8022 7648 8034
rect 7702 8032 7729 8034
rect 7738 8032 7959 8042
rect 7994 8039 8000 8042
rect 7702 8028 7959 8032
rect 7597 8014 7648 8022
rect 7695 8014 7959 8028
rect 8003 8034 8038 8042
rect 7549 7966 7568 8000
rect 7613 8006 7642 8014
rect 7613 8000 7630 8006
rect 7613 7998 7647 8000
rect 7695 7998 7711 8014
rect 7712 8004 7920 8014
rect 7921 8004 7937 8014
rect 7985 8010 8000 8025
rect 8003 8022 8004 8034
rect 8011 8022 8038 8034
rect 8003 8014 8038 8022
rect 8003 8013 8032 8014
rect 7723 8000 7937 8004
rect 7738 7998 7937 8000
rect 7972 8000 7985 8010
rect 8003 8000 8020 8013
rect 7972 7998 8020 8000
rect 7614 7994 7647 7998
rect 7610 7992 7647 7994
rect 7610 7991 7677 7992
rect 7610 7986 7641 7991
rect 7647 7986 7677 7991
rect 7610 7982 7677 7986
rect 7583 7979 7677 7982
rect 7583 7972 7632 7979
rect 7583 7966 7613 7972
rect 7632 7967 7637 7972
rect 7549 7950 7629 7966
rect 7641 7958 7677 7979
rect 7738 7974 7927 7998
rect 7972 7997 8019 7998
rect 7985 7992 8019 7997
rect 7753 7971 7927 7974
rect 7746 7968 7927 7971
rect 7955 7991 8019 7992
rect 7549 7948 7568 7950
rect 7583 7948 7617 7950
rect 7549 7932 7629 7948
rect 7549 7926 7568 7932
rect 7265 7900 7368 7910
rect 7219 7898 7368 7900
rect 7389 7898 7424 7910
rect 7058 7896 7220 7898
rect 7070 7876 7089 7896
rect 7104 7894 7134 7896
rect 6953 7868 6994 7876
rect 7076 7872 7089 7876
rect 7141 7880 7220 7896
rect 7252 7896 7424 7898
rect 7252 7880 7331 7896
rect 7338 7894 7368 7896
rect 6916 7858 6945 7868
rect 6959 7858 6988 7868
rect 7003 7858 7033 7872
rect 7076 7858 7119 7872
rect 7141 7868 7331 7880
rect 7396 7876 7402 7896
rect 7126 7858 7156 7868
rect 7157 7858 7315 7868
rect 7319 7858 7349 7868
rect 7353 7858 7383 7872
rect 7411 7858 7424 7896
rect 7496 7910 7525 7926
rect 7539 7910 7568 7926
rect 7583 7916 7613 7932
rect 7641 7910 7647 7958
rect 7650 7952 7669 7958
rect 7684 7952 7714 7960
rect 7650 7944 7714 7952
rect 7650 7928 7730 7944
rect 7746 7937 7808 7968
rect 7824 7937 7886 7968
rect 7955 7966 8004 7991
rect 8019 7966 8049 7982
rect 7918 7952 7948 7960
rect 7955 7958 8065 7966
rect 7918 7944 7963 7952
rect 7650 7926 7669 7928
rect 7684 7926 7730 7928
rect 7650 7910 7730 7926
rect 7757 7924 7792 7937
rect 7833 7934 7870 7937
rect 7833 7932 7875 7934
rect 7762 7921 7792 7924
rect 7771 7917 7778 7921
rect 7778 7916 7779 7917
rect 7737 7910 7747 7916
rect 7496 7902 7531 7910
rect 7496 7876 7497 7902
rect 7504 7876 7531 7902
rect 7439 7858 7469 7872
rect 7496 7868 7531 7876
rect 7533 7902 7574 7910
rect 7533 7876 7548 7902
rect 7555 7876 7574 7902
rect 7638 7898 7669 7910
rect 7684 7898 7787 7910
rect 7799 7900 7825 7926
rect 7840 7921 7870 7932
rect 7902 7928 7964 7944
rect 7902 7926 7948 7928
rect 7902 7910 7964 7926
rect 7976 7910 7982 7958
rect 7985 7950 8065 7958
rect 7985 7948 8004 7950
rect 8019 7948 8053 7950
rect 7985 7932 8065 7948
rect 7985 7910 8004 7932
rect 8019 7916 8049 7932
rect 8077 7926 8083 8000
rect 8086 7926 8105 8070
rect 8120 7926 8126 8070
rect 8135 8000 8148 8070
rect 8200 8066 8222 8070
rect 8193 8044 8222 8058
rect 8275 8044 8291 8058
rect 8329 8054 8335 8056
rect 8342 8054 8450 8070
rect 8457 8054 8463 8056
rect 8471 8054 8486 8070
rect 8552 8064 8571 8067
rect 8193 8042 8291 8044
rect 8318 8042 8486 8054
rect 8501 8044 8517 8058
rect 8552 8045 8574 8064
rect 8584 8058 8600 8059
rect 8583 8056 8600 8058
rect 8584 8051 8600 8056
rect 8574 8044 8580 8045
rect 8583 8044 8612 8051
rect 8501 8043 8612 8044
rect 8501 8042 8618 8043
rect 8177 8034 8228 8042
rect 8275 8034 8309 8042
rect 8177 8022 8202 8034
rect 8209 8022 8228 8034
rect 8282 8032 8309 8034
rect 8318 8032 8539 8042
rect 8574 8039 8580 8042
rect 8282 8028 8539 8032
rect 8177 8014 8228 8022
rect 8275 8014 8539 8028
rect 8583 8034 8618 8042
rect 8129 7966 8148 8000
rect 8193 8006 8222 8014
rect 8193 8000 8210 8006
rect 8193 7998 8227 8000
rect 8275 7998 8291 8014
rect 8292 8004 8500 8014
rect 8501 8004 8517 8014
rect 8565 8010 8580 8025
rect 8583 8022 8584 8034
rect 8591 8022 8618 8034
rect 8583 8014 8618 8022
rect 8583 8013 8612 8014
rect 8303 8000 8517 8004
rect 8318 7998 8517 8000
rect 8552 8000 8565 8010
rect 8583 8000 8600 8013
rect 8552 7998 8600 8000
rect 8194 7994 8227 7998
rect 8190 7992 8227 7994
rect 8190 7991 8257 7992
rect 8190 7986 8221 7991
rect 8227 7986 8257 7991
rect 8190 7982 8257 7986
rect 8163 7979 8257 7982
rect 8163 7972 8212 7979
rect 8163 7966 8193 7972
rect 8212 7967 8217 7972
rect 8129 7950 8209 7966
rect 8221 7958 8257 7979
rect 8318 7974 8507 7998
rect 8552 7997 8599 7998
rect 8565 7992 8599 7997
rect 8333 7971 8507 7974
rect 8326 7968 8507 7971
rect 8535 7991 8599 7992
rect 8129 7948 8148 7950
rect 8163 7948 8197 7950
rect 8129 7932 8209 7948
rect 8129 7926 8148 7932
rect 7845 7900 7948 7910
rect 7799 7898 7948 7900
rect 7969 7898 8004 7910
rect 7638 7896 7800 7898
rect 7650 7876 7669 7896
rect 7684 7894 7714 7896
rect 7533 7868 7574 7876
rect 7656 7872 7669 7876
rect 7721 7880 7800 7896
rect 7832 7896 8004 7898
rect 7832 7880 7911 7896
rect 7918 7894 7948 7896
rect 7496 7858 7525 7868
rect 7539 7858 7568 7868
rect 7583 7858 7613 7872
rect 7656 7858 7699 7872
rect 7721 7868 7911 7880
rect 7976 7876 7982 7896
rect 7706 7858 7736 7868
rect 7737 7858 7895 7868
rect 7899 7858 7929 7868
rect 7933 7858 7963 7872
rect 7991 7858 8004 7896
rect 8076 7910 8105 7926
rect 8119 7910 8148 7926
rect 8163 7916 8193 7932
rect 8221 7910 8227 7958
rect 8230 7952 8249 7958
rect 8264 7952 8294 7960
rect 8230 7944 8294 7952
rect 8230 7928 8310 7944
rect 8326 7937 8388 7968
rect 8404 7937 8466 7968
rect 8535 7966 8584 7991
rect 8599 7966 8629 7982
rect 8498 7952 8528 7960
rect 8535 7958 8645 7966
rect 8498 7944 8543 7952
rect 8230 7926 8249 7928
rect 8264 7926 8310 7928
rect 8230 7910 8310 7926
rect 8337 7924 8372 7937
rect 8413 7934 8450 7937
rect 8413 7932 8455 7934
rect 8342 7921 8372 7924
rect 8351 7917 8358 7921
rect 8358 7916 8359 7917
rect 8317 7910 8327 7916
rect 8076 7902 8111 7910
rect 8076 7876 8077 7902
rect 8084 7876 8111 7902
rect 8019 7858 8049 7872
rect 8076 7868 8111 7876
rect 8113 7902 8154 7910
rect 8113 7876 8128 7902
rect 8135 7876 8154 7902
rect 8218 7898 8249 7910
rect 8264 7898 8367 7910
rect 8379 7900 8405 7926
rect 8420 7921 8450 7932
rect 8482 7928 8544 7944
rect 8482 7926 8528 7928
rect 8482 7910 8544 7926
rect 8556 7910 8562 7958
rect 8565 7950 8645 7958
rect 8565 7948 8584 7950
rect 8599 7948 8633 7950
rect 8565 7932 8645 7948
rect 8565 7910 8584 7932
rect 8599 7916 8629 7932
rect 8657 7926 8663 8000
rect 8666 7926 8685 8070
rect 8700 7926 8706 8070
rect 8715 8000 8728 8070
rect 8780 8066 8802 8070
rect 8773 8044 8802 8058
rect 8855 8044 8871 8058
rect 8909 8054 8915 8056
rect 8922 8054 9030 8070
rect 9037 8054 9043 8056
rect 9051 8054 9066 8070
rect 9132 8064 9151 8067
rect 8773 8042 8871 8044
rect 8898 8042 9066 8054
rect 9081 8044 9097 8058
rect 9132 8045 9154 8064
rect 9164 8058 9180 8059
rect 9163 8056 9180 8058
rect 9164 8051 9180 8056
rect 9154 8044 9160 8045
rect 9163 8044 9192 8051
rect 9081 8043 9192 8044
rect 9081 8042 9198 8043
rect 8757 8034 8808 8042
rect 8855 8034 8889 8042
rect 8757 8022 8782 8034
rect 8789 8022 8808 8034
rect 8862 8032 8889 8034
rect 8898 8032 9119 8042
rect 9154 8039 9160 8042
rect 8862 8028 9119 8032
rect 8757 8014 8808 8022
rect 8855 8014 9119 8028
rect 9163 8034 9198 8042
rect 8709 7966 8728 8000
rect 8773 8006 8802 8014
rect 8773 8000 8790 8006
rect 8773 7998 8807 8000
rect 8855 7998 8871 8014
rect 8872 8004 9080 8014
rect 9081 8004 9097 8014
rect 9145 8010 9160 8025
rect 9163 8022 9164 8034
rect 9171 8022 9198 8034
rect 9163 8014 9198 8022
rect 9163 8013 9192 8014
rect 8883 8000 9097 8004
rect 8898 7998 9097 8000
rect 9132 8000 9145 8010
rect 9163 8000 9180 8013
rect 9132 7998 9180 8000
rect 8774 7994 8807 7998
rect 8770 7992 8807 7994
rect 8770 7991 8837 7992
rect 8770 7986 8801 7991
rect 8807 7986 8837 7991
rect 8770 7982 8837 7986
rect 8743 7979 8837 7982
rect 8743 7972 8792 7979
rect 8743 7966 8773 7972
rect 8792 7967 8797 7972
rect 8709 7950 8789 7966
rect 8801 7958 8837 7979
rect 8898 7974 9087 7998
rect 9132 7997 9179 7998
rect 9145 7992 9179 7997
rect 8913 7971 9087 7974
rect 8906 7968 9087 7971
rect 9115 7991 9179 7992
rect 8709 7948 8728 7950
rect 8743 7948 8777 7950
rect 8709 7932 8789 7948
rect 8709 7926 8728 7932
rect 8425 7900 8528 7910
rect 8379 7898 8528 7900
rect 8549 7898 8584 7910
rect 8218 7896 8380 7898
rect 8230 7876 8249 7896
rect 8264 7894 8294 7896
rect 8113 7868 8154 7876
rect 8236 7872 8249 7876
rect 8301 7880 8380 7896
rect 8412 7896 8584 7898
rect 8412 7880 8491 7896
rect 8498 7894 8528 7896
rect 8076 7858 8105 7868
rect 8119 7858 8148 7868
rect 8163 7858 8193 7872
rect 8236 7858 8279 7872
rect 8301 7868 8491 7880
rect 8556 7876 8562 7896
rect 8286 7858 8316 7868
rect 8317 7858 8475 7868
rect 8479 7858 8509 7868
rect 8513 7858 8543 7872
rect 8571 7858 8584 7896
rect 8656 7910 8685 7926
rect 8699 7910 8728 7926
rect 8743 7916 8773 7932
rect 8801 7910 8807 7958
rect 8810 7952 8829 7958
rect 8844 7952 8874 7960
rect 8810 7944 8874 7952
rect 8810 7928 8890 7944
rect 8906 7937 8968 7968
rect 8984 7937 9046 7968
rect 9115 7966 9164 7991
rect 9179 7966 9209 7982
rect 9078 7952 9108 7960
rect 9115 7958 9225 7966
rect 9078 7944 9123 7952
rect 8810 7926 8829 7928
rect 8844 7926 8890 7928
rect 8810 7910 8890 7926
rect 8917 7924 8952 7937
rect 8993 7934 9030 7937
rect 8993 7932 9035 7934
rect 8922 7921 8952 7924
rect 8931 7917 8938 7921
rect 8938 7916 8939 7917
rect 8897 7910 8907 7916
rect 8656 7902 8691 7910
rect 8656 7876 8657 7902
rect 8664 7876 8691 7902
rect 8599 7858 8629 7872
rect 8656 7868 8691 7876
rect 8693 7902 8734 7910
rect 8693 7876 8708 7902
rect 8715 7876 8734 7902
rect 8798 7898 8829 7910
rect 8844 7898 8947 7910
rect 8959 7900 8985 7926
rect 9000 7921 9030 7932
rect 9062 7928 9124 7944
rect 9062 7926 9108 7928
rect 9062 7910 9124 7926
rect 9136 7910 9142 7958
rect 9145 7950 9225 7958
rect 9145 7948 9164 7950
rect 9179 7948 9213 7950
rect 9145 7932 9225 7948
rect 9145 7910 9164 7932
rect 9179 7916 9209 7932
rect 9237 7926 9243 8000
rect 9246 7926 9265 8070
rect 9280 7926 9286 8070
rect 9295 8000 9308 8070
rect 9360 8066 9382 8070
rect 9353 8044 9382 8058
rect 9435 8044 9451 8058
rect 9489 8054 9495 8056
rect 9502 8054 9610 8070
rect 9617 8054 9623 8056
rect 9631 8054 9646 8070
rect 9712 8064 9731 8067
rect 9353 8042 9451 8044
rect 9478 8042 9646 8054
rect 9661 8044 9677 8058
rect 9712 8045 9734 8064
rect 9744 8058 9760 8059
rect 9743 8056 9760 8058
rect 9744 8051 9760 8056
rect 9734 8044 9740 8045
rect 9743 8044 9772 8051
rect 9661 8043 9772 8044
rect 9661 8042 9778 8043
rect 9337 8034 9388 8042
rect 9435 8034 9469 8042
rect 9337 8022 9362 8034
rect 9369 8022 9388 8034
rect 9442 8032 9469 8034
rect 9478 8032 9699 8042
rect 9734 8039 9740 8042
rect 9442 8028 9699 8032
rect 9337 8014 9388 8022
rect 9435 8014 9699 8028
rect 9743 8034 9778 8042
rect 9289 7966 9308 8000
rect 9353 8006 9382 8014
rect 9353 8000 9370 8006
rect 9353 7998 9387 8000
rect 9435 7998 9451 8014
rect 9452 8004 9660 8014
rect 9661 8004 9677 8014
rect 9725 8010 9740 8025
rect 9743 8022 9744 8034
rect 9751 8022 9778 8034
rect 9743 8014 9778 8022
rect 9743 8013 9772 8014
rect 9463 8000 9677 8004
rect 9478 7998 9677 8000
rect 9712 8000 9725 8010
rect 9743 8000 9760 8013
rect 9712 7998 9760 8000
rect 9354 7994 9387 7998
rect 9350 7992 9387 7994
rect 9350 7991 9417 7992
rect 9350 7986 9381 7991
rect 9387 7986 9417 7991
rect 9350 7982 9417 7986
rect 9323 7979 9417 7982
rect 9323 7972 9372 7979
rect 9323 7966 9353 7972
rect 9372 7967 9377 7972
rect 9289 7950 9369 7966
rect 9381 7958 9417 7979
rect 9478 7974 9667 7998
rect 9712 7997 9759 7998
rect 9725 7992 9759 7997
rect 9493 7971 9667 7974
rect 9486 7968 9667 7971
rect 9695 7991 9759 7992
rect 9289 7948 9308 7950
rect 9323 7948 9357 7950
rect 9289 7932 9369 7948
rect 9289 7926 9308 7932
rect 9005 7900 9108 7910
rect 8959 7898 9108 7900
rect 9129 7898 9164 7910
rect 8798 7896 8960 7898
rect 8810 7876 8829 7896
rect 8844 7894 8874 7896
rect 8693 7868 8734 7876
rect 8816 7872 8829 7876
rect 8881 7880 8960 7896
rect 8992 7896 9164 7898
rect 8992 7880 9071 7896
rect 9078 7894 9108 7896
rect 8656 7858 8685 7868
rect 8699 7858 8728 7868
rect 8743 7858 8773 7872
rect 8816 7858 8859 7872
rect 8881 7868 9071 7880
rect 9136 7876 9142 7896
rect 8866 7858 8896 7868
rect 8897 7858 9055 7868
rect 9059 7858 9089 7868
rect 9093 7858 9123 7872
rect 9151 7858 9164 7896
rect 9236 7910 9265 7926
rect 9279 7910 9308 7926
rect 9323 7916 9353 7932
rect 9381 7910 9387 7958
rect 9390 7952 9409 7958
rect 9424 7952 9454 7960
rect 9390 7944 9454 7952
rect 9390 7928 9470 7944
rect 9486 7937 9548 7968
rect 9564 7937 9626 7968
rect 9695 7966 9744 7991
rect 9759 7966 9789 7982
rect 9658 7952 9688 7960
rect 9695 7958 9805 7966
rect 9658 7944 9703 7952
rect 9390 7926 9409 7928
rect 9424 7926 9470 7928
rect 9390 7910 9470 7926
rect 9497 7924 9532 7937
rect 9573 7934 9610 7937
rect 9573 7932 9615 7934
rect 9502 7921 9532 7924
rect 9511 7917 9518 7921
rect 9518 7916 9519 7917
rect 9477 7910 9487 7916
rect 9236 7902 9271 7910
rect 9236 7876 9237 7902
rect 9244 7876 9271 7902
rect 9179 7858 9209 7872
rect 9236 7868 9271 7876
rect 9273 7902 9314 7910
rect 9273 7876 9288 7902
rect 9295 7876 9314 7902
rect 9378 7898 9409 7910
rect 9424 7898 9527 7910
rect 9539 7900 9565 7926
rect 9580 7921 9610 7932
rect 9642 7928 9704 7944
rect 9642 7926 9688 7928
rect 9642 7910 9704 7926
rect 9716 7910 9722 7958
rect 9725 7950 9805 7958
rect 9725 7948 9744 7950
rect 9759 7948 9793 7950
rect 9725 7932 9805 7948
rect 9725 7910 9744 7932
rect 9759 7916 9789 7932
rect 9817 7926 9823 8000
rect 9826 7926 9845 8070
rect 9860 7926 9866 8070
rect 9875 8000 9888 8070
rect 9940 8066 9962 8070
rect 9933 8044 9962 8058
rect 10015 8044 10031 8058
rect 10069 8054 10075 8056
rect 10082 8054 10190 8070
rect 10197 8054 10203 8056
rect 10211 8054 10226 8070
rect 10292 8064 10311 8067
rect 9933 8042 10031 8044
rect 10058 8042 10226 8054
rect 10241 8044 10257 8058
rect 10292 8045 10314 8064
rect 10324 8058 10340 8059
rect 10323 8056 10340 8058
rect 10324 8051 10340 8056
rect 10314 8044 10320 8045
rect 10323 8044 10352 8051
rect 10241 8043 10352 8044
rect 10241 8042 10358 8043
rect 9917 8034 9968 8042
rect 10015 8034 10049 8042
rect 9917 8022 9942 8034
rect 9949 8022 9968 8034
rect 10022 8032 10049 8034
rect 10058 8032 10279 8042
rect 10314 8039 10320 8042
rect 10022 8028 10279 8032
rect 9917 8014 9968 8022
rect 10015 8014 10279 8028
rect 10323 8034 10358 8042
rect 9869 7966 9888 8000
rect 9933 8006 9962 8014
rect 9933 8000 9950 8006
rect 9933 7998 9967 8000
rect 10015 7998 10031 8014
rect 10032 8004 10240 8014
rect 10241 8004 10257 8014
rect 10305 8010 10320 8025
rect 10323 8022 10324 8034
rect 10331 8022 10358 8034
rect 10323 8014 10358 8022
rect 10323 8013 10352 8014
rect 10043 8000 10257 8004
rect 10058 7998 10257 8000
rect 10292 8000 10305 8010
rect 10323 8000 10340 8013
rect 10292 7998 10340 8000
rect 9934 7994 9967 7998
rect 9930 7992 9967 7994
rect 9930 7991 9997 7992
rect 9930 7986 9961 7991
rect 9967 7986 9997 7991
rect 9930 7982 9997 7986
rect 9903 7979 9997 7982
rect 9903 7972 9952 7979
rect 9903 7966 9933 7972
rect 9952 7967 9957 7972
rect 9869 7950 9949 7966
rect 9961 7958 9997 7979
rect 10058 7974 10247 7998
rect 10292 7997 10339 7998
rect 10305 7992 10339 7997
rect 10073 7971 10247 7974
rect 10066 7968 10247 7971
rect 10275 7991 10339 7992
rect 9869 7948 9888 7950
rect 9903 7948 9937 7950
rect 9869 7932 9949 7948
rect 9869 7926 9888 7932
rect 9585 7900 9688 7910
rect 9539 7898 9688 7900
rect 9709 7898 9744 7910
rect 9378 7896 9540 7898
rect 9390 7876 9409 7896
rect 9424 7894 9454 7896
rect 9273 7868 9314 7876
rect 9396 7872 9409 7876
rect 9461 7880 9540 7896
rect 9572 7896 9744 7898
rect 9572 7880 9651 7896
rect 9658 7894 9688 7896
rect 9236 7858 9265 7868
rect 9279 7858 9308 7868
rect 9323 7858 9353 7872
rect 9396 7858 9439 7872
rect 9461 7868 9651 7880
rect 9716 7876 9722 7896
rect 9446 7858 9476 7868
rect 9477 7858 9635 7868
rect 9639 7858 9669 7868
rect 9673 7858 9703 7872
rect 9731 7858 9744 7896
rect 9816 7910 9845 7926
rect 9859 7910 9888 7926
rect 9903 7916 9933 7932
rect 9961 7910 9967 7958
rect 9970 7952 9989 7958
rect 10004 7952 10034 7960
rect 9970 7944 10034 7952
rect 9970 7928 10050 7944
rect 10066 7937 10128 7968
rect 10144 7937 10206 7968
rect 10275 7966 10324 7991
rect 10339 7966 10369 7982
rect 10238 7952 10268 7960
rect 10275 7958 10385 7966
rect 10238 7944 10283 7952
rect 9970 7926 9989 7928
rect 10004 7926 10050 7928
rect 9970 7910 10050 7926
rect 10077 7924 10112 7937
rect 10153 7934 10190 7937
rect 10153 7932 10195 7934
rect 10082 7921 10112 7924
rect 10091 7917 10098 7921
rect 10098 7916 10099 7917
rect 10057 7910 10067 7916
rect 9816 7902 9851 7910
rect 9816 7876 9817 7902
rect 9824 7876 9851 7902
rect 9759 7858 9789 7872
rect 9816 7868 9851 7876
rect 9853 7902 9894 7910
rect 9853 7876 9868 7902
rect 9875 7876 9894 7902
rect 9958 7898 9989 7910
rect 10004 7898 10107 7910
rect 10119 7900 10145 7926
rect 10160 7921 10190 7932
rect 10222 7928 10284 7944
rect 10222 7926 10268 7928
rect 10222 7910 10284 7926
rect 10296 7910 10302 7958
rect 10305 7950 10385 7958
rect 10305 7948 10324 7950
rect 10339 7948 10373 7950
rect 10305 7932 10385 7948
rect 10305 7910 10324 7932
rect 10339 7916 10369 7932
rect 10397 7926 10403 8000
rect 10406 7926 10425 8070
rect 10440 7926 10446 8070
rect 10455 8000 10468 8070
rect 10520 8066 10542 8070
rect 10513 8044 10542 8058
rect 10595 8044 10611 8058
rect 10649 8054 10655 8056
rect 10662 8054 10770 8070
rect 10777 8054 10783 8056
rect 10791 8054 10806 8070
rect 10872 8064 10891 8067
rect 10513 8042 10611 8044
rect 10638 8042 10806 8054
rect 10821 8044 10837 8058
rect 10872 8045 10894 8064
rect 10904 8058 10920 8059
rect 10903 8056 10920 8058
rect 10904 8051 10920 8056
rect 10894 8044 10900 8045
rect 10903 8044 10932 8051
rect 10821 8043 10932 8044
rect 10821 8042 10938 8043
rect 10497 8034 10548 8042
rect 10595 8034 10629 8042
rect 10497 8022 10522 8034
rect 10529 8022 10548 8034
rect 10602 8032 10629 8034
rect 10638 8032 10859 8042
rect 10894 8039 10900 8042
rect 10602 8028 10859 8032
rect 10497 8014 10548 8022
rect 10595 8014 10859 8028
rect 10903 8034 10938 8042
rect 10449 7966 10468 8000
rect 10513 8006 10542 8014
rect 10513 8000 10530 8006
rect 10513 7998 10547 8000
rect 10595 7998 10611 8014
rect 10612 8004 10820 8014
rect 10821 8004 10837 8014
rect 10885 8010 10900 8025
rect 10903 8022 10904 8034
rect 10911 8022 10938 8034
rect 10903 8014 10938 8022
rect 10903 8013 10932 8014
rect 10623 8000 10837 8004
rect 10638 7998 10837 8000
rect 10872 8000 10885 8010
rect 10903 8000 10920 8013
rect 10872 7998 10920 8000
rect 10514 7994 10547 7998
rect 10510 7992 10547 7994
rect 10510 7991 10577 7992
rect 10510 7986 10541 7991
rect 10547 7986 10577 7991
rect 10510 7982 10577 7986
rect 10483 7979 10577 7982
rect 10483 7972 10532 7979
rect 10483 7966 10513 7972
rect 10532 7967 10537 7972
rect 10449 7950 10529 7966
rect 10541 7958 10577 7979
rect 10638 7974 10827 7998
rect 10872 7997 10919 7998
rect 10885 7992 10919 7997
rect 10653 7971 10827 7974
rect 10646 7968 10827 7971
rect 10855 7991 10919 7992
rect 10449 7948 10468 7950
rect 10483 7948 10517 7950
rect 10449 7932 10529 7948
rect 10449 7926 10468 7932
rect 10165 7900 10268 7910
rect 10119 7898 10268 7900
rect 10289 7898 10324 7910
rect 9958 7896 10120 7898
rect 9970 7876 9989 7896
rect 10004 7894 10034 7896
rect 9853 7868 9894 7876
rect 9976 7872 9989 7876
rect 10041 7880 10120 7896
rect 10152 7896 10324 7898
rect 10152 7880 10231 7896
rect 10238 7894 10268 7896
rect 9816 7858 9845 7868
rect 9859 7858 9888 7868
rect 9903 7858 9933 7872
rect 9976 7858 10019 7872
rect 10041 7868 10231 7880
rect 10296 7876 10302 7896
rect 10026 7858 10056 7868
rect 10057 7858 10215 7868
rect 10219 7858 10249 7868
rect 10253 7858 10283 7872
rect 10311 7858 10324 7896
rect 10396 7910 10425 7926
rect 10439 7910 10468 7926
rect 10483 7916 10513 7932
rect 10541 7910 10547 7958
rect 10550 7952 10569 7958
rect 10584 7952 10614 7960
rect 10550 7944 10614 7952
rect 10550 7928 10630 7944
rect 10646 7937 10708 7968
rect 10724 7937 10786 7968
rect 10855 7966 10904 7991
rect 10919 7966 10949 7982
rect 10818 7952 10848 7960
rect 10855 7958 10965 7966
rect 10818 7944 10863 7952
rect 10550 7926 10569 7928
rect 10584 7926 10630 7928
rect 10550 7910 10630 7926
rect 10657 7924 10692 7937
rect 10733 7934 10770 7937
rect 10733 7932 10775 7934
rect 10662 7921 10692 7924
rect 10671 7917 10678 7921
rect 10678 7916 10679 7917
rect 10637 7910 10647 7916
rect 10396 7902 10431 7910
rect 10396 7876 10397 7902
rect 10404 7876 10431 7902
rect 10339 7858 10369 7872
rect 10396 7868 10431 7876
rect 10433 7902 10474 7910
rect 10433 7876 10448 7902
rect 10455 7876 10474 7902
rect 10538 7898 10569 7910
rect 10584 7898 10687 7910
rect 10699 7900 10725 7926
rect 10740 7921 10770 7932
rect 10802 7928 10864 7944
rect 10802 7926 10848 7928
rect 10802 7910 10864 7926
rect 10876 7910 10882 7958
rect 10885 7950 10965 7958
rect 10885 7948 10904 7950
rect 10919 7948 10953 7950
rect 10885 7932 10965 7948
rect 10885 7910 10904 7932
rect 10919 7916 10949 7932
rect 10977 7926 10983 8000
rect 10986 7926 11005 8070
rect 11020 7926 11026 8070
rect 11035 8000 11048 8070
rect 11100 8066 11122 8070
rect 11093 8044 11122 8058
rect 11175 8044 11191 8058
rect 11229 8054 11235 8056
rect 11242 8054 11350 8070
rect 11357 8054 11363 8056
rect 11371 8054 11386 8070
rect 11452 8064 11471 8067
rect 11093 8042 11191 8044
rect 11218 8042 11386 8054
rect 11401 8044 11417 8058
rect 11452 8045 11474 8064
rect 11484 8058 11500 8059
rect 11483 8056 11500 8058
rect 11484 8051 11500 8056
rect 11474 8044 11480 8045
rect 11483 8044 11512 8051
rect 11401 8043 11512 8044
rect 11401 8042 11518 8043
rect 11077 8034 11128 8042
rect 11175 8034 11209 8042
rect 11077 8022 11102 8034
rect 11109 8022 11128 8034
rect 11182 8032 11209 8034
rect 11218 8032 11439 8042
rect 11474 8039 11480 8042
rect 11182 8028 11439 8032
rect 11077 8014 11128 8022
rect 11175 8014 11439 8028
rect 11483 8034 11518 8042
rect 11029 7966 11048 8000
rect 11093 8006 11122 8014
rect 11093 8000 11110 8006
rect 11093 7998 11127 8000
rect 11175 7998 11191 8014
rect 11192 8004 11400 8014
rect 11401 8004 11417 8014
rect 11465 8010 11480 8025
rect 11483 8022 11484 8034
rect 11491 8022 11518 8034
rect 11483 8014 11518 8022
rect 11483 8013 11512 8014
rect 11203 8000 11417 8004
rect 11218 7998 11417 8000
rect 11452 8000 11465 8010
rect 11483 8000 11500 8013
rect 11452 7998 11500 8000
rect 11094 7994 11127 7998
rect 11090 7992 11127 7994
rect 11090 7991 11157 7992
rect 11090 7986 11121 7991
rect 11127 7986 11157 7991
rect 11090 7982 11157 7986
rect 11063 7979 11157 7982
rect 11063 7972 11112 7979
rect 11063 7966 11093 7972
rect 11112 7967 11117 7972
rect 11029 7950 11109 7966
rect 11121 7958 11157 7979
rect 11218 7974 11407 7998
rect 11452 7997 11499 7998
rect 11465 7992 11499 7997
rect 11233 7971 11407 7974
rect 11226 7968 11407 7971
rect 11435 7991 11499 7992
rect 11029 7948 11048 7950
rect 11063 7948 11097 7950
rect 11029 7932 11109 7948
rect 11029 7926 11048 7932
rect 10745 7900 10848 7910
rect 10699 7898 10848 7900
rect 10869 7898 10904 7910
rect 10538 7896 10700 7898
rect 10550 7876 10569 7896
rect 10584 7894 10614 7896
rect 10433 7868 10474 7876
rect 10556 7872 10569 7876
rect 10621 7880 10700 7896
rect 10732 7896 10904 7898
rect 10732 7880 10811 7896
rect 10818 7894 10848 7896
rect 10396 7858 10425 7868
rect 10439 7858 10468 7868
rect 10483 7858 10513 7872
rect 10556 7858 10599 7872
rect 10621 7868 10811 7880
rect 10876 7876 10882 7896
rect 10606 7858 10636 7868
rect 10637 7858 10795 7868
rect 10799 7858 10829 7868
rect 10833 7858 10863 7872
rect 10891 7858 10904 7896
rect 10976 7910 11005 7926
rect 11019 7910 11048 7926
rect 11063 7916 11093 7932
rect 11121 7910 11127 7958
rect 11130 7952 11149 7958
rect 11164 7952 11194 7960
rect 11130 7944 11194 7952
rect 11130 7928 11210 7944
rect 11226 7937 11288 7968
rect 11304 7937 11366 7968
rect 11435 7966 11484 7991
rect 11499 7966 11529 7982
rect 11398 7952 11428 7960
rect 11435 7958 11545 7966
rect 11398 7944 11443 7952
rect 11130 7926 11149 7928
rect 11164 7926 11210 7928
rect 11130 7910 11210 7926
rect 11237 7924 11272 7937
rect 11313 7934 11350 7937
rect 11313 7932 11355 7934
rect 11242 7921 11272 7924
rect 11251 7917 11258 7921
rect 11258 7916 11259 7917
rect 11217 7910 11227 7916
rect 10976 7902 11011 7910
rect 10976 7876 10977 7902
rect 10984 7876 11011 7902
rect 10919 7858 10949 7872
rect 10976 7868 11011 7876
rect 11013 7902 11054 7910
rect 11013 7876 11028 7902
rect 11035 7876 11054 7902
rect 11118 7898 11149 7910
rect 11164 7898 11267 7910
rect 11279 7900 11305 7926
rect 11320 7921 11350 7932
rect 11382 7928 11444 7944
rect 11382 7926 11428 7928
rect 11382 7910 11444 7926
rect 11456 7910 11462 7958
rect 11465 7950 11545 7958
rect 11465 7948 11484 7950
rect 11499 7948 11533 7950
rect 11465 7932 11545 7948
rect 11465 7910 11484 7932
rect 11499 7916 11529 7932
rect 11557 7926 11563 8000
rect 11566 7926 11585 8070
rect 11600 7926 11606 8070
rect 11615 8000 11628 8070
rect 11680 8066 11702 8070
rect 11673 8044 11702 8058
rect 11755 8044 11771 8058
rect 11809 8054 11815 8056
rect 11822 8054 11930 8070
rect 11937 8054 11943 8056
rect 11951 8054 11966 8070
rect 12032 8064 12051 8067
rect 11673 8042 11771 8044
rect 11798 8042 11966 8054
rect 11981 8044 11997 8058
rect 12032 8045 12054 8064
rect 12064 8058 12080 8059
rect 12063 8056 12080 8058
rect 12064 8051 12080 8056
rect 12054 8044 12060 8045
rect 12063 8044 12092 8051
rect 11981 8043 12092 8044
rect 11981 8042 12098 8043
rect 11657 8034 11708 8042
rect 11755 8034 11789 8042
rect 11657 8022 11682 8034
rect 11689 8022 11708 8034
rect 11762 8032 11789 8034
rect 11798 8032 12019 8042
rect 12054 8039 12060 8042
rect 11762 8028 12019 8032
rect 11657 8014 11708 8022
rect 11755 8014 12019 8028
rect 12063 8034 12098 8042
rect 11609 7966 11628 8000
rect 11673 8006 11702 8014
rect 11673 8000 11690 8006
rect 11673 7998 11707 8000
rect 11755 7998 11771 8014
rect 11772 8004 11980 8014
rect 11981 8004 11997 8014
rect 12045 8010 12060 8025
rect 12063 8022 12064 8034
rect 12071 8022 12098 8034
rect 12063 8014 12098 8022
rect 12063 8013 12092 8014
rect 11783 8000 11997 8004
rect 11798 7998 11997 8000
rect 12032 8000 12045 8010
rect 12063 8000 12080 8013
rect 12032 7998 12080 8000
rect 11674 7994 11707 7998
rect 11670 7992 11707 7994
rect 11670 7991 11737 7992
rect 11670 7986 11701 7991
rect 11707 7986 11737 7991
rect 11670 7982 11737 7986
rect 11643 7979 11737 7982
rect 11643 7972 11692 7979
rect 11643 7966 11673 7972
rect 11692 7967 11697 7972
rect 11609 7950 11689 7966
rect 11701 7958 11737 7979
rect 11798 7974 11987 7998
rect 12032 7997 12079 7998
rect 12045 7992 12079 7997
rect 11813 7971 11987 7974
rect 11806 7968 11987 7971
rect 12015 7991 12079 7992
rect 11609 7948 11628 7950
rect 11643 7948 11677 7950
rect 11609 7932 11689 7948
rect 11609 7926 11628 7932
rect 11325 7900 11428 7910
rect 11279 7898 11428 7900
rect 11449 7898 11484 7910
rect 11118 7896 11280 7898
rect 11130 7876 11149 7896
rect 11164 7894 11194 7896
rect 11013 7868 11054 7876
rect 11136 7872 11149 7876
rect 11201 7880 11280 7896
rect 11312 7896 11484 7898
rect 11312 7880 11391 7896
rect 11398 7894 11428 7896
rect 10976 7858 11005 7868
rect 11019 7858 11048 7868
rect 11063 7858 11093 7872
rect 11136 7858 11179 7872
rect 11201 7868 11391 7880
rect 11456 7876 11462 7896
rect 11186 7858 11216 7868
rect 11217 7858 11375 7868
rect 11379 7858 11409 7868
rect 11413 7858 11443 7872
rect 11471 7858 11484 7896
rect 11556 7910 11585 7926
rect 11599 7910 11628 7926
rect 11643 7916 11673 7932
rect 11701 7910 11707 7958
rect 11710 7952 11729 7958
rect 11744 7952 11774 7960
rect 11710 7944 11774 7952
rect 11710 7928 11790 7944
rect 11806 7937 11868 7968
rect 11884 7937 11946 7968
rect 12015 7966 12064 7991
rect 12079 7966 12109 7982
rect 11978 7952 12008 7960
rect 12015 7958 12125 7966
rect 11978 7944 12023 7952
rect 11710 7926 11729 7928
rect 11744 7926 11790 7928
rect 11710 7910 11790 7926
rect 11817 7924 11852 7937
rect 11893 7934 11930 7937
rect 11893 7932 11935 7934
rect 11822 7921 11852 7924
rect 11831 7917 11838 7921
rect 11838 7916 11839 7917
rect 11797 7910 11807 7916
rect 11556 7902 11591 7910
rect 11556 7876 11557 7902
rect 11564 7876 11591 7902
rect 11499 7858 11529 7872
rect 11556 7868 11591 7876
rect 11593 7902 11634 7910
rect 11593 7876 11608 7902
rect 11615 7876 11634 7902
rect 11698 7898 11729 7910
rect 11744 7898 11847 7910
rect 11859 7900 11885 7926
rect 11900 7921 11930 7932
rect 11962 7928 12024 7944
rect 11962 7926 12008 7928
rect 11962 7910 12024 7926
rect 12036 7910 12042 7958
rect 12045 7950 12125 7958
rect 12045 7948 12064 7950
rect 12079 7948 12113 7950
rect 12045 7932 12125 7948
rect 12045 7910 12064 7932
rect 12079 7916 12109 7932
rect 12137 7926 12143 8000
rect 12146 7926 12165 8070
rect 12180 7926 12186 8070
rect 12195 8000 12208 8070
rect 12260 8066 12282 8070
rect 12253 8044 12282 8058
rect 12335 8044 12351 8058
rect 12389 8054 12395 8056
rect 12402 8054 12510 8070
rect 12517 8054 12523 8056
rect 12531 8054 12546 8070
rect 12612 8064 12631 8067
rect 12253 8042 12351 8044
rect 12378 8042 12546 8054
rect 12561 8044 12577 8058
rect 12612 8045 12634 8064
rect 12644 8058 12660 8059
rect 12643 8056 12660 8058
rect 12644 8051 12660 8056
rect 12634 8044 12640 8045
rect 12643 8044 12672 8051
rect 12561 8043 12672 8044
rect 12561 8042 12678 8043
rect 12237 8034 12288 8042
rect 12335 8034 12369 8042
rect 12237 8022 12262 8034
rect 12269 8022 12288 8034
rect 12342 8032 12369 8034
rect 12378 8032 12599 8042
rect 12634 8039 12640 8042
rect 12342 8028 12599 8032
rect 12237 8014 12288 8022
rect 12335 8014 12599 8028
rect 12643 8034 12678 8042
rect 12189 7966 12208 8000
rect 12253 8006 12282 8014
rect 12253 8000 12270 8006
rect 12253 7998 12287 8000
rect 12335 7998 12351 8014
rect 12352 8004 12560 8014
rect 12561 8004 12577 8014
rect 12625 8010 12640 8025
rect 12643 8022 12644 8034
rect 12651 8022 12678 8034
rect 12643 8014 12678 8022
rect 12643 8013 12672 8014
rect 12363 8000 12577 8004
rect 12378 7998 12577 8000
rect 12612 8000 12625 8010
rect 12643 8000 12660 8013
rect 12612 7998 12660 8000
rect 12254 7994 12287 7998
rect 12250 7992 12287 7994
rect 12250 7991 12317 7992
rect 12250 7986 12281 7991
rect 12287 7986 12317 7991
rect 12250 7982 12317 7986
rect 12223 7979 12317 7982
rect 12223 7972 12272 7979
rect 12223 7966 12253 7972
rect 12272 7967 12277 7972
rect 12189 7950 12269 7966
rect 12281 7958 12317 7979
rect 12378 7974 12567 7998
rect 12612 7997 12659 7998
rect 12625 7992 12659 7997
rect 12393 7971 12567 7974
rect 12386 7968 12567 7971
rect 12595 7991 12659 7992
rect 12189 7948 12208 7950
rect 12223 7948 12257 7950
rect 12189 7932 12269 7948
rect 12189 7926 12208 7932
rect 11905 7900 12008 7910
rect 11859 7898 12008 7900
rect 12029 7898 12064 7910
rect 11698 7896 11860 7898
rect 11710 7876 11729 7896
rect 11744 7894 11774 7896
rect 11593 7868 11634 7876
rect 11716 7872 11729 7876
rect 11781 7880 11860 7896
rect 11892 7896 12064 7898
rect 11892 7880 11971 7896
rect 11978 7894 12008 7896
rect 11556 7858 11585 7868
rect 11599 7858 11628 7868
rect 11643 7858 11673 7872
rect 11716 7858 11759 7872
rect 11781 7868 11971 7880
rect 12036 7876 12042 7896
rect 11766 7858 11796 7868
rect 11797 7858 11955 7868
rect 11959 7858 11989 7868
rect 11993 7858 12023 7872
rect 12051 7858 12064 7896
rect 12136 7910 12165 7926
rect 12179 7910 12208 7926
rect 12223 7916 12253 7932
rect 12281 7910 12287 7958
rect 12290 7952 12309 7958
rect 12324 7952 12354 7960
rect 12290 7944 12354 7952
rect 12290 7928 12370 7944
rect 12386 7937 12448 7968
rect 12464 7937 12526 7968
rect 12595 7966 12644 7991
rect 12659 7966 12689 7982
rect 12558 7952 12588 7960
rect 12595 7958 12705 7966
rect 12558 7944 12603 7952
rect 12290 7926 12309 7928
rect 12324 7926 12370 7928
rect 12290 7910 12370 7926
rect 12397 7924 12432 7937
rect 12473 7934 12510 7937
rect 12473 7932 12515 7934
rect 12402 7921 12432 7924
rect 12411 7917 12418 7921
rect 12418 7916 12419 7917
rect 12377 7910 12387 7916
rect 12136 7902 12171 7910
rect 12136 7876 12137 7902
rect 12144 7876 12171 7902
rect 12079 7858 12109 7872
rect 12136 7868 12171 7876
rect 12173 7902 12214 7910
rect 12173 7876 12188 7902
rect 12195 7876 12214 7902
rect 12278 7898 12309 7910
rect 12324 7898 12427 7910
rect 12439 7900 12465 7926
rect 12480 7921 12510 7932
rect 12542 7928 12604 7944
rect 12542 7926 12588 7928
rect 12542 7910 12604 7926
rect 12616 7910 12622 7958
rect 12625 7950 12705 7958
rect 12625 7948 12644 7950
rect 12659 7948 12693 7950
rect 12625 7932 12705 7948
rect 12625 7910 12644 7932
rect 12659 7916 12689 7932
rect 12717 7926 12723 8000
rect 12726 7926 12745 8070
rect 12760 7926 12766 8070
rect 12775 8000 12788 8070
rect 12840 8066 12862 8070
rect 12833 8044 12862 8058
rect 12915 8044 12931 8058
rect 12969 8054 12975 8056
rect 12982 8054 13090 8070
rect 13097 8054 13103 8056
rect 13111 8054 13126 8070
rect 13192 8064 13211 8067
rect 12833 8042 12931 8044
rect 12958 8042 13126 8054
rect 13141 8044 13157 8058
rect 13192 8045 13214 8064
rect 13224 8058 13240 8059
rect 13223 8056 13240 8058
rect 13224 8051 13240 8056
rect 13214 8044 13220 8045
rect 13223 8044 13252 8051
rect 13141 8043 13252 8044
rect 13141 8042 13258 8043
rect 12817 8034 12868 8042
rect 12915 8034 12949 8042
rect 12817 8022 12842 8034
rect 12849 8022 12868 8034
rect 12922 8032 12949 8034
rect 12958 8032 13179 8042
rect 13214 8039 13220 8042
rect 12922 8028 13179 8032
rect 12817 8014 12868 8022
rect 12915 8014 13179 8028
rect 13223 8034 13258 8042
rect 12769 7966 12788 8000
rect 12833 8006 12862 8014
rect 12833 8000 12850 8006
rect 12833 7998 12867 8000
rect 12915 7998 12931 8014
rect 12932 8004 13140 8014
rect 13141 8004 13157 8014
rect 13205 8010 13220 8025
rect 13223 8022 13224 8034
rect 13231 8022 13258 8034
rect 13223 8014 13258 8022
rect 13223 8013 13252 8014
rect 12943 8000 13157 8004
rect 12958 7998 13157 8000
rect 13192 8000 13205 8010
rect 13223 8000 13240 8013
rect 13192 7998 13240 8000
rect 12834 7994 12867 7998
rect 12830 7992 12867 7994
rect 12830 7991 12897 7992
rect 12830 7986 12861 7991
rect 12867 7986 12897 7991
rect 12830 7982 12897 7986
rect 12803 7979 12897 7982
rect 12803 7972 12852 7979
rect 12803 7966 12833 7972
rect 12852 7967 12857 7972
rect 12769 7950 12849 7966
rect 12861 7958 12897 7979
rect 12958 7974 13147 7998
rect 13192 7997 13239 7998
rect 13205 7992 13239 7997
rect 12973 7971 13147 7974
rect 12966 7968 13147 7971
rect 13175 7991 13239 7992
rect 12769 7948 12788 7950
rect 12803 7948 12837 7950
rect 12769 7932 12849 7948
rect 12769 7926 12788 7932
rect 12485 7900 12588 7910
rect 12439 7898 12588 7900
rect 12609 7898 12644 7910
rect 12278 7896 12440 7898
rect 12290 7876 12309 7896
rect 12324 7894 12354 7896
rect 12173 7868 12214 7876
rect 12296 7872 12309 7876
rect 12361 7880 12440 7896
rect 12472 7896 12644 7898
rect 12472 7880 12551 7896
rect 12558 7894 12588 7896
rect 12136 7858 12165 7868
rect 12179 7858 12208 7868
rect 12223 7858 12253 7872
rect 12296 7858 12339 7872
rect 12361 7868 12551 7880
rect 12616 7876 12622 7896
rect 12346 7858 12376 7868
rect 12377 7858 12535 7868
rect 12539 7858 12569 7868
rect 12573 7858 12603 7872
rect 12631 7858 12644 7896
rect 12716 7910 12745 7926
rect 12759 7910 12788 7926
rect 12803 7916 12833 7932
rect 12861 7910 12867 7958
rect 12870 7952 12889 7958
rect 12904 7952 12934 7960
rect 12870 7944 12934 7952
rect 12870 7928 12950 7944
rect 12966 7937 13028 7968
rect 13044 7937 13106 7968
rect 13175 7966 13224 7991
rect 13239 7966 13269 7982
rect 13138 7952 13168 7960
rect 13175 7958 13285 7966
rect 13138 7944 13183 7952
rect 12870 7926 12889 7928
rect 12904 7926 12950 7928
rect 12870 7910 12950 7926
rect 12977 7924 13012 7937
rect 13053 7934 13090 7937
rect 13053 7932 13095 7934
rect 12982 7921 13012 7924
rect 12991 7917 12998 7921
rect 12998 7916 12999 7917
rect 12957 7910 12967 7916
rect 12716 7902 12751 7910
rect 12716 7876 12717 7902
rect 12724 7876 12751 7902
rect 12659 7858 12689 7872
rect 12716 7868 12751 7876
rect 12753 7902 12794 7910
rect 12753 7876 12768 7902
rect 12775 7876 12794 7902
rect 12858 7898 12889 7910
rect 12904 7898 13007 7910
rect 13019 7900 13045 7926
rect 13060 7921 13090 7932
rect 13122 7928 13184 7944
rect 13122 7926 13168 7928
rect 13122 7910 13184 7926
rect 13196 7910 13202 7958
rect 13205 7950 13285 7958
rect 13205 7948 13224 7950
rect 13239 7948 13273 7950
rect 13205 7932 13285 7948
rect 13205 7910 13224 7932
rect 13239 7916 13269 7932
rect 13297 7926 13303 8000
rect 13306 7926 13325 8070
rect 13340 7926 13346 8070
rect 13355 8000 13368 8070
rect 13420 8066 13442 8070
rect 13413 8044 13442 8058
rect 13495 8044 13511 8058
rect 13549 8054 13555 8056
rect 13562 8054 13670 8070
rect 13677 8054 13683 8056
rect 13691 8054 13706 8070
rect 13772 8064 13791 8067
rect 13413 8042 13511 8044
rect 13538 8042 13706 8054
rect 13721 8044 13737 8058
rect 13772 8045 13794 8064
rect 13804 8058 13820 8059
rect 13803 8056 13820 8058
rect 13804 8051 13820 8056
rect 13794 8044 13800 8045
rect 13803 8044 13832 8051
rect 13721 8043 13832 8044
rect 13721 8042 13838 8043
rect 13397 8034 13448 8042
rect 13495 8034 13529 8042
rect 13397 8022 13422 8034
rect 13429 8022 13448 8034
rect 13502 8032 13529 8034
rect 13538 8032 13759 8042
rect 13794 8039 13800 8042
rect 13502 8028 13759 8032
rect 13397 8014 13448 8022
rect 13495 8014 13759 8028
rect 13803 8034 13838 8042
rect 13349 7966 13368 8000
rect 13413 8006 13442 8014
rect 13413 8000 13430 8006
rect 13413 7998 13447 8000
rect 13495 7998 13511 8014
rect 13512 8004 13720 8014
rect 13721 8004 13737 8014
rect 13785 8010 13800 8025
rect 13803 8022 13804 8034
rect 13811 8022 13838 8034
rect 13803 8014 13838 8022
rect 13803 8013 13832 8014
rect 13523 8000 13737 8004
rect 13538 7998 13737 8000
rect 13772 8000 13785 8010
rect 13803 8000 13820 8013
rect 13772 7998 13820 8000
rect 13414 7994 13447 7998
rect 13410 7992 13447 7994
rect 13410 7991 13477 7992
rect 13410 7986 13441 7991
rect 13447 7986 13477 7991
rect 13410 7982 13477 7986
rect 13383 7979 13477 7982
rect 13383 7972 13432 7979
rect 13383 7966 13413 7972
rect 13432 7967 13437 7972
rect 13349 7950 13429 7966
rect 13441 7958 13477 7979
rect 13538 7974 13727 7998
rect 13772 7997 13819 7998
rect 13785 7992 13819 7997
rect 13553 7971 13727 7974
rect 13546 7968 13727 7971
rect 13755 7991 13819 7992
rect 13349 7948 13368 7950
rect 13383 7948 13417 7950
rect 13349 7932 13429 7948
rect 13349 7926 13368 7932
rect 13065 7900 13168 7910
rect 13019 7898 13168 7900
rect 13189 7898 13224 7910
rect 12858 7896 13020 7898
rect 12870 7876 12889 7896
rect 12904 7894 12934 7896
rect 12753 7868 12794 7876
rect 12876 7872 12889 7876
rect 12941 7880 13020 7896
rect 13052 7896 13224 7898
rect 13052 7880 13131 7896
rect 13138 7894 13168 7896
rect 12716 7858 12745 7868
rect 12759 7858 12788 7868
rect 12803 7858 12833 7872
rect 12876 7858 12919 7872
rect 12941 7868 13131 7880
rect 13196 7876 13202 7896
rect 12926 7858 12956 7868
rect 12957 7858 13115 7868
rect 13119 7858 13149 7868
rect 13153 7858 13183 7872
rect 13211 7858 13224 7896
rect 13296 7910 13325 7926
rect 13339 7910 13368 7926
rect 13383 7916 13413 7932
rect 13441 7910 13447 7958
rect 13450 7952 13469 7958
rect 13484 7952 13514 7960
rect 13450 7944 13514 7952
rect 13450 7928 13530 7944
rect 13546 7937 13608 7968
rect 13624 7937 13686 7968
rect 13755 7966 13804 7991
rect 13819 7966 13849 7982
rect 13718 7952 13748 7960
rect 13755 7958 13865 7966
rect 13718 7944 13763 7952
rect 13450 7926 13469 7928
rect 13484 7926 13530 7928
rect 13450 7910 13530 7926
rect 13557 7924 13592 7937
rect 13633 7934 13670 7937
rect 13633 7932 13675 7934
rect 13562 7921 13592 7924
rect 13571 7917 13578 7921
rect 13578 7916 13579 7917
rect 13537 7910 13547 7916
rect 13296 7902 13331 7910
rect 13296 7876 13297 7902
rect 13304 7876 13331 7902
rect 13239 7858 13269 7872
rect 13296 7868 13331 7876
rect 13333 7902 13374 7910
rect 13333 7876 13348 7902
rect 13355 7876 13374 7902
rect 13438 7898 13469 7910
rect 13484 7898 13587 7910
rect 13599 7900 13625 7926
rect 13640 7921 13670 7932
rect 13702 7928 13764 7944
rect 13702 7926 13748 7928
rect 13702 7910 13764 7926
rect 13776 7910 13782 7958
rect 13785 7950 13865 7958
rect 13785 7948 13804 7950
rect 13819 7948 13853 7950
rect 13785 7932 13865 7948
rect 13785 7910 13804 7932
rect 13819 7916 13849 7932
rect 13877 7926 13883 8000
rect 13886 7926 13905 8070
rect 13920 7926 13926 8070
rect 13935 8000 13948 8070
rect 14000 8066 14022 8070
rect 13993 8044 14022 8058
rect 14075 8044 14091 8058
rect 14129 8054 14135 8056
rect 14142 8054 14250 8070
rect 14257 8054 14263 8056
rect 14271 8054 14286 8070
rect 14352 8064 14371 8067
rect 13993 8042 14091 8044
rect 14118 8042 14286 8054
rect 14301 8044 14317 8058
rect 14352 8045 14374 8064
rect 14384 8058 14400 8059
rect 14383 8056 14400 8058
rect 14384 8051 14400 8056
rect 14374 8044 14380 8045
rect 14383 8044 14412 8051
rect 14301 8043 14412 8044
rect 14301 8042 14418 8043
rect 13977 8034 14028 8042
rect 14075 8034 14109 8042
rect 13977 8022 14002 8034
rect 14009 8022 14028 8034
rect 14082 8032 14109 8034
rect 14118 8032 14339 8042
rect 14374 8039 14380 8042
rect 14082 8028 14339 8032
rect 13977 8014 14028 8022
rect 14075 8014 14339 8028
rect 14383 8034 14418 8042
rect 13929 7966 13948 8000
rect 13993 8006 14022 8014
rect 13993 8000 14010 8006
rect 13993 7998 14027 8000
rect 14075 7998 14091 8014
rect 14092 8004 14300 8014
rect 14301 8004 14317 8014
rect 14365 8010 14380 8025
rect 14383 8022 14384 8034
rect 14391 8022 14418 8034
rect 14383 8014 14418 8022
rect 14383 8013 14412 8014
rect 14103 8000 14317 8004
rect 14118 7998 14317 8000
rect 14352 8000 14365 8010
rect 14383 8000 14400 8013
rect 14352 7998 14400 8000
rect 13994 7994 14027 7998
rect 13990 7992 14027 7994
rect 13990 7991 14057 7992
rect 13990 7986 14021 7991
rect 14027 7986 14057 7991
rect 13990 7982 14057 7986
rect 13963 7979 14057 7982
rect 13963 7972 14012 7979
rect 13963 7966 13993 7972
rect 14012 7967 14017 7972
rect 13929 7950 14009 7966
rect 14021 7958 14057 7979
rect 14118 7974 14307 7998
rect 14352 7997 14399 7998
rect 14365 7992 14399 7997
rect 14133 7971 14307 7974
rect 14126 7968 14307 7971
rect 14335 7991 14399 7992
rect 13929 7948 13948 7950
rect 13963 7948 13997 7950
rect 13929 7932 14009 7948
rect 13929 7926 13948 7932
rect 13645 7900 13748 7910
rect 13599 7898 13748 7900
rect 13769 7898 13804 7910
rect 13438 7896 13600 7898
rect 13450 7876 13469 7896
rect 13484 7894 13514 7896
rect 13333 7868 13374 7876
rect 13456 7872 13469 7876
rect 13521 7880 13600 7896
rect 13632 7896 13804 7898
rect 13632 7880 13711 7896
rect 13718 7894 13748 7896
rect 13296 7858 13325 7868
rect 13339 7858 13368 7868
rect 13383 7858 13413 7872
rect 13456 7858 13499 7872
rect 13521 7868 13711 7880
rect 13776 7876 13782 7896
rect 13506 7858 13536 7868
rect 13537 7858 13695 7868
rect 13699 7858 13729 7868
rect 13733 7858 13763 7872
rect 13791 7858 13804 7896
rect 13876 7910 13905 7926
rect 13919 7910 13948 7926
rect 13963 7916 13993 7932
rect 14021 7910 14027 7958
rect 14030 7952 14049 7958
rect 14064 7952 14094 7960
rect 14030 7944 14094 7952
rect 14030 7928 14110 7944
rect 14126 7937 14188 7968
rect 14204 7937 14266 7968
rect 14335 7966 14384 7991
rect 14399 7966 14429 7982
rect 14298 7952 14328 7960
rect 14335 7958 14445 7966
rect 14298 7944 14343 7952
rect 14030 7926 14049 7928
rect 14064 7926 14110 7928
rect 14030 7910 14110 7926
rect 14137 7924 14172 7937
rect 14213 7934 14250 7937
rect 14213 7932 14255 7934
rect 14142 7921 14172 7924
rect 14151 7917 14158 7921
rect 14158 7916 14159 7917
rect 14117 7910 14127 7916
rect 13876 7902 13911 7910
rect 13876 7876 13877 7902
rect 13884 7876 13911 7902
rect 13819 7858 13849 7872
rect 13876 7868 13911 7876
rect 13913 7902 13954 7910
rect 13913 7876 13928 7902
rect 13935 7876 13954 7902
rect 14018 7898 14049 7910
rect 14064 7898 14167 7910
rect 14179 7900 14205 7926
rect 14220 7921 14250 7932
rect 14282 7928 14344 7944
rect 14282 7926 14328 7928
rect 14282 7910 14344 7926
rect 14356 7910 14362 7958
rect 14365 7950 14445 7958
rect 14365 7948 14384 7950
rect 14399 7948 14433 7950
rect 14365 7932 14445 7948
rect 14365 7910 14384 7932
rect 14399 7916 14429 7932
rect 14457 7926 14463 8000
rect 14466 7926 14485 8070
rect 14500 7926 14506 8070
rect 14515 8000 14528 8070
rect 14580 8066 14602 8070
rect 14573 8044 14602 8058
rect 14655 8044 14671 8058
rect 14709 8054 14715 8056
rect 14722 8054 14830 8070
rect 14837 8054 14843 8056
rect 14851 8054 14866 8070
rect 14932 8064 14951 8067
rect 14573 8042 14671 8044
rect 14698 8042 14866 8054
rect 14881 8044 14897 8058
rect 14932 8045 14954 8064
rect 14964 8058 14980 8059
rect 14963 8056 14980 8058
rect 14964 8051 14980 8056
rect 14954 8044 14960 8045
rect 14963 8044 14992 8051
rect 14881 8043 14992 8044
rect 14881 8042 14998 8043
rect 14557 8034 14608 8042
rect 14655 8034 14689 8042
rect 14557 8022 14582 8034
rect 14589 8022 14608 8034
rect 14662 8032 14689 8034
rect 14698 8032 14919 8042
rect 14954 8039 14960 8042
rect 14662 8028 14919 8032
rect 14557 8014 14608 8022
rect 14655 8014 14919 8028
rect 14963 8034 14998 8042
rect 14509 7966 14528 8000
rect 14573 8006 14602 8014
rect 14573 8000 14590 8006
rect 14573 7998 14607 8000
rect 14655 7998 14671 8014
rect 14672 8004 14880 8014
rect 14881 8004 14897 8014
rect 14945 8010 14960 8025
rect 14963 8022 14964 8034
rect 14971 8022 14998 8034
rect 14963 8014 14998 8022
rect 14963 8013 14992 8014
rect 14683 8000 14897 8004
rect 14698 7998 14897 8000
rect 14932 8000 14945 8010
rect 14963 8000 14980 8013
rect 14932 7998 14980 8000
rect 14574 7994 14607 7998
rect 14570 7992 14607 7994
rect 14570 7991 14637 7992
rect 14570 7986 14601 7991
rect 14607 7986 14637 7991
rect 14570 7982 14637 7986
rect 14543 7979 14637 7982
rect 14543 7972 14592 7979
rect 14543 7966 14573 7972
rect 14592 7967 14597 7972
rect 14509 7950 14589 7966
rect 14601 7958 14637 7979
rect 14698 7974 14887 7998
rect 14932 7997 14979 7998
rect 14945 7992 14979 7997
rect 14713 7971 14887 7974
rect 14706 7968 14887 7971
rect 14915 7991 14979 7992
rect 14509 7948 14528 7950
rect 14543 7948 14577 7950
rect 14509 7932 14589 7948
rect 14509 7926 14528 7932
rect 14225 7900 14328 7910
rect 14179 7898 14328 7900
rect 14349 7898 14384 7910
rect 14018 7896 14180 7898
rect 14030 7876 14049 7896
rect 14064 7894 14094 7896
rect 13913 7868 13954 7876
rect 14036 7872 14049 7876
rect 14101 7880 14180 7896
rect 14212 7896 14384 7898
rect 14212 7880 14291 7896
rect 14298 7894 14328 7896
rect 13876 7858 13905 7868
rect 13919 7858 13948 7868
rect 13963 7858 13993 7872
rect 14036 7858 14079 7872
rect 14101 7868 14291 7880
rect 14356 7876 14362 7896
rect 14086 7858 14116 7868
rect 14117 7858 14275 7868
rect 14279 7858 14309 7868
rect 14313 7858 14343 7872
rect 14371 7858 14384 7896
rect 14456 7910 14485 7926
rect 14499 7910 14528 7926
rect 14543 7916 14573 7932
rect 14601 7910 14607 7958
rect 14610 7952 14629 7958
rect 14644 7952 14674 7960
rect 14610 7944 14674 7952
rect 14610 7928 14690 7944
rect 14706 7937 14768 7968
rect 14784 7937 14846 7968
rect 14915 7966 14964 7991
rect 14979 7966 15009 7982
rect 14878 7952 14908 7960
rect 14915 7958 15025 7966
rect 14878 7944 14923 7952
rect 14610 7926 14629 7928
rect 14644 7926 14690 7928
rect 14610 7910 14690 7926
rect 14717 7924 14752 7937
rect 14793 7934 14830 7937
rect 14793 7932 14835 7934
rect 14722 7921 14752 7924
rect 14731 7917 14738 7921
rect 14738 7916 14739 7917
rect 14697 7910 14707 7916
rect 14456 7902 14491 7910
rect 14456 7876 14457 7902
rect 14464 7876 14491 7902
rect 14399 7858 14429 7872
rect 14456 7868 14491 7876
rect 14493 7902 14534 7910
rect 14493 7876 14508 7902
rect 14515 7876 14534 7902
rect 14598 7898 14629 7910
rect 14644 7898 14747 7910
rect 14759 7900 14785 7926
rect 14800 7921 14830 7932
rect 14862 7928 14924 7944
rect 14862 7926 14908 7928
rect 14862 7910 14924 7926
rect 14936 7910 14942 7958
rect 14945 7950 15025 7958
rect 14945 7948 14964 7950
rect 14979 7948 15013 7950
rect 14945 7932 15025 7948
rect 14945 7910 14964 7932
rect 14979 7916 15009 7932
rect 15037 7926 15043 8000
rect 15046 7926 15065 8070
rect 15080 7926 15086 8070
rect 15095 8000 15108 8070
rect 15160 8066 15182 8070
rect 15153 8044 15182 8058
rect 15235 8044 15251 8058
rect 15289 8054 15295 8056
rect 15302 8054 15410 8070
rect 15417 8054 15423 8056
rect 15431 8054 15446 8070
rect 15512 8064 15531 8067
rect 15153 8042 15251 8044
rect 15278 8042 15446 8054
rect 15461 8044 15477 8058
rect 15512 8045 15534 8064
rect 15544 8058 15560 8059
rect 15543 8056 15560 8058
rect 15544 8051 15560 8056
rect 15534 8044 15540 8045
rect 15543 8044 15572 8051
rect 15461 8043 15572 8044
rect 15461 8042 15578 8043
rect 15137 8034 15188 8042
rect 15235 8034 15269 8042
rect 15137 8022 15162 8034
rect 15169 8022 15188 8034
rect 15242 8032 15269 8034
rect 15278 8032 15499 8042
rect 15534 8039 15540 8042
rect 15242 8028 15499 8032
rect 15137 8014 15188 8022
rect 15235 8014 15499 8028
rect 15543 8034 15578 8042
rect 15089 7966 15108 8000
rect 15153 8006 15182 8014
rect 15153 8000 15170 8006
rect 15153 7998 15187 8000
rect 15235 7998 15251 8014
rect 15252 8004 15460 8014
rect 15461 8004 15477 8014
rect 15525 8010 15540 8025
rect 15543 8022 15544 8034
rect 15551 8022 15578 8034
rect 15543 8014 15578 8022
rect 15543 8013 15572 8014
rect 15263 8000 15477 8004
rect 15278 7998 15477 8000
rect 15512 8000 15525 8010
rect 15543 8000 15560 8013
rect 15512 7998 15560 8000
rect 15154 7994 15187 7998
rect 15150 7992 15187 7994
rect 15150 7991 15217 7992
rect 15150 7986 15181 7991
rect 15187 7986 15217 7991
rect 15150 7982 15217 7986
rect 15123 7979 15217 7982
rect 15123 7972 15172 7979
rect 15123 7966 15153 7972
rect 15172 7967 15177 7972
rect 15089 7950 15169 7966
rect 15181 7958 15217 7979
rect 15278 7974 15467 7998
rect 15512 7997 15559 7998
rect 15525 7992 15559 7997
rect 15293 7971 15467 7974
rect 15286 7968 15467 7971
rect 15495 7991 15559 7992
rect 15089 7948 15108 7950
rect 15123 7948 15157 7950
rect 15089 7932 15169 7948
rect 15089 7926 15108 7932
rect 14805 7900 14908 7910
rect 14759 7898 14908 7900
rect 14929 7898 14964 7910
rect 14598 7896 14760 7898
rect 14610 7876 14629 7896
rect 14644 7894 14674 7896
rect 14493 7868 14534 7876
rect 14616 7872 14629 7876
rect 14681 7880 14760 7896
rect 14792 7896 14964 7898
rect 14792 7880 14871 7896
rect 14878 7894 14908 7896
rect 14456 7858 14485 7868
rect 14499 7858 14528 7868
rect 14543 7858 14573 7872
rect 14616 7858 14659 7872
rect 14681 7868 14871 7880
rect 14936 7876 14942 7896
rect 14666 7858 14696 7868
rect 14697 7858 14855 7868
rect 14859 7858 14889 7868
rect 14893 7858 14923 7872
rect 14951 7858 14964 7896
rect 15036 7910 15065 7926
rect 15079 7910 15108 7926
rect 15123 7916 15153 7932
rect 15181 7910 15187 7958
rect 15190 7952 15209 7958
rect 15224 7952 15254 7960
rect 15190 7944 15254 7952
rect 15190 7928 15270 7944
rect 15286 7937 15348 7968
rect 15364 7937 15426 7968
rect 15495 7966 15544 7991
rect 15559 7966 15589 7982
rect 15458 7952 15488 7960
rect 15495 7958 15605 7966
rect 15458 7944 15503 7952
rect 15190 7926 15209 7928
rect 15224 7926 15270 7928
rect 15190 7910 15270 7926
rect 15297 7924 15332 7937
rect 15373 7934 15410 7937
rect 15373 7932 15415 7934
rect 15302 7921 15332 7924
rect 15311 7917 15318 7921
rect 15318 7916 15319 7917
rect 15277 7910 15287 7916
rect 15036 7902 15071 7910
rect 15036 7876 15037 7902
rect 15044 7876 15071 7902
rect 14979 7858 15009 7872
rect 15036 7868 15071 7876
rect 15073 7902 15114 7910
rect 15073 7876 15088 7902
rect 15095 7876 15114 7902
rect 15178 7898 15209 7910
rect 15224 7898 15327 7910
rect 15339 7900 15365 7926
rect 15380 7921 15410 7932
rect 15442 7928 15504 7944
rect 15442 7926 15488 7928
rect 15442 7910 15504 7926
rect 15516 7910 15522 7958
rect 15525 7950 15605 7958
rect 15525 7948 15544 7950
rect 15559 7948 15593 7950
rect 15525 7932 15605 7948
rect 15525 7910 15544 7932
rect 15559 7916 15589 7932
rect 15617 7926 15623 8000
rect 15626 7926 15645 8070
rect 15660 7926 15666 8070
rect 15675 8000 15688 8070
rect 15740 8066 15762 8070
rect 15733 8044 15762 8058
rect 15815 8044 15831 8058
rect 15869 8054 15875 8056
rect 15882 8054 15990 8070
rect 15997 8054 16003 8056
rect 16011 8054 16026 8070
rect 16092 8064 16111 8067
rect 15733 8042 15831 8044
rect 15858 8042 16026 8054
rect 16041 8044 16057 8058
rect 16092 8045 16114 8064
rect 16124 8058 16140 8059
rect 16123 8056 16140 8058
rect 16124 8051 16140 8056
rect 16114 8044 16120 8045
rect 16123 8044 16152 8051
rect 16041 8043 16152 8044
rect 16041 8042 16158 8043
rect 15717 8034 15768 8042
rect 15815 8034 15849 8042
rect 15717 8022 15742 8034
rect 15749 8022 15768 8034
rect 15822 8032 15849 8034
rect 15858 8032 16079 8042
rect 16114 8039 16120 8042
rect 15822 8028 16079 8032
rect 15717 8014 15768 8022
rect 15815 8014 16079 8028
rect 16123 8034 16158 8042
rect 15669 7966 15688 8000
rect 15733 8006 15762 8014
rect 15733 8000 15750 8006
rect 15733 7998 15767 8000
rect 15815 7998 15831 8014
rect 15832 8004 16040 8014
rect 16041 8004 16057 8014
rect 16105 8010 16120 8025
rect 16123 8022 16124 8034
rect 16131 8022 16158 8034
rect 16123 8014 16158 8022
rect 16123 8013 16152 8014
rect 15843 8000 16057 8004
rect 15858 7998 16057 8000
rect 16092 8000 16105 8010
rect 16123 8000 16140 8013
rect 16092 7998 16140 8000
rect 15734 7994 15767 7998
rect 15730 7992 15767 7994
rect 15730 7991 15797 7992
rect 15730 7986 15761 7991
rect 15767 7986 15797 7991
rect 15730 7982 15797 7986
rect 15703 7979 15797 7982
rect 15703 7972 15752 7979
rect 15703 7966 15733 7972
rect 15752 7967 15757 7972
rect 15669 7950 15749 7966
rect 15761 7958 15797 7979
rect 15858 7974 16047 7998
rect 16092 7997 16139 7998
rect 16105 7992 16139 7997
rect 15873 7971 16047 7974
rect 15866 7968 16047 7971
rect 16075 7991 16139 7992
rect 15669 7948 15688 7950
rect 15703 7948 15737 7950
rect 15669 7932 15749 7948
rect 15669 7926 15688 7932
rect 15385 7900 15488 7910
rect 15339 7898 15488 7900
rect 15509 7898 15544 7910
rect 15178 7896 15340 7898
rect 15190 7876 15209 7896
rect 15224 7894 15254 7896
rect 15073 7868 15114 7876
rect 15196 7872 15209 7876
rect 15261 7880 15340 7896
rect 15372 7896 15544 7898
rect 15372 7880 15451 7896
rect 15458 7894 15488 7896
rect 15036 7858 15065 7868
rect 15079 7858 15108 7868
rect 15123 7858 15153 7872
rect 15196 7858 15239 7872
rect 15261 7868 15451 7880
rect 15516 7876 15522 7896
rect 15246 7858 15276 7868
rect 15277 7858 15435 7868
rect 15439 7858 15469 7868
rect 15473 7858 15503 7872
rect 15531 7858 15544 7896
rect 15616 7910 15645 7926
rect 15659 7910 15688 7926
rect 15703 7916 15733 7932
rect 15761 7910 15767 7958
rect 15770 7952 15789 7958
rect 15804 7952 15834 7960
rect 15770 7944 15834 7952
rect 15770 7928 15850 7944
rect 15866 7937 15928 7968
rect 15944 7937 16006 7968
rect 16075 7966 16124 7991
rect 16139 7966 16169 7982
rect 16038 7952 16068 7960
rect 16075 7958 16185 7966
rect 16038 7944 16083 7952
rect 15770 7926 15789 7928
rect 15804 7926 15850 7928
rect 15770 7910 15850 7926
rect 15877 7924 15912 7937
rect 15953 7934 15990 7937
rect 15953 7932 15995 7934
rect 15882 7921 15912 7924
rect 15891 7917 15898 7921
rect 15898 7916 15899 7917
rect 15857 7910 15867 7916
rect 15616 7902 15651 7910
rect 15616 7876 15617 7902
rect 15624 7876 15651 7902
rect 15559 7858 15589 7872
rect 15616 7868 15651 7876
rect 15653 7902 15694 7910
rect 15653 7876 15668 7902
rect 15675 7876 15694 7902
rect 15758 7898 15789 7910
rect 15804 7898 15907 7910
rect 15919 7900 15945 7926
rect 15960 7921 15990 7932
rect 16022 7928 16084 7944
rect 16022 7926 16068 7928
rect 16022 7910 16084 7926
rect 16096 7910 16102 7958
rect 16105 7950 16185 7958
rect 16105 7948 16124 7950
rect 16139 7948 16173 7950
rect 16105 7932 16185 7948
rect 16105 7910 16124 7932
rect 16139 7916 16169 7932
rect 16197 7926 16203 8000
rect 16206 7926 16225 8070
rect 16240 7926 16246 8070
rect 16255 8000 16268 8070
rect 16320 8066 16342 8070
rect 16313 8044 16342 8058
rect 16395 8044 16411 8058
rect 16449 8054 16455 8056
rect 16462 8054 16570 8070
rect 16577 8054 16583 8056
rect 16591 8054 16606 8070
rect 16672 8064 16691 8067
rect 16313 8042 16411 8044
rect 16438 8042 16606 8054
rect 16621 8044 16637 8058
rect 16672 8045 16694 8064
rect 16704 8058 16720 8059
rect 16703 8056 16720 8058
rect 16704 8051 16720 8056
rect 16694 8044 16700 8045
rect 16703 8044 16732 8051
rect 16621 8043 16732 8044
rect 16621 8042 16738 8043
rect 16297 8034 16348 8042
rect 16395 8034 16429 8042
rect 16297 8022 16322 8034
rect 16329 8022 16348 8034
rect 16402 8032 16429 8034
rect 16438 8032 16659 8042
rect 16694 8039 16700 8042
rect 16402 8028 16659 8032
rect 16297 8014 16348 8022
rect 16395 8014 16659 8028
rect 16703 8034 16738 8042
rect 16249 7966 16268 8000
rect 16313 8006 16342 8014
rect 16313 8000 16330 8006
rect 16313 7998 16347 8000
rect 16395 7998 16411 8014
rect 16412 8004 16620 8014
rect 16621 8004 16637 8014
rect 16685 8010 16700 8025
rect 16703 8022 16704 8034
rect 16711 8022 16738 8034
rect 16703 8014 16738 8022
rect 16703 8013 16732 8014
rect 16423 8000 16637 8004
rect 16438 7998 16637 8000
rect 16672 8000 16685 8010
rect 16703 8000 16720 8013
rect 16672 7998 16720 8000
rect 16314 7994 16347 7998
rect 16310 7992 16347 7994
rect 16310 7991 16377 7992
rect 16310 7986 16341 7991
rect 16347 7986 16377 7991
rect 16310 7982 16377 7986
rect 16283 7979 16377 7982
rect 16283 7972 16332 7979
rect 16283 7966 16313 7972
rect 16332 7967 16337 7972
rect 16249 7950 16329 7966
rect 16341 7958 16377 7979
rect 16438 7974 16627 7998
rect 16672 7997 16719 7998
rect 16685 7992 16719 7997
rect 16453 7971 16627 7974
rect 16446 7968 16627 7971
rect 16655 7991 16719 7992
rect 16249 7948 16268 7950
rect 16283 7948 16317 7950
rect 16249 7932 16329 7948
rect 16249 7926 16268 7932
rect 15965 7900 16068 7910
rect 15919 7898 16068 7900
rect 16089 7898 16124 7910
rect 15758 7896 15920 7898
rect 15770 7876 15789 7896
rect 15804 7894 15834 7896
rect 15653 7868 15694 7876
rect 15776 7872 15789 7876
rect 15841 7880 15920 7896
rect 15952 7896 16124 7898
rect 15952 7880 16031 7896
rect 16038 7894 16068 7896
rect 15616 7858 15645 7868
rect 15659 7858 15688 7868
rect 15703 7858 15733 7872
rect 15776 7858 15819 7872
rect 15841 7868 16031 7880
rect 16096 7876 16102 7896
rect 15826 7858 15856 7868
rect 15857 7858 16015 7868
rect 16019 7858 16049 7868
rect 16053 7858 16083 7872
rect 16111 7858 16124 7896
rect 16196 7910 16225 7926
rect 16239 7910 16268 7926
rect 16283 7916 16313 7932
rect 16341 7910 16347 7958
rect 16350 7952 16369 7958
rect 16384 7952 16414 7960
rect 16350 7944 16414 7952
rect 16350 7928 16430 7944
rect 16446 7937 16508 7968
rect 16524 7937 16586 7968
rect 16655 7966 16704 7991
rect 16719 7966 16749 7982
rect 16618 7952 16648 7960
rect 16655 7958 16765 7966
rect 16618 7944 16663 7952
rect 16350 7926 16369 7928
rect 16384 7926 16430 7928
rect 16350 7910 16430 7926
rect 16457 7924 16492 7937
rect 16533 7934 16570 7937
rect 16533 7932 16575 7934
rect 16462 7921 16492 7924
rect 16471 7917 16478 7921
rect 16478 7916 16479 7917
rect 16437 7910 16447 7916
rect 16196 7902 16231 7910
rect 16196 7876 16197 7902
rect 16204 7876 16231 7902
rect 16139 7858 16169 7872
rect 16196 7868 16231 7876
rect 16233 7902 16274 7910
rect 16233 7876 16248 7902
rect 16255 7876 16274 7902
rect 16338 7898 16369 7910
rect 16384 7898 16487 7910
rect 16499 7900 16525 7926
rect 16540 7921 16570 7932
rect 16602 7928 16664 7944
rect 16602 7926 16648 7928
rect 16602 7910 16664 7926
rect 16676 7910 16682 7958
rect 16685 7950 16765 7958
rect 16685 7948 16704 7950
rect 16719 7948 16753 7950
rect 16685 7932 16765 7948
rect 16685 7910 16704 7932
rect 16719 7916 16749 7932
rect 16777 7926 16783 8000
rect 16786 7926 16805 8070
rect 16820 7926 16826 8070
rect 16835 8000 16848 8070
rect 16900 8066 16922 8070
rect 16893 8044 16922 8058
rect 16975 8044 16991 8058
rect 17029 8054 17035 8056
rect 17042 8054 17150 8070
rect 17157 8054 17163 8056
rect 17171 8054 17186 8070
rect 17252 8064 17271 8067
rect 16893 8042 16991 8044
rect 17018 8042 17186 8054
rect 17201 8044 17217 8058
rect 17252 8045 17274 8064
rect 17284 8058 17300 8059
rect 17283 8056 17300 8058
rect 17284 8051 17300 8056
rect 17274 8044 17280 8045
rect 17283 8044 17312 8051
rect 17201 8043 17312 8044
rect 17201 8042 17318 8043
rect 16877 8034 16928 8042
rect 16975 8034 17009 8042
rect 16877 8022 16902 8034
rect 16909 8022 16928 8034
rect 16982 8032 17009 8034
rect 17018 8032 17239 8042
rect 17274 8039 17280 8042
rect 16982 8028 17239 8032
rect 16877 8014 16928 8022
rect 16975 8014 17239 8028
rect 17283 8034 17318 8042
rect 16829 7966 16848 8000
rect 16893 8006 16922 8014
rect 16893 8000 16910 8006
rect 16893 7998 16927 8000
rect 16975 7998 16991 8014
rect 16992 8004 17200 8014
rect 17201 8004 17217 8014
rect 17265 8010 17280 8025
rect 17283 8022 17284 8034
rect 17291 8022 17318 8034
rect 17283 8014 17318 8022
rect 17283 8013 17312 8014
rect 17003 8000 17217 8004
rect 17018 7998 17217 8000
rect 17252 8000 17265 8010
rect 17283 8000 17300 8013
rect 17252 7998 17300 8000
rect 16894 7994 16927 7998
rect 16890 7992 16927 7994
rect 16890 7991 16957 7992
rect 16890 7986 16921 7991
rect 16927 7986 16957 7991
rect 16890 7982 16957 7986
rect 16863 7979 16957 7982
rect 16863 7972 16912 7979
rect 16863 7966 16893 7972
rect 16912 7967 16917 7972
rect 16829 7950 16909 7966
rect 16921 7958 16957 7979
rect 17018 7974 17207 7998
rect 17252 7997 17299 7998
rect 17265 7992 17299 7997
rect 17033 7971 17207 7974
rect 17026 7968 17207 7971
rect 17235 7991 17299 7992
rect 16829 7948 16848 7950
rect 16863 7948 16897 7950
rect 16829 7932 16909 7948
rect 16829 7926 16848 7932
rect 16545 7900 16648 7910
rect 16499 7898 16648 7900
rect 16669 7898 16704 7910
rect 16338 7896 16500 7898
rect 16350 7876 16369 7896
rect 16384 7894 16414 7896
rect 16233 7868 16274 7876
rect 16356 7872 16369 7876
rect 16421 7880 16500 7896
rect 16532 7896 16704 7898
rect 16532 7880 16611 7896
rect 16618 7894 16648 7896
rect 16196 7858 16225 7868
rect 16239 7858 16268 7868
rect 16283 7858 16313 7872
rect 16356 7858 16399 7872
rect 16421 7868 16611 7880
rect 16676 7876 16682 7896
rect 16406 7858 16436 7868
rect 16437 7858 16595 7868
rect 16599 7858 16629 7868
rect 16633 7858 16663 7872
rect 16691 7858 16704 7896
rect 16776 7910 16805 7926
rect 16819 7910 16848 7926
rect 16863 7916 16893 7932
rect 16921 7910 16927 7958
rect 16930 7952 16949 7958
rect 16964 7952 16994 7960
rect 16930 7944 16994 7952
rect 16930 7928 17010 7944
rect 17026 7937 17088 7968
rect 17104 7937 17166 7968
rect 17235 7966 17284 7991
rect 17299 7966 17329 7982
rect 17198 7952 17228 7960
rect 17235 7958 17345 7966
rect 17198 7944 17243 7952
rect 16930 7926 16949 7928
rect 16964 7926 17010 7928
rect 16930 7910 17010 7926
rect 17037 7924 17072 7937
rect 17113 7934 17150 7937
rect 17113 7932 17155 7934
rect 17042 7921 17072 7924
rect 17051 7917 17058 7921
rect 17058 7916 17059 7917
rect 17017 7910 17027 7916
rect 16776 7902 16811 7910
rect 16776 7876 16777 7902
rect 16784 7876 16811 7902
rect 16719 7858 16749 7872
rect 16776 7868 16811 7876
rect 16813 7902 16854 7910
rect 16813 7876 16828 7902
rect 16835 7876 16854 7902
rect 16918 7898 16949 7910
rect 16964 7898 17067 7910
rect 17079 7900 17105 7926
rect 17120 7921 17150 7932
rect 17182 7928 17244 7944
rect 17182 7926 17228 7928
rect 17182 7910 17244 7926
rect 17256 7910 17262 7958
rect 17265 7950 17345 7958
rect 17265 7948 17284 7950
rect 17299 7948 17333 7950
rect 17265 7932 17345 7948
rect 17265 7910 17284 7932
rect 17299 7916 17329 7932
rect 17357 7926 17363 8000
rect 17366 7926 17385 8070
rect 17400 7926 17406 8070
rect 17415 8000 17428 8070
rect 17480 8066 17502 8070
rect 17473 8044 17502 8058
rect 17555 8044 17571 8058
rect 17609 8054 17615 8056
rect 17622 8054 17730 8070
rect 17737 8054 17743 8056
rect 17751 8054 17766 8070
rect 17832 8064 17851 8067
rect 17473 8042 17571 8044
rect 17598 8042 17766 8054
rect 17781 8044 17797 8058
rect 17832 8045 17854 8064
rect 17864 8058 17880 8059
rect 17863 8056 17880 8058
rect 17864 8051 17880 8056
rect 17854 8044 17860 8045
rect 17863 8044 17892 8051
rect 17781 8043 17892 8044
rect 17781 8042 17898 8043
rect 17457 8034 17508 8042
rect 17555 8034 17589 8042
rect 17457 8022 17482 8034
rect 17489 8022 17508 8034
rect 17562 8032 17589 8034
rect 17598 8032 17819 8042
rect 17854 8039 17860 8042
rect 17562 8028 17819 8032
rect 17457 8014 17508 8022
rect 17555 8014 17819 8028
rect 17863 8034 17898 8042
rect 17409 7966 17428 8000
rect 17473 8006 17502 8014
rect 17473 8000 17490 8006
rect 17473 7998 17507 8000
rect 17555 7998 17571 8014
rect 17572 8004 17780 8014
rect 17781 8004 17797 8014
rect 17845 8010 17860 8025
rect 17863 8022 17864 8034
rect 17871 8022 17898 8034
rect 17863 8014 17898 8022
rect 17863 8013 17892 8014
rect 17583 8000 17797 8004
rect 17598 7998 17797 8000
rect 17832 8000 17845 8010
rect 17863 8000 17880 8013
rect 17832 7998 17880 8000
rect 17474 7994 17507 7998
rect 17470 7992 17507 7994
rect 17470 7991 17537 7992
rect 17470 7986 17501 7991
rect 17507 7986 17537 7991
rect 17470 7982 17537 7986
rect 17443 7979 17537 7982
rect 17443 7972 17492 7979
rect 17443 7966 17473 7972
rect 17492 7967 17497 7972
rect 17409 7950 17489 7966
rect 17501 7958 17537 7979
rect 17598 7974 17787 7998
rect 17832 7997 17879 7998
rect 17845 7992 17879 7997
rect 17613 7971 17787 7974
rect 17606 7968 17787 7971
rect 17815 7991 17879 7992
rect 17409 7948 17428 7950
rect 17443 7948 17477 7950
rect 17409 7932 17489 7948
rect 17409 7926 17428 7932
rect 17125 7900 17228 7910
rect 17079 7898 17228 7900
rect 17249 7898 17284 7910
rect 16918 7896 17080 7898
rect 16930 7876 16949 7896
rect 16964 7894 16994 7896
rect 16813 7868 16854 7876
rect 16936 7872 16949 7876
rect 17001 7880 17080 7896
rect 17112 7896 17284 7898
rect 17112 7880 17191 7896
rect 17198 7894 17228 7896
rect 16776 7858 16805 7868
rect 16819 7858 16848 7868
rect 16863 7858 16893 7872
rect 16936 7858 16979 7872
rect 17001 7868 17191 7880
rect 17256 7876 17262 7896
rect 16986 7858 17016 7868
rect 17017 7858 17175 7868
rect 17179 7858 17209 7868
rect 17213 7858 17243 7872
rect 17271 7858 17284 7896
rect 17356 7910 17385 7926
rect 17399 7910 17428 7926
rect 17443 7916 17473 7932
rect 17501 7910 17507 7958
rect 17510 7952 17529 7958
rect 17544 7952 17574 7960
rect 17510 7944 17574 7952
rect 17510 7928 17590 7944
rect 17606 7937 17668 7968
rect 17684 7937 17746 7968
rect 17815 7966 17864 7991
rect 17879 7966 17909 7982
rect 17778 7952 17808 7960
rect 17815 7958 17925 7966
rect 17778 7944 17823 7952
rect 17510 7926 17529 7928
rect 17544 7926 17590 7928
rect 17510 7910 17590 7926
rect 17617 7924 17652 7937
rect 17693 7934 17730 7937
rect 17693 7932 17735 7934
rect 17622 7921 17652 7924
rect 17631 7917 17638 7921
rect 17638 7916 17639 7917
rect 17597 7910 17607 7916
rect 17356 7902 17391 7910
rect 17356 7876 17357 7902
rect 17364 7876 17391 7902
rect 17299 7858 17329 7872
rect 17356 7868 17391 7876
rect 17393 7902 17434 7910
rect 17393 7876 17408 7902
rect 17415 7876 17434 7902
rect 17498 7898 17529 7910
rect 17544 7898 17647 7910
rect 17659 7900 17685 7926
rect 17700 7921 17730 7932
rect 17762 7928 17824 7944
rect 17762 7926 17808 7928
rect 17762 7910 17824 7926
rect 17836 7910 17842 7958
rect 17845 7950 17925 7958
rect 17845 7948 17864 7950
rect 17879 7948 17913 7950
rect 17845 7932 17925 7948
rect 17845 7910 17864 7932
rect 17879 7916 17909 7932
rect 17937 7926 17943 8000
rect 17946 7926 17965 8070
rect 17980 7926 17986 8070
rect 17995 8000 18008 8070
rect 18060 8066 18082 8070
rect 18053 8044 18082 8058
rect 18135 8044 18151 8058
rect 18189 8054 18195 8056
rect 18202 8054 18310 8070
rect 18317 8054 18323 8056
rect 18331 8054 18346 8070
rect 18412 8064 18431 8067
rect 18053 8042 18151 8044
rect 18178 8042 18346 8054
rect 18361 8044 18377 8058
rect 18412 8045 18434 8064
rect 18444 8058 18460 8059
rect 18443 8056 18460 8058
rect 18444 8051 18460 8056
rect 18434 8044 18440 8045
rect 18443 8044 18472 8051
rect 18361 8043 18472 8044
rect 18361 8042 18478 8043
rect 18037 8034 18088 8042
rect 18135 8034 18169 8042
rect 18037 8022 18062 8034
rect 18069 8022 18088 8034
rect 18142 8032 18169 8034
rect 18178 8032 18399 8042
rect 18434 8039 18440 8042
rect 18142 8028 18399 8032
rect 18037 8014 18088 8022
rect 18135 8014 18399 8028
rect 18443 8034 18478 8042
rect 17989 7966 18008 8000
rect 18053 8006 18082 8014
rect 18053 8000 18070 8006
rect 18053 7998 18087 8000
rect 18135 7998 18151 8014
rect 18152 8004 18360 8014
rect 18361 8004 18377 8014
rect 18425 8010 18440 8025
rect 18443 8022 18444 8034
rect 18451 8022 18478 8034
rect 18443 8014 18478 8022
rect 18443 8013 18472 8014
rect 18163 8000 18377 8004
rect 18178 7998 18377 8000
rect 18412 8000 18425 8010
rect 18443 8000 18460 8013
rect 18412 7998 18460 8000
rect 18054 7994 18087 7998
rect 18050 7992 18087 7994
rect 18050 7991 18117 7992
rect 18050 7986 18081 7991
rect 18087 7986 18117 7991
rect 18050 7982 18117 7986
rect 18023 7979 18117 7982
rect 18023 7972 18072 7979
rect 18023 7966 18053 7972
rect 18072 7967 18077 7972
rect 17989 7950 18069 7966
rect 18081 7958 18117 7979
rect 18178 7974 18367 7998
rect 18412 7997 18459 7998
rect 18425 7992 18459 7997
rect 18193 7971 18367 7974
rect 18186 7968 18367 7971
rect 18395 7991 18459 7992
rect 17989 7948 18008 7950
rect 18023 7948 18057 7950
rect 17989 7932 18069 7948
rect 17989 7926 18008 7932
rect 17705 7900 17808 7910
rect 17659 7898 17808 7900
rect 17829 7898 17864 7910
rect 17498 7896 17660 7898
rect 17510 7876 17529 7896
rect 17544 7894 17574 7896
rect 17393 7868 17434 7876
rect 17516 7872 17529 7876
rect 17581 7880 17660 7896
rect 17692 7896 17864 7898
rect 17692 7880 17771 7896
rect 17778 7894 17808 7896
rect 17356 7858 17385 7868
rect 17399 7858 17428 7868
rect 17443 7858 17473 7872
rect 17516 7858 17559 7872
rect 17581 7868 17771 7880
rect 17836 7876 17842 7896
rect 17566 7858 17596 7868
rect 17597 7858 17755 7868
rect 17759 7858 17789 7868
rect 17793 7858 17823 7872
rect 17851 7858 17864 7896
rect 17936 7910 17965 7926
rect 17979 7910 18008 7926
rect 18023 7916 18053 7932
rect 18081 7910 18087 7958
rect 18090 7952 18109 7958
rect 18124 7952 18154 7960
rect 18090 7944 18154 7952
rect 18090 7928 18170 7944
rect 18186 7937 18248 7968
rect 18264 7937 18326 7968
rect 18395 7966 18444 7991
rect 18459 7966 18489 7982
rect 18358 7952 18388 7960
rect 18395 7958 18505 7966
rect 18358 7944 18403 7952
rect 18090 7926 18109 7928
rect 18124 7926 18170 7928
rect 18090 7910 18170 7926
rect 18197 7924 18232 7937
rect 18273 7934 18310 7937
rect 18273 7932 18315 7934
rect 18202 7921 18232 7924
rect 18211 7917 18218 7921
rect 18218 7916 18219 7917
rect 18177 7910 18187 7916
rect 17936 7902 17971 7910
rect 17936 7876 17937 7902
rect 17944 7876 17971 7902
rect 17879 7858 17909 7872
rect 17936 7868 17971 7876
rect 17973 7902 18014 7910
rect 17973 7876 17988 7902
rect 17995 7876 18014 7902
rect 18078 7898 18109 7910
rect 18124 7898 18227 7910
rect 18239 7900 18265 7926
rect 18280 7921 18310 7932
rect 18342 7928 18404 7944
rect 18342 7926 18388 7928
rect 18342 7910 18404 7926
rect 18416 7910 18422 7958
rect 18425 7950 18505 7958
rect 18425 7948 18444 7950
rect 18459 7948 18493 7950
rect 18425 7932 18505 7948
rect 18425 7910 18444 7932
rect 18459 7916 18489 7932
rect 18517 7926 18523 8000
rect 18532 7926 18545 8070
rect 18285 7900 18388 7910
rect 18239 7898 18388 7900
rect 18409 7898 18444 7910
rect 18078 7896 18240 7898
rect 18090 7876 18109 7896
rect 18124 7894 18154 7896
rect 17973 7868 18014 7876
rect 18096 7872 18109 7876
rect 18161 7880 18240 7896
rect 18272 7896 18444 7898
rect 18272 7880 18351 7896
rect 18358 7894 18388 7896
rect 17936 7858 17965 7868
rect 17979 7858 18008 7868
rect 18023 7858 18053 7872
rect 18096 7858 18139 7872
rect 18161 7868 18351 7880
rect 18416 7876 18422 7896
rect 18146 7858 18176 7868
rect 18177 7858 18335 7868
rect 18339 7858 18369 7868
rect 18373 7858 18403 7872
rect 18431 7858 18444 7896
rect 18516 7910 18545 7926
rect 18516 7902 18551 7910
rect 18516 7876 18517 7902
rect 18524 7876 18551 7902
rect 18459 7858 18489 7872
rect 18516 7868 18551 7876
rect 18516 7858 18545 7868
rect -1 7852 18545 7858
rect 0 7844 18545 7852
rect 15 7814 28 7844
rect 43 7830 73 7844
rect 116 7830 159 7844
rect 166 7830 386 7844
rect 393 7830 423 7844
rect 83 7816 98 7828
rect 117 7816 130 7830
rect 198 7826 351 7830
rect 80 7814 102 7816
rect 180 7814 372 7826
rect 451 7814 464 7844
rect 479 7830 509 7844
rect 546 7814 565 7844
rect 580 7814 586 7844
rect 595 7814 608 7844
rect 623 7830 653 7844
rect 696 7830 739 7844
rect 746 7830 966 7844
rect 973 7830 1003 7844
rect 663 7816 678 7828
rect 697 7816 710 7830
rect 778 7826 931 7830
rect 660 7814 682 7816
rect 760 7814 952 7826
rect 1031 7814 1044 7844
rect 1059 7830 1089 7844
rect 1126 7814 1145 7844
rect 1160 7814 1166 7844
rect 1175 7814 1188 7844
rect 1203 7830 1233 7844
rect 1276 7830 1319 7844
rect 1326 7830 1546 7844
rect 1553 7830 1583 7844
rect 1243 7816 1258 7828
rect 1277 7816 1290 7830
rect 1358 7826 1511 7830
rect 1240 7814 1262 7816
rect 1340 7814 1532 7826
rect 1611 7814 1624 7844
rect 1639 7830 1669 7844
rect 1706 7814 1725 7844
rect 1740 7814 1746 7844
rect 1755 7814 1768 7844
rect 1783 7830 1813 7844
rect 1856 7830 1899 7844
rect 1906 7830 2126 7844
rect 2133 7830 2163 7844
rect 1823 7816 1838 7828
rect 1857 7816 1870 7830
rect 1938 7826 2091 7830
rect 1820 7814 1842 7816
rect 1920 7814 2112 7826
rect 2191 7814 2204 7844
rect 2219 7830 2249 7844
rect 2286 7814 2305 7844
rect 2320 7814 2326 7844
rect 2335 7814 2348 7844
rect 2363 7830 2393 7844
rect 2436 7830 2479 7844
rect 2486 7830 2706 7844
rect 2713 7830 2743 7844
rect 2403 7816 2418 7828
rect 2437 7816 2450 7830
rect 2518 7826 2671 7830
rect 2400 7814 2422 7816
rect 2500 7814 2692 7826
rect 2771 7814 2784 7844
rect 2799 7830 2829 7844
rect 2866 7814 2885 7844
rect 2900 7814 2906 7844
rect 2915 7814 2928 7844
rect 2943 7830 2973 7844
rect 3016 7830 3059 7844
rect 3066 7830 3286 7844
rect 3293 7830 3323 7844
rect 2983 7816 2998 7828
rect 3017 7816 3030 7830
rect 3098 7826 3251 7830
rect 2980 7814 3002 7816
rect 3080 7814 3272 7826
rect 3351 7814 3364 7844
rect 3379 7830 3409 7844
rect 3446 7814 3465 7844
rect 3480 7814 3486 7844
rect 3495 7814 3508 7844
rect 3523 7830 3553 7844
rect 3596 7830 3639 7844
rect 3646 7830 3866 7844
rect 3873 7830 3903 7844
rect 3563 7816 3578 7828
rect 3597 7816 3610 7830
rect 3678 7826 3831 7830
rect 3560 7814 3582 7816
rect 3660 7814 3852 7826
rect 3931 7814 3944 7844
rect 3959 7830 3989 7844
rect 4026 7814 4045 7844
rect 4060 7814 4066 7844
rect 4075 7814 4088 7844
rect 4103 7830 4133 7844
rect 4176 7830 4219 7844
rect 4226 7830 4446 7844
rect 4453 7830 4483 7844
rect 4143 7816 4158 7828
rect 4177 7816 4190 7830
rect 4258 7826 4411 7830
rect 4140 7814 4162 7816
rect 4240 7814 4432 7826
rect 4511 7814 4524 7844
rect 4539 7830 4569 7844
rect 4606 7814 4625 7844
rect 4640 7814 4646 7844
rect 4655 7814 4668 7844
rect 4683 7830 4713 7844
rect 4756 7830 4799 7844
rect 4806 7830 5026 7844
rect 5033 7830 5063 7844
rect 4723 7816 4738 7828
rect 4757 7816 4770 7830
rect 4838 7826 4991 7830
rect 4720 7814 4742 7816
rect 4820 7814 5012 7826
rect 5091 7814 5104 7844
rect 5119 7830 5149 7844
rect 5186 7814 5205 7844
rect 5220 7814 5226 7844
rect 5235 7814 5248 7844
rect 5263 7830 5293 7844
rect 5336 7830 5379 7844
rect 5386 7830 5606 7844
rect 5613 7830 5643 7844
rect 5303 7816 5318 7828
rect 5337 7816 5350 7830
rect 5418 7826 5571 7830
rect 5300 7814 5322 7816
rect 5400 7814 5592 7826
rect 5671 7814 5684 7844
rect 5699 7830 5729 7844
rect 5766 7814 5785 7844
rect 5800 7814 5806 7844
rect 5815 7814 5828 7844
rect 5843 7830 5873 7844
rect 5916 7830 5959 7844
rect 5966 7830 6186 7844
rect 6193 7830 6223 7844
rect 5883 7816 5898 7828
rect 5917 7816 5930 7830
rect 5998 7826 6151 7830
rect 5880 7814 5902 7816
rect 5980 7814 6172 7826
rect 6251 7814 6264 7844
rect 6279 7830 6309 7844
rect 6346 7814 6365 7844
rect 6380 7814 6386 7844
rect 6395 7814 6408 7844
rect 6423 7830 6453 7844
rect 6496 7830 6539 7844
rect 6546 7830 6766 7844
rect 6773 7830 6803 7844
rect 6463 7816 6478 7828
rect 6497 7816 6510 7830
rect 6578 7826 6731 7830
rect 6460 7814 6482 7816
rect 6560 7814 6752 7826
rect 6831 7814 6844 7844
rect 6859 7830 6889 7844
rect 6926 7814 6945 7844
rect 6960 7814 6966 7844
rect 6975 7814 6988 7844
rect 7003 7830 7033 7844
rect 7076 7830 7119 7844
rect 7126 7830 7346 7844
rect 7353 7830 7383 7844
rect 7043 7816 7058 7828
rect 7077 7816 7090 7830
rect 7158 7826 7311 7830
rect 7040 7814 7062 7816
rect 7140 7814 7332 7826
rect 7411 7814 7424 7844
rect 7439 7830 7469 7844
rect 7506 7814 7525 7844
rect 7540 7814 7546 7844
rect 7555 7814 7568 7844
rect 7583 7830 7613 7844
rect 7656 7830 7699 7844
rect 7706 7830 7926 7844
rect 7933 7830 7963 7844
rect 7623 7816 7638 7828
rect 7657 7816 7670 7830
rect 7738 7826 7891 7830
rect 7620 7814 7642 7816
rect 7720 7814 7912 7826
rect 7991 7814 8004 7844
rect 8019 7830 8049 7844
rect 8086 7814 8105 7844
rect 8120 7814 8126 7844
rect 8135 7814 8148 7844
rect 8163 7830 8193 7844
rect 8236 7830 8279 7844
rect 8286 7830 8506 7844
rect 8513 7830 8543 7844
rect 8203 7816 8218 7828
rect 8237 7816 8250 7830
rect 8318 7826 8471 7830
rect 8200 7814 8222 7816
rect 8300 7814 8492 7826
rect 8571 7814 8584 7844
rect 8599 7830 8629 7844
rect 8666 7814 8685 7844
rect 8700 7814 8706 7844
rect 8715 7814 8728 7844
rect 8743 7830 8773 7844
rect 8816 7830 8859 7844
rect 8866 7830 9086 7844
rect 9093 7830 9123 7844
rect 8783 7816 8798 7828
rect 8817 7816 8830 7830
rect 8898 7826 9051 7830
rect 8780 7814 8802 7816
rect 8880 7814 9072 7826
rect 9151 7814 9164 7844
rect 9179 7830 9209 7844
rect 9246 7814 9265 7844
rect 9280 7814 9286 7844
rect 9295 7814 9308 7844
rect 9323 7830 9353 7844
rect 9396 7830 9439 7844
rect 9446 7830 9666 7844
rect 9673 7830 9703 7844
rect 9363 7816 9378 7828
rect 9397 7816 9410 7830
rect 9478 7826 9631 7830
rect 9360 7814 9382 7816
rect 9460 7814 9652 7826
rect 9731 7814 9744 7844
rect 9759 7830 9789 7844
rect 9826 7814 9845 7844
rect 9860 7814 9866 7844
rect 9875 7814 9888 7844
rect 9903 7830 9933 7844
rect 9976 7830 10019 7844
rect 10026 7830 10246 7844
rect 10253 7830 10283 7844
rect 9943 7816 9958 7828
rect 9977 7816 9990 7830
rect 10058 7826 10211 7830
rect 9940 7814 9962 7816
rect 10040 7814 10232 7826
rect 10311 7814 10324 7844
rect 10339 7830 10369 7844
rect 10406 7814 10425 7844
rect 10440 7814 10446 7844
rect 10455 7814 10468 7844
rect 10483 7830 10513 7844
rect 10556 7830 10599 7844
rect 10606 7830 10826 7844
rect 10833 7830 10863 7844
rect 10523 7816 10538 7828
rect 10557 7816 10570 7830
rect 10638 7826 10791 7830
rect 10520 7814 10542 7816
rect 10620 7814 10812 7826
rect 10891 7814 10904 7844
rect 10919 7830 10949 7844
rect 10986 7814 11005 7844
rect 11020 7814 11026 7844
rect 11035 7814 11048 7844
rect 11063 7830 11093 7844
rect 11136 7830 11179 7844
rect 11186 7830 11406 7844
rect 11413 7830 11443 7844
rect 11103 7816 11118 7828
rect 11137 7816 11150 7830
rect 11218 7826 11371 7830
rect 11100 7814 11122 7816
rect 11200 7814 11392 7826
rect 11471 7814 11484 7844
rect 11499 7830 11529 7844
rect 11566 7814 11585 7844
rect 11600 7814 11606 7844
rect 11615 7814 11628 7844
rect 11643 7830 11673 7844
rect 11716 7830 11759 7844
rect 11766 7830 11986 7844
rect 11993 7830 12023 7844
rect 11683 7816 11698 7828
rect 11717 7816 11730 7830
rect 11798 7826 11951 7830
rect 11680 7814 11702 7816
rect 11780 7814 11972 7826
rect 12051 7814 12064 7844
rect 12079 7830 12109 7844
rect 12146 7814 12165 7844
rect 12180 7814 12186 7844
rect 12195 7814 12208 7844
rect 12223 7830 12253 7844
rect 12296 7830 12339 7844
rect 12346 7830 12566 7844
rect 12573 7830 12603 7844
rect 12263 7816 12278 7828
rect 12297 7816 12310 7830
rect 12378 7826 12531 7830
rect 12260 7814 12282 7816
rect 12360 7814 12552 7826
rect 12631 7814 12644 7844
rect 12659 7830 12689 7844
rect 12726 7814 12745 7844
rect 12760 7814 12766 7844
rect 12775 7814 12788 7844
rect 12803 7830 12833 7844
rect 12876 7830 12919 7844
rect 12926 7830 13146 7844
rect 13153 7830 13183 7844
rect 12843 7816 12858 7828
rect 12877 7816 12890 7830
rect 12958 7826 13111 7830
rect 12840 7814 12862 7816
rect 12940 7814 13132 7826
rect 13211 7814 13224 7844
rect 13239 7830 13269 7844
rect 13306 7814 13325 7844
rect 13340 7814 13346 7844
rect 13355 7814 13368 7844
rect 13383 7830 13413 7844
rect 13456 7830 13499 7844
rect 13506 7830 13726 7844
rect 13733 7830 13763 7844
rect 13423 7816 13438 7828
rect 13457 7816 13470 7830
rect 13538 7826 13691 7830
rect 13420 7814 13442 7816
rect 13520 7814 13712 7826
rect 13791 7814 13804 7844
rect 13819 7830 13849 7844
rect 13886 7814 13905 7844
rect 13920 7814 13926 7844
rect 13935 7814 13948 7844
rect 13963 7830 13993 7844
rect 14036 7830 14079 7844
rect 14086 7830 14306 7844
rect 14313 7830 14343 7844
rect 14003 7816 14018 7828
rect 14037 7816 14050 7830
rect 14118 7826 14271 7830
rect 14000 7814 14022 7816
rect 14100 7814 14292 7826
rect 14371 7814 14384 7844
rect 14399 7830 14429 7844
rect 14466 7814 14485 7844
rect 14500 7814 14506 7844
rect 14515 7814 14528 7844
rect 14543 7830 14573 7844
rect 14616 7830 14659 7844
rect 14666 7830 14886 7844
rect 14893 7830 14923 7844
rect 14583 7816 14598 7828
rect 14617 7816 14630 7830
rect 14698 7826 14851 7830
rect 14580 7814 14602 7816
rect 14680 7814 14872 7826
rect 14951 7814 14964 7844
rect 14979 7830 15009 7844
rect 15046 7814 15065 7844
rect 15080 7814 15086 7844
rect 15095 7814 15108 7844
rect 15123 7830 15153 7844
rect 15196 7830 15239 7844
rect 15246 7830 15466 7844
rect 15473 7830 15503 7844
rect 15163 7816 15178 7828
rect 15197 7816 15210 7830
rect 15278 7826 15431 7830
rect 15160 7814 15182 7816
rect 15260 7814 15452 7826
rect 15531 7814 15544 7844
rect 15559 7830 15589 7844
rect 15626 7814 15645 7844
rect 15660 7814 15666 7844
rect 15675 7814 15688 7844
rect 15703 7830 15733 7844
rect 15776 7830 15819 7844
rect 15826 7830 16046 7844
rect 16053 7830 16083 7844
rect 15743 7816 15758 7828
rect 15777 7816 15790 7830
rect 15858 7826 16011 7830
rect 15740 7814 15762 7816
rect 15840 7814 16032 7826
rect 16111 7814 16124 7844
rect 16139 7830 16169 7844
rect 16206 7814 16225 7844
rect 16240 7814 16246 7844
rect 16255 7814 16268 7844
rect 16283 7830 16313 7844
rect 16356 7830 16399 7844
rect 16406 7830 16626 7844
rect 16633 7830 16663 7844
rect 16323 7816 16338 7828
rect 16357 7816 16370 7830
rect 16438 7826 16591 7830
rect 16320 7814 16342 7816
rect 16420 7814 16612 7826
rect 16691 7814 16704 7844
rect 16719 7830 16749 7844
rect 16786 7814 16805 7844
rect 16820 7814 16826 7844
rect 16835 7814 16848 7844
rect 16863 7830 16893 7844
rect 16936 7830 16979 7844
rect 16986 7830 17206 7844
rect 17213 7830 17243 7844
rect 16903 7816 16918 7828
rect 16937 7816 16950 7830
rect 17018 7826 17171 7830
rect 16900 7814 16922 7816
rect 17000 7814 17192 7826
rect 17271 7814 17284 7844
rect 17299 7830 17329 7844
rect 17366 7814 17385 7844
rect 17400 7814 17406 7844
rect 17415 7814 17428 7844
rect 17443 7830 17473 7844
rect 17516 7830 17559 7844
rect 17566 7830 17786 7844
rect 17793 7830 17823 7844
rect 17483 7816 17498 7828
rect 17517 7816 17530 7830
rect 17598 7826 17751 7830
rect 17480 7814 17502 7816
rect 17580 7814 17772 7826
rect 17851 7814 17864 7844
rect 17879 7830 17909 7844
rect 17946 7814 17965 7844
rect 17980 7814 17986 7844
rect 17995 7814 18008 7844
rect 18023 7830 18053 7844
rect 18096 7830 18139 7844
rect 18146 7830 18366 7844
rect 18373 7830 18403 7844
rect 18063 7816 18078 7828
rect 18097 7816 18110 7830
rect 18178 7826 18331 7830
rect 18060 7814 18082 7816
rect 18160 7814 18352 7826
rect 18431 7814 18444 7844
rect 18459 7830 18489 7844
rect 18532 7814 18545 7844
rect 0 7800 18545 7814
rect 15 7730 28 7800
rect 80 7796 102 7800
rect 73 7774 102 7788
rect 155 7774 171 7788
rect 209 7784 215 7786
rect 222 7784 330 7800
rect 337 7784 343 7786
rect 351 7784 366 7800
rect 432 7794 451 7797
rect 73 7772 171 7774
rect 198 7772 366 7784
rect 381 7774 397 7788
rect 432 7775 454 7794
rect 464 7788 480 7789
rect 463 7786 480 7788
rect 464 7781 480 7786
rect 454 7774 460 7775
rect 463 7774 492 7781
rect 381 7773 492 7774
rect 381 7772 498 7773
rect 57 7764 108 7772
rect 155 7764 189 7772
rect 57 7752 82 7764
rect 89 7752 108 7764
rect 162 7762 189 7764
rect 198 7762 419 7772
rect 454 7769 460 7772
rect 162 7758 419 7762
rect 57 7744 108 7752
rect 155 7744 419 7758
rect 463 7764 498 7772
rect 9 7696 28 7730
rect 73 7736 102 7744
rect 73 7730 90 7736
rect 73 7728 107 7730
rect 155 7728 171 7744
rect 172 7734 380 7744
rect 381 7734 397 7744
rect 445 7740 460 7755
rect 463 7752 464 7764
rect 471 7752 498 7764
rect 463 7744 498 7752
rect 463 7743 492 7744
rect 183 7730 397 7734
rect 198 7728 397 7730
rect 432 7730 445 7740
rect 463 7730 480 7743
rect 432 7728 480 7730
rect 74 7724 107 7728
rect 70 7722 107 7724
rect 70 7721 137 7722
rect 70 7716 101 7721
rect 107 7716 137 7721
rect 70 7712 137 7716
rect 43 7709 137 7712
rect 43 7702 92 7709
rect 43 7696 73 7702
rect 92 7697 97 7702
rect 9 7680 89 7696
rect 101 7688 137 7709
rect 198 7704 387 7728
rect 432 7727 479 7728
rect 445 7722 479 7727
rect 213 7701 387 7704
rect 206 7698 387 7701
rect 415 7721 479 7722
rect 9 7678 28 7680
rect 43 7678 77 7680
rect 9 7662 89 7678
rect 9 7656 28 7662
rect -1 7640 28 7656
rect 43 7646 73 7662
rect 101 7640 107 7688
rect 110 7682 129 7688
rect 144 7682 174 7690
rect 110 7674 174 7682
rect 110 7658 190 7674
rect 206 7667 268 7698
rect 284 7667 346 7698
rect 415 7696 464 7721
rect 479 7696 509 7712
rect 378 7682 408 7690
rect 415 7688 525 7696
rect 378 7674 423 7682
rect 110 7656 129 7658
rect 144 7656 190 7658
rect 110 7640 190 7656
rect 217 7654 252 7667
rect 293 7664 330 7667
rect 293 7662 335 7664
rect 222 7651 252 7654
rect 231 7647 238 7651
rect 238 7646 239 7647
rect 197 7640 207 7646
rect -7 7632 34 7640
rect -7 7606 8 7632
rect 15 7606 34 7632
rect 98 7628 129 7640
rect 144 7628 247 7640
rect 259 7630 285 7656
rect 300 7651 330 7662
rect 362 7658 424 7674
rect 362 7656 408 7658
rect 362 7640 424 7656
rect 436 7640 442 7688
rect 445 7680 525 7688
rect 445 7678 464 7680
rect 479 7678 513 7680
rect 445 7662 525 7678
rect 445 7640 464 7662
rect 479 7646 509 7662
rect 537 7656 543 7730
rect 546 7656 565 7800
rect 580 7656 586 7800
rect 595 7730 608 7800
rect 660 7796 682 7800
rect 653 7774 682 7788
rect 735 7774 751 7788
rect 789 7784 795 7786
rect 802 7784 910 7800
rect 917 7784 923 7786
rect 931 7784 946 7800
rect 1012 7794 1031 7797
rect 653 7772 751 7774
rect 778 7772 946 7784
rect 961 7774 977 7788
rect 1012 7775 1034 7794
rect 1044 7788 1060 7789
rect 1043 7786 1060 7788
rect 1044 7781 1060 7786
rect 1034 7774 1040 7775
rect 1043 7774 1072 7781
rect 961 7773 1072 7774
rect 961 7772 1078 7773
rect 637 7764 688 7772
rect 735 7764 769 7772
rect 637 7752 662 7764
rect 669 7752 688 7764
rect 742 7762 769 7764
rect 778 7762 999 7772
rect 1034 7769 1040 7772
rect 742 7758 999 7762
rect 637 7744 688 7752
rect 735 7744 999 7758
rect 1043 7764 1078 7772
rect 589 7696 608 7730
rect 653 7736 682 7744
rect 653 7730 670 7736
rect 653 7728 687 7730
rect 735 7728 751 7744
rect 752 7734 960 7744
rect 961 7734 977 7744
rect 1025 7740 1040 7755
rect 1043 7752 1044 7764
rect 1051 7752 1078 7764
rect 1043 7744 1078 7752
rect 1043 7743 1072 7744
rect 763 7730 977 7734
rect 778 7728 977 7730
rect 1012 7730 1025 7740
rect 1043 7730 1060 7743
rect 1012 7728 1060 7730
rect 654 7724 687 7728
rect 650 7722 687 7724
rect 650 7721 717 7722
rect 650 7716 681 7721
rect 687 7716 717 7721
rect 650 7712 717 7716
rect 623 7709 717 7712
rect 623 7702 672 7709
rect 623 7696 653 7702
rect 672 7697 677 7702
rect 589 7680 669 7696
rect 681 7688 717 7709
rect 778 7704 967 7728
rect 1012 7727 1059 7728
rect 1025 7722 1059 7727
rect 793 7701 967 7704
rect 786 7698 967 7701
rect 995 7721 1059 7722
rect 589 7678 608 7680
rect 623 7678 657 7680
rect 589 7662 669 7678
rect 589 7656 608 7662
rect 305 7630 408 7640
rect 259 7628 408 7630
rect 429 7628 464 7640
rect 98 7626 260 7628
rect 110 7606 129 7626
rect 144 7624 174 7626
rect -7 7598 34 7606
rect 116 7602 129 7606
rect 181 7610 260 7626
rect 292 7626 464 7628
rect 292 7610 371 7626
rect 378 7624 408 7626
rect -1 7588 28 7598
rect 43 7588 73 7602
rect 116 7588 159 7602
rect 181 7598 371 7610
rect 436 7606 442 7626
rect 166 7588 196 7598
rect 197 7588 355 7598
rect 359 7588 389 7598
rect 393 7588 423 7602
rect 451 7588 464 7626
rect 536 7640 565 7656
rect 579 7640 608 7656
rect 623 7646 653 7662
rect 681 7640 687 7688
rect 690 7682 709 7688
rect 724 7682 754 7690
rect 690 7674 754 7682
rect 690 7658 770 7674
rect 786 7667 848 7698
rect 864 7667 926 7698
rect 995 7696 1044 7721
rect 1059 7696 1089 7712
rect 958 7682 988 7690
rect 995 7688 1105 7696
rect 958 7674 1003 7682
rect 690 7656 709 7658
rect 724 7656 770 7658
rect 690 7640 770 7656
rect 797 7654 832 7667
rect 873 7664 910 7667
rect 873 7662 915 7664
rect 802 7651 832 7654
rect 811 7647 818 7651
rect 818 7646 819 7647
rect 777 7640 787 7646
rect 536 7632 571 7640
rect 536 7606 537 7632
rect 544 7606 571 7632
rect 479 7588 509 7602
rect 536 7598 571 7606
rect 573 7632 614 7640
rect 573 7606 588 7632
rect 595 7606 614 7632
rect 678 7628 709 7640
rect 724 7628 827 7640
rect 839 7630 865 7656
rect 880 7651 910 7662
rect 942 7658 1004 7674
rect 942 7656 988 7658
rect 942 7640 1004 7656
rect 1016 7640 1022 7688
rect 1025 7680 1105 7688
rect 1025 7678 1044 7680
rect 1059 7678 1093 7680
rect 1025 7662 1105 7678
rect 1025 7640 1044 7662
rect 1059 7646 1089 7662
rect 1117 7656 1123 7730
rect 1126 7656 1145 7800
rect 1160 7656 1166 7800
rect 1175 7730 1188 7800
rect 1240 7796 1262 7800
rect 1233 7774 1262 7788
rect 1315 7774 1331 7788
rect 1369 7784 1375 7786
rect 1382 7784 1490 7800
rect 1497 7784 1503 7786
rect 1511 7784 1526 7800
rect 1592 7794 1611 7797
rect 1233 7772 1331 7774
rect 1358 7772 1526 7784
rect 1541 7774 1557 7788
rect 1592 7775 1614 7794
rect 1624 7788 1640 7789
rect 1623 7786 1640 7788
rect 1624 7781 1640 7786
rect 1614 7774 1620 7775
rect 1623 7774 1652 7781
rect 1541 7773 1652 7774
rect 1541 7772 1658 7773
rect 1217 7764 1268 7772
rect 1315 7764 1349 7772
rect 1217 7752 1242 7764
rect 1249 7752 1268 7764
rect 1322 7762 1349 7764
rect 1358 7762 1579 7772
rect 1614 7769 1620 7772
rect 1322 7758 1579 7762
rect 1217 7744 1268 7752
rect 1315 7744 1579 7758
rect 1623 7764 1658 7772
rect 1169 7696 1188 7730
rect 1233 7736 1262 7744
rect 1233 7730 1250 7736
rect 1233 7728 1267 7730
rect 1315 7728 1331 7744
rect 1332 7734 1540 7744
rect 1541 7734 1557 7744
rect 1605 7740 1620 7755
rect 1623 7752 1624 7764
rect 1631 7752 1658 7764
rect 1623 7744 1658 7752
rect 1623 7743 1652 7744
rect 1343 7730 1557 7734
rect 1358 7728 1557 7730
rect 1592 7730 1605 7740
rect 1623 7730 1640 7743
rect 1592 7728 1640 7730
rect 1234 7724 1267 7728
rect 1230 7722 1267 7724
rect 1230 7721 1297 7722
rect 1230 7716 1261 7721
rect 1267 7716 1297 7721
rect 1230 7712 1297 7716
rect 1203 7709 1297 7712
rect 1203 7702 1252 7709
rect 1203 7696 1233 7702
rect 1252 7697 1257 7702
rect 1169 7680 1249 7696
rect 1261 7688 1297 7709
rect 1358 7704 1547 7728
rect 1592 7727 1639 7728
rect 1605 7722 1639 7727
rect 1373 7701 1547 7704
rect 1366 7698 1547 7701
rect 1575 7721 1639 7722
rect 1169 7678 1188 7680
rect 1203 7678 1237 7680
rect 1169 7662 1249 7678
rect 1169 7656 1188 7662
rect 885 7630 988 7640
rect 839 7628 988 7630
rect 1009 7628 1044 7640
rect 678 7626 840 7628
rect 690 7606 709 7626
rect 724 7624 754 7626
rect 573 7598 614 7606
rect 696 7602 709 7606
rect 761 7610 840 7626
rect 872 7626 1044 7628
rect 872 7610 951 7626
rect 958 7624 988 7626
rect 536 7588 565 7598
rect 579 7588 608 7598
rect 623 7588 653 7602
rect 696 7588 739 7602
rect 761 7598 951 7610
rect 1016 7606 1022 7626
rect 746 7588 776 7598
rect 777 7588 935 7598
rect 939 7588 969 7598
rect 973 7588 1003 7602
rect 1031 7588 1044 7626
rect 1116 7640 1145 7656
rect 1159 7640 1188 7656
rect 1203 7646 1233 7662
rect 1261 7640 1267 7688
rect 1270 7682 1289 7688
rect 1304 7682 1334 7690
rect 1270 7674 1334 7682
rect 1270 7658 1350 7674
rect 1366 7667 1428 7698
rect 1444 7667 1506 7698
rect 1575 7696 1624 7721
rect 1639 7696 1669 7712
rect 1538 7682 1568 7690
rect 1575 7688 1685 7696
rect 1538 7674 1583 7682
rect 1270 7656 1289 7658
rect 1304 7656 1350 7658
rect 1270 7640 1350 7656
rect 1377 7654 1412 7667
rect 1453 7664 1490 7667
rect 1453 7662 1495 7664
rect 1382 7651 1412 7654
rect 1391 7647 1398 7651
rect 1398 7646 1399 7647
rect 1357 7640 1367 7646
rect 1116 7632 1151 7640
rect 1116 7606 1117 7632
rect 1124 7606 1151 7632
rect 1059 7588 1089 7602
rect 1116 7598 1151 7606
rect 1153 7632 1194 7640
rect 1153 7606 1168 7632
rect 1175 7606 1194 7632
rect 1258 7628 1289 7640
rect 1304 7628 1407 7640
rect 1419 7630 1445 7656
rect 1460 7651 1490 7662
rect 1522 7658 1584 7674
rect 1522 7656 1568 7658
rect 1522 7640 1584 7656
rect 1596 7640 1602 7688
rect 1605 7680 1685 7688
rect 1605 7678 1624 7680
rect 1639 7678 1673 7680
rect 1605 7662 1685 7678
rect 1605 7640 1624 7662
rect 1639 7646 1669 7662
rect 1697 7656 1703 7730
rect 1706 7656 1725 7800
rect 1740 7656 1746 7800
rect 1755 7730 1768 7800
rect 1820 7796 1842 7800
rect 1813 7774 1842 7788
rect 1895 7774 1911 7788
rect 1949 7784 1955 7786
rect 1962 7784 2070 7800
rect 2077 7784 2083 7786
rect 2091 7784 2106 7800
rect 2172 7794 2191 7797
rect 1813 7772 1911 7774
rect 1938 7772 2106 7784
rect 2121 7774 2137 7788
rect 2172 7775 2194 7794
rect 2204 7788 2220 7789
rect 2203 7786 2220 7788
rect 2204 7781 2220 7786
rect 2194 7774 2200 7775
rect 2203 7774 2232 7781
rect 2121 7773 2232 7774
rect 2121 7772 2238 7773
rect 1797 7764 1848 7772
rect 1895 7764 1929 7772
rect 1797 7752 1822 7764
rect 1829 7752 1848 7764
rect 1902 7762 1929 7764
rect 1938 7762 2159 7772
rect 2194 7769 2200 7772
rect 1902 7758 2159 7762
rect 1797 7744 1848 7752
rect 1895 7744 2159 7758
rect 2203 7764 2238 7772
rect 1749 7696 1768 7730
rect 1813 7736 1842 7744
rect 1813 7730 1830 7736
rect 1813 7728 1847 7730
rect 1895 7728 1911 7744
rect 1912 7734 2120 7744
rect 2121 7734 2137 7744
rect 2185 7740 2200 7755
rect 2203 7752 2204 7764
rect 2211 7752 2238 7764
rect 2203 7744 2238 7752
rect 2203 7743 2232 7744
rect 1923 7730 2137 7734
rect 1938 7728 2137 7730
rect 2172 7730 2185 7740
rect 2203 7730 2220 7743
rect 2172 7728 2220 7730
rect 1814 7724 1847 7728
rect 1810 7722 1847 7724
rect 1810 7721 1877 7722
rect 1810 7716 1841 7721
rect 1847 7716 1877 7721
rect 1810 7712 1877 7716
rect 1783 7709 1877 7712
rect 1783 7702 1832 7709
rect 1783 7696 1813 7702
rect 1832 7697 1837 7702
rect 1749 7680 1829 7696
rect 1841 7688 1877 7709
rect 1938 7704 2127 7728
rect 2172 7727 2219 7728
rect 2185 7722 2219 7727
rect 1953 7701 2127 7704
rect 1946 7698 2127 7701
rect 2155 7721 2219 7722
rect 1749 7678 1768 7680
rect 1783 7678 1817 7680
rect 1749 7662 1829 7678
rect 1749 7656 1768 7662
rect 1465 7630 1568 7640
rect 1419 7628 1568 7630
rect 1589 7628 1624 7640
rect 1258 7626 1420 7628
rect 1270 7606 1289 7626
rect 1304 7624 1334 7626
rect 1153 7598 1194 7606
rect 1276 7602 1289 7606
rect 1341 7610 1420 7626
rect 1452 7626 1624 7628
rect 1452 7610 1531 7626
rect 1538 7624 1568 7626
rect 1116 7588 1145 7598
rect 1159 7588 1188 7598
rect 1203 7588 1233 7602
rect 1276 7588 1319 7602
rect 1341 7598 1531 7610
rect 1596 7606 1602 7626
rect 1326 7588 1356 7598
rect 1357 7588 1515 7598
rect 1519 7588 1549 7598
rect 1553 7588 1583 7602
rect 1611 7588 1624 7626
rect 1696 7640 1725 7656
rect 1739 7640 1768 7656
rect 1783 7646 1813 7662
rect 1841 7640 1847 7688
rect 1850 7682 1869 7688
rect 1884 7682 1914 7690
rect 1850 7674 1914 7682
rect 1850 7658 1930 7674
rect 1946 7667 2008 7698
rect 2024 7667 2086 7698
rect 2155 7696 2204 7721
rect 2219 7696 2249 7712
rect 2118 7682 2148 7690
rect 2155 7688 2265 7696
rect 2118 7674 2163 7682
rect 1850 7656 1869 7658
rect 1884 7656 1930 7658
rect 1850 7640 1930 7656
rect 1957 7654 1992 7667
rect 2033 7664 2070 7667
rect 2033 7662 2075 7664
rect 1962 7651 1992 7654
rect 1971 7647 1978 7651
rect 1978 7646 1979 7647
rect 1937 7640 1947 7646
rect 1696 7632 1731 7640
rect 1696 7606 1697 7632
rect 1704 7606 1731 7632
rect 1639 7588 1669 7602
rect 1696 7598 1731 7606
rect 1733 7632 1774 7640
rect 1733 7606 1748 7632
rect 1755 7606 1774 7632
rect 1838 7628 1869 7640
rect 1884 7628 1987 7640
rect 1999 7630 2025 7656
rect 2040 7651 2070 7662
rect 2102 7658 2164 7674
rect 2102 7656 2148 7658
rect 2102 7640 2164 7656
rect 2176 7640 2182 7688
rect 2185 7680 2265 7688
rect 2185 7678 2204 7680
rect 2219 7678 2253 7680
rect 2185 7662 2265 7678
rect 2185 7640 2204 7662
rect 2219 7646 2249 7662
rect 2277 7656 2283 7730
rect 2286 7656 2305 7800
rect 2320 7656 2326 7800
rect 2335 7730 2348 7800
rect 2400 7796 2422 7800
rect 2393 7774 2422 7788
rect 2475 7774 2491 7788
rect 2529 7784 2535 7786
rect 2542 7784 2650 7800
rect 2657 7784 2663 7786
rect 2671 7784 2686 7800
rect 2752 7794 2771 7797
rect 2393 7772 2491 7774
rect 2518 7772 2686 7784
rect 2701 7774 2717 7788
rect 2752 7775 2774 7794
rect 2784 7788 2800 7789
rect 2783 7786 2800 7788
rect 2784 7781 2800 7786
rect 2774 7774 2780 7775
rect 2783 7774 2812 7781
rect 2701 7773 2812 7774
rect 2701 7772 2818 7773
rect 2377 7764 2428 7772
rect 2475 7764 2509 7772
rect 2377 7752 2402 7764
rect 2409 7752 2428 7764
rect 2482 7762 2509 7764
rect 2518 7762 2739 7772
rect 2774 7769 2780 7772
rect 2482 7758 2739 7762
rect 2377 7744 2428 7752
rect 2475 7744 2739 7758
rect 2783 7764 2818 7772
rect 2329 7696 2348 7730
rect 2393 7736 2422 7744
rect 2393 7730 2410 7736
rect 2393 7728 2427 7730
rect 2475 7728 2491 7744
rect 2492 7734 2700 7744
rect 2701 7734 2717 7744
rect 2765 7740 2780 7755
rect 2783 7752 2784 7764
rect 2791 7752 2818 7764
rect 2783 7744 2818 7752
rect 2783 7743 2812 7744
rect 2503 7730 2717 7734
rect 2518 7728 2717 7730
rect 2752 7730 2765 7740
rect 2783 7730 2800 7743
rect 2752 7728 2800 7730
rect 2394 7724 2427 7728
rect 2390 7722 2427 7724
rect 2390 7721 2457 7722
rect 2390 7716 2421 7721
rect 2427 7716 2457 7721
rect 2390 7712 2457 7716
rect 2363 7709 2457 7712
rect 2363 7702 2412 7709
rect 2363 7696 2393 7702
rect 2412 7697 2417 7702
rect 2329 7680 2409 7696
rect 2421 7688 2457 7709
rect 2518 7704 2707 7728
rect 2752 7727 2799 7728
rect 2765 7722 2799 7727
rect 2533 7701 2707 7704
rect 2526 7698 2707 7701
rect 2735 7721 2799 7722
rect 2329 7678 2348 7680
rect 2363 7678 2397 7680
rect 2329 7662 2409 7678
rect 2329 7656 2348 7662
rect 2045 7630 2148 7640
rect 1999 7628 2148 7630
rect 2169 7628 2204 7640
rect 1838 7626 2000 7628
rect 1850 7606 1869 7626
rect 1884 7624 1914 7626
rect 1733 7598 1774 7606
rect 1856 7602 1869 7606
rect 1921 7610 2000 7626
rect 2032 7626 2204 7628
rect 2032 7610 2111 7626
rect 2118 7624 2148 7626
rect 1696 7588 1725 7598
rect 1739 7588 1768 7598
rect 1783 7588 1813 7602
rect 1856 7588 1899 7602
rect 1921 7598 2111 7610
rect 2176 7606 2182 7626
rect 1906 7588 1936 7598
rect 1937 7588 2095 7598
rect 2099 7588 2129 7598
rect 2133 7588 2163 7602
rect 2191 7588 2204 7626
rect 2276 7640 2305 7656
rect 2319 7640 2348 7656
rect 2363 7646 2393 7662
rect 2421 7640 2427 7688
rect 2430 7682 2449 7688
rect 2464 7682 2494 7690
rect 2430 7674 2494 7682
rect 2430 7658 2510 7674
rect 2526 7667 2588 7698
rect 2604 7667 2666 7698
rect 2735 7696 2784 7721
rect 2799 7696 2829 7712
rect 2698 7682 2728 7690
rect 2735 7688 2845 7696
rect 2698 7674 2743 7682
rect 2430 7656 2449 7658
rect 2464 7656 2510 7658
rect 2430 7640 2510 7656
rect 2537 7654 2572 7667
rect 2613 7664 2650 7667
rect 2613 7662 2655 7664
rect 2542 7651 2572 7654
rect 2551 7647 2558 7651
rect 2558 7646 2559 7647
rect 2517 7640 2527 7646
rect 2276 7632 2311 7640
rect 2276 7606 2277 7632
rect 2284 7606 2311 7632
rect 2219 7588 2249 7602
rect 2276 7598 2311 7606
rect 2313 7632 2354 7640
rect 2313 7606 2328 7632
rect 2335 7606 2354 7632
rect 2418 7628 2449 7640
rect 2464 7628 2567 7640
rect 2579 7630 2605 7656
rect 2620 7651 2650 7662
rect 2682 7658 2744 7674
rect 2682 7656 2728 7658
rect 2682 7640 2744 7656
rect 2756 7640 2762 7688
rect 2765 7680 2845 7688
rect 2765 7678 2784 7680
rect 2799 7678 2833 7680
rect 2765 7662 2845 7678
rect 2765 7640 2784 7662
rect 2799 7646 2829 7662
rect 2857 7656 2863 7730
rect 2866 7656 2885 7800
rect 2900 7656 2906 7800
rect 2915 7730 2928 7800
rect 2980 7796 3002 7800
rect 2973 7774 3002 7788
rect 3055 7774 3071 7788
rect 3109 7784 3115 7786
rect 3122 7784 3230 7800
rect 3237 7784 3243 7786
rect 3251 7784 3266 7800
rect 3332 7794 3351 7797
rect 2973 7772 3071 7774
rect 3098 7772 3266 7784
rect 3281 7774 3297 7788
rect 3332 7775 3354 7794
rect 3364 7788 3380 7789
rect 3363 7786 3380 7788
rect 3364 7781 3380 7786
rect 3354 7774 3360 7775
rect 3363 7774 3392 7781
rect 3281 7773 3392 7774
rect 3281 7772 3398 7773
rect 2957 7764 3008 7772
rect 3055 7764 3089 7772
rect 2957 7752 2982 7764
rect 2989 7752 3008 7764
rect 3062 7762 3089 7764
rect 3098 7762 3319 7772
rect 3354 7769 3360 7772
rect 3062 7758 3319 7762
rect 2957 7744 3008 7752
rect 3055 7744 3319 7758
rect 3363 7764 3398 7772
rect 2909 7696 2928 7730
rect 2973 7736 3002 7744
rect 2973 7730 2990 7736
rect 2973 7728 3007 7730
rect 3055 7728 3071 7744
rect 3072 7734 3280 7744
rect 3281 7734 3297 7744
rect 3345 7740 3360 7755
rect 3363 7752 3364 7764
rect 3371 7752 3398 7764
rect 3363 7744 3398 7752
rect 3363 7743 3392 7744
rect 3083 7730 3297 7734
rect 3098 7728 3297 7730
rect 3332 7730 3345 7740
rect 3363 7730 3380 7743
rect 3332 7728 3380 7730
rect 2974 7724 3007 7728
rect 2970 7722 3007 7724
rect 2970 7721 3037 7722
rect 2970 7716 3001 7721
rect 3007 7716 3037 7721
rect 2970 7712 3037 7716
rect 2943 7709 3037 7712
rect 2943 7702 2992 7709
rect 2943 7696 2973 7702
rect 2992 7697 2997 7702
rect 2909 7680 2989 7696
rect 3001 7688 3037 7709
rect 3098 7704 3287 7728
rect 3332 7727 3379 7728
rect 3345 7722 3379 7727
rect 3113 7701 3287 7704
rect 3106 7698 3287 7701
rect 3315 7721 3379 7722
rect 2909 7678 2928 7680
rect 2943 7678 2977 7680
rect 2909 7662 2989 7678
rect 2909 7656 2928 7662
rect 2625 7630 2728 7640
rect 2579 7628 2728 7630
rect 2749 7628 2784 7640
rect 2418 7626 2580 7628
rect 2430 7606 2449 7626
rect 2464 7624 2494 7626
rect 2313 7598 2354 7606
rect 2436 7602 2449 7606
rect 2501 7610 2580 7626
rect 2612 7626 2784 7628
rect 2612 7610 2691 7626
rect 2698 7624 2728 7626
rect 2276 7588 2305 7598
rect 2319 7588 2348 7598
rect 2363 7588 2393 7602
rect 2436 7588 2479 7602
rect 2501 7598 2691 7610
rect 2756 7606 2762 7626
rect 2486 7588 2516 7598
rect 2517 7588 2675 7598
rect 2679 7588 2709 7598
rect 2713 7588 2743 7602
rect 2771 7588 2784 7626
rect 2856 7640 2885 7656
rect 2899 7640 2928 7656
rect 2943 7646 2973 7662
rect 3001 7640 3007 7688
rect 3010 7682 3029 7688
rect 3044 7682 3074 7690
rect 3010 7674 3074 7682
rect 3010 7658 3090 7674
rect 3106 7667 3168 7698
rect 3184 7667 3246 7698
rect 3315 7696 3364 7721
rect 3379 7696 3409 7712
rect 3278 7682 3308 7690
rect 3315 7688 3425 7696
rect 3278 7674 3323 7682
rect 3010 7656 3029 7658
rect 3044 7656 3090 7658
rect 3010 7640 3090 7656
rect 3117 7654 3152 7667
rect 3193 7664 3230 7667
rect 3193 7662 3235 7664
rect 3122 7651 3152 7654
rect 3131 7647 3138 7651
rect 3138 7646 3139 7647
rect 3097 7640 3107 7646
rect 2856 7632 2891 7640
rect 2856 7606 2857 7632
rect 2864 7606 2891 7632
rect 2799 7588 2829 7602
rect 2856 7598 2891 7606
rect 2893 7632 2934 7640
rect 2893 7606 2908 7632
rect 2915 7606 2934 7632
rect 2998 7628 3029 7640
rect 3044 7628 3147 7640
rect 3159 7630 3185 7656
rect 3200 7651 3230 7662
rect 3262 7658 3324 7674
rect 3262 7656 3308 7658
rect 3262 7640 3324 7656
rect 3336 7640 3342 7688
rect 3345 7680 3425 7688
rect 3345 7678 3364 7680
rect 3379 7678 3413 7680
rect 3345 7662 3425 7678
rect 3345 7640 3364 7662
rect 3379 7646 3409 7662
rect 3437 7656 3443 7730
rect 3446 7656 3465 7800
rect 3480 7656 3486 7800
rect 3495 7730 3508 7800
rect 3560 7796 3582 7800
rect 3553 7774 3582 7788
rect 3635 7774 3651 7788
rect 3689 7784 3695 7786
rect 3702 7784 3810 7800
rect 3817 7784 3823 7786
rect 3831 7784 3846 7800
rect 3912 7794 3931 7797
rect 3553 7772 3651 7774
rect 3678 7772 3846 7784
rect 3861 7774 3877 7788
rect 3912 7775 3934 7794
rect 3944 7788 3960 7789
rect 3943 7786 3960 7788
rect 3944 7781 3960 7786
rect 3934 7774 3940 7775
rect 3943 7774 3972 7781
rect 3861 7773 3972 7774
rect 3861 7772 3978 7773
rect 3537 7764 3588 7772
rect 3635 7764 3669 7772
rect 3537 7752 3562 7764
rect 3569 7752 3588 7764
rect 3642 7762 3669 7764
rect 3678 7762 3899 7772
rect 3934 7769 3940 7772
rect 3642 7758 3899 7762
rect 3537 7744 3588 7752
rect 3635 7744 3899 7758
rect 3943 7764 3978 7772
rect 3489 7696 3508 7730
rect 3553 7736 3582 7744
rect 3553 7730 3570 7736
rect 3553 7728 3587 7730
rect 3635 7728 3651 7744
rect 3652 7734 3860 7744
rect 3861 7734 3877 7744
rect 3925 7740 3940 7755
rect 3943 7752 3944 7764
rect 3951 7752 3978 7764
rect 3943 7744 3978 7752
rect 3943 7743 3972 7744
rect 3663 7730 3877 7734
rect 3678 7728 3877 7730
rect 3912 7730 3925 7740
rect 3943 7730 3960 7743
rect 3912 7728 3960 7730
rect 3554 7724 3587 7728
rect 3550 7722 3587 7724
rect 3550 7721 3617 7722
rect 3550 7716 3581 7721
rect 3587 7716 3617 7721
rect 3550 7712 3617 7716
rect 3523 7709 3617 7712
rect 3523 7702 3572 7709
rect 3523 7696 3553 7702
rect 3572 7697 3577 7702
rect 3489 7680 3569 7696
rect 3581 7688 3617 7709
rect 3678 7704 3867 7728
rect 3912 7727 3959 7728
rect 3925 7722 3959 7727
rect 3693 7701 3867 7704
rect 3686 7698 3867 7701
rect 3895 7721 3959 7722
rect 3489 7678 3508 7680
rect 3523 7678 3557 7680
rect 3489 7662 3569 7678
rect 3489 7656 3508 7662
rect 3205 7630 3308 7640
rect 3159 7628 3308 7630
rect 3329 7628 3364 7640
rect 2998 7626 3160 7628
rect 3010 7606 3029 7626
rect 3044 7624 3074 7626
rect 2893 7598 2934 7606
rect 3016 7602 3029 7606
rect 3081 7610 3160 7626
rect 3192 7626 3364 7628
rect 3192 7610 3271 7626
rect 3278 7624 3308 7626
rect 2856 7588 2885 7598
rect 2899 7588 2928 7598
rect 2943 7588 2973 7602
rect 3016 7588 3059 7602
rect 3081 7598 3271 7610
rect 3336 7606 3342 7626
rect 3066 7588 3096 7598
rect 3097 7588 3255 7598
rect 3259 7588 3289 7598
rect 3293 7588 3323 7602
rect 3351 7588 3364 7626
rect 3436 7640 3465 7656
rect 3479 7640 3508 7656
rect 3523 7646 3553 7662
rect 3581 7640 3587 7688
rect 3590 7682 3609 7688
rect 3624 7682 3654 7690
rect 3590 7674 3654 7682
rect 3590 7658 3670 7674
rect 3686 7667 3748 7698
rect 3764 7667 3826 7698
rect 3895 7696 3944 7721
rect 3959 7696 3989 7712
rect 3858 7682 3888 7690
rect 3895 7688 4005 7696
rect 3858 7674 3903 7682
rect 3590 7656 3609 7658
rect 3624 7656 3670 7658
rect 3590 7640 3670 7656
rect 3697 7654 3732 7667
rect 3773 7664 3810 7667
rect 3773 7662 3815 7664
rect 3702 7651 3732 7654
rect 3711 7647 3718 7651
rect 3718 7646 3719 7647
rect 3677 7640 3687 7646
rect 3436 7632 3471 7640
rect 3436 7606 3437 7632
rect 3444 7606 3471 7632
rect 3379 7588 3409 7602
rect 3436 7598 3471 7606
rect 3473 7632 3514 7640
rect 3473 7606 3488 7632
rect 3495 7606 3514 7632
rect 3578 7628 3609 7640
rect 3624 7628 3727 7640
rect 3739 7630 3765 7656
rect 3780 7651 3810 7662
rect 3842 7658 3904 7674
rect 3842 7656 3888 7658
rect 3842 7640 3904 7656
rect 3916 7640 3922 7688
rect 3925 7680 4005 7688
rect 3925 7678 3944 7680
rect 3959 7678 3993 7680
rect 3925 7662 4005 7678
rect 3925 7640 3944 7662
rect 3959 7646 3989 7662
rect 4017 7656 4023 7730
rect 4026 7656 4045 7800
rect 4060 7656 4066 7800
rect 4075 7730 4088 7800
rect 4140 7796 4162 7800
rect 4133 7774 4162 7788
rect 4215 7774 4231 7788
rect 4269 7784 4275 7786
rect 4282 7784 4390 7800
rect 4397 7784 4403 7786
rect 4411 7784 4426 7800
rect 4492 7794 4511 7797
rect 4133 7772 4231 7774
rect 4258 7772 4426 7784
rect 4441 7774 4457 7788
rect 4492 7775 4514 7794
rect 4524 7788 4540 7789
rect 4523 7786 4540 7788
rect 4524 7781 4540 7786
rect 4514 7774 4520 7775
rect 4523 7774 4552 7781
rect 4441 7773 4552 7774
rect 4441 7772 4558 7773
rect 4117 7764 4168 7772
rect 4215 7764 4249 7772
rect 4117 7752 4142 7764
rect 4149 7752 4168 7764
rect 4222 7762 4249 7764
rect 4258 7762 4479 7772
rect 4514 7769 4520 7772
rect 4222 7758 4479 7762
rect 4117 7744 4168 7752
rect 4215 7744 4479 7758
rect 4523 7764 4558 7772
rect 4069 7696 4088 7730
rect 4133 7736 4162 7744
rect 4133 7730 4150 7736
rect 4133 7728 4167 7730
rect 4215 7728 4231 7744
rect 4232 7734 4440 7744
rect 4441 7734 4457 7744
rect 4505 7740 4520 7755
rect 4523 7752 4524 7764
rect 4531 7752 4558 7764
rect 4523 7744 4558 7752
rect 4523 7743 4552 7744
rect 4243 7730 4457 7734
rect 4258 7728 4457 7730
rect 4492 7730 4505 7740
rect 4523 7730 4540 7743
rect 4492 7728 4540 7730
rect 4134 7724 4167 7728
rect 4130 7722 4167 7724
rect 4130 7721 4197 7722
rect 4130 7716 4161 7721
rect 4167 7716 4197 7721
rect 4130 7712 4197 7716
rect 4103 7709 4197 7712
rect 4103 7702 4152 7709
rect 4103 7696 4133 7702
rect 4152 7697 4157 7702
rect 4069 7680 4149 7696
rect 4161 7688 4197 7709
rect 4258 7704 4447 7728
rect 4492 7727 4539 7728
rect 4505 7722 4539 7727
rect 4273 7701 4447 7704
rect 4266 7698 4447 7701
rect 4475 7721 4539 7722
rect 4069 7678 4088 7680
rect 4103 7678 4137 7680
rect 4069 7662 4149 7678
rect 4069 7656 4088 7662
rect 3785 7630 3888 7640
rect 3739 7628 3888 7630
rect 3909 7628 3944 7640
rect 3578 7626 3740 7628
rect 3590 7606 3609 7626
rect 3624 7624 3654 7626
rect 3473 7598 3514 7606
rect 3596 7602 3609 7606
rect 3661 7610 3740 7626
rect 3772 7626 3944 7628
rect 3772 7610 3851 7626
rect 3858 7624 3888 7626
rect 3436 7588 3465 7598
rect 3479 7588 3508 7598
rect 3523 7588 3553 7602
rect 3596 7588 3639 7602
rect 3661 7598 3851 7610
rect 3916 7606 3922 7626
rect 3646 7588 3676 7598
rect 3677 7588 3835 7598
rect 3839 7588 3869 7598
rect 3873 7588 3903 7602
rect 3931 7588 3944 7626
rect 4016 7640 4045 7656
rect 4059 7640 4088 7656
rect 4103 7646 4133 7662
rect 4161 7640 4167 7688
rect 4170 7682 4189 7688
rect 4204 7682 4234 7690
rect 4170 7674 4234 7682
rect 4170 7658 4250 7674
rect 4266 7667 4328 7698
rect 4344 7667 4406 7698
rect 4475 7696 4524 7721
rect 4539 7696 4569 7712
rect 4438 7682 4468 7690
rect 4475 7688 4585 7696
rect 4438 7674 4483 7682
rect 4170 7656 4189 7658
rect 4204 7656 4250 7658
rect 4170 7640 4250 7656
rect 4277 7654 4312 7667
rect 4353 7664 4390 7667
rect 4353 7662 4395 7664
rect 4282 7651 4312 7654
rect 4291 7647 4298 7651
rect 4298 7646 4299 7647
rect 4257 7640 4267 7646
rect 4016 7632 4051 7640
rect 4016 7606 4017 7632
rect 4024 7606 4051 7632
rect 3959 7588 3989 7602
rect 4016 7598 4051 7606
rect 4053 7632 4094 7640
rect 4053 7606 4068 7632
rect 4075 7606 4094 7632
rect 4158 7628 4189 7640
rect 4204 7628 4307 7640
rect 4319 7630 4345 7656
rect 4360 7651 4390 7662
rect 4422 7658 4484 7674
rect 4422 7656 4468 7658
rect 4422 7640 4484 7656
rect 4496 7640 4502 7688
rect 4505 7680 4585 7688
rect 4505 7678 4524 7680
rect 4539 7678 4573 7680
rect 4505 7662 4585 7678
rect 4505 7640 4524 7662
rect 4539 7646 4569 7662
rect 4597 7656 4603 7730
rect 4606 7656 4625 7800
rect 4640 7656 4646 7800
rect 4655 7730 4668 7800
rect 4720 7796 4742 7800
rect 4713 7774 4742 7788
rect 4795 7774 4811 7788
rect 4849 7784 4855 7786
rect 4862 7784 4970 7800
rect 4977 7784 4983 7786
rect 4991 7784 5006 7800
rect 5072 7794 5091 7797
rect 4713 7772 4811 7774
rect 4838 7772 5006 7784
rect 5021 7774 5037 7788
rect 5072 7775 5094 7794
rect 5104 7788 5120 7789
rect 5103 7786 5120 7788
rect 5104 7781 5120 7786
rect 5094 7774 5100 7775
rect 5103 7774 5132 7781
rect 5021 7773 5132 7774
rect 5021 7772 5138 7773
rect 4697 7764 4748 7772
rect 4795 7764 4829 7772
rect 4697 7752 4722 7764
rect 4729 7752 4748 7764
rect 4802 7762 4829 7764
rect 4838 7762 5059 7772
rect 5094 7769 5100 7772
rect 4802 7758 5059 7762
rect 4697 7744 4748 7752
rect 4795 7744 5059 7758
rect 5103 7764 5138 7772
rect 4649 7696 4668 7730
rect 4713 7736 4742 7744
rect 4713 7730 4730 7736
rect 4713 7728 4747 7730
rect 4795 7728 4811 7744
rect 4812 7734 5020 7744
rect 5021 7734 5037 7744
rect 5085 7740 5100 7755
rect 5103 7752 5104 7764
rect 5111 7752 5138 7764
rect 5103 7744 5138 7752
rect 5103 7743 5132 7744
rect 4823 7730 5037 7734
rect 4838 7728 5037 7730
rect 5072 7730 5085 7740
rect 5103 7730 5120 7743
rect 5072 7728 5120 7730
rect 4714 7724 4747 7728
rect 4710 7722 4747 7724
rect 4710 7721 4777 7722
rect 4710 7716 4741 7721
rect 4747 7716 4777 7721
rect 4710 7712 4777 7716
rect 4683 7709 4777 7712
rect 4683 7702 4732 7709
rect 4683 7696 4713 7702
rect 4732 7697 4737 7702
rect 4649 7680 4729 7696
rect 4741 7688 4777 7709
rect 4838 7704 5027 7728
rect 5072 7727 5119 7728
rect 5085 7722 5119 7727
rect 4853 7701 5027 7704
rect 4846 7698 5027 7701
rect 5055 7721 5119 7722
rect 4649 7678 4668 7680
rect 4683 7678 4717 7680
rect 4649 7662 4729 7678
rect 4649 7656 4668 7662
rect 4365 7630 4468 7640
rect 4319 7628 4468 7630
rect 4489 7628 4524 7640
rect 4158 7626 4320 7628
rect 4170 7606 4189 7626
rect 4204 7624 4234 7626
rect 4053 7598 4094 7606
rect 4176 7602 4189 7606
rect 4241 7610 4320 7626
rect 4352 7626 4524 7628
rect 4352 7610 4431 7626
rect 4438 7624 4468 7626
rect 4016 7588 4045 7598
rect 4059 7588 4088 7598
rect 4103 7588 4133 7602
rect 4176 7588 4219 7602
rect 4241 7598 4431 7610
rect 4496 7606 4502 7626
rect 4226 7588 4256 7598
rect 4257 7588 4415 7598
rect 4419 7588 4449 7598
rect 4453 7588 4483 7602
rect 4511 7588 4524 7626
rect 4596 7640 4625 7656
rect 4639 7640 4668 7656
rect 4683 7646 4713 7662
rect 4741 7640 4747 7688
rect 4750 7682 4769 7688
rect 4784 7682 4814 7690
rect 4750 7674 4814 7682
rect 4750 7658 4830 7674
rect 4846 7667 4908 7698
rect 4924 7667 4986 7698
rect 5055 7696 5104 7721
rect 5119 7696 5149 7712
rect 5018 7682 5048 7690
rect 5055 7688 5165 7696
rect 5018 7674 5063 7682
rect 4750 7656 4769 7658
rect 4784 7656 4830 7658
rect 4750 7640 4830 7656
rect 4857 7654 4892 7667
rect 4933 7664 4970 7667
rect 4933 7662 4975 7664
rect 4862 7651 4892 7654
rect 4871 7647 4878 7651
rect 4878 7646 4879 7647
rect 4837 7640 4847 7646
rect 4596 7632 4631 7640
rect 4596 7606 4597 7632
rect 4604 7606 4631 7632
rect 4539 7588 4569 7602
rect 4596 7598 4631 7606
rect 4633 7632 4674 7640
rect 4633 7606 4648 7632
rect 4655 7606 4674 7632
rect 4738 7628 4769 7640
rect 4784 7628 4887 7640
rect 4899 7630 4925 7656
rect 4940 7651 4970 7662
rect 5002 7658 5064 7674
rect 5002 7656 5048 7658
rect 5002 7640 5064 7656
rect 5076 7640 5082 7688
rect 5085 7680 5165 7688
rect 5085 7678 5104 7680
rect 5119 7678 5153 7680
rect 5085 7662 5165 7678
rect 5085 7640 5104 7662
rect 5119 7646 5149 7662
rect 5177 7656 5183 7730
rect 5186 7656 5205 7800
rect 5220 7656 5226 7800
rect 5235 7730 5248 7800
rect 5300 7796 5322 7800
rect 5293 7774 5322 7788
rect 5375 7774 5391 7788
rect 5429 7784 5435 7786
rect 5442 7784 5550 7800
rect 5557 7784 5563 7786
rect 5571 7784 5586 7800
rect 5652 7794 5671 7797
rect 5293 7772 5391 7774
rect 5418 7772 5586 7784
rect 5601 7774 5617 7788
rect 5652 7775 5674 7794
rect 5684 7788 5700 7789
rect 5683 7786 5700 7788
rect 5684 7781 5700 7786
rect 5674 7774 5680 7775
rect 5683 7774 5712 7781
rect 5601 7773 5712 7774
rect 5601 7772 5718 7773
rect 5277 7764 5328 7772
rect 5375 7764 5409 7772
rect 5277 7752 5302 7764
rect 5309 7752 5328 7764
rect 5382 7762 5409 7764
rect 5418 7762 5639 7772
rect 5674 7769 5680 7772
rect 5382 7758 5639 7762
rect 5277 7744 5328 7752
rect 5375 7744 5639 7758
rect 5683 7764 5718 7772
rect 5229 7696 5248 7730
rect 5293 7736 5322 7744
rect 5293 7730 5310 7736
rect 5293 7728 5327 7730
rect 5375 7728 5391 7744
rect 5392 7734 5600 7744
rect 5601 7734 5617 7744
rect 5665 7740 5680 7755
rect 5683 7752 5684 7764
rect 5691 7752 5718 7764
rect 5683 7744 5718 7752
rect 5683 7743 5712 7744
rect 5403 7730 5617 7734
rect 5418 7728 5617 7730
rect 5652 7730 5665 7740
rect 5683 7730 5700 7743
rect 5652 7728 5700 7730
rect 5294 7724 5327 7728
rect 5290 7722 5327 7724
rect 5290 7721 5357 7722
rect 5290 7716 5321 7721
rect 5327 7716 5357 7721
rect 5290 7712 5357 7716
rect 5263 7709 5357 7712
rect 5263 7702 5312 7709
rect 5263 7696 5293 7702
rect 5312 7697 5317 7702
rect 5229 7680 5309 7696
rect 5321 7688 5357 7709
rect 5418 7704 5607 7728
rect 5652 7727 5699 7728
rect 5665 7722 5699 7727
rect 5433 7701 5607 7704
rect 5426 7698 5607 7701
rect 5635 7721 5699 7722
rect 5229 7678 5248 7680
rect 5263 7678 5297 7680
rect 5229 7662 5309 7678
rect 5229 7656 5248 7662
rect 4945 7630 5048 7640
rect 4899 7628 5048 7630
rect 5069 7628 5104 7640
rect 4738 7626 4900 7628
rect 4750 7606 4769 7626
rect 4784 7624 4814 7626
rect 4633 7598 4674 7606
rect 4756 7602 4769 7606
rect 4821 7610 4900 7626
rect 4932 7626 5104 7628
rect 4932 7610 5011 7626
rect 5018 7624 5048 7626
rect 4596 7588 4625 7598
rect 4639 7588 4668 7598
rect 4683 7588 4713 7602
rect 4756 7588 4799 7602
rect 4821 7598 5011 7610
rect 5076 7606 5082 7626
rect 4806 7588 4836 7598
rect 4837 7588 4995 7598
rect 4999 7588 5029 7598
rect 5033 7588 5063 7602
rect 5091 7588 5104 7626
rect 5176 7640 5205 7656
rect 5219 7640 5248 7656
rect 5263 7646 5293 7662
rect 5321 7640 5327 7688
rect 5330 7682 5349 7688
rect 5364 7682 5394 7690
rect 5330 7674 5394 7682
rect 5330 7658 5410 7674
rect 5426 7667 5488 7698
rect 5504 7667 5566 7698
rect 5635 7696 5684 7721
rect 5699 7696 5729 7712
rect 5598 7682 5628 7690
rect 5635 7688 5745 7696
rect 5598 7674 5643 7682
rect 5330 7656 5349 7658
rect 5364 7656 5410 7658
rect 5330 7640 5410 7656
rect 5437 7654 5472 7667
rect 5513 7664 5550 7667
rect 5513 7662 5555 7664
rect 5442 7651 5472 7654
rect 5451 7647 5458 7651
rect 5458 7646 5459 7647
rect 5417 7640 5427 7646
rect 5176 7632 5211 7640
rect 5176 7606 5177 7632
rect 5184 7606 5211 7632
rect 5119 7588 5149 7602
rect 5176 7598 5211 7606
rect 5213 7632 5254 7640
rect 5213 7606 5228 7632
rect 5235 7606 5254 7632
rect 5318 7628 5349 7640
rect 5364 7628 5467 7640
rect 5479 7630 5505 7656
rect 5520 7651 5550 7662
rect 5582 7658 5644 7674
rect 5582 7656 5628 7658
rect 5582 7640 5644 7656
rect 5656 7640 5662 7688
rect 5665 7680 5745 7688
rect 5665 7678 5684 7680
rect 5699 7678 5733 7680
rect 5665 7662 5745 7678
rect 5665 7640 5684 7662
rect 5699 7646 5729 7662
rect 5757 7656 5763 7730
rect 5766 7656 5785 7800
rect 5800 7656 5806 7800
rect 5815 7730 5828 7800
rect 5880 7796 5902 7800
rect 5873 7774 5902 7788
rect 5955 7774 5971 7788
rect 6009 7784 6015 7786
rect 6022 7784 6130 7800
rect 6137 7784 6143 7786
rect 6151 7784 6166 7800
rect 6232 7794 6251 7797
rect 5873 7772 5971 7774
rect 5998 7772 6166 7784
rect 6181 7774 6197 7788
rect 6232 7775 6254 7794
rect 6264 7788 6280 7789
rect 6263 7786 6280 7788
rect 6264 7781 6280 7786
rect 6254 7774 6260 7775
rect 6263 7774 6292 7781
rect 6181 7773 6292 7774
rect 6181 7772 6298 7773
rect 5857 7764 5908 7772
rect 5955 7764 5989 7772
rect 5857 7752 5882 7764
rect 5889 7752 5908 7764
rect 5962 7762 5989 7764
rect 5998 7762 6219 7772
rect 6254 7769 6260 7772
rect 5962 7758 6219 7762
rect 5857 7744 5908 7752
rect 5955 7744 6219 7758
rect 6263 7764 6298 7772
rect 5809 7696 5828 7730
rect 5873 7736 5902 7744
rect 5873 7730 5890 7736
rect 5873 7728 5907 7730
rect 5955 7728 5971 7744
rect 5972 7734 6180 7744
rect 6181 7734 6197 7744
rect 6245 7740 6260 7755
rect 6263 7752 6264 7764
rect 6271 7752 6298 7764
rect 6263 7744 6298 7752
rect 6263 7743 6292 7744
rect 5983 7730 6197 7734
rect 5998 7728 6197 7730
rect 6232 7730 6245 7740
rect 6263 7730 6280 7743
rect 6232 7728 6280 7730
rect 5874 7724 5907 7728
rect 5870 7722 5907 7724
rect 5870 7721 5937 7722
rect 5870 7716 5901 7721
rect 5907 7716 5937 7721
rect 5870 7712 5937 7716
rect 5843 7709 5937 7712
rect 5843 7702 5892 7709
rect 5843 7696 5873 7702
rect 5892 7697 5897 7702
rect 5809 7680 5889 7696
rect 5901 7688 5937 7709
rect 5998 7704 6187 7728
rect 6232 7727 6279 7728
rect 6245 7722 6279 7727
rect 6013 7701 6187 7704
rect 6006 7698 6187 7701
rect 6215 7721 6279 7722
rect 5809 7678 5828 7680
rect 5843 7678 5877 7680
rect 5809 7662 5889 7678
rect 5809 7656 5828 7662
rect 5525 7630 5628 7640
rect 5479 7628 5628 7630
rect 5649 7628 5684 7640
rect 5318 7626 5480 7628
rect 5330 7606 5349 7626
rect 5364 7624 5394 7626
rect 5213 7598 5254 7606
rect 5336 7602 5349 7606
rect 5401 7610 5480 7626
rect 5512 7626 5684 7628
rect 5512 7610 5591 7626
rect 5598 7624 5628 7626
rect 5176 7588 5205 7598
rect 5219 7588 5248 7598
rect 5263 7588 5293 7602
rect 5336 7588 5379 7602
rect 5401 7598 5591 7610
rect 5656 7606 5662 7626
rect 5386 7588 5416 7598
rect 5417 7588 5575 7598
rect 5579 7588 5609 7598
rect 5613 7588 5643 7602
rect 5671 7588 5684 7626
rect 5756 7640 5785 7656
rect 5799 7640 5828 7656
rect 5843 7646 5873 7662
rect 5901 7640 5907 7688
rect 5910 7682 5929 7688
rect 5944 7682 5974 7690
rect 5910 7674 5974 7682
rect 5910 7658 5990 7674
rect 6006 7667 6068 7698
rect 6084 7667 6146 7698
rect 6215 7696 6264 7721
rect 6279 7696 6309 7712
rect 6178 7682 6208 7690
rect 6215 7688 6325 7696
rect 6178 7674 6223 7682
rect 5910 7656 5929 7658
rect 5944 7656 5990 7658
rect 5910 7640 5990 7656
rect 6017 7654 6052 7667
rect 6093 7664 6130 7667
rect 6093 7662 6135 7664
rect 6022 7651 6052 7654
rect 6031 7647 6038 7651
rect 6038 7646 6039 7647
rect 5997 7640 6007 7646
rect 5756 7632 5791 7640
rect 5756 7606 5757 7632
rect 5764 7606 5791 7632
rect 5699 7588 5729 7602
rect 5756 7598 5791 7606
rect 5793 7632 5834 7640
rect 5793 7606 5808 7632
rect 5815 7606 5834 7632
rect 5898 7628 5929 7640
rect 5944 7628 6047 7640
rect 6059 7630 6085 7656
rect 6100 7651 6130 7662
rect 6162 7658 6224 7674
rect 6162 7656 6208 7658
rect 6162 7640 6224 7656
rect 6236 7640 6242 7688
rect 6245 7680 6325 7688
rect 6245 7678 6264 7680
rect 6279 7678 6313 7680
rect 6245 7662 6325 7678
rect 6245 7640 6264 7662
rect 6279 7646 6309 7662
rect 6337 7656 6343 7730
rect 6346 7656 6365 7800
rect 6380 7656 6386 7800
rect 6395 7730 6408 7800
rect 6460 7796 6482 7800
rect 6453 7774 6482 7788
rect 6535 7774 6551 7788
rect 6589 7784 6595 7786
rect 6602 7784 6710 7800
rect 6717 7784 6723 7786
rect 6731 7784 6746 7800
rect 6812 7794 6831 7797
rect 6453 7772 6551 7774
rect 6578 7772 6746 7784
rect 6761 7774 6777 7788
rect 6812 7775 6834 7794
rect 6844 7788 6860 7789
rect 6843 7786 6860 7788
rect 6844 7781 6860 7786
rect 6834 7774 6840 7775
rect 6843 7774 6872 7781
rect 6761 7773 6872 7774
rect 6761 7772 6878 7773
rect 6437 7764 6488 7772
rect 6535 7764 6569 7772
rect 6437 7752 6462 7764
rect 6469 7752 6488 7764
rect 6542 7762 6569 7764
rect 6578 7762 6799 7772
rect 6834 7769 6840 7772
rect 6542 7758 6799 7762
rect 6437 7744 6488 7752
rect 6535 7744 6799 7758
rect 6843 7764 6878 7772
rect 6389 7696 6408 7730
rect 6453 7736 6482 7744
rect 6453 7730 6470 7736
rect 6453 7728 6487 7730
rect 6535 7728 6551 7744
rect 6552 7734 6760 7744
rect 6761 7734 6777 7744
rect 6825 7740 6840 7755
rect 6843 7752 6844 7764
rect 6851 7752 6878 7764
rect 6843 7744 6878 7752
rect 6843 7743 6872 7744
rect 6563 7730 6777 7734
rect 6578 7728 6777 7730
rect 6812 7730 6825 7740
rect 6843 7730 6860 7743
rect 6812 7728 6860 7730
rect 6454 7724 6487 7728
rect 6450 7722 6487 7724
rect 6450 7721 6517 7722
rect 6450 7716 6481 7721
rect 6487 7716 6517 7721
rect 6450 7712 6517 7716
rect 6423 7709 6517 7712
rect 6423 7702 6472 7709
rect 6423 7696 6453 7702
rect 6472 7697 6477 7702
rect 6389 7680 6469 7696
rect 6481 7688 6517 7709
rect 6578 7704 6767 7728
rect 6812 7727 6859 7728
rect 6825 7722 6859 7727
rect 6593 7701 6767 7704
rect 6586 7698 6767 7701
rect 6795 7721 6859 7722
rect 6389 7678 6408 7680
rect 6423 7678 6457 7680
rect 6389 7662 6469 7678
rect 6389 7656 6408 7662
rect 6105 7630 6208 7640
rect 6059 7628 6208 7630
rect 6229 7628 6264 7640
rect 5898 7626 6060 7628
rect 5910 7606 5929 7626
rect 5944 7624 5974 7626
rect 5793 7598 5834 7606
rect 5916 7602 5929 7606
rect 5981 7610 6060 7626
rect 6092 7626 6264 7628
rect 6092 7610 6171 7626
rect 6178 7624 6208 7626
rect 5756 7588 5785 7598
rect 5799 7588 5828 7598
rect 5843 7588 5873 7602
rect 5916 7588 5959 7602
rect 5981 7598 6171 7610
rect 6236 7606 6242 7626
rect 5966 7588 5996 7598
rect 5997 7588 6155 7598
rect 6159 7588 6189 7598
rect 6193 7588 6223 7602
rect 6251 7588 6264 7626
rect 6336 7640 6365 7656
rect 6379 7640 6408 7656
rect 6423 7646 6453 7662
rect 6481 7640 6487 7688
rect 6490 7682 6509 7688
rect 6524 7682 6554 7690
rect 6490 7674 6554 7682
rect 6490 7658 6570 7674
rect 6586 7667 6648 7698
rect 6664 7667 6726 7698
rect 6795 7696 6844 7721
rect 6859 7696 6889 7712
rect 6758 7682 6788 7690
rect 6795 7688 6905 7696
rect 6758 7674 6803 7682
rect 6490 7656 6509 7658
rect 6524 7656 6570 7658
rect 6490 7640 6570 7656
rect 6597 7654 6632 7667
rect 6673 7664 6710 7667
rect 6673 7662 6715 7664
rect 6602 7651 6632 7654
rect 6611 7647 6618 7651
rect 6618 7646 6619 7647
rect 6577 7640 6587 7646
rect 6336 7632 6371 7640
rect 6336 7606 6337 7632
rect 6344 7606 6371 7632
rect 6279 7588 6309 7602
rect 6336 7598 6371 7606
rect 6373 7632 6414 7640
rect 6373 7606 6388 7632
rect 6395 7606 6414 7632
rect 6478 7628 6509 7640
rect 6524 7628 6627 7640
rect 6639 7630 6665 7656
rect 6680 7651 6710 7662
rect 6742 7658 6804 7674
rect 6742 7656 6788 7658
rect 6742 7640 6804 7656
rect 6816 7640 6822 7688
rect 6825 7680 6905 7688
rect 6825 7678 6844 7680
rect 6859 7678 6893 7680
rect 6825 7662 6905 7678
rect 6825 7640 6844 7662
rect 6859 7646 6889 7662
rect 6917 7656 6923 7730
rect 6926 7656 6945 7800
rect 6960 7656 6966 7800
rect 6975 7730 6988 7800
rect 7040 7796 7062 7800
rect 7033 7774 7062 7788
rect 7115 7774 7131 7788
rect 7169 7784 7175 7786
rect 7182 7784 7290 7800
rect 7297 7784 7303 7786
rect 7311 7784 7326 7800
rect 7392 7794 7411 7797
rect 7033 7772 7131 7774
rect 7158 7772 7326 7784
rect 7341 7774 7357 7788
rect 7392 7775 7414 7794
rect 7424 7788 7440 7789
rect 7423 7786 7440 7788
rect 7424 7781 7440 7786
rect 7414 7774 7420 7775
rect 7423 7774 7452 7781
rect 7341 7773 7452 7774
rect 7341 7772 7458 7773
rect 7017 7764 7068 7772
rect 7115 7764 7149 7772
rect 7017 7752 7042 7764
rect 7049 7752 7068 7764
rect 7122 7762 7149 7764
rect 7158 7762 7379 7772
rect 7414 7769 7420 7772
rect 7122 7758 7379 7762
rect 7017 7744 7068 7752
rect 7115 7744 7379 7758
rect 7423 7764 7458 7772
rect 6969 7696 6988 7730
rect 7033 7736 7062 7744
rect 7033 7730 7050 7736
rect 7033 7728 7067 7730
rect 7115 7728 7131 7744
rect 7132 7734 7340 7744
rect 7341 7734 7357 7744
rect 7405 7740 7420 7755
rect 7423 7752 7424 7764
rect 7431 7752 7458 7764
rect 7423 7744 7458 7752
rect 7423 7743 7452 7744
rect 7143 7730 7357 7734
rect 7158 7728 7357 7730
rect 7392 7730 7405 7740
rect 7423 7730 7440 7743
rect 7392 7728 7440 7730
rect 7034 7724 7067 7728
rect 7030 7722 7067 7724
rect 7030 7721 7097 7722
rect 7030 7716 7061 7721
rect 7067 7716 7097 7721
rect 7030 7712 7097 7716
rect 7003 7709 7097 7712
rect 7003 7702 7052 7709
rect 7003 7696 7033 7702
rect 7052 7697 7057 7702
rect 6969 7680 7049 7696
rect 7061 7688 7097 7709
rect 7158 7704 7347 7728
rect 7392 7727 7439 7728
rect 7405 7722 7439 7727
rect 7173 7701 7347 7704
rect 7166 7698 7347 7701
rect 7375 7721 7439 7722
rect 6969 7678 6988 7680
rect 7003 7678 7037 7680
rect 6969 7662 7049 7678
rect 6969 7656 6988 7662
rect 6685 7630 6788 7640
rect 6639 7628 6788 7630
rect 6809 7628 6844 7640
rect 6478 7626 6640 7628
rect 6490 7606 6509 7626
rect 6524 7624 6554 7626
rect 6373 7598 6414 7606
rect 6496 7602 6509 7606
rect 6561 7610 6640 7626
rect 6672 7626 6844 7628
rect 6672 7610 6751 7626
rect 6758 7624 6788 7626
rect 6336 7588 6365 7598
rect 6379 7588 6408 7598
rect 6423 7588 6453 7602
rect 6496 7588 6539 7602
rect 6561 7598 6751 7610
rect 6816 7606 6822 7626
rect 6546 7588 6576 7598
rect 6577 7588 6735 7598
rect 6739 7588 6769 7598
rect 6773 7588 6803 7602
rect 6831 7588 6844 7626
rect 6916 7640 6945 7656
rect 6959 7640 6988 7656
rect 7003 7646 7033 7662
rect 7061 7640 7067 7688
rect 7070 7682 7089 7688
rect 7104 7682 7134 7690
rect 7070 7674 7134 7682
rect 7070 7658 7150 7674
rect 7166 7667 7228 7698
rect 7244 7667 7306 7698
rect 7375 7696 7424 7721
rect 7439 7696 7469 7712
rect 7338 7682 7368 7690
rect 7375 7688 7485 7696
rect 7338 7674 7383 7682
rect 7070 7656 7089 7658
rect 7104 7656 7150 7658
rect 7070 7640 7150 7656
rect 7177 7654 7212 7667
rect 7253 7664 7290 7667
rect 7253 7662 7295 7664
rect 7182 7651 7212 7654
rect 7191 7647 7198 7651
rect 7198 7646 7199 7647
rect 7157 7640 7167 7646
rect 6916 7632 6951 7640
rect 6916 7606 6917 7632
rect 6924 7606 6951 7632
rect 6859 7588 6889 7602
rect 6916 7598 6951 7606
rect 6953 7632 6994 7640
rect 6953 7606 6968 7632
rect 6975 7606 6994 7632
rect 7058 7628 7089 7640
rect 7104 7628 7207 7640
rect 7219 7630 7245 7656
rect 7260 7651 7290 7662
rect 7322 7658 7384 7674
rect 7322 7656 7368 7658
rect 7322 7640 7384 7656
rect 7396 7640 7402 7688
rect 7405 7680 7485 7688
rect 7405 7678 7424 7680
rect 7439 7678 7473 7680
rect 7405 7662 7485 7678
rect 7405 7640 7424 7662
rect 7439 7646 7469 7662
rect 7497 7656 7503 7730
rect 7506 7656 7525 7800
rect 7540 7656 7546 7800
rect 7555 7730 7568 7800
rect 7620 7796 7642 7800
rect 7613 7774 7642 7788
rect 7695 7774 7711 7788
rect 7749 7784 7755 7786
rect 7762 7784 7870 7800
rect 7877 7784 7883 7786
rect 7891 7784 7906 7800
rect 7972 7794 7991 7797
rect 7613 7772 7711 7774
rect 7738 7772 7906 7784
rect 7921 7774 7937 7788
rect 7972 7775 7994 7794
rect 8004 7788 8020 7789
rect 8003 7786 8020 7788
rect 8004 7781 8020 7786
rect 7994 7774 8000 7775
rect 8003 7774 8032 7781
rect 7921 7773 8032 7774
rect 7921 7772 8038 7773
rect 7597 7764 7648 7772
rect 7695 7764 7729 7772
rect 7597 7752 7622 7764
rect 7629 7752 7648 7764
rect 7702 7762 7729 7764
rect 7738 7762 7959 7772
rect 7994 7769 8000 7772
rect 7702 7758 7959 7762
rect 7597 7744 7648 7752
rect 7695 7744 7959 7758
rect 8003 7764 8038 7772
rect 7549 7696 7568 7730
rect 7613 7736 7642 7744
rect 7613 7730 7630 7736
rect 7613 7728 7647 7730
rect 7695 7728 7711 7744
rect 7712 7734 7920 7744
rect 7921 7734 7937 7744
rect 7985 7740 8000 7755
rect 8003 7752 8004 7764
rect 8011 7752 8038 7764
rect 8003 7744 8038 7752
rect 8003 7743 8032 7744
rect 7723 7730 7937 7734
rect 7738 7728 7937 7730
rect 7972 7730 7985 7740
rect 8003 7730 8020 7743
rect 7972 7728 8020 7730
rect 7614 7724 7647 7728
rect 7610 7722 7647 7724
rect 7610 7721 7677 7722
rect 7610 7716 7641 7721
rect 7647 7716 7677 7721
rect 7610 7712 7677 7716
rect 7583 7709 7677 7712
rect 7583 7702 7632 7709
rect 7583 7696 7613 7702
rect 7632 7697 7637 7702
rect 7549 7680 7629 7696
rect 7641 7688 7677 7709
rect 7738 7704 7927 7728
rect 7972 7727 8019 7728
rect 7985 7722 8019 7727
rect 7753 7701 7927 7704
rect 7746 7698 7927 7701
rect 7955 7721 8019 7722
rect 7549 7678 7568 7680
rect 7583 7678 7617 7680
rect 7549 7662 7629 7678
rect 7549 7656 7568 7662
rect 7265 7630 7368 7640
rect 7219 7628 7368 7630
rect 7389 7628 7424 7640
rect 7058 7626 7220 7628
rect 7070 7606 7089 7626
rect 7104 7624 7134 7626
rect 6953 7598 6994 7606
rect 7076 7602 7089 7606
rect 7141 7610 7220 7626
rect 7252 7626 7424 7628
rect 7252 7610 7331 7626
rect 7338 7624 7368 7626
rect 6916 7588 6945 7598
rect 6959 7588 6988 7598
rect 7003 7588 7033 7602
rect 7076 7588 7119 7602
rect 7141 7598 7331 7610
rect 7396 7606 7402 7626
rect 7126 7588 7156 7598
rect 7157 7588 7315 7598
rect 7319 7588 7349 7598
rect 7353 7588 7383 7602
rect 7411 7588 7424 7626
rect 7496 7640 7525 7656
rect 7539 7640 7568 7656
rect 7583 7646 7613 7662
rect 7641 7640 7647 7688
rect 7650 7682 7669 7688
rect 7684 7682 7714 7690
rect 7650 7674 7714 7682
rect 7650 7658 7730 7674
rect 7746 7667 7808 7698
rect 7824 7667 7886 7698
rect 7955 7696 8004 7721
rect 8019 7696 8049 7712
rect 7918 7682 7948 7690
rect 7955 7688 8065 7696
rect 7918 7674 7963 7682
rect 7650 7656 7669 7658
rect 7684 7656 7730 7658
rect 7650 7640 7730 7656
rect 7757 7654 7792 7667
rect 7833 7664 7870 7667
rect 7833 7662 7875 7664
rect 7762 7651 7792 7654
rect 7771 7647 7778 7651
rect 7778 7646 7779 7647
rect 7737 7640 7747 7646
rect 7496 7632 7531 7640
rect 7496 7606 7497 7632
rect 7504 7606 7531 7632
rect 7439 7588 7469 7602
rect 7496 7598 7531 7606
rect 7533 7632 7574 7640
rect 7533 7606 7548 7632
rect 7555 7606 7574 7632
rect 7638 7628 7669 7640
rect 7684 7628 7787 7640
rect 7799 7630 7825 7656
rect 7840 7651 7870 7662
rect 7902 7658 7964 7674
rect 7902 7656 7948 7658
rect 7902 7640 7964 7656
rect 7976 7640 7982 7688
rect 7985 7680 8065 7688
rect 7985 7678 8004 7680
rect 8019 7678 8053 7680
rect 7985 7662 8065 7678
rect 7985 7640 8004 7662
rect 8019 7646 8049 7662
rect 8077 7656 8083 7730
rect 8086 7656 8105 7800
rect 8120 7656 8126 7800
rect 8135 7730 8148 7800
rect 8200 7796 8222 7800
rect 8193 7774 8222 7788
rect 8275 7774 8291 7788
rect 8329 7784 8335 7786
rect 8342 7784 8450 7800
rect 8457 7784 8463 7786
rect 8471 7784 8486 7800
rect 8552 7794 8571 7797
rect 8193 7772 8291 7774
rect 8318 7772 8486 7784
rect 8501 7774 8517 7788
rect 8552 7775 8574 7794
rect 8584 7788 8600 7789
rect 8583 7786 8600 7788
rect 8584 7781 8600 7786
rect 8574 7774 8580 7775
rect 8583 7774 8612 7781
rect 8501 7773 8612 7774
rect 8501 7772 8618 7773
rect 8177 7764 8228 7772
rect 8275 7764 8309 7772
rect 8177 7752 8202 7764
rect 8209 7752 8228 7764
rect 8282 7762 8309 7764
rect 8318 7762 8539 7772
rect 8574 7769 8580 7772
rect 8282 7758 8539 7762
rect 8177 7744 8228 7752
rect 8275 7744 8539 7758
rect 8583 7764 8618 7772
rect 8129 7696 8148 7730
rect 8193 7736 8222 7744
rect 8193 7730 8210 7736
rect 8193 7728 8227 7730
rect 8275 7728 8291 7744
rect 8292 7734 8500 7744
rect 8501 7734 8517 7744
rect 8565 7740 8580 7755
rect 8583 7752 8584 7764
rect 8591 7752 8618 7764
rect 8583 7744 8618 7752
rect 8583 7743 8612 7744
rect 8303 7730 8517 7734
rect 8318 7728 8517 7730
rect 8552 7730 8565 7740
rect 8583 7730 8600 7743
rect 8552 7728 8600 7730
rect 8194 7724 8227 7728
rect 8190 7722 8227 7724
rect 8190 7721 8257 7722
rect 8190 7716 8221 7721
rect 8227 7716 8257 7721
rect 8190 7712 8257 7716
rect 8163 7709 8257 7712
rect 8163 7702 8212 7709
rect 8163 7696 8193 7702
rect 8212 7697 8217 7702
rect 8129 7680 8209 7696
rect 8221 7688 8257 7709
rect 8318 7704 8507 7728
rect 8552 7727 8599 7728
rect 8565 7722 8599 7727
rect 8333 7701 8507 7704
rect 8326 7698 8507 7701
rect 8535 7721 8599 7722
rect 8129 7678 8148 7680
rect 8163 7678 8197 7680
rect 8129 7662 8209 7678
rect 8129 7656 8148 7662
rect 7845 7630 7948 7640
rect 7799 7628 7948 7630
rect 7969 7628 8004 7640
rect 7638 7626 7800 7628
rect 7650 7606 7669 7626
rect 7684 7624 7714 7626
rect 7533 7598 7574 7606
rect 7656 7602 7669 7606
rect 7721 7610 7800 7626
rect 7832 7626 8004 7628
rect 7832 7610 7911 7626
rect 7918 7624 7948 7626
rect 7496 7588 7525 7598
rect 7539 7588 7568 7598
rect 7583 7588 7613 7602
rect 7656 7588 7699 7602
rect 7721 7598 7911 7610
rect 7976 7606 7982 7626
rect 7706 7588 7736 7598
rect 7737 7588 7895 7598
rect 7899 7588 7929 7598
rect 7933 7588 7963 7602
rect 7991 7588 8004 7626
rect 8076 7640 8105 7656
rect 8119 7640 8148 7656
rect 8163 7646 8193 7662
rect 8221 7640 8227 7688
rect 8230 7682 8249 7688
rect 8264 7682 8294 7690
rect 8230 7674 8294 7682
rect 8230 7658 8310 7674
rect 8326 7667 8388 7698
rect 8404 7667 8466 7698
rect 8535 7696 8584 7721
rect 8599 7696 8629 7712
rect 8498 7682 8528 7690
rect 8535 7688 8645 7696
rect 8498 7674 8543 7682
rect 8230 7656 8249 7658
rect 8264 7656 8310 7658
rect 8230 7640 8310 7656
rect 8337 7654 8372 7667
rect 8413 7664 8450 7667
rect 8413 7662 8455 7664
rect 8342 7651 8372 7654
rect 8351 7647 8358 7651
rect 8358 7646 8359 7647
rect 8317 7640 8327 7646
rect 8076 7632 8111 7640
rect 8076 7606 8077 7632
rect 8084 7606 8111 7632
rect 8019 7588 8049 7602
rect 8076 7598 8111 7606
rect 8113 7632 8154 7640
rect 8113 7606 8128 7632
rect 8135 7606 8154 7632
rect 8218 7628 8249 7640
rect 8264 7628 8367 7640
rect 8379 7630 8405 7656
rect 8420 7651 8450 7662
rect 8482 7658 8544 7674
rect 8482 7656 8528 7658
rect 8482 7640 8544 7656
rect 8556 7640 8562 7688
rect 8565 7680 8645 7688
rect 8565 7678 8584 7680
rect 8599 7678 8633 7680
rect 8565 7662 8645 7678
rect 8565 7640 8584 7662
rect 8599 7646 8629 7662
rect 8657 7656 8663 7730
rect 8666 7656 8685 7800
rect 8700 7656 8706 7800
rect 8715 7730 8728 7800
rect 8780 7796 8802 7800
rect 8773 7774 8802 7788
rect 8855 7774 8871 7788
rect 8909 7784 8915 7786
rect 8922 7784 9030 7800
rect 9037 7784 9043 7786
rect 9051 7784 9066 7800
rect 9132 7794 9151 7797
rect 8773 7772 8871 7774
rect 8898 7772 9066 7784
rect 9081 7774 9097 7788
rect 9132 7775 9154 7794
rect 9164 7788 9180 7789
rect 9163 7786 9180 7788
rect 9164 7781 9180 7786
rect 9154 7774 9160 7775
rect 9163 7774 9192 7781
rect 9081 7773 9192 7774
rect 9081 7772 9198 7773
rect 8757 7764 8808 7772
rect 8855 7764 8889 7772
rect 8757 7752 8782 7764
rect 8789 7752 8808 7764
rect 8862 7762 8889 7764
rect 8898 7762 9119 7772
rect 9154 7769 9160 7772
rect 8862 7758 9119 7762
rect 8757 7744 8808 7752
rect 8855 7744 9119 7758
rect 9163 7764 9198 7772
rect 8709 7696 8728 7730
rect 8773 7736 8802 7744
rect 8773 7730 8790 7736
rect 8773 7728 8807 7730
rect 8855 7728 8871 7744
rect 8872 7734 9080 7744
rect 9081 7734 9097 7744
rect 9145 7740 9160 7755
rect 9163 7752 9164 7764
rect 9171 7752 9198 7764
rect 9163 7744 9198 7752
rect 9163 7743 9192 7744
rect 8883 7730 9097 7734
rect 8898 7728 9097 7730
rect 9132 7730 9145 7740
rect 9163 7730 9180 7743
rect 9132 7728 9180 7730
rect 8774 7724 8807 7728
rect 8770 7722 8807 7724
rect 8770 7721 8837 7722
rect 8770 7716 8801 7721
rect 8807 7716 8837 7721
rect 8770 7712 8837 7716
rect 8743 7709 8837 7712
rect 8743 7702 8792 7709
rect 8743 7696 8773 7702
rect 8792 7697 8797 7702
rect 8709 7680 8789 7696
rect 8801 7688 8837 7709
rect 8898 7704 9087 7728
rect 9132 7727 9179 7728
rect 9145 7722 9179 7727
rect 8913 7701 9087 7704
rect 8906 7698 9087 7701
rect 9115 7721 9179 7722
rect 8709 7678 8728 7680
rect 8743 7678 8777 7680
rect 8709 7662 8789 7678
rect 8709 7656 8728 7662
rect 8425 7630 8528 7640
rect 8379 7628 8528 7630
rect 8549 7628 8584 7640
rect 8218 7626 8380 7628
rect 8230 7606 8249 7626
rect 8264 7624 8294 7626
rect 8113 7598 8154 7606
rect 8236 7602 8249 7606
rect 8301 7610 8380 7626
rect 8412 7626 8584 7628
rect 8412 7610 8491 7626
rect 8498 7624 8528 7626
rect 8076 7588 8105 7598
rect 8119 7588 8148 7598
rect 8163 7588 8193 7602
rect 8236 7588 8279 7602
rect 8301 7598 8491 7610
rect 8556 7606 8562 7626
rect 8286 7588 8316 7598
rect 8317 7588 8475 7598
rect 8479 7588 8509 7598
rect 8513 7588 8543 7602
rect 8571 7588 8584 7626
rect 8656 7640 8685 7656
rect 8699 7640 8728 7656
rect 8743 7646 8773 7662
rect 8801 7640 8807 7688
rect 8810 7682 8829 7688
rect 8844 7682 8874 7690
rect 8810 7674 8874 7682
rect 8810 7658 8890 7674
rect 8906 7667 8968 7698
rect 8984 7667 9046 7698
rect 9115 7696 9164 7721
rect 9179 7696 9209 7712
rect 9078 7682 9108 7690
rect 9115 7688 9225 7696
rect 9078 7674 9123 7682
rect 8810 7656 8829 7658
rect 8844 7656 8890 7658
rect 8810 7640 8890 7656
rect 8917 7654 8952 7667
rect 8993 7664 9030 7667
rect 8993 7662 9035 7664
rect 8922 7651 8952 7654
rect 8931 7647 8938 7651
rect 8938 7646 8939 7647
rect 8897 7640 8907 7646
rect 8656 7632 8691 7640
rect 8656 7606 8657 7632
rect 8664 7606 8691 7632
rect 8599 7588 8629 7602
rect 8656 7598 8691 7606
rect 8693 7632 8734 7640
rect 8693 7606 8708 7632
rect 8715 7606 8734 7632
rect 8798 7628 8829 7640
rect 8844 7628 8947 7640
rect 8959 7630 8985 7656
rect 9000 7651 9030 7662
rect 9062 7658 9124 7674
rect 9062 7656 9108 7658
rect 9062 7640 9124 7656
rect 9136 7640 9142 7688
rect 9145 7680 9225 7688
rect 9145 7678 9164 7680
rect 9179 7678 9213 7680
rect 9145 7662 9225 7678
rect 9145 7640 9164 7662
rect 9179 7646 9209 7662
rect 9237 7656 9243 7730
rect 9246 7656 9265 7800
rect 9280 7656 9286 7800
rect 9295 7730 9308 7800
rect 9360 7796 9382 7800
rect 9353 7774 9382 7788
rect 9435 7774 9451 7788
rect 9489 7784 9495 7786
rect 9502 7784 9610 7800
rect 9617 7784 9623 7786
rect 9631 7784 9646 7800
rect 9712 7794 9731 7797
rect 9353 7772 9451 7774
rect 9478 7772 9646 7784
rect 9661 7774 9677 7788
rect 9712 7775 9734 7794
rect 9744 7788 9760 7789
rect 9743 7786 9760 7788
rect 9744 7781 9760 7786
rect 9734 7774 9740 7775
rect 9743 7774 9772 7781
rect 9661 7773 9772 7774
rect 9661 7772 9778 7773
rect 9337 7764 9388 7772
rect 9435 7764 9469 7772
rect 9337 7752 9362 7764
rect 9369 7752 9388 7764
rect 9442 7762 9469 7764
rect 9478 7762 9699 7772
rect 9734 7769 9740 7772
rect 9442 7758 9699 7762
rect 9337 7744 9388 7752
rect 9435 7744 9699 7758
rect 9743 7764 9778 7772
rect 9289 7696 9308 7730
rect 9353 7736 9382 7744
rect 9353 7730 9370 7736
rect 9353 7728 9387 7730
rect 9435 7728 9451 7744
rect 9452 7734 9660 7744
rect 9661 7734 9677 7744
rect 9725 7740 9740 7755
rect 9743 7752 9744 7764
rect 9751 7752 9778 7764
rect 9743 7744 9778 7752
rect 9743 7743 9772 7744
rect 9463 7730 9677 7734
rect 9478 7728 9677 7730
rect 9712 7730 9725 7740
rect 9743 7730 9760 7743
rect 9712 7728 9760 7730
rect 9354 7724 9387 7728
rect 9350 7722 9387 7724
rect 9350 7721 9417 7722
rect 9350 7716 9381 7721
rect 9387 7716 9417 7721
rect 9350 7712 9417 7716
rect 9323 7709 9417 7712
rect 9323 7702 9372 7709
rect 9323 7696 9353 7702
rect 9372 7697 9377 7702
rect 9289 7680 9369 7696
rect 9381 7688 9417 7709
rect 9478 7704 9667 7728
rect 9712 7727 9759 7728
rect 9725 7722 9759 7727
rect 9493 7701 9667 7704
rect 9486 7698 9667 7701
rect 9695 7721 9759 7722
rect 9289 7678 9308 7680
rect 9323 7678 9357 7680
rect 9289 7662 9369 7678
rect 9289 7656 9308 7662
rect 9005 7630 9108 7640
rect 8959 7628 9108 7630
rect 9129 7628 9164 7640
rect 8798 7626 8960 7628
rect 8810 7606 8829 7626
rect 8844 7624 8874 7626
rect 8693 7598 8734 7606
rect 8816 7602 8829 7606
rect 8881 7610 8960 7626
rect 8992 7626 9164 7628
rect 8992 7610 9071 7626
rect 9078 7624 9108 7626
rect 8656 7588 8685 7598
rect 8699 7588 8728 7598
rect 8743 7588 8773 7602
rect 8816 7588 8859 7602
rect 8881 7598 9071 7610
rect 9136 7606 9142 7626
rect 8866 7588 8896 7598
rect 8897 7588 9055 7598
rect 9059 7588 9089 7598
rect 9093 7588 9123 7602
rect 9151 7588 9164 7626
rect 9236 7640 9265 7656
rect 9279 7640 9308 7656
rect 9323 7646 9353 7662
rect 9381 7640 9387 7688
rect 9390 7682 9409 7688
rect 9424 7682 9454 7690
rect 9390 7674 9454 7682
rect 9390 7658 9470 7674
rect 9486 7667 9548 7698
rect 9564 7667 9626 7698
rect 9695 7696 9744 7721
rect 9759 7696 9789 7712
rect 9658 7682 9688 7690
rect 9695 7688 9805 7696
rect 9658 7674 9703 7682
rect 9390 7656 9409 7658
rect 9424 7656 9470 7658
rect 9390 7640 9470 7656
rect 9497 7654 9532 7667
rect 9573 7664 9610 7667
rect 9573 7662 9615 7664
rect 9502 7651 9532 7654
rect 9511 7647 9518 7651
rect 9518 7646 9519 7647
rect 9477 7640 9487 7646
rect 9236 7632 9271 7640
rect 9236 7606 9237 7632
rect 9244 7606 9271 7632
rect 9179 7588 9209 7602
rect 9236 7598 9271 7606
rect 9273 7632 9314 7640
rect 9273 7606 9288 7632
rect 9295 7606 9314 7632
rect 9378 7628 9409 7640
rect 9424 7628 9527 7640
rect 9539 7630 9565 7656
rect 9580 7651 9610 7662
rect 9642 7658 9704 7674
rect 9642 7656 9688 7658
rect 9642 7640 9704 7656
rect 9716 7640 9722 7688
rect 9725 7680 9805 7688
rect 9725 7678 9744 7680
rect 9759 7678 9793 7680
rect 9725 7662 9805 7678
rect 9725 7640 9744 7662
rect 9759 7646 9789 7662
rect 9817 7656 9823 7730
rect 9826 7656 9845 7800
rect 9860 7656 9866 7800
rect 9875 7730 9888 7800
rect 9940 7796 9962 7800
rect 9933 7774 9962 7788
rect 10015 7774 10031 7788
rect 10069 7784 10075 7786
rect 10082 7784 10190 7800
rect 10197 7784 10203 7786
rect 10211 7784 10226 7800
rect 10292 7794 10311 7797
rect 9933 7772 10031 7774
rect 10058 7772 10226 7784
rect 10241 7774 10257 7788
rect 10292 7775 10314 7794
rect 10324 7788 10340 7789
rect 10323 7786 10340 7788
rect 10324 7781 10340 7786
rect 10314 7774 10320 7775
rect 10323 7774 10352 7781
rect 10241 7773 10352 7774
rect 10241 7772 10358 7773
rect 9917 7764 9968 7772
rect 10015 7764 10049 7772
rect 9917 7752 9942 7764
rect 9949 7752 9968 7764
rect 10022 7762 10049 7764
rect 10058 7762 10279 7772
rect 10314 7769 10320 7772
rect 10022 7758 10279 7762
rect 9917 7744 9968 7752
rect 10015 7744 10279 7758
rect 10323 7764 10358 7772
rect 9869 7696 9888 7730
rect 9933 7736 9962 7744
rect 9933 7730 9950 7736
rect 9933 7728 9967 7730
rect 10015 7728 10031 7744
rect 10032 7734 10240 7744
rect 10241 7734 10257 7744
rect 10305 7740 10320 7755
rect 10323 7752 10324 7764
rect 10331 7752 10358 7764
rect 10323 7744 10358 7752
rect 10323 7743 10352 7744
rect 10043 7730 10257 7734
rect 10058 7728 10257 7730
rect 10292 7730 10305 7740
rect 10323 7730 10340 7743
rect 10292 7728 10340 7730
rect 9934 7724 9967 7728
rect 9930 7722 9967 7724
rect 9930 7721 9997 7722
rect 9930 7716 9961 7721
rect 9967 7716 9997 7721
rect 9930 7712 9997 7716
rect 9903 7709 9997 7712
rect 9903 7702 9952 7709
rect 9903 7696 9933 7702
rect 9952 7697 9957 7702
rect 9869 7680 9949 7696
rect 9961 7688 9997 7709
rect 10058 7704 10247 7728
rect 10292 7727 10339 7728
rect 10305 7722 10339 7727
rect 10073 7701 10247 7704
rect 10066 7698 10247 7701
rect 10275 7721 10339 7722
rect 9869 7678 9888 7680
rect 9903 7678 9937 7680
rect 9869 7662 9949 7678
rect 9869 7656 9888 7662
rect 9585 7630 9688 7640
rect 9539 7628 9688 7630
rect 9709 7628 9744 7640
rect 9378 7626 9540 7628
rect 9390 7606 9409 7626
rect 9424 7624 9454 7626
rect 9273 7598 9314 7606
rect 9396 7602 9409 7606
rect 9461 7610 9540 7626
rect 9572 7626 9744 7628
rect 9572 7610 9651 7626
rect 9658 7624 9688 7626
rect 9236 7588 9265 7598
rect 9279 7588 9308 7598
rect 9323 7588 9353 7602
rect 9396 7588 9439 7602
rect 9461 7598 9651 7610
rect 9716 7606 9722 7626
rect 9446 7588 9476 7598
rect 9477 7588 9635 7598
rect 9639 7588 9669 7598
rect 9673 7588 9703 7602
rect 9731 7588 9744 7626
rect 9816 7640 9845 7656
rect 9859 7640 9888 7656
rect 9903 7646 9933 7662
rect 9961 7640 9967 7688
rect 9970 7682 9989 7688
rect 10004 7682 10034 7690
rect 9970 7674 10034 7682
rect 9970 7658 10050 7674
rect 10066 7667 10128 7698
rect 10144 7667 10206 7698
rect 10275 7696 10324 7721
rect 10339 7696 10369 7712
rect 10238 7682 10268 7690
rect 10275 7688 10385 7696
rect 10238 7674 10283 7682
rect 9970 7656 9989 7658
rect 10004 7656 10050 7658
rect 9970 7640 10050 7656
rect 10077 7654 10112 7667
rect 10153 7664 10190 7667
rect 10153 7662 10195 7664
rect 10082 7651 10112 7654
rect 10091 7647 10098 7651
rect 10098 7646 10099 7647
rect 10057 7640 10067 7646
rect 9816 7632 9851 7640
rect 9816 7606 9817 7632
rect 9824 7606 9851 7632
rect 9759 7588 9789 7602
rect 9816 7598 9851 7606
rect 9853 7632 9894 7640
rect 9853 7606 9868 7632
rect 9875 7606 9894 7632
rect 9958 7628 9989 7640
rect 10004 7628 10107 7640
rect 10119 7630 10145 7656
rect 10160 7651 10190 7662
rect 10222 7658 10284 7674
rect 10222 7656 10268 7658
rect 10222 7640 10284 7656
rect 10296 7640 10302 7688
rect 10305 7680 10385 7688
rect 10305 7678 10324 7680
rect 10339 7678 10373 7680
rect 10305 7662 10385 7678
rect 10305 7640 10324 7662
rect 10339 7646 10369 7662
rect 10397 7656 10403 7730
rect 10406 7656 10425 7800
rect 10440 7656 10446 7800
rect 10455 7730 10468 7800
rect 10520 7796 10542 7800
rect 10513 7774 10542 7788
rect 10595 7774 10611 7788
rect 10649 7784 10655 7786
rect 10662 7784 10770 7800
rect 10777 7784 10783 7786
rect 10791 7784 10806 7800
rect 10872 7794 10891 7797
rect 10513 7772 10611 7774
rect 10638 7772 10806 7784
rect 10821 7774 10837 7788
rect 10872 7775 10894 7794
rect 10904 7788 10920 7789
rect 10903 7786 10920 7788
rect 10904 7781 10920 7786
rect 10894 7774 10900 7775
rect 10903 7774 10932 7781
rect 10821 7773 10932 7774
rect 10821 7772 10938 7773
rect 10497 7764 10548 7772
rect 10595 7764 10629 7772
rect 10497 7752 10522 7764
rect 10529 7752 10548 7764
rect 10602 7762 10629 7764
rect 10638 7762 10859 7772
rect 10894 7769 10900 7772
rect 10602 7758 10859 7762
rect 10497 7744 10548 7752
rect 10595 7744 10859 7758
rect 10903 7764 10938 7772
rect 10449 7696 10468 7730
rect 10513 7736 10542 7744
rect 10513 7730 10530 7736
rect 10513 7728 10547 7730
rect 10595 7728 10611 7744
rect 10612 7734 10820 7744
rect 10821 7734 10837 7744
rect 10885 7740 10900 7755
rect 10903 7752 10904 7764
rect 10911 7752 10938 7764
rect 10903 7744 10938 7752
rect 10903 7743 10932 7744
rect 10623 7730 10837 7734
rect 10638 7728 10837 7730
rect 10872 7730 10885 7740
rect 10903 7730 10920 7743
rect 10872 7728 10920 7730
rect 10514 7724 10547 7728
rect 10510 7722 10547 7724
rect 10510 7721 10577 7722
rect 10510 7716 10541 7721
rect 10547 7716 10577 7721
rect 10510 7712 10577 7716
rect 10483 7709 10577 7712
rect 10483 7702 10532 7709
rect 10483 7696 10513 7702
rect 10532 7697 10537 7702
rect 10449 7680 10529 7696
rect 10541 7688 10577 7709
rect 10638 7704 10827 7728
rect 10872 7727 10919 7728
rect 10885 7722 10919 7727
rect 10653 7701 10827 7704
rect 10646 7698 10827 7701
rect 10855 7721 10919 7722
rect 10449 7678 10468 7680
rect 10483 7678 10517 7680
rect 10449 7662 10529 7678
rect 10449 7656 10468 7662
rect 10165 7630 10268 7640
rect 10119 7628 10268 7630
rect 10289 7628 10324 7640
rect 9958 7626 10120 7628
rect 9970 7606 9989 7626
rect 10004 7624 10034 7626
rect 9853 7598 9894 7606
rect 9976 7602 9989 7606
rect 10041 7610 10120 7626
rect 10152 7626 10324 7628
rect 10152 7610 10231 7626
rect 10238 7624 10268 7626
rect 9816 7588 9845 7598
rect 9859 7588 9888 7598
rect 9903 7588 9933 7602
rect 9976 7588 10019 7602
rect 10041 7598 10231 7610
rect 10296 7606 10302 7626
rect 10026 7588 10056 7598
rect 10057 7588 10215 7598
rect 10219 7588 10249 7598
rect 10253 7588 10283 7602
rect 10311 7588 10324 7626
rect 10396 7640 10425 7656
rect 10439 7640 10468 7656
rect 10483 7646 10513 7662
rect 10541 7640 10547 7688
rect 10550 7682 10569 7688
rect 10584 7682 10614 7690
rect 10550 7674 10614 7682
rect 10550 7658 10630 7674
rect 10646 7667 10708 7698
rect 10724 7667 10786 7698
rect 10855 7696 10904 7721
rect 10919 7696 10949 7712
rect 10818 7682 10848 7690
rect 10855 7688 10965 7696
rect 10818 7674 10863 7682
rect 10550 7656 10569 7658
rect 10584 7656 10630 7658
rect 10550 7640 10630 7656
rect 10657 7654 10692 7667
rect 10733 7664 10770 7667
rect 10733 7662 10775 7664
rect 10662 7651 10692 7654
rect 10671 7647 10678 7651
rect 10678 7646 10679 7647
rect 10637 7640 10647 7646
rect 10396 7632 10431 7640
rect 10396 7606 10397 7632
rect 10404 7606 10431 7632
rect 10339 7588 10369 7602
rect 10396 7598 10431 7606
rect 10433 7632 10474 7640
rect 10433 7606 10448 7632
rect 10455 7606 10474 7632
rect 10538 7628 10569 7640
rect 10584 7628 10687 7640
rect 10699 7630 10725 7656
rect 10740 7651 10770 7662
rect 10802 7658 10864 7674
rect 10802 7656 10848 7658
rect 10802 7640 10864 7656
rect 10876 7640 10882 7688
rect 10885 7680 10965 7688
rect 10885 7678 10904 7680
rect 10919 7678 10953 7680
rect 10885 7662 10965 7678
rect 10885 7640 10904 7662
rect 10919 7646 10949 7662
rect 10977 7656 10983 7730
rect 10986 7656 11005 7800
rect 11020 7656 11026 7800
rect 11035 7730 11048 7800
rect 11100 7796 11122 7800
rect 11093 7774 11122 7788
rect 11175 7774 11191 7788
rect 11229 7784 11235 7786
rect 11242 7784 11350 7800
rect 11357 7784 11363 7786
rect 11371 7784 11386 7800
rect 11452 7794 11471 7797
rect 11093 7772 11191 7774
rect 11218 7772 11386 7784
rect 11401 7774 11417 7788
rect 11452 7775 11474 7794
rect 11484 7788 11500 7789
rect 11483 7786 11500 7788
rect 11484 7781 11500 7786
rect 11474 7774 11480 7775
rect 11483 7774 11512 7781
rect 11401 7773 11512 7774
rect 11401 7772 11518 7773
rect 11077 7764 11128 7772
rect 11175 7764 11209 7772
rect 11077 7752 11102 7764
rect 11109 7752 11128 7764
rect 11182 7762 11209 7764
rect 11218 7762 11439 7772
rect 11474 7769 11480 7772
rect 11182 7758 11439 7762
rect 11077 7744 11128 7752
rect 11175 7744 11439 7758
rect 11483 7764 11518 7772
rect 11029 7696 11048 7730
rect 11093 7736 11122 7744
rect 11093 7730 11110 7736
rect 11093 7728 11127 7730
rect 11175 7728 11191 7744
rect 11192 7734 11400 7744
rect 11401 7734 11417 7744
rect 11465 7740 11480 7755
rect 11483 7752 11484 7764
rect 11491 7752 11518 7764
rect 11483 7744 11518 7752
rect 11483 7743 11512 7744
rect 11203 7730 11417 7734
rect 11218 7728 11417 7730
rect 11452 7730 11465 7740
rect 11483 7730 11500 7743
rect 11452 7728 11500 7730
rect 11094 7724 11127 7728
rect 11090 7722 11127 7724
rect 11090 7721 11157 7722
rect 11090 7716 11121 7721
rect 11127 7716 11157 7721
rect 11090 7712 11157 7716
rect 11063 7709 11157 7712
rect 11063 7702 11112 7709
rect 11063 7696 11093 7702
rect 11112 7697 11117 7702
rect 11029 7680 11109 7696
rect 11121 7688 11157 7709
rect 11218 7704 11407 7728
rect 11452 7727 11499 7728
rect 11465 7722 11499 7727
rect 11233 7701 11407 7704
rect 11226 7698 11407 7701
rect 11435 7721 11499 7722
rect 11029 7678 11048 7680
rect 11063 7678 11097 7680
rect 11029 7662 11109 7678
rect 11029 7656 11048 7662
rect 10745 7630 10848 7640
rect 10699 7628 10848 7630
rect 10869 7628 10904 7640
rect 10538 7626 10700 7628
rect 10550 7606 10569 7626
rect 10584 7624 10614 7626
rect 10433 7598 10474 7606
rect 10556 7602 10569 7606
rect 10621 7610 10700 7626
rect 10732 7626 10904 7628
rect 10732 7610 10811 7626
rect 10818 7624 10848 7626
rect 10396 7588 10425 7598
rect 10439 7588 10468 7598
rect 10483 7588 10513 7602
rect 10556 7588 10599 7602
rect 10621 7598 10811 7610
rect 10876 7606 10882 7626
rect 10606 7588 10636 7598
rect 10637 7588 10795 7598
rect 10799 7588 10829 7598
rect 10833 7588 10863 7602
rect 10891 7588 10904 7626
rect 10976 7640 11005 7656
rect 11019 7640 11048 7656
rect 11063 7646 11093 7662
rect 11121 7640 11127 7688
rect 11130 7682 11149 7688
rect 11164 7682 11194 7690
rect 11130 7674 11194 7682
rect 11130 7658 11210 7674
rect 11226 7667 11288 7698
rect 11304 7667 11366 7698
rect 11435 7696 11484 7721
rect 11499 7696 11529 7712
rect 11398 7682 11428 7690
rect 11435 7688 11545 7696
rect 11398 7674 11443 7682
rect 11130 7656 11149 7658
rect 11164 7656 11210 7658
rect 11130 7640 11210 7656
rect 11237 7654 11272 7667
rect 11313 7664 11350 7667
rect 11313 7662 11355 7664
rect 11242 7651 11272 7654
rect 11251 7647 11258 7651
rect 11258 7646 11259 7647
rect 11217 7640 11227 7646
rect 10976 7632 11011 7640
rect 10976 7606 10977 7632
rect 10984 7606 11011 7632
rect 10919 7588 10949 7602
rect 10976 7598 11011 7606
rect 11013 7632 11054 7640
rect 11013 7606 11028 7632
rect 11035 7606 11054 7632
rect 11118 7628 11149 7640
rect 11164 7628 11267 7640
rect 11279 7630 11305 7656
rect 11320 7651 11350 7662
rect 11382 7658 11444 7674
rect 11382 7656 11428 7658
rect 11382 7640 11444 7656
rect 11456 7640 11462 7688
rect 11465 7680 11545 7688
rect 11465 7678 11484 7680
rect 11499 7678 11533 7680
rect 11465 7662 11545 7678
rect 11465 7640 11484 7662
rect 11499 7646 11529 7662
rect 11557 7656 11563 7730
rect 11566 7656 11585 7800
rect 11600 7656 11606 7800
rect 11615 7730 11628 7800
rect 11680 7796 11702 7800
rect 11673 7774 11702 7788
rect 11755 7774 11771 7788
rect 11809 7784 11815 7786
rect 11822 7784 11930 7800
rect 11937 7784 11943 7786
rect 11951 7784 11966 7800
rect 12032 7794 12051 7797
rect 11673 7772 11771 7774
rect 11798 7772 11966 7784
rect 11981 7774 11997 7788
rect 12032 7775 12054 7794
rect 12064 7788 12080 7789
rect 12063 7786 12080 7788
rect 12064 7781 12080 7786
rect 12054 7774 12060 7775
rect 12063 7774 12092 7781
rect 11981 7773 12092 7774
rect 11981 7772 12098 7773
rect 11657 7764 11708 7772
rect 11755 7764 11789 7772
rect 11657 7752 11682 7764
rect 11689 7752 11708 7764
rect 11762 7762 11789 7764
rect 11798 7762 12019 7772
rect 12054 7769 12060 7772
rect 11762 7758 12019 7762
rect 11657 7744 11708 7752
rect 11755 7744 12019 7758
rect 12063 7764 12098 7772
rect 11609 7696 11628 7730
rect 11673 7736 11702 7744
rect 11673 7730 11690 7736
rect 11673 7728 11707 7730
rect 11755 7728 11771 7744
rect 11772 7734 11980 7744
rect 11981 7734 11997 7744
rect 12045 7740 12060 7755
rect 12063 7752 12064 7764
rect 12071 7752 12098 7764
rect 12063 7744 12098 7752
rect 12063 7743 12092 7744
rect 11783 7730 11997 7734
rect 11798 7728 11997 7730
rect 12032 7730 12045 7740
rect 12063 7730 12080 7743
rect 12032 7728 12080 7730
rect 11674 7724 11707 7728
rect 11670 7722 11707 7724
rect 11670 7721 11737 7722
rect 11670 7716 11701 7721
rect 11707 7716 11737 7721
rect 11670 7712 11737 7716
rect 11643 7709 11737 7712
rect 11643 7702 11692 7709
rect 11643 7696 11673 7702
rect 11692 7697 11697 7702
rect 11609 7680 11689 7696
rect 11701 7688 11737 7709
rect 11798 7704 11987 7728
rect 12032 7727 12079 7728
rect 12045 7722 12079 7727
rect 11813 7701 11987 7704
rect 11806 7698 11987 7701
rect 12015 7721 12079 7722
rect 11609 7678 11628 7680
rect 11643 7678 11677 7680
rect 11609 7662 11689 7678
rect 11609 7656 11628 7662
rect 11325 7630 11428 7640
rect 11279 7628 11428 7630
rect 11449 7628 11484 7640
rect 11118 7626 11280 7628
rect 11130 7606 11149 7626
rect 11164 7624 11194 7626
rect 11013 7598 11054 7606
rect 11136 7602 11149 7606
rect 11201 7610 11280 7626
rect 11312 7626 11484 7628
rect 11312 7610 11391 7626
rect 11398 7624 11428 7626
rect 10976 7588 11005 7598
rect 11019 7588 11048 7598
rect 11063 7588 11093 7602
rect 11136 7588 11179 7602
rect 11201 7598 11391 7610
rect 11456 7606 11462 7626
rect 11186 7588 11216 7598
rect 11217 7588 11375 7598
rect 11379 7588 11409 7598
rect 11413 7588 11443 7602
rect 11471 7588 11484 7626
rect 11556 7640 11585 7656
rect 11599 7640 11628 7656
rect 11643 7646 11673 7662
rect 11701 7640 11707 7688
rect 11710 7682 11729 7688
rect 11744 7682 11774 7690
rect 11710 7674 11774 7682
rect 11710 7658 11790 7674
rect 11806 7667 11868 7698
rect 11884 7667 11946 7698
rect 12015 7696 12064 7721
rect 12079 7696 12109 7712
rect 11978 7682 12008 7690
rect 12015 7688 12125 7696
rect 11978 7674 12023 7682
rect 11710 7656 11729 7658
rect 11744 7656 11790 7658
rect 11710 7640 11790 7656
rect 11817 7654 11852 7667
rect 11893 7664 11930 7667
rect 11893 7662 11935 7664
rect 11822 7651 11852 7654
rect 11831 7647 11838 7651
rect 11838 7646 11839 7647
rect 11797 7640 11807 7646
rect 11556 7632 11591 7640
rect 11556 7606 11557 7632
rect 11564 7606 11591 7632
rect 11499 7588 11529 7602
rect 11556 7598 11591 7606
rect 11593 7632 11634 7640
rect 11593 7606 11608 7632
rect 11615 7606 11634 7632
rect 11698 7628 11729 7640
rect 11744 7628 11847 7640
rect 11859 7630 11885 7656
rect 11900 7651 11930 7662
rect 11962 7658 12024 7674
rect 11962 7656 12008 7658
rect 11962 7640 12024 7656
rect 12036 7640 12042 7688
rect 12045 7680 12125 7688
rect 12045 7678 12064 7680
rect 12079 7678 12113 7680
rect 12045 7662 12125 7678
rect 12045 7640 12064 7662
rect 12079 7646 12109 7662
rect 12137 7656 12143 7730
rect 12146 7656 12165 7800
rect 12180 7656 12186 7800
rect 12195 7730 12208 7800
rect 12260 7796 12282 7800
rect 12253 7774 12282 7788
rect 12335 7774 12351 7788
rect 12389 7784 12395 7786
rect 12402 7784 12510 7800
rect 12517 7784 12523 7786
rect 12531 7784 12546 7800
rect 12612 7794 12631 7797
rect 12253 7772 12351 7774
rect 12378 7772 12546 7784
rect 12561 7774 12577 7788
rect 12612 7775 12634 7794
rect 12644 7788 12660 7789
rect 12643 7786 12660 7788
rect 12644 7781 12660 7786
rect 12634 7774 12640 7775
rect 12643 7774 12672 7781
rect 12561 7773 12672 7774
rect 12561 7772 12678 7773
rect 12237 7764 12288 7772
rect 12335 7764 12369 7772
rect 12237 7752 12262 7764
rect 12269 7752 12288 7764
rect 12342 7762 12369 7764
rect 12378 7762 12599 7772
rect 12634 7769 12640 7772
rect 12342 7758 12599 7762
rect 12237 7744 12288 7752
rect 12335 7744 12599 7758
rect 12643 7764 12678 7772
rect 12189 7696 12208 7730
rect 12253 7736 12282 7744
rect 12253 7730 12270 7736
rect 12253 7728 12287 7730
rect 12335 7728 12351 7744
rect 12352 7734 12560 7744
rect 12561 7734 12577 7744
rect 12625 7740 12640 7755
rect 12643 7752 12644 7764
rect 12651 7752 12678 7764
rect 12643 7744 12678 7752
rect 12643 7743 12672 7744
rect 12363 7730 12577 7734
rect 12378 7728 12577 7730
rect 12612 7730 12625 7740
rect 12643 7730 12660 7743
rect 12612 7728 12660 7730
rect 12254 7724 12287 7728
rect 12250 7722 12287 7724
rect 12250 7721 12317 7722
rect 12250 7716 12281 7721
rect 12287 7716 12317 7721
rect 12250 7712 12317 7716
rect 12223 7709 12317 7712
rect 12223 7702 12272 7709
rect 12223 7696 12253 7702
rect 12272 7697 12277 7702
rect 12189 7680 12269 7696
rect 12281 7688 12317 7709
rect 12378 7704 12567 7728
rect 12612 7727 12659 7728
rect 12625 7722 12659 7727
rect 12393 7701 12567 7704
rect 12386 7698 12567 7701
rect 12595 7721 12659 7722
rect 12189 7678 12208 7680
rect 12223 7678 12257 7680
rect 12189 7662 12269 7678
rect 12189 7656 12208 7662
rect 11905 7630 12008 7640
rect 11859 7628 12008 7630
rect 12029 7628 12064 7640
rect 11698 7626 11860 7628
rect 11710 7606 11729 7626
rect 11744 7624 11774 7626
rect 11593 7598 11634 7606
rect 11716 7602 11729 7606
rect 11781 7610 11860 7626
rect 11892 7626 12064 7628
rect 11892 7610 11971 7626
rect 11978 7624 12008 7626
rect 11556 7588 11585 7598
rect 11599 7588 11628 7598
rect 11643 7588 11673 7602
rect 11716 7588 11759 7602
rect 11781 7598 11971 7610
rect 12036 7606 12042 7626
rect 11766 7588 11796 7598
rect 11797 7588 11955 7598
rect 11959 7588 11989 7598
rect 11993 7588 12023 7602
rect 12051 7588 12064 7626
rect 12136 7640 12165 7656
rect 12179 7640 12208 7656
rect 12223 7646 12253 7662
rect 12281 7640 12287 7688
rect 12290 7682 12309 7688
rect 12324 7682 12354 7690
rect 12290 7674 12354 7682
rect 12290 7658 12370 7674
rect 12386 7667 12448 7698
rect 12464 7667 12526 7698
rect 12595 7696 12644 7721
rect 12659 7696 12689 7712
rect 12558 7682 12588 7690
rect 12595 7688 12705 7696
rect 12558 7674 12603 7682
rect 12290 7656 12309 7658
rect 12324 7656 12370 7658
rect 12290 7640 12370 7656
rect 12397 7654 12432 7667
rect 12473 7664 12510 7667
rect 12473 7662 12515 7664
rect 12402 7651 12432 7654
rect 12411 7647 12418 7651
rect 12418 7646 12419 7647
rect 12377 7640 12387 7646
rect 12136 7632 12171 7640
rect 12136 7606 12137 7632
rect 12144 7606 12171 7632
rect 12079 7588 12109 7602
rect 12136 7598 12171 7606
rect 12173 7632 12214 7640
rect 12173 7606 12188 7632
rect 12195 7606 12214 7632
rect 12278 7628 12309 7640
rect 12324 7628 12427 7640
rect 12439 7630 12465 7656
rect 12480 7651 12510 7662
rect 12542 7658 12604 7674
rect 12542 7656 12588 7658
rect 12542 7640 12604 7656
rect 12616 7640 12622 7688
rect 12625 7680 12705 7688
rect 12625 7678 12644 7680
rect 12659 7678 12693 7680
rect 12625 7662 12705 7678
rect 12625 7640 12644 7662
rect 12659 7646 12689 7662
rect 12717 7656 12723 7730
rect 12726 7656 12745 7800
rect 12760 7656 12766 7800
rect 12775 7730 12788 7800
rect 12840 7796 12862 7800
rect 12833 7774 12862 7788
rect 12915 7774 12931 7788
rect 12969 7784 12975 7786
rect 12982 7784 13090 7800
rect 13097 7784 13103 7786
rect 13111 7784 13126 7800
rect 13192 7794 13211 7797
rect 12833 7772 12931 7774
rect 12958 7772 13126 7784
rect 13141 7774 13157 7788
rect 13192 7775 13214 7794
rect 13224 7788 13240 7789
rect 13223 7786 13240 7788
rect 13224 7781 13240 7786
rect 13214 7774 13220 7775
rect 13223 7774 13252 7781
rect 13141 7773 13252 7774
rect 13141 7772 13258 7773
rect 12817 7764 12868 7772
rect 12915 7764 12949 7772
rect 12817 7752 12842 7764
rect 12849 7752 12868 7764
rect 12922 7762 12949 7764
rect 12958 7762 13179 7772
rect 13214 7769 13220 7772
rect 12922 7758 13179 7762
rect 12817 7744 12868 7752
rect 12915 7744 13179 7758
rect 13223 7764 13258 7772
rect 12769 7696 12788 7730
rect 12833 7736 12862 7744
rect 12833 7730 12850 7736
rect 12833 7728 12867 7730
rect 12915 7728 12931 7744
rect 12932 7734 13140 7744
rect 13141 7734 13157 7744
rect 13205 7740 13220 7755
rect 13223 7752 13224 7764
rect 13231 7752 13258 7764
rect 13223 7744 13258 7752
rect 13223 7743 13252 7744
rect 12943 7730 13157 7734
rect 12958 7728 13157 7730
rect 13192 7730 13205 7740
rect 13223 7730 13240 7743
rect 13192 7728 13240 7730
rect 12834 7724 12867 7728
rect 12830 7722 12867 7724
rect 12830 7721 12897 7722
rect 12830 7716 12861 7721
rect 12867 7716 12897 7721
rect 12830 7712 12897 7716
rect 12803 7709 12897 7712
rect 12803 7702 12852 7709
rect 12803 7696 12833 7702
rect 12852 7697 12857 7702
rect 12769 7680 12849 7696
rect 12861 7688 12897 7709
rect 12958 7704 13147 7728
rect 13192 7727 13239 7728
rect 13205 7722 13239 7727
rect 12973 7701 13147 7704
rect 12966 7698 13147 7701
rect 13175 7721 13239 7722
rect 12769 7678 12788 7680
rect 12803 7678 12837 7680
rect 12769 7662 12849 7678
rect 12769 7656 12788 7662
rect 12485 7630 12588 7640
rect 12439 7628 12588 7630
rect 12609 7628 12644 7640
rect 12278 7626 12440 7628
rect 12290 7606 12309 7626
rect 12324 7624 12354 7626
rect 12173 7598 12214 7606
rect 12296 7602 12309 7606
rect 12361 7610 12440 7626
rect 12472 7626 12644 7628
rect 12472 7610 12551 7626
rect 12558 7624 12588 7626
rect 12136 7588 12165 7598
rect 12179 7588 12208 7598
rect 12223 7588 12253 7602
rect 12296 7588 12339 7602
rect 12361 7598 12551 7610
rect 12616 7606 12622 7626
rect 12346 7588 12376 7598
rect 12377 7588 12535 7598
rect 12539 7588 12569 7598
rect 12573 7588 12603 7602
rect 12631 7588 12644 7626
rect 12716 7640 12745 7656
rect 12759 7640 12788 7656
rect 12803 7646 12833 7662
rect 12861 7640 12867 7688
rect 12870 7682 12889 7688
rect 12904 7682 12934 7690
rect 12870 7674 12934 7682
rect 12870 7658 12950 7674
rect 12966 7667 13028 7698
rect 13044 7667 13106 7698
rect 13175 7696 13224 7721
rect 13239 7696 13269 7712
rect 13138 7682 13168 7690
rect 13175 7688 13285 7696
rect 13138 7674 13183 7682
rect 12870 7656 12889 7658
rect 12904 7656 12950 7658
rect 12870 7640 12950 7656
rect 12977 7654 13012 7667
rect 13053 7664 13090 7667
rect 13053 7662 13095 7664
rect 12982 7651 13012 7654
rect 12991 7647 12998 7651
rect 12998 7646 12999 7647
rect 12957 7640 12967 7646
rect 12716 7632 12751 7640
rect 12716 7606 12717 7632
rect 12724 7606 12751 7632
rect 12659 7588 12689 7602
rect 12716 7598 12751 7606
rect 12753 7632 12794 7640
rect 12753 7606 12768 7632
rect 12775 7606 12794 7632
rect 12858 7628 12889 7640
rect 12904 7628 13007 7640
rect 13019 7630 13045 7656
rect 13060 7651 13090 7662
rect 13122 7658 13184 7674
rect 13122 7656 13168 7658
rect 13122 7640 13184 7656
rect 13196 7640 13202 7688
rect 13205 7680 13285 7688
rect 13205 7678 13224 7680
rect 13239 7678 13273 7680
rect 13205 7662 13285 7678
rect 13205 7640 13224 7662
rect 13239 7646 13269 7662
rect 13297 7656 13303 7730
rect 13306 7656 13325 7800
rect 13340 7656 13346 7800
rect 13355 7730 13368 7800
rect 13420 7796 13442 7800
rect 13413 7774 13442 7788
rect 13495 7774 13511 7788
rect 13549 7784 13555 7786
rect 13562 7784 13670 7800
rect 13677 7784 13683 7786
rect 13691 7784 13706 7800
rect 13772 7794 13791 7797
rect 13413 7772 13511 7774
rect 13538 7772 13706 7784
rect 13721 7774 13737 7788
rect 13772 7775 13794 7794
rect 13804 7788 13820 7789
rect 13803 7786 13820 7788
rect 13804 7781 13820 7786
rect 13794 7774 13800 7775
rect 13803 7774 13832 7781
rect 13721 7773 13832 7774
rect 13721 7772 13838 7773
rect 13397 7764 13448 7772
rect 13495 7764 13529 7772
rect 13397 7752 13422 7764
rect 13429 7752 13448 7764
rect 13502 7762 13529 7764
rect 13538 7762 13759 7772
rect 13794 7769 13800 7772
rect 13502 7758 13759 7762
rect 13397 7744 13448 7752
rect 13495 7744 13759 7758
rect 13803 7764 13838 7772
rect 13349 7696 13368 7730
rect 13413 7736 13442 7744
rect 13413 7730 13430 7736
rect 13413 7728 13447 7730
rect 13495 7728 13511 7744
rect 13512 7734 13720 7744
rect 13721 7734 13737 7744
rect 13785 7740 13800 7755
rect 13803 7752 13804 7764
rect 13811 7752 13838 7764
rect 13803 7744 13838 7752
rect 13803 7743 13832 7744
rect 13523 7730 13737 7734
rect 13538 7728 13737 7730
rect 13772 7730 13785 7740
rect 13803 7730 13820 7743
rect 13772 7728 13820 7730
rect 13414 7724 13447 7728
rect 13410 7722 13447 7724
rect 13410 7721 13477 7722
rect 13410 7716 13441 7721
rect 13447 7716 13477 7721
rect 13410 7712 13477 7716
rect 13383 7709 13477 7712
rect 13383 7702 13432 7709
rect 13383 7696 13413 7702
rect 13432 7697 13437 7702
rect 13349 7680 13429 7696
rect 13441 7688 13477 7709
rect 13538 7704 13727 7728
rect 13772 7727 13819 7728
rect 13785 7722 13819 7727
rect 13553 7701 13727 7704
rect 13546 7698 13727 7701
rect 13755 7721 13819 7722
rect 13349 7678 13368 7680
rect 13383 7678 13417 7680
rect 13349 7662 13429 7678
rect 13349 7656 13368 7662
rect 13065 7630 13168 7640
rect 13019 7628 13168 7630
rect 13189 7628 13224 7640
rect 12858 7626 13020 7628
rect 12870 7606 12889 7626
rect 12904 7624 12934 7626
rect 12753 7598 12794 7606
rect 12876 7602 12889 7606
rect 12941 7610 13020 7626
rect 13052 7626 13224 7628
rect 13052 7610 13131 7626
rect 13138 7624 13168 7626
rect 12716 7588 12745 7598
rect 12759 7588 12788 7598
rect 12803 7588 12833 7602
rect 12876 7588 12919 7602
rect 12941 7598 13131 7610
rect 13196 7606 13202 7626
rect 12926 7588 12956 7598
rect 12957 7588 13115 7598
rect 13119 7588 13149 7598
rect 13153 7588 13183 7602
rect 13211 7588 13224 7626
rect 13296 7640 13325 7656
rect 13339 7640 13368 7656
rect 13383 7646 13413 7662
rect 13441 7640 13447 7688
rect 13450 7682 13469 7688
rect 13484 7682 13514 7690
rect 13450 7674 13514 7682
rect 13450 7658 13530 7674
rect 13546 7667 13608 7698
rect 13624 7667 13686 7698
rect 13755 7696 13804 7721
rect 13819 7696 13849 7712
rect 13718 7682 13748 7690
rect 13755 7688 13865 7696
rect 13718 7674 13763 7682
rect 13450 7656 13469 7658
rect 13484 7656 13530 7658
rect 13450 7640 13530 7656
rect 13557 7654 13592 7667
rect 13633 7664 13670 7667
rect 13633 7662 13675 7664
rect 13562 7651 13592 7654
rect 13571 7647 13578 7651
rect 13578 7646 13579 7647
rect 13537 7640 13547 7646
rect 13296 7632 13331 7640
rect 13296 7606 13297 7632
rect 13304 7606 13331 7632
rect 13239 7588 13269 7602
rect 13296 7598 13331 7606
rect 13333 7632 13374 7640
rect 13333 7606 13348 7632
rect 13355 7606 13374 7632
rect 13438 7628 13469 7640
rect 13484 7628 13587 7640
rect 13599 7630 13625 7656
rect 13640 7651 13670 7662
rect 13702 7658 13764 7674
rect 13702 7656 13748 7658
rect 13702 7640 13764 7656
rect 13776 7640 13782 7688
rect 13785 7680 13865 7688
rect 13785 7678 13804 7680
rect 13819 7678 13853 7680
rect 13785 7662 13865 7678
rect 13785 7640 13804 7662
rect 13819 7646 13849 7662
rect 13877 7656 13883 7730
rect 13886 7656 13905 7800
rect 13920 7656 13926 7800
rect 13935 7730 13948 7800
rect 14000 7796 14022 7800
rect 13993 7774 14022 7788
rect 14075 7774 14091 7788
rect 14129 7784 14135 7786
rect 14142 7784 14250 7800
rect 14257 7784 14263 7786
rect 14271 7784 14286 7800
rect 14352 7794 14371 7797
rect 13993 7772 14091 7774
rect 14118 7772 14286 7784
rect 14301 7774 14317 7788
rect 14352 7775 14374 7794
rect 14384 7788 14400 7789
rect 14383 7786 14400 7788
rect 14384 7781 14400 7786
rect 14374 7774 14380 7775
rect 14383 7774 14412 7781
rect 14301 7773 14412 7774
rect 14301 7772 14418 7773
rect 13977 7764 14028 7772
rect 14075 7764 14109 7772
rect 13977 7752 14002 7764
rect 14009 7752 14028 7764
rect 14082 7762 14109 7764
rect 14118 7762 14339 7772
rect 14374 7769 14380 7772
rect 14082 7758 14339 7762
rect 13977 7744 14028 7752
rect 14075 7744 14339 7758
rect 14383 7764 14418 7772
rect 13929 7696 13948 7730
rect 13993 7736 14022 7744
rect 13993 7730 14010 7736
rect 13993 7728 14027 7730
rect 14075 7728 14091 7744
rect 14092 7734 14300 7744
rect 14301 7734 14317 7744
rect 14365 7740 14380 7755
rect 14383 7752 14384 7764
rect 14391 7752 14418 7764
rect 14383 7744 14418 7752
rect 14383 7743 14412 7744
rect 14103 7730 14317 7734
rect 14118 7728 14317 7730
rect 14352 7730 14365 7740
rect 14383 7730 14400 7743
rect 14352 7728 14400 7730
rect 13994 7724 14027 7728
rect 13990 7722 14027 7724
rect 13990 7721 14057 7722
rect 13990 7716 14021 7721
rect 14027 7716 14057 7721
rect 13990 7712 14057 7716
rect 13963 7709 14057 7712
rect 13963 7702 14012 7709
rect 13963 7696 13993 7702
rect 14012 7697 14017 7702
rect 13929 7680 14009 7696
rect 14021 7688 14057 7709
rect 14118 7704 14307 7728
rect 14352 7727 14399 7728
rect 14365 7722 14399 7727
rect 14133 7701 14307 7704
rect 14126 7698 14307 7701
rect 14335 7721 14399 7722
rect 13929 7678 13948 7680
rect 13963 7678 13997 7680
rect 13929 7662 14009 7678
rect 13929 7656 13948 7662
rect 13645 7630 13748 7640
rect 13599 7628 13748 7630
rect 13769 7628 13804 7640
rect 13438 7626 13600 7628
rect 13450 7606 13469 7626
rect 13484 7624 13514 7626
rect 13333 7598 13374 7606
rect 13456 7602 13469 7606
rect 13521 7610 13600 7626
rect 13632 7626 13804 7628
rect 13632 7610 13711 7626
rect 13718 7624 13748 7626
rect 13296 7588 13325 7598
rect 13339 7588 13368 7598
rect 13383 7588 13413 7602
rect 13456 7588 13499 7602
rect 13521 7598 13711 7610
rect 13776 7606 13782 7626
rect 13506 7588 13536 7598
rect 13537 7588 13695 7598
rect 13699 7588 13729 7598
rect 13733 7588 13763 7602
rect 13791 7588 13804 7626
rect 13876 7640 13905 7656
rect 13919 7640 13948 7656
rect 13963 7646 13993 7662
rect 14021 7640 14027 7688
rect 14030 7682 14049 7688
rect 14064 7682 14094 7690
rect 14030 7674 14094 7682
rect 14030 7658 14110 7674
rect 14126 7667 14188 7698
rect 14204 7667 14266 7698
rect 14335 7696 14384 7721
rect 14399 7696 14429 7712
rect 14298 7682 14328 7690
rect 14335 7688 14445 7696
rect 14298 7674 14343 7682
rect 14030 7656 14049 7658
rect 14064 7656 14110 7658
rect 14030 7640 14110 7656
rect 14137 7654 14172 7667
rect 14213 7664 14250 7667
rect 14213 7662 14255 7664
rect 14142 7651 14172 7654
rect 14151 7647 14158 7651
rect 14158 7646 14159 7647
rect 14117 7640 14127 7646
rect 13876 7632 13911 7640
rect 13876 7606 13877 7632
rect 13884 7606 13911 7632
rect 13819 7588 13849 7602
rect 13876 7598 13911 7606
rect 13913 7632 13954 7640
rect 13913 7606 13928 7632
rect 13935 7606 13954 7632
rect 14018 7628 14049 7640
rect 14064 7628 14167 7640
rect 14179 7630 14205 7656
rect 14220 7651 14250 7662
rect 14282 7658 14344 7674
rect 14282 7656 14328 7658
rect 14282 7640 14344 7656
rect 14356 7640 14362 7688
rect 14365 7680 14445 7688
rect 14365 7678 14384 7680
rect 14399 7678 14433 7680
rect 14365 7662 14445 7678
rect 14365 7640 14384 7662
rect 14399 7646 14429 7662
rect 14457 7656 14463 7730
rect 14466 7656 14485 7800
rect 14500 7656 14506 7800
rect 14515 7730 14528 7800
rect 14580 7796 14602 7800
rect 14573 7774 14602 7788
rect 14655 7774 14671 7788
rect 14709 7784 14715 7786
rect 14722 7784 14830 7800
rect 14837 7784 14843 7786
rect 14851 7784 14866 7800
rect 14932 7794 14951 7797
rect 14573 7772 14671 7774
rect 14698 7772 14866 7784
rect 14881 7774 14897 7788
rect 14932 7775 14954 7794
rect 14964 7788 14980 7789
rect 14963 7786 14980 7788
rect 14964 7781 14980 7786
rect 14954 7774 14960 7775
rect 14963 7774 14992 7781
rect 14881 7773 14992 7774
rect 14881 7772 14998 7773
rect 14557 7764 14608 7772
rect 14655 7764 14689 7772
rect 14557 7752 14582 7764
rect 14589 7752 14608 7764
rect 14662 7762 14689 7764
rect 14698 7762 14919 7772
rect 14954 7769 14960 7772
rect 14662 7758 14919 7762
rect 14557 7744 14608 7752
rect 14655 7744 14919 7758
rect 14963 7764 14998 7772
rect 14509 7696 14528 7730
rect 14573 7736 14602 7744
rect 14573 7730 14590 7736
rect 14573 7728 14607 7730
rect 14655 7728 14671 7744
rect 14672 7734 14880 7744
rect 14881 7734 14897 7744
rect 14945 7740 14960 7755
rect 14963 7752 14964 7764
rect 14971 7752 14998 7764
rect 14963 7744 14998 7752
rect 14963 7743 14992 7744
rect 14683 7730 14897 7734
rect 14698 7728 14897 7730
rect 14932 7730 14945 7740
rect 14963 7730 14980 7743
rect 14932 7728 14980 7730
rect 14574 7724 14607 7728
rect 14570 7722 14607 7724
rect 14570 7721 14637 7722
rect 14570 7716 14601 7721
rect 14607 7716 14637 7721
rect 14570 7712 14637 7716
rect 14543 7709 14637 7712
rect 14543 7702 14592 7709
rect 14543 7696 14573 7702
rect 14592 7697 14597 7702
rect 14509 7680 14589 7696
rect 14601 7688 14637 7709
rect 14698 7704 14887 7728
rect 14932 7727 14979 7728
rect 14945 7722 14979 7727
rect 14713 7701 14887 7704
rect 14706 7698 14887 7701
rect 14915 7721 14979 7722
rect 14509 7678 14528 7680
rect 14543 7678 14577 7680
rect 14509 7662 14589 7678
rect 14509 7656 14528 7662
rect 14225 7630 14328 7640
rect 14179 7628 14328 7630
rect 14349 7628 14384 7640
rect 14018 7626 14180 7628
rect 14030 7606 14049 7626
rect 14064 7624 14094 7626
rect 13913 7598 13954 7606
rect 14036 7602 14049 7606
rect 14101 7610 14180 7626
rect 14212 7626 14384 7628
rect 14212 7610 14291 7626
rect 14298 7624 14328 7626
rect 13876 7588 13905 7598
rect 13919 7588 13948 7598
rect 13963 7588 13993 7602
rect 14036 7588 14079 7602
rect 14101 7598 14291 7610
rect 14356 7606 14362 7626
rect 14086 7588 14116 7598
rect 14117 7588 14275 7598
rect 14279 7588 14309 7598
rect 14313 7588 14343 7602
rect 14371 7588 14384 7626
rect 14456 7640 14485 7656
rect 14499 7640 14528 7656
rect 14543 7646 14573 7662
rect 14601 7640 14607 7688
rect 14610 7682 14629 7688
rect 14644 7682 14674 7690
rect 14610 7674 14674 7682
rect 14610 7658 14690 7674
rect 14706 7667 14768 7698
rect 14784 7667 14846 7698
rect 14915 7696 14964 7721
rect 14979 7696 15009 7712
rect 14878 7682 14908 7690
rect 14915 7688 15025 7696
rect 14878 7674 14923 7682
rect 14610 7656 14629 7658
rect 14644 7656 14690 7658
rect 14610 7640 14690 7656
rect 14717 7654 14752 7667
rect 14793 7664 14830 7667
rect 14793 7662 14835 7664
rect 14722 7651 14752 7654
rect 14731 7647 14738 7651
rect 14738 7646 14739 7647
rect 14697 7640 14707 7646
rect 14456 7632 14491 7640
rect 14456 7606 14457 7632
rect 14464 7606 14491 7632
rect 14399 7588 14429 7602
rect 14456 7598 14491 7606
rect 14493 7632 14534 7640
rect 14493 7606 14508 7632
rect 14515 7606 14534 7632
rect 14598 7628 14629 7640
rect 14644 7628 14747 7640
rect 14759 7630 14785 7656
rect 14800 7651 14830 7662
rect 14862 7658 14924 7674
rect 14862 7656 14908 7658
rect 14862 7640 14924 7656
rect 14936 7640 14942 7688
rect 14945 7680 15025 7688
rect 14945 7678 14964 7680
rect 14979 7678 15013 7680
rect 14945 7662 15025 7678
rect 14945 7640 14964 7662
rect 14979 7646 15009 7662
rect 15037 7656 15043 7730
rect 15046 7656 15065 7800
rect 15080 7656 15086 7800
rect 15095 7730 15108 7800
rect 15160 7796 15182 7800
rect 15153 7774 15182 7788
rect 15235 7774 15251 7788
rect 15289 7784 15295 7786
rect 15302 7784 15410 7800
rect 15417 7784 15423 7786
rect 15431 7784 15446 7800
rect 15512 7794 15531 7797
rect 15153 7772 15251 7774
rect 15278 7772 15446 7784
rect 15461 7774 15477 7788
rect 15512 7775 15534 7794
rect 15544 7788 15560 7789
rect 15543 7786 15560 7788
rect 15544 7781 15560 7786
rect 15534 7774 15540 7775
rect 15543 7774 15572 7781
rect 15461 7773 15572 7774
rect 15461 7772 15578 7773
rect 15137 7764 15188 7772
rect 15235 7764 15269 7772
rect 15137 7752 15162 7764
rect 15169 7752 15188 7764
rect 15242 7762 15269 7764
rect 15278 7762 15499 7772
rect 15534 7769 15540 7772
rect 15242 7758 15499 7762
rect 15137 7744 15188 7752
rect 15235 7744 15499 7758
rect 15543 7764 15578 7772
rect 15089 7696 15108 7730
rect 15153 7736 15182 7744
rect 15153 7730 15170 7736
rect 15153 7728 15187 7730
rect 15235 7728 15251 7744
rect 15252 7734 15460 7744
rect 15461 7734 15477 7744
rect 15525 7740 15540 7755
rect 15543 7752 15544 7764
rect 15551 7752 15578 7764
rect 15543 7744 15578 7752
rect 15543 7743 15572 7744
rect 15263 7730 15477 7734
rect 15278 7728 15477 7730
rect 15512 7730 15525 7740
rect 15543 7730 15560 7743
rect 15512 7728 15560 7730
rect 15154 7724 15187 7728
rect 15150 7722 15187 7724
rect 15150 7721 15217 7722
rect 15150 7716 15181 7721
rect 15187 7716 15217 7721
rect 15150 7712 15217 7716
rect 15123 7709 15217 7712
rect 15123 7702 15172 7709
rect 15123 7696 15153 7702
rect 15172 7697 15177 7702
rect 15089 7680 15169 7696
rect 15181 7688 15217 7709
rect 15278 7704 15467 7728
rect 15512 7727 15559 7728
rect 15525 7722 15559 7727
rect 15293 7701 15467 7704
rect 15286 7698 15467 7701
rect 15495 7721 15559 7722
rect 15089 7678 15108 7680
rect 15123 7678 15157 7680
rect 15089 7662 15169 7678
rect 15089 7656 15108 7662
rect 14805 7630 14908 7640
rect 14759 7628 14908 7630
rect 14929 7628 14964 7640
rect 14598 7626 14760 7628
rect 14610 7606 14629 7626
rect 14644 7624 14674 7626
rect 14493 7598 14534 7606
rect 14616 7602 14629 7606
rect 14681 7610 14760 7626
rect 14792 7626 14964 7628
rect 14792 7610 14871 7626
rect 14878 7624 14908 7626
rect 14456 7588 14485 7598
rect 14499 7588 14528 7598
rect 14543 7588 14573 7602
rect 14616 7588 14659 7602
rect 14681 7598 14871 7610
rect 14936 7606 14942 7626
rect 14666 7588 14696 7598
rect 14697 7588 14855 7598
rect 14859 7588 14889 7598
rect 14893 7588 14923 7602
rect 14951 7588 14964 7626
rect 15036 7640 15065 7656
rect 15079 7640 15108 7656
rect 15123 7646 15153 7662
rect 15181 7640 15187 7688
rect 15190 7682 15209 7688
rect 15224 7682 15254 7690
rect 15190 7674 15254 7682
rect 15190 7658 15270 7674
rect 15286 7667 15348 7698
rect 15364 7667 15426 7698
rect 15495 7696 15544 7721
rect 15559 7696 15589 7712
rect 15458 7682 15488 7690
rect 15495 7688 15605 7696
rect 15458 7674 15503 7682
rect 15190 7656 15209 7658
rect 15224 7656 15270 7658
rect 15190 7640 15270 7656
rect 15297 7654 15332 7667
rect 15373 7664 15410 7667
rect 15373 7662 15415 7664
rect 15302 7651 15332 7654
rect 15311 7647 15318 7651
rect 15318 7646 15319 7647
rect 15277 7640 15287 7646
rect 15036 7632 15071 7640
rect 15036 7606 15037 7632
rect 15044 7606 15071 7632
rect 14979 7588 15009 7602
rect 15036 7598 15071 7606
rect 15073 7632 15114 7640
rect 15073 7606 15088 7632
rect 15095 7606 15114 7632
rect 15178 7628 15209 7640
rect 15224 7628 15327 7640
rect 15339 7630 15365 7656
rect 15380 7651 15410 7662
rect 15442 7658 15504 7674
rect 15442 7656 15488 7658
rect 15442 7640 15504 7656
rect 15516 7640 15522 7688
rect 15525 7680 15605 7688
rect 15525 7678 15544 7680
rect 15559 7678 15593 7680
rect 15525 7662 15605 7678
rect 15525 7640 15544 7662
rect 15559 7646 15589 7662
rect 15617 7656 15623 7730
rect 15626 7656 15645 7800
rect 15660 7656 15666 7800
rect 15675 7730 15688 7800
rect 15740 7796 15762 7800
rect 15733 7774 15762 7788
rect 15815 7774 15831 7788
rect 15869 7784 15875 7786
rect 15882 7784 15990 7800
rect 15997 7784 16003 7786
rect 16011 7784 16026 7800
rect 16092 7794 16111 7797
rect 15733 7772 15831 7774
rect 15858 7772 16026 7784
rect 16041 7774 16057 7788
rect 16092 7775 16114 7794
rect 16124 7788 16140 7789
rect 16123 7786 16140 7788
rect 16124 7781 16140 7786
rect 16114 7774 16120 7775
rect 16123 7774 16152 7781
rect 16041 7773 16152 7774
rect 16041 7772 16158 7773
rect 15717 7764 15768 7772
rect 15815 7764 15849 7772
rect 15717 7752 15742 7764
rect 15749 7752 15768 7764
rect 15822 7762 15849 7764
rect 15858 7762 16079 7772
rect 16114 7769 16120 7772
rect 15822 7758 16079 7762
rect 15717 7744 15768 7752
rect 15815 7744 16079 7758
rect 16123 7764 16158 7772
rect 15669 7696 15688 7730
rect 15733 7736 15762 7744
rect 15733 7730 15750 7736
rect 15733 7728 15767 7730
rect 15815 7728 15831 7744
rect 15832 7734 16040 7744
rect 16041 7734 16057 7744
rect 16105 7740 16120 7755
rect 16123 7752 16124 7764
rect 16131 7752 16158 7764
rect 16123 7744 16158 7752
rect 16123 7743 16152 7744
rect 15843 7730 16057 7734
rect 15858 7728 16057 7730
rect 16092 7730 16105 7740
rect 16123 7730 16140 7743
rect 16092 7728 16140 7730
rect 15734 7724 15767 7728
rect 15730 7722 15767 7724
rect 15730 7721 15797 7722
rect 15730 7716 15761 7721
rect 15767 7716 15797 7721
rect 15730 7712 15797 7716
rect 15703 7709 15797 7712
rect 15703 7702 15752 7709
rect 15703 7696 15733 7702
rect 15752 7697 15757 7702
rect 15669 7680 15749 7696
rect 15761 7688 15797 7709
rect 15858 7704 16047 7728
rect 16092 7727 16139 7728
rect 16105 7722 16139 7727
rect 15873 7701 16047 7704
rect 15866 7698 16047 7701
rect 16075 7721 16139 7722
rect 15669 7678 15688 7680
rect 15703 7678 15737 7680
rect 15669 7662 15749 7678
rect 15669 7656 15688 7662
rect 15385 7630 15488 7640
rect 15339 7628 15488 7630
rect 15509 7628 15544 7640
rect 15178 7626 15340 7628
rect 15190 7606 15209 7626
rect 15224 7624 15254 7626
rect 15073 7598 15114 7606
rect 15196 7602 15209 7606
rect 15261 7610 15340 7626
rect 15372 7626 15544 7628
rect 15372 7610 15451 7626
rect 15458 7624 15488 7626
rect 15036 7588 15065 7598
rect 15079 7588 15108 7598
rect 15123 7588 15153 7602
rect 15196 7588 15239 7602
rect 15261 7598 15451 7610
rect 15516 7606 15522 7626
rect 15246 7588 15276 7598
rect 15277 7588 15435 7598
rect 15439 7588 15469 7598
rect 15473 7588 15503 7602
rect 15531 7588 15544 7626
rect 15616 7640 15645 7656
rect 15659 7640 15688 7656
rect 15703 7646 15733 7662
rect 15761 7640 15767 7688
rect 15770 7682 15789 7688
rect 15804 7682 15834 7690
rect 15770 7674 15834 7682
rect 15770 7658 15850 7674
rect 15866 7667 15928 7698
rect 15944 7667 16006 7698
rect 16075 7696 16124 7721
rect 16139 7696 16169 7712
rect 16038 7682 16068 7690
rect 16075 7688 16185 7696
rect 16038 7674 16083 7682
rect 15770 7656 15789 7658
rect 15804 7656 15850 7658
rect 15770 7640 15850 7656
rect 15877 7654 15912 7667
rect 15953 7664 15990 7667
rect 15953 7662 15995 7664
rect 15882 7651 15912 7654
rect 15891 7647 15898 7651
rect 15898 7646 15899 7647
rect 15857 7640 15867 7646
rect 15616 7632 15651 7640
rect 15616 7606 15617 7632
rect 15624 7606 15651 7632
rect 15559 7588 15589 7602
rect 15616 7598 15651 7606
rect 15653 7632 15694 7640
rect 15653 7606 15668 7632
rect 15675 7606 15694 7632
rect 15758 7628 15789 7640
rect 15804 7628 15907 7640
rect 15919 7630 15945 7656
rect 15960 7651 15990 7662
rect 16022 7658 16084 7674
rect 16022 7656 16068 7658
rect 16022 7640 16084 7656
rect 16096 7640 16102 7688
rect 16105 7680 16185 7688
rect 16105 7678 16124 7680
rect 16139 7678 16173 7680
rect 16105 7662 16185 7678
rect 16105 7640 16124 7662
rect 16139 7646 16169 7662
rect 16197 7656 16203 7730
rect 16206 7656 16225 7800
rect 16240 7656 16246 7800
rect 16255 7730 16268 7800
rect 16320 7796 16342 7800
rect 16313 7774 16342 7788
rect 16395 7774 16411 7788
rect 16449 7784 16455 7786
rect 16462 7784 16570 7800
rect 16577 7784 16583 7786
rect 16591 7784 16606 7800
rect 16672 7794 16691 7797
rect 16313 7772 16411 7774
rect 16438 7772 16606 7784
rect 16621 7774 16637 7788
rect 16672 7775 16694 7794
rect 16704 7788 16720 7789
rect 16703 7786 16720 7788
rect 16704 7781 16720 7786
rect 16694 7774 16700 7775
rect 16703 7774 16732 7781
rect 16621 7773 16732 7774
rect 16621 7772 16738 7773
rect 16297 7764 16348 7772
rect 16395 7764 16429 7772
rect 16297 7752 16322 7764
rect 16329 7752 16348 7764
rect 16402 7762 16429 7764
rect 16438 7762 16659 7772
rect 16694 7769 16700 7772
rect 16402 7758 16659 7762
rect 16297 7744 16348 7752
rect 16395 7744 16659 7758
rect 16703 7764 16738 7772
rect 16249 7696 16268 7730
rect 16313 7736 16342 7744
rect 16313 7730 16330 7736
rect 16313 7728 16347 7730
rect 16395 7728 16411 7744
rect 16412 7734 16620 7744
rect 16621 7734 16637 7744
rect 16685 7740 16700 7755
rect 16703 7752 16704 7764
rect 16711 7752 16738 7764
rect 16703 7744 16738 7752
rect 16703 7743 16732 7744
rect 16423 7730 16637 7734
rect 16438 7728 16637 7730
rect 16672 7730 16685 7740
rect 16703 7730 16720 7743
rect 16672 7728 16720 7730
rect 16314 7724 16347 7728
rect 16310 7722 16347 7724
rect 16310 7721 16377 7722
rect 16310 7716 16341 7721
rect 16347 7716 16377 7721
rect 16310 7712 16377 7716
rect 16283 7709 16377 7712
rect 16283 7702 16332 7709
rect 16283 7696 16313 7702
rect 16332 7697 16337 7702
rect 16249 7680 16329 7696
rect 16341 7688 16377 7709
rect 16438 7704 16627 7728
rect 16672 7727 16719 7728
rect 16685 7722 16719 7727
rect 16453 7701 16627 7704
rect 16446 7698 16627 7701
rect 16655 7721 16719 7722
rect 16249 7678 16268 7680
rect 16283 7678 16317 7680
rect 16249 7662 16329 7678
rect 16249 7656 16268 7662
rect 15965 7630 16068 7640
rect 15919 7628 16068 7630
rect 16089 7628 16124 7640
rect 15758 7626 15920 7628
rect 15770 7606 15789 7626
rect 15804 7624 15834 7626
rect 15653 7598 15694 7606
rect 15776 7602 15789 7606
rect 15841 7610 15920 7626
rect 15952 7626 16124 7628
rect 15952 7610 16031 7626
rect 16038 7624 16068 7626
rect 15616 7588 15645 7598
rect 15659 7588 15688 7598
rect 15703 7588 15733 7602
rect 15776 7588 15819 7602
rect 15841 7598 16031 7610
rect 16096 7606 16102 7626
rect 15826 7588 15856 7598
rect 15857 7588 16015 7598
rect 16019 7588 16049 7598
rect 16053 7588 16083 7602
rect 16111 7588 16124 7626
rect 16196 7640 16225 7656
rect 16239 7640 16268 7656
rect 16283 7646 16313 7662
rect 16341 7640 16347 7688
rect 16350 7682 16369 7688
rect 16384 7682 16414 7690
rect 16350 7674 16414 7682
rect 16350 7658 16430 7674
rect 16446 7667 16508 7698
rect 16524 7667 16586 7698
rect 16655 7696 16704 7721
rect 16719 7696 16749 7712
rect 16618 7682 16648 7690
rect 16655 7688 16765 7696
rect 16618 7674 16663 7682
rect 16350 7656 16369 7658
rect 16384 7656 16430 7658
rect 16350 7640 16430 7656
rect 16457 7654 16492 7667
rect 16533 7664 16570 7667
rect 16533 7662 16575 7664
rect 16462 7651 16492 7654
rect 16471 7647 16478 7651
rect 16478 7646 16479 7647
rect 16437 7640 16447 7646
rect 16196 7632 16231 7640
rect 16196 7606 16197 7632
rect 16204 7606 16231 7632
rect 16139 7588 16169 7602
rect 16196 7598 16231 7606
rect 16233 7632 16274 7640
rect 16233 7606 16248 7632
rect 16255 7606 16274 7632
rect 16338 7628 16369 7640
rect 16384 7628 16487 7640
rect 16499 7630 16525 7656
rect 16540 7651 16570 7662
rect 16602 7658 16664 7674
rect 16602 7656 16648 7658
rect 16602 7640 16664 7656
rect 16676 7640 16682 7688
rect 16685 7680 16765 7688
rect 16685 7678 16704 7680
rect 16719 7678 16753 7680
rect 16685 7662 16765 7678
rect 16685 7640 16704 7662
rect 16719 7646 16749 7662
rect 16777 7656 16783 7730
rect 16786 7656 16805 7800
rect 16820 7656 16826 7800
rect 16835 7730 16848 7800
rect 16900 7796 16922 7800
rect 16893 7774 16922 7788
rect 16975 7774 16991 7788
rect 17029 7784 17035 7786
rect 17042 7784 17150 7800
rect 17157 7784 17163 7786
rect 17171 7784 17186 7800
rect 17252 7794 17271 7797
rect 16893 7772 16991 7774
rect 17018 7772 17186 7784
rect 17201 7774 17217 7788
rect 17252 7775 17274 7794
rect 17284 7788 17300 7789
rect 17283 7786 17300 7788
rect 17284 7781 17300 7786
rect 17274 7774 17280 7775
rect 17283 7774 17312 7781
rect 17201 7773 17312 7774
rect 17201 7772 17318 7773
rect 16877 7764 16928 7772
rect 16975 7764 17009 7772
rect 16877 7752 16902 7764
rect 16909 7752 16928 7764
rect 16982 7762 17009 7764
rect 17018 7762 17239 7772
rect 17274 7769 17280 7772
rect 16982 7758 17239 7762
rect 16877 7744 16928 7752
rect 16975 7744 17239 7758
rect 17283 7764 17318 7772
rect 16829 7696 16848 7730
rect 16893 7736 16922 7744
rect 16893 7730 16910 7736
rect 16893 7728 16927 7730
rect 16975 7728 16991 7744
rect 16992 7734 17200 7744
rect 17201 7734 17217 7744
rect 17265 7740 17280 7755
rect 17283 7752 17284 7764
rect 17291 7752 17318 7764
rect 17283 7744 17318 7752
rect 17283 7743 17312 7744
rect 17003 7730 17217 7734
rect 17018 7728 17217 7730
rect 17252 7730 17265 7740
rect 17283 7730 17300 7743
rect 17252 7728 17300 7730
rect 16894 7724 16927 7728
rect 16890 7722 16927 7724
rect 16890 7721 16957 7722
rect 16890 7716 16921 7721
rect 16927 7716 16957 7721
rect 16890 7712 16957 7716
rect 16863 7709 16957 7712
rect 16863 7702 16912 7709
rect 16863 7696 16893 7702
rect 16912 7697 16917 7702
rect 16829 7680 16909 7696
rect 16921 7688 16957 7709
rect 17018 7704 17207 7728
rect 17252 7727 17299 7728
rect 17265 7722 17299 7727
rect 17033 7701 17207 7704
rect 17026 7698 17207 7701
rect 17235 7721 17299 7722
rect 16829 7678 16848 7680
rect 16863 7678 16897 7680
rect 16829 7662 16909 7678
rect 16829 7656 16848 7662
rect 16545 7630 16648 7640
rect 16499 7628 16648 7630
rect 16669 7628 16704 7640
rect 16338 7626 16500 7628
rect 16350 7606 16369 7626
rect 16384 7624 16414 7626
rect 16233 7598 16274 7606
rect 16356 7602 16369 7606
rect 16421 7610 16500 7626
rect 16532 7626 16704 7628
rect 16532 7610 16611 7626
rect 16618 7624 16648 7626
rect 16196 7588 16225 7598
rect 16239 7588 16268 7598
rect 16283 7588 16313 7602
rect 16356 7588 16399 7602
rect 16421 7598 16611 7610
rect 16676 7606 16682 7626
rect 16406 7588 16436 7598
rect 16437 7588 16595 7598
rect 16599 7588 16629 7598
rect 16633 7588 16663 7602
rect 16691 7588 16704 7626
rect 16776 7640 16805 7656
rect 16819 7640 16848 7656
rect 16863 7646 16893 7662
rect 16921 7640 16927 7688
rect 16930 7682 16949 7688
rect 16964 7682 16994 7690
rect 16930 7674 16994 7682
rect 16930 7658 17010 7674
rect 17026 7667 17088 7698
rect 17104 7667 17166 7698
rect 17235 7696 17284 7721
rect 17299 7696 17329 7712
rect 17198 7682 17228 7690
rect 17235 7688 17345 7696
rect 17198 7674 17243 7682
rect 16930 7656 16949 7658
rect 16964 7656 17010 7658
rect 16930 7640 17010 7656
rect 17037 7654 17072 7667
rect 17113 7664 17150 7667
rect 17113 7662 17155 7664
rect 17042 7651 17072 7654
rect 17051 7647 17058 7651
rect 17058 7646 17059 7647
rect 17017 7640 17027 7646
rect 16776 7632 16811 7640
rect 16776 7606 16777 7632
rect 16784 7606 16811 7632
rect 16719 7588 16749 7602
rect 16776 7598 16811 7606
rect 16813 7632 16854 7640
rect 16813 7606 16828 7632
rect 16835 7606 16854 7632
rect 16918 7628 16949 7640
rect 16964 7628 17067 7640
rect 17079 7630 17105 7656
rect 17120 7651 17150 7662
rect 17182 7658 17244 7674
rect 17182 7656 17228 7658
rect 17182 7640 17244 7656
rect 17256 7640 17262 7688
rect 17265 7680 17345 7688
rect 17265 7678 17284 7680
rect 17299 7678 17333 7680
rect 17265 7662 17345 7678
rect 17265 7640 17284 7662
rect 17299 7646 17329 7662
rect 17357 7656 17363 7730
rect 17366 7656 17385 7800
rect 17400 7656 17406 7800
rect 17415 7730 17428 7800
rect 17480 7796 17502 7800
rect 17473 7774 17502 7788
rect 17555 7774 17571 7788
rect 17609 7784 17615 7786
rect 17622 7784 17730 7800
rect 17737 7784 17743 7786
rect 17751 7784 17766 7800
rect 17832 7794 17851 7797
rect 17473 7772 17571 7774
rect 17598 7772 17766 7784
rect 17781 7774 17797 7788
rect 17832 7775 17854 7794
rect 17864 7788 17880 7789
rect 17863 7786 17880 7788
rect 17864 7781 17880 7786
rect 17854 7774 17860 7775
rect 17863 7774 17892 7781
rect 17781 7773 17892 7774
rect 17781 7772 17898 7773
rect 17457 7764 17508 7772
rect 17555 7764 17589 7772
rect 17457 7752 17482 7764
rect 17489 7752 17508 7764
rect 17562 7762 17589 7764
rect 17598 7762 17819 7772
rect 17854 7769 17860 7772
rect 17562 7758 17819 7762
rect 17457 7744 17508 7752
rect 17555 7744 17819 7758
rect 17863 7764 17898 7772
rect 17409 7696 17428 7730
rect 17473 7736 17502 7744
rect 17473 7730 17490 7736
rect 17473 7728 17507 7730
rect 17555 7728 17571 7744
rect 17572 7734 17780 7744
rect 17781 7734 17797 7744
rect 17845 7740 17860 7755
rect 17863 7752 17864 7764
rect 17871 7752 17898 7764
rect 17863 7744 17898 7752
rect 17863 7743 17892 7744
rect 17583 7730 17797 7734
rect 17598 7728 17797 7730
rect 17832 7730 17845 7740
rect 17863 7730 17880 7743
rect 17832 7728 17880 7730
rect 17474 7724 17507 7728
rect 17470 7722 17507 7724
rect 17470 7721 17537 7722
rect 17470 7716 17501 7721
rect 17507 7716 17537 7721
rect 17470 7712 17537 7716
rect 17443 7709 17537 7712
rect 17443 7702 17492 7709
rect 17443 7696 17473 7702
rect 17492 7697 17497 7702
rect 17409 7680 17489 7696
rect 17501 7688 17537 7709
rect 17598 7704 17787 7728
rect 17832 7727 17879 7728
rect 17845 7722 17879 7727
rect 17613 7701 17787 7704
rect 17606 7698 17787 7701
rect 17815 7721 17879 7722
rect 17409 7678 17428 7680
rect 17443 7678 17477 7680
rect 17409 7662 17489 7678
rect 17409 7656 17428 7662
rect 17125 7630 17228 7640
rect 17079 7628 17228 7630
rect 17249 7628 17284 7640
rect 16918 7626 17080 7628
rect 16930 7606 16949 7626
rect 16964 7624 16994 7626
rect 16813 7598 16854 7606
rect 16936 7602 16949 7606
rect 17001 7610 17080 7626
rect 17112 7626 17284 7628
rect 17112 7610 17191 7626
rect 17198 7624 17228 7626
rect 16776 7588 16805 7598
rect 16819 7588 16848 7598
rect 16863 7588 16893 7602
rect 16936 7588 16979 7602
rect 17001 7598 17191 7610
rect 17256 7606 17262 7626
rect 16986 7588 17016 7598
rect 17017 7588 17175 7598
rect 17179 7588 17209 7598
rect 17213 7588 17243 7602
rect 17271 7588 17284 7626
rect 17356 7640 17385 7656
rect 17399 7640 17428 7656
rect 17443 7646 17473 7662
rect 17501 7640 17507 7688
rect 17510 7682 17529 7688
rect 17544 7682 17574 7690
rect 17510 7674 17574 7682
rect 17510 7658 17590 7674
rect 17606 7667 17668 7698
rect 17684 7667 17746 7698
rect 17815 7696 17864 7721
rect 17879 7696 17909 7712
rect 17778 7682 17808 7690
rect 17815 7688 17925 7696
rect 17778 7674 17823 7682
rect 17510 7656 17529 7658
rect 17544 7656 17590 7658
rect 17510 7640 17590 7656
rect 17617 7654 17652 7667
rect 17693 7664 17730 7667
rect 17693 7662 17735 7664
rect 17622 7651 17652 7654
rect 17631 7647 17638 7651
rect 17638 7646 17639 7647
rect 17597 7640 17607 7646
rect 17356 7632 17391 7640
rect 17356 7606 17357 7632
rect 17364 7606 17391 7632
rect 17299 7588 17329 7602
rect 17356 7598 17391 7606
rect 17393 7632 17434 7640
rect 17393 7606 17408 7632
rect 17415 7606 17434 7632
rect 17498 7628 17529 7640
rect 17544 7628 17647 7640
rect 17659 7630 17685 7656
rect 17700 7651 17730 7662
rect 17762 7658 17824 7674
rect 17762 7656 17808 7658
rect 17762 7640 17824 7656
rect 17836 7640 17842 7688
rect 17845 7680 17925 7688
rect 17845 7678 17864 7680
rect 17879 7678 17913 7680
rect 17845 7662 17925 7678
rect 17845 7640 17864 7662
rect 17879 7646 17909 7662
rect 17937 7656 17943 7730
rect 17946 7656 17965 7800
rect 17980 7656 17986 7800
rect 17995 7730 18008 7800
rect 18060 7796 18082 7800
rect 18053 7774 18082 7788
rect 18135 7774 18151 7788
rect 18189 7784 18195 7786
rect 18202 7784 18310 7800
rect 18317 7784 18323 7786
rect 18331 7784 18346 7800
rect 18412 7794 18431 7797
rect 18053 7772 18151 7774
rect 18178 7772 18346 7784
rect 18361 7774 18377 7788
rect 18412 7775 18434 7794
rect 18444 7788 18460 7789
rect 18443 7786 18460 7788
rect 18444 7781 18460 7786
rect 18434 7774 18440 7775
rect 18443 7774 18472 7781
rect 18361 7773 18472 7774
rect 18361 7772 18478 7773
rect 18037 7764 18088 7772
rect 18135 7764 18169 7772
rect 18037 7752 18062 7764
rect 18069 7752 18088 7764
rect 18142 7762 18169 7764
rect 18178 7762 18399 7772
rect 18434 7769 18440 7772
rect 18142 7758 18399 7762
rect 18037 7744 18088 7752
rect 18135 7744 18399 7758
rect 18443 7764 18478 7772
rect 17989 7696 18008 7730
rect 18053 7736 18082 7744
rect 18053 7730 18070 7736
rect 18053 7728 18087 7730
rect 18135 7728 18151 7744
rect 18152 7734 18360 7744
rect 18361 7734 18377 7744
rect 18425 7740 18440 7755
rect 18443 7752 18444 7764
rect 18451 7752 18478 7764
rect 18443 7744 18478 7752
rect 18443 7743 18472 7744
rect 18163 7730 18377 7734
rect 18178 7728 18377 7730
rect 18412 7730 18425 7740
rect 18443 7730 18460 7743
rect 18412 7728 18460 7730
rect 18054 7724 18087 7728
rect 18050 7722 18087 7724
rect 18050 7721 18117 7722
rect 18050 7716 18081 7721
rect 18087 7716 18117 7721
rect 18050 7712 18117 7716
rect 18023 7709 18117 7712
rect 18023 7702 18072 7709
rect 18023 7696 18053 7702
rect 18072 7697 18077 7702
rect 17989 7680 18069 7696
rect 18081 7688 18117 7709
rect 18178 7704 18367 7728
rect 18412 7727 18459 7728
rect 18425 7722 18459 7727
rect 18193 7701 18367 7704
rect 18186 7698 18367 7701
rect 18395 7721 18459 7722
rect 17989 7678 18008 7680
rect 18023 7678 18057 7680
rect 17989 7662 18069 7678
rect 17989 7656 18008 7662
rect 17705 7630 17808 7640
rect 17659 7628 17808 7630
rect 17829 7628 17864 7640
rect 17498 7626 17660 7628
rect 17510 7606 17529 7626
rect 17544 7624 17574 7626
rect 17393 7598 17434 7606
rect 17516 7602 17529 7606
rect 17581 7610 17660 7626
rect 17692 7626 17864 7628
rect 17692 7610 17771 7626
rect 17778 7624 17808 7626
rect 17356 7588 17385 7598
rect 17399 7588 17428 7598
rect 17443 7588 17473 7602
rect 17516 7588 17559 7602
rect 17581 7598 17771 7610
rect 17836 7606 17842 7626
rect 17566 7588 17596 7598
rect 17597 7588 17755 7598
rect 17759 7588 17789 7598
rect 17793 7588 17823 7602
rect 17851 7588 17864 7626
rect 17936 7640 17965 7656
rect 17979 7640 18008 7656
rect 18023 7646 18053 7662
rect 18081 7640 18087 7688
rect 18090 7682 18109 7688
rect 18124 7682 18154 7690
rect 18090 7674 18154 7682
rect 18090 7658 18170 7674
rect 18186 7667 18248 7698
rect 18264 7667 18326 7698
rect 18395 7696 18444 7721
rect 18459 7696 18489 7712
rect 18358 7682 18388 7690
rect 18395 7688 18505 7696
rect 18358 7674 18403 7682
rect 18090 7656 18109 7658
rect 18124 7656 18170 7658
rect 18090 7640 18170 7656
rect 18197 7654 18232 7667
rect 18273 7664 18310 7667
rect 18273 7662 18315 7664
rect 18202 7651 18232 7654
rect 18211 7647 18218 7651
rect 18218 7646 18219 7647
rect 18177 7640 18187 7646
rect 17936 7632 17971 7640
rect 17936 7606 17937 7632
rect 17944 7606 17971 7632
rect 17879 7588 17909 7602
rect 17936 7598 17971 7606
rect 17973 7632 18014 7640
rect 17973 7606 17988 7632
rect 17995 7606 18014 7632
rect 18078 7628 18109 7640
rect 18124 7628 18227 7640
rect 18239 7630 18265 7656
rect 18280 7651 18310 7662
rect 18342 7658 18404 7674
rect 18342 7656 18388 7658
rect 18342 7640 18404 7656
rect 18416 7640 18422 7688
rect 18425 7680 18505 7688
rect 18425 7678 18444 7680
rect 18459 7678 18493 7680
rect 18425 7662 18505 7678
rect 18425 7640 18444 7662
rect 18459 7646 18489 7662
rect 18517 7656 18523 7730
rect 18532 7656 18545 7800
rect 18285 7630 18388 7640
rect 18239 7628 18388 7630
rect 18409 7628 18444 7640
rect 18078 7626 18240 7628
rect 18090 7606 18109 7626
rect 18124 7624 18154 7626
rect 17973 7598 18014 7606
rect 18096 7602 18109 7606
rect 18161 7610 18240 7626
rect 18272 7626 18444 7628
rect 18272 7610 18351 7626
rect 18358 7624 18388 7626
rect 17936 7588 17965 7598
rect 17979 7588 18008 7598
rect 18023 7588 18053 7602
rect 18096 7588 18139 7602
rect 18161 7598 18351 7610
rect 18416 7606 18422 7626
rect 18146 7588 18176 7598
rect 18177 7588 18335 7598
rect 18339 7588 18369 7598
rect 18373 7588 18403 7602
rect 18431 7588 18444 7626
rect 18516 7640 18545 7656
rect 18516 7632 18551 7640
rect 18516 7606 18517 7632
rect 18524 7606 18551 7632
rect 18459 7588 18489 7602
rect 18516 7598 18551 7606
rect 18516 7588 18545 7598
rect -1 7582 18545 7588
rect 0 7574 18545 7582
rect 15 7544 28 7574
rect 43 7560 73 7574
rect 116 7560 159 7574
rect 166 7560 386 7574
rect 393 7560 423 7574
rect 83 7546 98 7558
rect 117 7546 130 7560
rect 198 7556 351 7560
rect 80 7544 102 7546
rect 180 7544 372 7556
rect 451 7544 464 7574
rect 479 7560 509 7574
rect 546 7544 565 7574
rect 580 7544 586 7574
rect 595 7544 608 7574
rect 623 7560 653 7574
rect 696 7560 739 7574
rect 746 7560 966 7574
rect 973 7560 1003 7574
rect 663 7546 678 7558
rect 697 7546 710 7560
rect 778 7556 931 7560
rect 660 7544 682 7546
rect 760 7544 952 7556
rect 1031 7544 1044 7574
rect 1059 7560 1089 7574
rect 1126 7544 1145 7574
rect 1160 7544 1166 7574
rect 1175 7544 1188 7574
rect 1203 7560 1233 7574
rect 1276 7560 1319 7574
rect 1326 7560 1546 7574
rect 1553 7560 1583 7574
rect 1243 7546 1258 7558
rect 1277 7546 1290 7560
rect 1358 7556 1511 7560
rect 1240 7544 1262 7546
rect 1340 7544 1532 7556
rect 1611 7544 1624 7574
rect 1639 7560 1669 7574
rect 1706 7544 1725 7574
rect 1740 7544 1746 7574
rect 1755 7544 1768 7574
rect 1783 7560 1813 7574
rect 1856 7560 1899 7574
rect 1906 7560 2126 7574
rect 2133 7560 2163 7574
rect 1823 7546 1838 7558
rect 1857 7546 1870 7560
rect 1938 7556 2091 7560
rect 1820 7544 1842 7546
rect 1920 7544 2112 7556
rect 2191 7544 2204 7574
rect 2219 7560 2249 7574
rect 2286 7544 2305 7574
rect 2320 7544 2326 7574
rect 2335 7544 2348 7574
rect 2363 7560 2393 7574
rect 2436 7560 2479 7574
rect 2486 7560 2706 7574
rect 2713 7560 2743 7574
rect 2403 7546 2418 7558
rect 2437 7546 2450 7560
rect 2518 7556 2671 7560
rect 2400 7544 2422 7546
rect 2500 7544 2692 7556
rect 2771 7544 2784 7574
rect 2799 7560 2829 7574
rect 2866 7544 2885 7574
rect 2900 7544 2906 7574
rect 2915 7544 2928 7574
rect 2943 7560 2973 7574
rect 3016 7560 3059 7574
rect 3066 7560 3286 7574
rect 3293 7560 3323 7574
rect 2983 7546 2998 7558
rect 3017 7546 3030 7560
rect 3098 7556 3251 7560
rect 2980 7544 3002 7546
rect 3080 7544 3272 7556
rect 3351 7544 3364 7574
rect 3379 7560 3409 7574
rect 3446 7544 3465 7574
rect 3480 7544 3486 7574
rect 3495 7544 3508 7574
rect 3523 7560 3553 7574
rect 3596 7560 3639 7574
rect 3646 7560 3866 7574
rect 3873 7560 3903 7574
rect 3563 7546 3578 7558
rect 3597 7546 3610 7560
rect 3678 7556 3831 7560
rect 3560 7544 3582 7546
rect 3660 7544 3852 7556
rect 3931 7544 3944 7574
rect 3959 7560 3989 7574
rect 4026 7544 4045 7574
rect 4060 7544 4066 7574
rect 4075 7544 4088 7574
rect 4103 7560 4133 7574
rect 4176 7560 4219 7574
rect 4226 7560 4446 7574
rect 4453 7560 4483 7574
rect 4143 7546 4158 7558
rect 4177 7546 4190 7560
rect 4258 7556 4411 7560
rect 4140 7544 4162 7546
rect 4240 7544 4432 7556
rect 4511 7544 4524 7574
rect 4539 7560 4569 7574
rect 4606 7544 4625 7574
rect 4640 7544 4646 7574
rect 4655 7544 4668 7574
rect 4683 7560 4713 7574
rect 4756 7560 4799 7574
rect 4806 7560 5026 7574
rect 5033 7560 5063 7574
rect 4723 7546 4738 7558
rect 4757 7546 4770 7560
rect 4838 7556 4991 7560
rect 4720 7544 4742 7546
rect 4820 7544 5012 7556
rect 5091 7544 5104 7574
rect 5119 7560 5149 7574
rect 5186 7544 5205 7574
rect 5220 7544 5226 7574
rect 5235 7544 5248 7574
rect 5263 7560 5293 7574
rect 5336 7560 5379 7574
rect 5386 7560 5606 7574
rect 5613 7560 5643 7574
rect 5303 7546 5318 7558
rect 5337 7546 5350 7560
rect 5418 7556 5571 7560
rect 5300 7544 5322 7546
rect 5400 7544 5592 7556
rect 5671 7544 5684 7574
rect 5699 7560 5729 7574
rect 5766 7544 5785 7574
rect 5800 7544 5806 7574
rect 5815 7544 5828 7574
rect 5843 7560 5873 7574
rect 5916 7560 5959 7574
rect 5966 7560 6186 7574
rect 6193 7560 6223 7574
rect 5883 7546 5898 7558
rect 5917 7546 5930 7560
rect 5998 7556 6151 7560
rect 5880 7544 5902 7546
rect 5980 7544 6172 7556
rect 6251 7544 6264 7574
rect 6279 7560 6309 7574
rect 6346 7544 6365 7574
rect 6380 7544 6386 7574
rect 6395 7544 6408 7574
rect 6423 7560 6453 7574
rect 6496 7560 6539 7574
rect 6546 7560 6766 7574
rect 6773 7560 6803 7574
rect 6463 7546 6478 7558
rect 6497 7546 6510 7560
rect 6578 7556 6731 7560
rect 6460 7544 6482 7546
rect 6560 7544 6752 7556
rect 6831 7544 6844 7574
rect 6859 7560 6889 7574
rect 6926 7544 6945 7574
rect 6960 7544 6966 7574
rect 6975 7544 6988 7574
rect 7003 7560 7033 7574
rect 7076 7560 7119 7574
rect 7126 7560 7346 7574
rect 7353 7560 7383 7574
rect 7043 7546 7058 7558
rect 7077 7546 7090 7560
rect 7158 7556 7311 7560
rect 7040 7544 7062 7546
rect 7140 7544 7332 7556
rect 7411 7544 7424 7574
rect 7439 7560 7469 7574
rect 7506 7544 7525 7574
rect 7540 7544 7546 7574
rect 7555 7544 7568 7574
rect 7583 7560 7613 7574
rect 7656 7560 7699 7574
rect 7706 7560 7926 7574
rect 7933 7560 7963 7574
rect 7623 7546 7638 7558
rect 7657 7546 7670 7560
rect 7738 7556 7891 7560
rect 7620 7544 7642 7546
rect 7720 7544 7912 7556
rect 7991 7544 8004 7574
rect 8019 7560 8049 7574
rect 8086 7544 8105 7574
rect 8120 7544 8126 7574
rect 8135 7544 8148 7574
rect 8163 7560 8193 7574
rect 8236 7560 8279 7574
rect 8286 7560 8506 7574
rect 8513 7560 8543 7574
rect 8203 7546 8218 7558
rect 8237 7546 8250 7560
rect 8318 7556 8471 7560
rect 8200 7544 8222 7546
rect 8300 7544 8492 7556
rect 8571 7544 8584 7574
rect 8599 7560 8629 7574
rect 8666 7544 8685 7574
rect 8700 7544 8706 7574
rect 8715 7544 8728 7574
rect 8743 7560 8773 7574
rect 8816 7560 8859 7574
rect 8866 7560 9086 7574
rect 9093 7560 9123 7574
rect 8783 7546 8798 7558
rect 8817 7546 8830 7560
rect 8898 7556 9051 7560
rect 8780 7544 8802 7546
rect 8880 7544 9072 7556
rect 9151 7544 9164 7574
rect 9179 7560 9209 7574
rect 9246 7544 9265 7574
rect 9280 7544 9286 7574
rect 9295 7544 9308 7574
rect 9323 7560 9353 7574
rect 9396 7560 9439 7574
rect 9446 7560 9666 7574
rect 9673 7560 9703 7574
rect 9363 7546 9378 7558
rect 9397 7546 9410 7560
rect 9478 7556 9631 7560
rect 9360 7544 9382 7546
rect 9460 7544 9652 7556
rect 9731 7544 9744 7574
rect 9759 7560 9789 7574
rect 9826 7544 9845 7574
rect 9860 7544 9866 7574
rect 9875 7544 9888 7574
rect 9903 7560 9933 7574
rect 9976 7560 10019 7574
rect 10026 7560 10246 7574
rect 10253 7560 10283 7574
rect 9943 7546 9958 7558
rect 9977 7546 9990 7560
rect 10058 7556 10211 7560
rect 9940 7544 9962 7546
rect 10040 7544 10232 7556
rect 10311 7544 10324 7574
rect 10339 7560 10369 7574
rect 10406 7544 10425 7574
rect 10440 7544 10446 7574
rect 10455 7544 10468 7574
rect 10483 7560 10513 7574
rect 10556 7560 10599 7574
rect 10606 7560 10826 7574
rect 10833 7560 10863 7574
rect 10523 7546 10538 7558
rect 10557 7546 10570 7560
rect 10638 7556 10791 7560
rect 10520 7544 10542 7546
rect 10620 7544 10812 7556
rect 10891 7544 10904 7574
rect 10919 7560 10949 7574
rect 10986 7544 11005 7574
rect 11020 7544 11026 7574
rect 11035 7544 11048 7574
rect 11063 7560 11093 7574
rect 11136 7560 11179 7574
rect 11186 7560 11406 7574
rect 11413 7560 11443 7574
rect 11103 7546 11118 7558
rect 11137 7546 11150 7560
rect 11218 7556 11371 7560
rect 11100 7544 11122 7546
rect 11200 7544 11392 7556
rect 11471 7544 11484 7574
rect 11499 7560 11529 7574
rect 11566 7544 11585 7574
rect 11600 7544 11606 7574
rect 11615 7544 11628 7574
rect 11643 7560 11673 7574
rect 11716 7560 11759 7574
rect 11766 7560 11986 7574
rect 11993 7560 12023 7574
rect 11683 7546 11698 7558
rect 11717 7546 11730 7560
rect 11798 7556 11951 7560
rect 11680 7544 11702 7546
rect 11780 7544 11972 7556
rect 12051 7544 12064 7574
rect 12079 7560 12109 7574
rect 12146 7544 12165 7574
rect 12180 7544 12186 7574
rect 12195 7544 12208 7574
rect 12223 7560 12253 7574
rect 12296 7560 12339 7574
rect 12346 7560 12566 7574
rect 12573 7560 12603 7574
rect 12263 7546 12278 7558
rect 12297 7546 12310 7560
rect 12378 7556 12531 7560
rect 12260 7544 12282 7546
rect 12360 7544 12552 7556
rect 12631 7544 12644 7574
rect 12659 7560 12689 7574
rect 12726 7544 12745 7574
rect 12760 7544 12766 7574
rect 12775 7544 12788 7574
rect 12803 7560 12833 7574
rect 12876 7560 12919 7574
rect 12926 7560 13146 7574
rect 13153 7560 13183 7574
rect 12843 7546 12858 7558
rect 12877 7546 12890 7560
rect 12958 7556 13111 7560
rect 12840 7544 12862 7546
rect 12940 7544 13132 7556
rect 13211 7544 13224 7574
rect 13239 7560 13269 7574
rect 13306 7544 13325 7574
rect 13340 7544 13346 7574
rect 13355 7544 13368 7574
rect 13383 7560 13413 7574
rect 13456 7560 13499 7574
rect 13506 7560 13726 7574
rect 13733 7560 13763 7574
rect 13423 7546 13438 7558
rect 13457 7546 13470 7560
rect 13538 7556 13691 7560
rect 13420 7544 13442 7546
rect 13520 7544 13712 7556
rect 13791 7544 13804 7574
rect 13819 7560 13849 7574
rect 13886 7544 13905 7574
rect 13920 7544 13926 7574
rect 13935 7544 13948 7574
rect 13963 7560 13993 7574
rect 14036 7560 14079 7574
rect 14086 7560 14306 7574
rect 14313 7560 14343 7574
rect 14003 7546 14018 7558
rect 14037 7546 14050 7560
rect 14118 7556 14271 7560
rect 14000 7544 14022 7546
rect 14100 7544 14292 7556
rect 14371 7544 14384 7574
rect 14399 7560 14429 7574
rect 14466 7544 14485 7574
rect 14500 7544 14506 7574
rect 14515 7544 14528 7574
rect 14543 7560 14573 7574
rect 14616 7560 14659 7574
rect 14666 7560 14886 7574
rect 14893 7560 14923 7574
rect 14583 7546 14598 7558
rect 14617 7546 14630 7560
rect 14698 7556 14851 7560
rect 14580 7544 14602 7546
rect 14680 7544 14872 7556
rect 14951 7544 14964 7574
rect 14979 7560 15009 7574
rect 15046 7544 15065 7574
rect 15080 7544 15086 7574
rect 15095 7544 15108 7574
rect 15123 7560 15153 7574
rect 15196 7560 15239 7574
rect 15246 7560 15466 7574
rect 15473 7560 15503 7574
rect 15163 7546 15178 7558
rect 15197 7546 15210 7560
rect 15278 7556 15431 7560
rect 15160 7544 15182 7546
rect 15260 7544 15452 7556
rect 15531 7544 15544 7574
rect 15559 7560 15589 7574
rect 15626 7544 15645 7574
rect 15660 7544 15666 7574
rect 15675 7544 15688 7574
rect 15703 7560 15733 7574
rect 15776 7560 15819 7574
rect 15826 7560 16046 7574
rect 16053 7560 16083 7574
rect 15743 7546 15758 7558
rect 15777 7546 15790 7560
rect 15858 7556 16011 7560
rect 15740 7544 15762 7546
rect 15840 7544 16032 7556
rect 16111 7544 16124 7574
rect 16139 7560 16169 7574
rect 16206 7544 16225 7574
rect 16240 7544 16246 7574
rect 16255 7544 16268 7574
rect 16283 7560 16313 7574
rect 16356 7560 16399 7574
rect 16406 7560 16626 7574
rect 16633 7560 16663 7574
rect 16323 7546 16338 7558
rect 16357 7546 16370 7560
rect 16438 7556 16591 7560
rect 16320 7544 16342 7546
rect 16420 7544 16612 7556
rect 16691 7544 16704 7574
rect 16719 7560 16749 7574
rect 16786 7544 16805 7574
rect 16820 7544 16826 7574
rect 16835 7544 16848 7574
rect 16863 7560 16893 7574
rect 16936 7560 16979 7574
rect 16986 7560 17206 7574
rect 17213 7560 17243 7574
rect 16903 7546 16918 7558
rect 16937 7546 16950 7560
rect 17018 7556 17171 7560
rect 16900 7544 16922 7546
rect 17000 7544 17192 7556
rect 17271 7544 17284 7574
rect 17299 7560 17329 7574
rect 17366 7544 17385 7574
rect 17400 7544 17406 7574
rect 17415 7544 17428 7574
rect 17443 7560 17473 7574
rect 17516 7560 17559 7574
rect 17566 7560 17786 7574
rect 17793 7560 17823 7574
rect 17483 7546 17498 7558
rect 17517 7546 17530 7560
rect 17598 7556 17751 7560
rect 17480 7544 17502 7546
rect 17580 7544 17772 7556
rect 17851 7544 17864 7574
rect 17879 7560 17909 7574
rect 17946 7544 17965 7574
rect 17980 7544 17986 7574
rect 17995 7544 18008 7574
rect 18023 7560 18053 7574
rect 18096 7560 18139 7574
rect 18146 7560 18366 7574
rect 18373 7560 18403 7574
rect 18063 7546 18078 7558
rect 18097 7546 18110 7560
rect 18178 7556 18331 7560
rect 18060 7544 18082 7546
rect 18160 7544 18352 7556
rect 18431 7544 18444 7574
rect 18459 7560 18489 7574
rect 18532 7544 18545 7574
rect 0 7530 18545 7544
rect 15 7460 28 7530
rect 80 7526 102 7530
rect 73 7504 102 7518
rect 155 7504 171 7518
rect 209 7514 215 7516
rect 222 7514 330 7530
rect 337 7514 343 7516
rect 351 7514 366 7530
rect 432 7524 451 7527
rect 73 7502 171 7504
rect 198 7502 366 7514
rect 381 7504 397 7518
rect 432 7505 454 7524
rect 464 7518 480 7519
rect 463 7516 480 7518
rect 464 7511 480 7516
rect 454 7504 460 7505
rect 463 7504 492 7511
rect 381 7503 492 7504
rect 381 7502 498 7503
rect 57 7494 108 7502
rect 155 7494 189 7502
rect 57 7482 82 7494
rect 89 7482 108 7494
rect 162 7492 189 7494
rect 198 7492 419 7502
rect 454 7499 460 7502
rect 162 7488 419 7492
rect 57 7474 108 7482
rect 155 7474 419 7488
rect 463 7494 498 7502
rect 9 7426 28 7460
rect 73 7466 102 7474
rect 73 7460 90 7466
rect 73 7458 107 7460
rect 155 7458 171 7474
rect 172 7464 380 7474
rect 381 7464 397 7474
rect 445 7470 460 7485
rect 463 7482 464 7494
rect 471 7482 498 7494
rect 463 7474 498 7482
rect 463 7473 492 7474
rect 183 7460 397 7464
rect 198 7458 397 7460
rect 432 7460 445 7470
rect 463 7460 480 7473
rect 432 7458 480 7460
rect 74 7454 107 7458
rect 70 7452 107 7454
rect 70 7451 137 7452
rect 70 7446 101 7451
rect 107 7446 137 7451
rect 70 7442 137 7446
rect 43 7439 137 7442
rect 43 7432 92 7439
rect 43 7426 73 7432
rect 92 7427 97 7432
rect 9 7410 89 7426
rect 101 7418 137 7439
rect 198 7434 387 7458
rect 432 7457 479 7458
rect 445 7452 479 7457
rect 213 7431 387 7434
rect 206 7428 387 7431
rect 415 7451 479 7452
rect 9 7408 28 7410
rect 43 7408 77 7410
rect 9 7392 89 7408
rect 9 7386 28 7392
rect -1 7370 28 7386
rect 43 7376 73 7392
rect 101 7370 107 7418
rect 110 7412 129 7418
rect 144 7412 174 7420
rect 110 7404 174 7412
rect 110 7388 190 7404
rect 206 7397 268 7428
rect 284 7397 346 7428
rect 415 7426 464 7451
rect 479 7426 509 7442
rect 378 7412 408 7420
rect 415 7418 525 7426
rect 378 7404 423 7412
rect 110 7386 129 7388
rect 144 7386 190 7388
rect 110 7370 190 7386
rect 217 7384 252 7397
rect 293 7394 330 7397
rect 293 7392 335 7394
rect 222 7381 252 7384
rect 231 7377 238 7381
rect 238 7376 239 7377
rect 197 7370 207 7376
rect -7 7362 34 7370
rect -7 7336 8 7362
rect 15 7336 34 7362
rect 98 7358 129 7370
rect 144 7358 247 7370
rect 259 7360 285 7386
rect 300 7381 330 7392
rect 362 7388 424 7404
rect 362 7386 408 7388
rect 362 7370 424 7386
rect 436 7370 442 7418
rect 445 7410 525 7418
rect 445 7408 464 7410
rect 479 7408 513 7410
rect 445 7392 525 7408
rect 445 7370 464 7392
rect 479 7376 509 7392
rect 537 7386 543 7460
rect 546 7386 565 7530
rect 580 7386 586 7530
rect 595 7460 608 7530
rect 660 7526 682 7530
rect 653 7504 682 7518
rect 735 7504 751 7518
rect 789 7514 795 7516
rect 802 7514 910 7530
rect 917 7514 923 7516
rect 931 7514 946 7530
rect 1012 7524 1031 7527
rect 653 7502 751 7504
rect 778 7502 946 7514
rect 961 7504 977 7518
rect 1012 7505 1034 7524
rect 1044 7518 1060 7519
rect 1043 7516 1060 7518
rect 1044 7511 1060 7516
rect 1034 7504 1040 7505
rect 1043 7504 1072 7511
rect 961 7503 1072 7504
rect 961 7502 1078 7503
rect 637 7494 688 7502
rect 735 7494 769 7502
rect 637 7482 662 7494
rect 669 7482 688 7494
rect 742 7492 769 7494
rect 778 7492 999 7502
rect 1034 7499 1040 7502
rect 742 7488 999 7492
rect 637 7474 688 7482
rect 735 7474 999 7488
rect 1043 7494 1078 7502
rect 589 7426 608 7460
rect 653 7466 682 7474
rect 653 7460 670 7466
rect 653 7458 687 7460
rect 735 7458 751 7474
rect 752 7464 960 7474
rect 961 7464 977 7474
rect 1025 7470 1040 7485
rect 1043 7482 1044 7494
rect 1051 7482 1078 7494
rect 1043 7474 1078 7482
rect 1043 7473 1072 7474
rect 763 7460 977 7464
rect 778 7458 977 7460
rect 1012 7460 1025 7470
rect 1043 7460 1060 7473
rect 1012 7458 1060 7460
rect 654 7454 687 7458
rect 650 7452 687 7454
rect 650 7451 717 7452
rect 650 7446 681 7451
rect 687 7446 717 7451
rect 650 7442 717 7446
rect 623 7439 717 7442
rect 623 7432 672 7439
rect 623 7426 653 7432
rect 672 7427 677 7432
rect 589 7410 669 7426
rect 681 7418 717 7439
rect 778 7434 967 7458
rect 1012 7457 1059 7458
rect 1025 7452 1059 7457
rect 793 7431 967 7434
rect 786 7428 967 7431
rect 995 7451 1059 7452
rect 589 7408 608 7410
rect 623 7408 657 7410
rect 589 7392 669 7408
rect 589 7386 608 7392
rect 305 7360 408 7370
rect 259 7358 408 7360
rect 429 7358 464 7370
rect 98 7356 260 7358
rect 110 7336 129 7356
rect 144 7354 174 7356
rect -7 7328 34 7336
rect 116 7332 129 7336
rect 181 7340 260 7356
rect 292 7356 464 7358
rect 292 7340 371 7356
rect 378 7354 408 7356
rect -1 7318 28 7328
rect 43 7318 73 7332
rect 116 7318 159 7332
rect 181 7328 371 7340
rect 436 7336 442 7356
rect 166 7318 196 7328
rect 197 7318 355 7328
rect 359 7318 389 7328
rect 393 7318 423 7332
rect 451 7318 464 7356
rect 536 7370 565 7386
rect 579 7370 608 7386
rect 623 7376 653 7392
rect 681 7370 687 7418
rect 690 7412 709 7418
rect 724 7412 754 7420
rect 690 7404 754 7412
rect 690 7388 770 7404
rect 786 7397 848 7428
rect 864 7397 926 7428
rect 995 7426 1044 7451
rect 1059 7426 1089 7442
rect 958 7412 988 7420
rect 995 7418 1105 7426
rect 958 7404 1003 7412
rect 690 7386 709 7388
rect 724 7386 770 7388
rect 690 7370 770 7386
rect 797 7384 832 7397
rect 873 7394 910 7397
rect 873 7392 915 7394
rect 802 7381 832 7384
rect 811 7377 818 7381
rect 818 7376 819 7377
rect 777 7370 787 7376
rect 536 7362 571 7370
rect 536 7336 537 7362
rect 544 7336 571 7362
rect 479 7318 509 7332
rect 536 7328 571 7336
rect 573 7362 614 7370
rect 573 7336 588 7362
rect 595 7336 614 7362
rect 678 7358 709 7370
rect 724 7358 827 7370
rect 839 7360 865 7386
rect 880 7381 910 7392
rect 942 7388 1004 7404
rect 942 7386 988 7388
rect 942 7370 1004 7386
rect 1016 7370 1022 7418
rect 1025 7410 1105 7418
rect 1025 7408 1044 7410
rect 1059 7408 1093 7410
rect 1025 7392 1105 7408
rect 1025 7370 1044 7392
rect 1059 7376 1089 7392
rect 1117 7386 1123 7460
rect 1126 7386 1145 7530
rect 1160 7386 1166 7530
rect 1175 7460 1188 7530
rect 1240 7526 1262 7530
rect 1233 7504 1262 7518
rect 1315 7504 1331 7518
rect 1369 7514 1375 7516
rect 1382 7514 1490 7530
rect 1497 7514 1503 7516
rect 1511 7514 1526 7530
rect 1592 7524 1611 7527
rect 1233 7502 1331 7504
rect 1358 7502 1526 7514
rect 1541 7504 1557 7518
rect 1592 7505 1614 7524
rect 1624 7518 1640 7519
rect 1623 7516 1640 7518
rect 1624 7511 1640 7516
rect 1614 7504 1620 7505
rect 1623 7504 1652 7511
rect 1541 7503 1652 7504
rect 1541 7502 1658 7503
rect 1217 7494 1268 7502
rect 1315 7494 1349 7502
rect 1217 7482 1242 7494
rect 1249 7482 1268 7494
rect 1322 7492 1349 7494
rect 1358 7492 1579 7502
rect 1614 7499 1620 7502
rect 1322 7488 1579 7492
rect 1217 7474 1268 7482
rect 1315 7474 1579 7488
rect 1623 7494 1658 7502
rect 1169 7426 1188 7460
rect 1233 7466 1262 7474
rect 1233 7460 1250 7466
rect 1233 7458 1267 7460
rect 1315 7458 1331 7474
rect 1332 7464 1540 7474
rect 1541 7464 1557 7474
rect 1605 7470 1620 7485
rect 1623 7482 1624 7494
rect 1631 7482 1658 7494
rect 1623 7474 1658 7482
rect 1623 7473 1652 7474
rect 1343 7460 1557 7464
rect 1358 7458 1557 7460
rect 1592 7460 1605 7470
rect 1623 7460 1640 7473
rect 1592 7458 1640 7460
rect 1234 7454 1267 7458
rect 1230 7452 1267 7454
rect 1230 7451 1297 7452
rect 1230 7446 1261 7451
rect 1267 7446 1297 7451
rect 1230 7442 1297 7446
rect 1203 7439 1297 7442
rect 1203 7432 1252 7439
rect 1203 7426 1233 7432
rect 1252 7427 1257 7432
rect 1169 7410 1249 7426
rect 1261 7418 1297 7439
rect 1358 7434 1547 7458
rect 1592 7457 1639 7458
rect 1605 7452 1639 7457
rect 1373 7431 1547 7434
rect 1366 7428 1547 7431
rect 1575 7451 1639 7452
rect 1169 7408 1188 7410
rect 1203 7408 1237 7410
rect 1169 7392 1249 7408
rect 1169 7386 1188 7392
rect 885 7360 988 7370
rect 839 7358 988 7360
rect 1009 7358 1044 7370
rect 678 7356 840 7358
rect 690 7336 709 7356
rect 724 7354 754 7356
rect 573 7328 614 7336
rect 696 7332 709 7336
rect 761 7340 840 7356
rect 872 7356 1044 7358
rect 872 7340 951 7356
rect 958 7354 988 7356
rect 536 7318 565 7328
rect 579 7318 608 7328
rect 623 7318 653 7332
rect 696 7318 739 7332
rect 761 7328 951 7340
rect 1016 7336 1022 7356
rect 746 7318 776 7328
rect 777 7318 935 7328
rect 939 7318 969 7328
rect 973 7318 1003 7332
rect 1031 7318 1044 7356
rect 1116 7370 1145 7386
rect 1159 7370 1188 7386
rect 1203 7376 1233 7392
rect 1261 7370 1267 7418
rect 1270 7412 1289 7418
rect 1304 7412 1334 7420
rect 1270 7404 1334 7412
rect 1270 7388 1350 7404
rect 1366 7397 1428 7428
rect 1444 7397 1506 7428
rect 1575 7426 1624 7451
rect 1639 7426 1669 7442
rect 1538 7412 1568 7420
rect 1575 7418 1685 7426
rect 1538 7404 1583 7412
rect 1270 7386 1289 7388
rect 1304 7386 1350 7388
rect 1270 7370 1350 7386
rect 1377 7384 1412 7397
rect 1453 7394 1490 7397
rect 1453 7392 1495 7394
rect 1382 7381 1412 7384
rect 1391 7377 1398 7381
rect 1398 7376 1399 7377
rect 1357 7370 1367 7376
rect 1116 7362 1151 7370
rect 1116 7336 1117 7362
rect 1124 7336 1151 7362
rect 1059 7318 1089 7332
rect 1116 7328 1151 7336
rect 1153 7362 1194 7370
rect 1153 7336 1168 7362
rect 1175 7336 1194 7362
rect 1258 7358 1289 7370
rect 1304 7358 1407 7370
rect 1419 7360 1445 7386
rect 1460 7381 1490 7392
rect 1522 7388 1584 7404
rect 1522 7386 1568 7388
rect 1522 7370 1584 7386
rect 1596 7370 1602 7418
rect 1605 7410 1685 7418
rect 1605 7408 1624 7410
rect 1639 7408 1673 7410
rect 1605 7392 1685 7408
rect 1605 7370 1624 7392
rect 1639 7376 1669 7392
rect 1697 7386 1703 7460
rect 1706 7386 1725 7530
rect 1740 7386 1746 7530
rect 1755 7460 1768 7530
rect 1820 7526 1842 7530
rect 1813 7504 1842 7518
rect 1895 7504 1911 7518
rect 1949 7514 1955 7516
rect 1962 7514 2070 7530
rect 2077 7514 2083 7516
rect 2091 7514 2106 7530
rect 2172 7524 2191 7527
rect 1813 7502 1911 7504
rect 1938 7502 2106 7514
rect 2121 7504 2137 7518
rect 2172 7505 2194 7524
rect 2204 7518 2220 7519
rect 2203 7516 2220 7518
rect 2204 7511 2220 7516
rect 2194 7504 2200 7505
rect 2203 7504 2232 7511
rect 2121 7503 2232 7504
rect 2121 7502 2238 7503
rect 1797 7494 1848 7502
rect 1895 7494 1929 7502
rect 1797 7482 1822 7494
rect 1829 7482 1848 7494
rect 1902 7492 1929 7494
rect 1938 7492 2159 7502
rect 2194 7499 2200 7502
rect 1902 7488 2159 7492
rect 1797 7474 1848 7482
rect 1895 7474 2159 7488
rect 2203 7494 2238 7502
rect 1749 7426 1768 7460
rect 1813 7466 1842 7474
rect 1813 7460 1830 7466
rect 1813 7458 1847 7460
rect 1895 7458 1911 7474
rect 1912 7464 2120 7474
rect 2121 7464 2137 7474
rect 2185 7470 2200 7485
rect 2203 7482 2204 7494
rect 2211 7482 2238 7494
rect 2203 7474 2238 7482
rect 2203 7473 2232 7474
rect 1923 7460 2137 7464
rect 1938 7458 2137 7460
rect 2172 7460 2185 7470
rect 2203 7460 2220 7473
rect 2172 7458 2220 7460
rect 1814 7454 1847 7458
rect 1810 7452 1847 7454
rect 1810 7451 1877 7452
rect 1810 7446 1841 7451
rect 1847 7446 1877 7451
rect 1810 7442 1877 7446
rect 1783 7439 1877 7442
rect 1783 7432 1832 7439
rect 1783 7426 1813 7432
rect 1832 7427 1837 7432
rect 1749 7410 1829 7426
rect 1841 7418 1877 7439
rect 1938 7434 2127 7458
rect 2172 7457 2219 7458
rect 2185 7452 2219 7457
rect 1953 7431 2127 7434
rect 1946 7428 2127 7431
rect 2155 7451 2219 7452
rect 1749 7408 1768 7410
rect 1783 7408 1817 7410
rect 1749 7392 1829 7408
rect 1749 7386 1768 7392
rect 1465 7360 1568 7370
rect 1419 7358 1568 7360
rect 1589 7358 1624 7370
rect 1258 7356 1420 7358
rect 1270 7336 1289 7356
rect 1304 7354 1334 7356
rect 1153 7328 1194 7336
rect 1276 7332 1289 7336
rect 1341 7340 1420 7356
rect 1452 7356 1624 7358
rect 1452 7340 1531 7356
rect 1538 7354 1568 7356
rect 1116 7318 1145 7328
rect 1159 7318 1188 7328
rect 1203 7318 1233 7332
rect 1276 7318 1319 7332
rect 1341 7328 1531 7340
rect 1596 7336 1602 7356
rect 1326 7318 1356 7328
rect 1357 7318 1515 7328
rect 1519 7318 1549 7328
rect 1553 7318 1583 7332
rect 1611 7318 1624 7356
rect 1696 7370 1725 7386
rect 1739 7370 1768 7386
rect 1783 7376 1813 7392
rect 1841 7370 1847 7418
rect 1850 7412 1869 7418
rect 1884 7412 1914 7420
rect 1850 7404 1914 7412
rect 1850 7388 1930 7404
rect 1946 7397 2008 7428
rect 2024 7397 2086 7428
rect 2155 7426 2204 7451
rect 2219 7426 2249 7442
rect 2118 7412 2148 7420
rect 2155 7418 2265 7426
rect 2118 7404 2163 7412
rect 1850 7386 1869 7388
rect 1884 7386 1930 7388
rect 1850 7370 1930 7386
rect 1957 7384 1992 7397
rect 2033 7394 2070 7397
rect 2033 7392 2075 7394
rect 1962 7381 1992 7384
rect 1971 7377 1978 7381
rect 1978 7376 1979 7377
rect 1937 7370 1947 7376
rect 1696 7362 1731 7370
rect 1696 7336 1697 7362
rect 1704 7336 1731 7362
rect 1639 7318 1669 7332
rect 1696 7328 1731 7336
rect 1733 7362 1774 7370
rect 1733 7336 1748 7362
rect 1755 7336 1774 7362
rect 1838 7358 1869 7370
rect 1884 7358 1987 7370
rect 1999 7360 2025 7386
rect 2040 7381 2070 7392
rect 2102 7388 2164 7404
rect 2102 7386 2148 7388
rect 2102 7370 2164 7386
rect 2176 7370 2182 7418
rect 2185 7410 2265 7418
rect 2185 7408 2204 7410
rect 2219 7408 2253 7410
rect 2185 7392 2265 7408
rect 2185 7370 2204 7392
rect 2219 7376 2249 7392
rect 2277 7386 2283 7460
rect 2286 7386 2305 7530
rect 2320 7386 2326 7530
rect 2335 7460 2348 7530
rect 2400 7526 2422 7530
rect 2393 7504 2422 7518
rect 2475 7504 2491 7518
rect 2529 7514 2535 7516
rect 2542 7514 2650 7530
rect 2657 7514 2663 7516
rect 2671 7514 2686 7530
rect 2752 7524 2771 7527
rect 2393 7502 2491 7504
rect 2518 7502 2686 7514
rect 2701 7504 2717 7518
rect 2752 7505 2774 7524
rect 2784 7518 2800 7519
rect 2783 7516 2800 7518
rect 2784 7511 2800 7516
rect 2774 7504 2780 7505
rect 2783 7504 2812 7511
rect 2701 7503 2812 7504
rect 2701 7502 2818 7503
rect 2377 7494 2428 7502
rect 2475 7494 2509 7502
rect 2377 7482 2402 7494
rect 2409 7482 2428 7494
rect 2482 7492 2509 7494
rect 2518 7492 2739 7502
rect 2774 7499 2780 7502
rect 2482 7488 2739 7492
rect 2377 7474 2428 7482
rect 2475 7474 2739 7488
rect 2783 7494 2818 7502
rect 2329 7426 2348 7460
rect 2393 7466 2422 7474
rect 2393 7460 2410 7466
rect 2393 7458 2427 7460
rect 2475 7458 2491 7474
rect 2492 7464 2700 7474
rect 2701 7464 2717 7474
rect 2765 7470 2780 7485
rect 2783 7482 2784 7494
rect 2791 7482 2818 7494
rect 2783 7474 2818 7482
rect 2783 7473 2812 7474
rect 2503 7460 2717 7464
rect 2518 7458 2717 7460
rect 2752 7460 2765 7470
rect 2783 7460 2800 7473
rect 2752 7458 2800 7460
rect 2394 7454 2427 7458
rect 2390 7452 2427 7454
rect 2390 7451 2457 7452
rect 2390 7446 2421 7451
rect 2427 7446 2457 7451
rect 2390 7442 2457 7446
rect 2363 7439 2457 7442
rect 2363 7432 2412 7439
rect 2363 7426 2393 7432
rect 2412 7427 2417 7432
rect 2329 7410 2409 7426
rect 2421 7418 2457 7439
rect 2518 7434 2707 7458
rect 2752 7457 2799 7458
rect 2765 7452 2799 7457
rect 2533 7431 2707 7434
rect 2526 7428 2707 7431
rect 2735 7451 2799 7452
rect 2329 7408 2348 7410
rect 2363 7408 2397 7410
rect 2329 7392 2409 7408
rect 2329 7386 2348 7392
rect 2045 7360 2148 7370
rect 1999 7358 2148 7360
rect 2169 7358 2204 7370
rect 1838 7356 2000 7358
rect 1850 7336 1869 7356
rect 1884 7354 1914 7356
rect 1733 7328 1774 7336
rect 1856 7332 1869 7336
rect 1921 7340 2000 7356
rect 2032 7356 2204 7358
rect 2032 7340 2111 7356
rect 2118 7354 2148 7356
rect 1696 7318 1725 7328
rect 1739 7318 1768 7328
rect 1783 7318 1813 7332
rect 1856 7318 1899 7332
rect 1921 7328 2111 7340
rect 2176 7336 2182 7356
rect 1906 7318 1936 7328
rect 1937 7318 2095 7328
rect 2099 7318 2129 7328
rect 2133 7318 2163 7332
rect 2191 7318 2204 7356
rect 2276 7370 2305 7386
rect 2319 7370 2348 7386
rect 2363 7376 2393 7392
rect 2421 7370 2427 7418
rect 2430 7412 2449 7418
rect 2464 7412 2494 7420
rect 2430 7404 2494 7412
rect 2430 7388 2510 7404
rect 2526 7397 2588 7428
rect 2604 7397 2666 7428
rect 2735 7426 2784 7451
rect 2799 7426 2829 7442
rect 2698 7412 2728 7420
rect 2735 7418 2845 7426
rect 2698 7404 2743 7412
rect 2430 7386 2449 7388
rect 2464 7386 2510 7388
rect 2430 7370 2510 7386
rect 2537 7384 2572 7397
rect 2613 7394 2650 7397
rect 2613 7392 2655 7394
rect 2542 7381 2572 7384
rect 2551 7377 2558 7381
rect 2558 7376 2559 7377
rect 2517 7370 2527 7376
rect 2276 7362 2311 7370
rect 2276 7336 2277 7362
rect 2284 7336 2311 7362
rect 2219 7318 2249 7332
rect 2276 7328 2311 7336
rect 2313 7362 2354 7370
rect 2313 7336 2328 7362
rect 2335 7336 2354 7362
rect 2418 7358 2449 7370
rect 2464 7358 2567 7370
rect 2579 7360 2605 7386
rect 2620 7381 2650 7392
rect 2682 7388 2744 7404
rect 2682 7386 2728 7388
rect 2682 7370 2744 7386
rect 2756 7370 2762 7418
rect 2765 7410 2845 7418
rect 2765 7408 2784 7410
rect 2799 7408 2833 7410
rect 2765 7392 2845 7408
rect 2765 7370 2784 7392
rect 2799 7376 2829 7392
rect 2857 7386 2863 7460
rect 2866 7386 2885 7530
rect 2900 7386 2906 7530
rect 2915 7460 2928 7530
rect 2980 7526 3002 7530
rect 2973 7504 3002 7518
rect 3055 7504 3071 7518
rect 3109 7514 3115 7516
rect 3122 7514 3230 7530
rect 3237 7514 3243 7516
rect 3251 7514 3266 7530
rect 3332 7524 3351 7527
rect 2973 7502 3071 7504
rect 3098 7502 3266 7514
rect 3281 7504 3297 7518
rect 3332 7505 3354 7524
rect 3364 7518 3380 7519
rect 3363 7516 3380 7518
rect 3364 7511 3380 7516
rect 3354 7504 3360 7505
rect 3363 7504 3392 7511
rect 3281 7503 3392 7504
rect 3281 7502 3398 7503
rect 2957 7494 3008 7502
rect 3055 7494 3089 7502
rect 2957 7482 2982 7494
rect 2989 7482 3008 7494
rect 3062 7492 3089 7494
rect 3098 7492 3319 7502
rect 3354 7499 3360 7502
rect 3062 7488 3319 7492
rect 2957 7474 3008 7482
rect 3055 7474 3319 7488
rect 3363 7494 3398 7502
rect 2909 7426 2928 7460
rect 2973 7466 3002 7474
rect 2973 7460 2990 7466
rect 2973 7458 3007 7460
rect 3055 7458 3071 7474
rect 3072 7464 3280 7474
rect 3281 7464 3297 7474
rect 3345 7470 3360 7485
rect 3363 7482 3364 7494
rect 3371 7482 3398 7494
rect 3363 7474 3398 7482
rect 3363 7473 3392 7474
rect 3083 7460 3297 7464
rect 3098 7458 3297 7460
rect 3332 7460 3345 7470
rect 3363 7460 3380 7473
rect 3332 7458 3380 7460
rect 2974 7454 3007 7458
rect 2970 7452 3007 7454
rect 2970 7451 3037 7452
rect 2970 7446 3001 7451
rect 3007 7446 3037 7451
rect 2970 7442 3037 7446
rect 2943 7439 3037 7442
rect 2943 7432 2992 7439
rect 2943 7426 2973 7432
rect 2992 7427 2997 7432
rect 2909 7410 2989 7426
rect 3001 7418 3037 7439
rect 3098 7434 3287 7458
rect 3332 7457 3379 7458
rect 3345 7452 3379 7457
rect 3113 7431 3287 7434
rect 3106 7428 3287 7431
rect 3315 7451 3379 7452
rect 2909 7408 2928 7410
rect 2943 7408 2977 7410
rect 2909 7392 2989 7408
rect 2909 7386 2928 7392
rect 2625 7360 2728 7370
rect 2579 7358 2728 7360
rect 2749 7358 2784 7370
rect 2418 7356 2580 7358
rect 2430 7336 2449 7356
rect 2464 7354 2494 7356
rect 2313 7328 2354 7336
rect 2436 7332 2449 7336
rect 2501 7340 2580 7356
rect 2612 7356 2784 7358
rect 2612 7340 2691 7356
rect 2698 7354 2728 7356
rect 2276 7318 2305 7328
rect 2319 7318 2348 7328
rect 2363 7318 2393 7332
rect 2436 7318 2479 7332
rect 2501 7328 2691 7340
rect 2756 7336 2762 7356
rect 2486 7318 2516 7328
rect 2517 7318 2675 7328
rect 2679 7318 2709 7328
rect 2713 7318 2743 7332
rect 2771 7318 2784 7356
rect 2856 7370 2885 7386
rect 2899 7370 2928 7386
rect 2943 7376 2973 7392
rect 3001 7370 3007 7418
rect 3010 7412 3029 7418
rect 3044 7412 3074 7420
rect 3010 7404 3074 7412
rect 3010 7388 3090 7404
rect 3106 7397 3168 7428
rect 3184 7397 3246 7428
rect 3315 7426 3364 7451
rect 3379 7426 3409 7442
rect 3278 7412 3308 7420
rect 3315 7418 3425 7426
rect 3278 7404 3323 7412
rect 3010 7386 3029 7388
rect 3044 7386 3090 7388
rect 3010 7370 3090 7386
rect 3117 7384 3152 7397
rect 3193 7394 3230 7397
rect 3193 7392 3235 7394
rect 3122 7381 3152 7384
rect 3131 7377 3138 7381
rect 3138 7376 3139 7377
rect 3097 7370 3107 7376
rect 2856 7362 2891 7370
rect 2856 7336 2857 7362
rect 2864 7336 2891 7362
rect 2799 7318 2829 7332
rect 2856 7328 2891 7336
rect 2893 7362 2934 7370
rect 2893 7336 2908 7362
rect 2915 7336 2934 7362
rect 2998 7358 3029 7370
rect 3044 7358 3147 7370
rect 3159 7360 3185 7386
rect 3200 7381 3230 7392
rect 3262 7388 3324 7404
rect 3262 7386 3308 7388
rect 3262 7370 3324 7386
rect 3336 7370 3342 7418
rect 3345 7410 3425 7418
rect 3345 7408 3364 7410
rect 3379 7408 3413 7410
rect 3345 7392 3425 7408
rect 3345 7370 3364 7392
rect 3379 7376 3409 7392
rect 3437 7386 3443 7460
rect 3446 7386 3465 7530
rect 3480 7386 3486 7530
rect 3495 7460 3508 7530
rect 3560 7526 3582 7530
rect 3553 7504 3582 7518
rect 3635 7504 3651 7518
rect 3689 7514 3695 7516
rect 3702 7514 3810 7530
rect 3817 7514 3823 7516
rect 3831 7514 3846 7530
rect 3912 7524 3931 7527
rect 3553 7502 3651 7504
rect 3678 7502 3846 7514
rect 3861 7504 3877 7518
rect 3912 7505 3934 7524
rect 3944 7518 3960 7519
rect 3943 7516 3960 7518
rect 3944 7511 3960 7516
rect 3934 7504 3940 7505
rect 3943 7504 3972 7511
rect 3861 7503 3972 7504
rect 3861 7502 3978 7503
rect 3537 7494 3588 7502
rect 3635 7494 3669 7502
rect 3537 7482 3562 7494
rect 3569 7482 3588 7494
rect 3642 7492 3669 7494
rect 3678 7492 3899 7502
rect 3934 7499 3940 7502
rect 3642 7488 3899 7492
rect 3537 7474 3588 7482
rect 3635 7474 3899 7488
rect 3943 7494 3978 7502
rect 3489 7426 3508 7460
rect 3553 7466 3582 7474
rect 3553 7460 3570 7466
rect 3553 7458 3587 7460
rect 3635 7458 3651 7474
rect 3652 7464 3860 7474
rect 3861 7464 3877 7474
rect 3925 7470 3940 7485
rect 3943 7482 3944 7494
rect 3951 7482 3978 7494
rect 3943 7474 3978 7482
rect 3943 7473 3972 7474
rect 3663 7460 3877 7464
rect 3678 7458 3877 7460
rect 3912 7460 3925 7470
rect 3943 7460 3960 7473
rect 3912 7458 3960 7460
rect 3554 7454 3587 7458
rect 3550 7452 3587 7454
rect 3550 7451 3617 7452
rect 3550 7446 3581 7451
rect 3587 7446 3617 7451
rect 3550 7442 3617 7446
rect 3523 7439 3617 7442
rect 3523 7432 3572 7439
rect 3523 7426 3553 7432
rect 3572 7427 3577 7432
rect 3489 7410 3569 7426
rect 3581 7418 3617 7439
rect 3678 7434 3867 7458
rect 3912 7457 3959 7458
rect 3925 7452 3959 7457
rect 3693 7431 3867 7434
rect 3686 7428 3867 7431
rect 3895 7451 3959 7452
rect 3489 7408 3508 7410
rect 3523 7408 3557 7410
rect 3489 7392 3569 7408
rect 3489 7386 3508 7392
rect 3205 7360 3308 7370
rect 3159 7358 3308 7360
rect 3329 7358 3364 7370
rect 2998 7356 3160 7358
rect 3010 7336 3029 7356
rect 3044 7354 3074 7356
rect 2893 7328 2934 7336
rect 3016 7332 3029 7336
rect 3081 7340 3160 7356
rect 3192 7356 3364 7358
rect 3192 7340 3271 7356
rect 3278 7354 3308 7356
rect 2856 7318 2885 7328
rect 2899 7318 2928 7328
rect 2943 7318 2973 7332
rect 3016 7318 3059 7332
rect 3081 7328 3271 7340
rect 3336 7336 3342 7356
rect 3066 7318 3096 7328
rect 3097 7318 3255 7328
rect 3259 7318 3289 7328
rect 3293 7318 3323 7332
rect 3351 7318 3364 7356
rect 3436 7370 3465 7386
rect 3479 7370 3508 7386
rect 3523 7376 3553 7392
rect 3581 7370 3587 7418
rect 3590 7412 3609 7418
rect 3624 7412 3654 7420
rect 3590 7404 3654 7412
rect 3590 7388 3670 7404
rect 3686 7397 3748 7428
rect 3764 7397 3826 7428
rect 3895 7426 3944 7451
rect 3959 7426 3989 7442
rect 3858 7412 3888 7420
rect 3895 7418 4005 7426
rect 3858 7404 3903 7412
rect 3590 7386 3609 7388
rect 3624 7386 3670 7388
rect 3590 7370 3670 7386
rect 3697 7384 3732 7397
rect 3773 7394 3810 7397
rect 3773 7392 3815 7394
rect 3702 7381 3732 7384
rect 3711 7377 3718 7381
rect 3718 7376 3719 7377
rect 3677 7370 3687 7376
rect 3436 7362 3471 7370
rect 3436 7336 3437 7362
rect 3444 7336 3471 7362
rect 3379 7318 3409 7332
rect 3436 7328 3471 7336
rect 3473 7362 3514 7370
rect 3473 7336 3488 7362
rect 3495 7336 3514 7362
rect 3578 7358 3609 7370
rect 3624 7358 3727 7370
rect 3739 7360 3765 7386
rect 3780 7381 3810 7392
rect 3842 7388 3904 7404
rect 3842 7386 3888 7388
rect 3842 7370 3904 7386
rect 3916 7370 3922 7418
rect 3925 7410 4005 7418
rect 3925 7408 3944 7410
rect 3959 7408 3993 7410
rect 3925 7392 4005 7408
rect 3925 7370 3944 7392
rect 3959 7376 3989 7392
rect 4017 7386 4023 7460
rect 4026 7386 4045 7530
rect 4060 7386 4066 7530
rect 4075 7460 4088 7530
rect 4140 7526 4162 7530
rect 4133 7504 4162 7518
rect 4215 7504 4231 7518
rect 4269 7514 4275 7516
rect 4282 7514 4390 7530
rect 4397 7514 4403 7516
rect 4411 7514 4426 7530
rect 4492 7524 4511 7527
rect 4133 7502 4231 7504
rect 4258 7502 4426 7514
rect 4441 7504 4457 7518
rect 4492 7505 4514 7524
rect 4524 7518 4540 7519
rect 4523 7516 4540 7518
rect 4524 7511 4540 7516
rect 4514 7504 4520 7505
rect 4523 7504 4552 7511
rect 4441 7503 4552 7504
rect 4441 7502 4558 7503
rect 4117 7494 4168 7502
rect 4215 7494 4249 7502
rect 4117 7482 4142 7494
rect 4149 7482 4168 7494
rect 4222 7492 4249 7494
rect 4258 7492 4479 7502
rect 4514 7499 4520 7502
rect 4222 7488 4479 7492
rect 4117 7474 4168 7482
rect 4215 7474 4479 7488
rect 4523 7494 4558 7502
rect 4069 7426 4088 7460
rect 4133 7466 4162 7474
rect 4133 7460 4150 7466
rect 4133 7458 4167 7460
rect 4215 7458 4231 7474
rect 4232 7464 4440 7474
rect 4441 7464 4457 7474
rect 4505 7470 4520 7485
rect 4523 7482 4524 7494
rect 4531 7482 4558 7494
rect 4523 7474 4558 7482
rect 4523 7473 4552 7474
rect 4243 7460 4457 7464
rect 4258 7458 4457 7460
rect 4492 7460 4505 7470
rect 4523 7460 4540 7473
rect 4492 7458 4540 7460
rect 4134 7454 4167 7458
rect 4130 7452 4167 7454
rect 4130 7451 4197 7452
rect 4130 7446 4161 7451
rect 4167 7446 4197 7451
rect 4130 7442 4197 7446
rect 4103 7439 4197 7442
rect 4103 7432 4152 7439
rect 4103 7426 4133 7432
rect 4152 7427 4157 7432
rect 4069 7410 4149 7426
rect 4161 7418 4197 7439
rect 4258 7434 4447 7458
rect 4492 7457 4539 7458
rect 4505 7452 4539 7457
rect 4273 7431 4447 7434
rect 4266 7428 4447 7431
rect 4475 7451 4539 7452
rect 4069 7408 4088 7410
rect 4103 7408 4137 7410
rect 4069 7392 4149 7408
rect 4069 7386 4088 7392
rect 3785 7360 3888 7370
rect 3739 7358 3888 7360
rect 3909 7358 3944 7370
rect 3578 7356 3740 7358
rect 3590 7336 3609 7356
rect 3624 7354 3654 7356
rect 3473 7328 3514 7336
rect 3596 7332 3609 7336
rect 3661 7340 3740 7356
rect 3772 7356 3944 7358
rect 3772 7340 3851 7356
rect 3858 7354 3888 7356
rect 3436 7318 3465 7328
rect 3479 7318 3508 7328
rect 3523 7318 3553 7332
rect 3596 7318 3639 7332
rect 3661 7328 3851 7340
rect 3916 7336 3922 7356
rect 3646 7318 3676 7328
rect 3677 7318 3835 7328
rect 3839 7318 3869 7328
rect 3873 7318 3903 7332
rect 3931 7318 3944 7356
rect 4016 7370 4045 7386
rect 4059 7370 4088 7386
rect 4103 7376 4133 7392
rect 4161 7370 4167 7418
rect 4170 7412 4189 7418
rect 4204 7412 4234 7420
rect 4170 7404 4234 7412
rect 4170 7388 4250 7404
rect 4266 7397 4328 7428
rect 4344 7397 4406 7428
rect 4475 7426 4524 7451
rect 4539 7426 4569 7442
rect 4438 7412 4468 7420
rect 4475 7418 4585 7426
rect 4438 7404 4483 7412
rect 4170 7386 4189 7388
rect 4204 7386 4250 7388
rect 4170 7370 4250 7386
rect 4277 7384 4312 7397
rect 4353 7394 4390 7397
rect 4353 7392 4395 7394
rect 4282 7381 4312 7384
rect 4291 7377 4298 7381
rect 4298 7376 4299 7377
rect 4257 7370 4267 7376
rect 4016 7362 4051 7370
rect 4016 7336 4017 7362
rect 4024 7336 4051 7362
rect 3959 7318 3989 7332
rect 4016 7328 4051 7336
rect 4053 7362 4094 7370
rect 4053 7336 4068 7362
rect 4075 7336 4094 7362
rect 4158 7358 4189 7370
rect 4204 7358 4307 7370
rect 4319 7360 4345 7386
rect 4360 7381 4390 7392
rect 4422 7388 4484 7404
rect 4422 7386 4468 7388
rect 4422 7370 4484 7386
rect 4496 7370 4502 7418
rect 4505 7410 4585 7418
rect 4505 7408 4524 7410
rect 4539 7408 4573 7410
rect 4505 7392 4585 7408
rect 4505 7370 4524 7392
rect 4539 7376 4569 7392
rect 4597 7386 4603 7460
rect 4606 7386 4625 7530
rect 4640 7386 4646 7530
rect 4655 7460 4668 7530
rect 4720 7526 4742 7530
rect 4713 7504 4742 7518
rect 4795 7504 4811 7518
rect 4849 7514 4855 7516
rect 4862 7514 4970 7530
rect 4977 7514 4983 7516
rect 4991 7514 5006 7530
rect 5072 7524 5091 7527
rect 4713 7502 4811 7504
rect 4838 7502 5006 7514
rect 5021 7504 5037 7518
rect 5072 7505 5094 7524
rect 5104 7518 5120 7519
rect 5103 7516 5120 7518
rect 5104 7511 5120 7516
rect 5094 7504 5100 7505
rect 5103 7504 5132 7511
rect 5021 7503 5132 7504
rect 5021 7502 5138 7503
rect 4697 7494 4748 7502
rect 4795 7494 4829 7502
rect 4697 7482 4722 7494
rect 4729 7482 4748 7494
rect 4802 7492 4829 7494
rect 4838 7492 5059 7502
rect 5094 7499 5100 7502
rect 4802 7488 5059 7492
rect 4697 7474 4748 7482
rect 4795 7474 5059 7488
rect 5103 7494 5138 7502
rect 4649 7426 4668 7460
rect 4713 7466 4742 7474
rect 4713 7460 4730 7466
rect 4713 7458 4747 7460
rect 4795 7458 4811 7474
rect 4812 7464 5020 7474
rect 5021 7464 5037 7474
rect 5085 7470 5100 7485
rect 5103 7482 5104 7494
rect 5111 7482 5138 7494
rect 5103 7474 5138 7482
rect 5103 7473 5132 7474
rect 4823 7460 5037 7464
rect 4838 7458 5037 7460
rect 5072 7460 5085 7470
rect 5103 7460 5120 7473
rect 5072 7458 5120 7460
rect 4714 7454 4747 7458
rect 4710 7452 4747 7454
rect 4710 7451 4777 7452
rect 4710 7446 4741 7451
rect 4747 7446 4777 7451
rect 4710 7442 4777 7446
rect 4683 7439 4777 7442
rect 4683 7432 4732 7439
rect 4683 7426 4713 7432
rect 4732 7427 4737 7432
rect 4649 7410 4729 7426
rect 4741 7418 4777 7439
rect 4838 7434 5027 7458
rect 5072 7457 5119 7458
rect 5085 7452 5119 7457
rect 4853 7431 5027 7434
rect 4846 7428 5027 7431
rect 5055 7451 5119 7452
rect 4649 7408 4668 7410
rect 4683 7408 4717 7410
rect 4649 7392 4729 7408
rect 4649 7386 4668 7392
rect 4365 7360 4468 7370
rect 4319 7358 4468 7360
rect 4489 7358 4524 7370
rect 4158 7356 4320 7358
rect 4170 7336 4189 7356
rect 4204 7354 4234 7356
rect 4053 7328 4094 7336
rect 4176 7332 4189 7336
rect 4241 7340 4320 7356
rect 4352 7356 4524 7358
rect 4352 7340 4431 7356
rect 4438 7354 4468 7356
rect 4016 7318 4045 7328
rect 4059 7318 4088 7328
rect 4103 7318 4133 7332
rect 4176 7318 4219 7332
rect 4241 7328 4431 7340
rect 4496 7336 4502 7356
rect 4226 7318 4256 7328
rect 4257 7318 4415 7328
rect 4419 7318 4449 7328
rect 4453 7318 4483 7332
rect 4511 7318 4524 7356
rect 4596 7370 4625 7386
rect 4639 7370 4668 7386
rect 4683 7376 4713 7392
rect 4741 7370 4747 7418
rect 4750 7412 4769 7418
rect 4784 7412 4814 7420
rect 4750 7404 4814 7412
rect 4750 7388 4830 7404
rect 4846 7397 4908 7428
rect 4924 7397 4986 7428
rect 5055 7426 5104 7451
rect 5119 7426 5149 7442
rect 5018 7412 5048 7420
rect 5055 7418 5165 7426
rect 5018 7404 5063 7412
rect 4750 7386 4769 7388
rect 4784 7386 4830 7388
rect 4750 7370 4830 7386
rect 4857 7384 4892 7397
rect 4933 7394 4970 7397
rect 4933 7392 4975 7394
rect 4862 7381 4892 7384
rect 4871 7377 4878 7381
rect 4878 7376 4879 7377
rect 4837 7370 4847 7376
rect 4596 7362 4631 7370
rect 4596 7336 4597 7362
rect 4604 7336 4631 7362
rect 4539 7318 4569 7332
rect 4596 7328 4631 7336
rect 4633 7362 4674 7370
rect 4633 7336 4648 7362
rect 4655 7336 4674 7362
rect 4738 7358 4769 7370
rect 4784 7358 4887 7370
rect 4899 7360 4925 7386
rect 4940 7381 4970 7392
rect 5002 7388 5064 7404
rect 5002 7386 5048 7388
rect 5002 7370 5064 7386
rect 5076 7370 5082 7418
rect 5085 7410 5165 7418
rect 5085 7408 5104 7410
rect 5119 7408 5153 7410
rect 5085 7392 5165 7408
rect 5085 7370 5104 7392
rect 5119 7376 5149 7392
rect 5177 7386 5183 7460
rect 5186 7386 5205 7530
rect 5220 7386 5226 7530
rect 5235 7460 5248 7530
rect 5300 7526 5322 7530
rect 5293 7504 5322 7518
rect 5375 7504 5391 7518
rect 5429 7514 5435 7516
rect 5442 7514 5550 7530
rect 5557 7514 5563 7516
rect 5571 7514 5586 7530
rect 5652 7524 5671 7527
rect 5293 7502 5391 7504
rect 5418 7502 5586 7514
rect 5601 7504 5617 7518
rect 5652 7505 5674 7524
rect 5684 7518 5700 7519
rect 5683 7516 5700 7518
rect 5684 7511 5700 7516
rect 5674 7504 5680 7505
rect 5683 7504 5712 7511
rect 5601 7503 5712 7504
rect 5601 7502 5718 7503
rect 5277 7494 5328 7502
rect 5375 7494 5409 7502
rect 5277 7482 5302 7494
rect 5309 7482 5328 7494
rect 5382 7492 5409 7494
rect 5418 7492 5639 7502
rect 5674 7499 5680 7502
rect 5382 7488 5639 7492
rect 5277 7474 5328 7482
rect 5375 7474 5639 7488
rect 5683 7494 5718 7502
rect 5229 7426 5248 7460
rect 5293 7466 5322 7474
rect 5293 7460 5310 7466
rect 5293 7458 5327 7460
rect 5375 7458 5391 7474
rect 5392 7464 5600 7474
rect 5601 7464 5617 7474
rect 5665 7470 5680 7485
rect 5683 7482 5684 7494
rect 5691 7482 5718 7494
rect 5683 7474 5718 7482
rect 5683 7473 5712 7474
rect 5403 7460 5617 7464
rect 5418 7458 5617 7460
rect 5652 7460 5665 7470
rect 5683 7460 5700 7473
rect 5652 7458 5700 7460
rect 5294 7454 5327 7458
rect 5290 7452 5327 7454
rect 5290 7451 5357 7452
rect 5290 7446 5321 7451
rect 5327 7446 5357 7451
rect 5290 7442 5357 7446
rect 5263 7439 5357 7442
rect 5263 7432 5312 7439
rect 5263 7426 5293 7432
rect 5312 7427 5317 7432
rect 5229 7410 5309 7426
rect 5321 7418 5357 7439
rect 5418 7434 5607 7458
rect 5652 7457 5699 7458
rect 5665 7452 5699 7457
rect 5433 7431 5607 7434
rect 5426 7428 5607 7431
rect 5635 7451 5699 7452
rect 5229 7408 5248 7410
rect 5263 7408 5297 7410
rect 5229 7392 5309 7408
rect 5229 7386 5248 7392
rect 4945 7360 5048 7370
rect 4899 7358 5048 7360
rect 5069 7358 5104 7370
rect 4738 7356 4900 7358
rect 4750 7336 4769 7356
rect 4784 7354 4814 7356
rect 4633 7328 4674 7336
rect 4756 7332 4769 7336
rect 4821 7340 4900 7356
rect 4932 7356 5104 7358
rect 4932 7340 5011 7356
rect 5018 7354 5048 7356
rect 4596 7318 4625 7328
rect 4639 7318 4668 7328
rect 4683 7318 4713 7332
rect 4756 7318 4799 7332
rect 4821 7328 5011 7340
rect 5076 7336 5082 7356
rect 4806 7318 4836 7328
rect 4837 7318 4995 7328
rect 4999 7318 5029 7328
rect 5033 7318 5063 7332
rect 5091 7318 5104 7356
rect 5176 7370 5205 7386
rect 5219 7370 5248 7386
rect 5263 7376 5293 7392
rect 5321 7370 5327 7418
rect 5330 7412 5349 7418
rect 5364 7412 5394 7420
rect 5330 7404 5394 7412
rect 5330 7388 5410 7404
rect 5426 7397 5488 7428
rect 5504 7397 5566 7428
rect 5635 7426 5684 7451
rect 5699 7426 5729 7442
rect 5598 7412 5628 7420
rect 5635 7418 5745 7426
rect 5598 7404 5643 7412
rect 5330 7386 5349 7388
rect 5364 7386 5410 7388
rect 5330 7370 5410 7386
rect 5437 7384 5472 7397
rect 5513 7394 5550 7397
rect 5513 7392 5555 7394
rect 5442 7381 5472 7384
rect 5451 7377 5458 7381
rect 5458 7376 5459 7377
rect 5417 7370 5427 7376
rect 5176 7362 5211 7370
rect 5176 7336 5177 7362
rect 5184 7336 5211 7362
rect 5119 7318 5149 7332
rect 5176 7328 5211 7336
rect 5213 7362 5254 7370
rect 5213 7336 5228 7362
rect 5235 7336 5254 7362
rect 5318 7358 5349 7370
rect 5364 7358 5467 7370
rect 5479 7360 5505 7386
rect 5520 7381 5550 7392
rect 5582 7388 5644 7404
rect 5582 7386 5628 7388
rect 5582 7370 5644 7386
rect 5656 7370 5662 7418
rect 5665 7410 5745 7418
rect 5665 7408 5684 7410
rect 5699 7408 5733 7410
rect 5665 7392 5745 7408
rect 5665 7370 5684 7392
rect 5699 7376 5729 7392
rect 5757 7386 5763 7460
rect 5766 7386 5785 7530
rect 5800 7386 5806 7530
rect 5815 7460 5828 7530
rect 5880 7526 5902 7530
rect 5873 7504 5902 7518
rect 5955 7504 5971 7518
rect 6009 7514 6015 7516
rect 6022 7514 6130 7530
rect 6137 7514 6143 7516
rect 6151 7514 6166 7530
rect 6232 7524 6251 7527
rect 5873 7502 5971 7504
rect 5998 7502 6166 7514
rect 6181 7504 6197 7518
rect 6232 7505 6254 7524
rect 6264 7518 6280 7519
rect 6263 7516 6280 7518
rect 6264 7511 6280 7516
rect 6254 7504 6260 7505
rect 6263 7504 6292 7511
rect 6181 7503 6292 7504
rect 6181 7502 6298 7503
rect 5857 7494 5908 7502
rect 5955 7494 5989 7502
rect 5857 7482 5882 7494
rect 5889 7482 5908 7494
rect 5962 7492 5989 7494
rect 5998 7492 6219 7502
rect 6254 7499 6260 7502
rect 5962 7488 6219 7492
rect 5857 7474 5908 7482
rect 5955 7474 6219 7488
rect 6263 7494 6298 7502
rect 5809 7426 5828 7460
rect 5873 7466 5902 7474
rect 5873 7460 5890 7466
rect 5873 7458 5907 7460
rect 5955 7458 5971 7474
rect 5972 7464 6180 7474
rect 6181 7464 6197 7474
rect 6245 7470 6260 7485
rect 6263 7482 6264 7494
rect 6271 7482 6298 7494
rect 6263 7474 6298 7482
rect 6263 7473 6292 7474
rect 5983 7460 6197 7464
rect 5998 7458 6197 7460
rect 6232 7460 6245 7470
rect 6263 7460 6280 7473
rect 6232 7458 6280 7460
rect 5874 7454 5907 7458
rect 5870 7452 5907 7454
rect 5870 7451 5937 7452
rect 5870 7446 5901 7451
rect 5907 7446 5937 7451
rect 5870 7442 5937 7446
rect 5843 7439 5937 7442
rect 5843 7432 5892 7439
rect 5843 7426 5873 7432
rect 5892 7427 5897 7432
rect 5809 7410 5889 7426
rect 5901 7418 5937 7439
rect 5998 7434 6187 7458
rect 6232 7457 6279 7458
rect 6245 7452 6279 7457
rect 6013 7431 6187 7434
rect 6006 7428 6187 7431
rect 6215 7451 6279 7452
rect 5809 7408 5828 7410
rect 5843 7408 5877 7410
rect 5809 7392 5889 7408
rect 5809 7386 5828 7392
rect 5525 7360 5628 7370
rect 5479 7358 5628 7360
rect 5649 7358 5684 7370
rect 5318 7356 5480 7358
rect 5330 7336 5349 7356
rect 5364 7354 5394 7356
rect 5213 7328 5254 7336
rect 5336 7332 5349 7336
rect 5401 7340 5480 7356
rect 5512 7356 5684 7358
rect 5512 7340 5591 7356
rect 5598 7354 5628 7356
rect 5176 7318 5205 7328
rect 5219 7318 5248 7328
rect 5263 7318 5293 7332
rect 5336 7318 5379 7332
rect 5401 7328 5591 7340
rect 5656 7336 5662 7356
rect 5386 7318 5416 7328
rect 5417 7318 5575 7328
rect 5579 7318 5609 7328
rect 5613 7318 5643 7332
rect 5671 7318 5684 7356
rect 5756 7370 5785 7386
rect 5799 7370 5828 7386
rect 5843 7376 5873 7392
rect 5901 7370 5907 7418
rect 5910 7412 5929 7418
rect 5944 7412 5974 7420
rect 5910 7404 5974 7412
rect 5910 7388 5990 7404
rect 6006 7397 6068 7428
rect 6084 7397 6146 7428
rect 6215 7426 6264 7451
rect 6279 7426 6309 7442
rect 6178 7412 6208 7420
rect 6215 7418 6325 7426
rect 6178 7404 6223 7412
rect 5910 7386 5929 7388
rect 5944 7386 5990 7388
rect 5910 7370 5990 7386
rect 6017 7384 6052 7397
rect 6093 7394 6130 7397
rect 6093 7392 6135 7394
rect 6022 7381 6052 7384
rect 6031 7377 6038 7381
rect 6038 7376 6039 7377
rect 5997 7370 6007 7376
rect 5756 7362 5791 7370
rect 5756 7336 5757 7362
rect 5764 7336 5791 7362
rect 5699 7318 5729 7332
rect 5756 7328 5791 7336
rect 5793 7362 5834 7370
rect 5793 7336 5808 7362
rect 5815 7336 5834 7362
rect 5898 7358 5929 7370
rect 5944 7358 6047 7370
rect 6059 7360 6085 7386
rect 6100 7381 6130 7392
rect 6162 7388 6224 7404
rect 6162 7386 6208 7388
rect 6162 7370 6224 7386
rect 6236 7370 6242 7418
rect 6245 7410 6325 7418
rect 6245 7408 6264 7410
rect 6279 7408 6313 7410
rect 6245 7392 6325 7408
rect 6245 7370 6264 7392
rect 6279 7376 6309 7392
rect 6337 7386 6343 7460
rect 6346 7386 6365 7530
rect 6380 7386 6386 7530
rect 6395 7460 6408 7530
rect 6460 7526 6482 7530
rect 6453 7504 6482 7518
rect 6535 7504 6551 7518
rect 6589 7514 6595 7516
rect 6602 7514 6710 7530
rect 6717 7514 6723 7516
rect 6731 7514 6746 7530
rect 6812 7524 6831 7527
rect 6453 7502 6551 7504
rect 6578 7502 6746 7514
rect 6761 7504 6777 7518
rect 6812 7505 6834 7524
rect 6844 7518 6860 7519
rect 6843 7516 6860 7518
rect 6844 7511 6860 7516
rect 6834 7504 6840 7505
rect 6843 7504 6872 7511
rect 6761 7503 6872 7504
rect 6761 7502 6878 7503
rect 6437 7494 6488 7502
rect 6535 7494 6569 7502
rect 6437 7482 6462 7494
rect 6469 7482 6488 7494
rect 6542 7492 6569 7494
rect 6578 7492 6799 7502
rect 6834 7499 6840 7502
rect 6542 7488 6799 7492
rect 6437 7474 6488 7482
rect 6535 7474 6799 7488
rect 6843 7494 6878 7502
rect 6389 7426 6408 7460
rect 6453 7466 6482 7474
rect 6453 7460 6470 7466
rect 6453 7458 6487 7460
rect 6535 7458 6551 7474
rect 6552 7464 6760 7474
rect 6761 7464 6777 7474
rect 6825 7470 6840 7485
rect 6843 7482 6844 7494
rect 6851 7482 6878 7494
rect 6843 7474 6878 7482
rect 6843 7473 6872 7474
rect 6563 7460 6777 7464
rect 6578 7458 6777 7460
rect 6812 7460 6825 7470
rect 6843 7460 6860 7473
rect 6812 7458 6860 7460
rect 6454 7454 6487 7458
rect 6450 7452 6487 7454
rect 6450 7451 6517 7452
rect 6450 7446 6481 7451
rect 6487 7446 6517 7451
rect 6450 7442 6517 7446
rect 6423 7439 6517 7442
rect 6423 7432 6472 7439
rect 6423 7426 6453 7432
rect 6472 7427 6477 7432
rect 6389 7410 6469 7426
rect 6481 7418 6517 7439
rect 6578 7434 6767 7458
rect 6812 7457 6859 7458
rect 6825 7452 6859 7457
rect 6593 7431 6767 7434
rect 6586 7428 6767 7431
rect 6795 7451 6859 7452
rect 6389 7408 6408 7410
rect 6423 7408 6457 7410
rect 6389 7392 6469 7408
rect 6389 7386 6408 7392
rect 6105 7360 6208 7370
rect 6059 7358 6208 7360
rect 6229 7358 6264 7370
rect 5898 7356 6060 7358
rect 5910 7336 5929 7356
rect 5944 7354 5974 7356
rect 5793 7328 5834 7336
rect 5916 7332 5929 7336
rect 5981 7340 6060 7356
rect 6092 7356 6264 7358
rect 6092 7340 6171 7356
rect 6178 7354 6208 7356
rect 5756 7318 5785 7328
rect 5799 7318 5828 7328
rect 5843 7318 5873 7332
rect 5916 7318 5959 7332
rect 5981 7328 6171 7340
rect 6236 7336 6242 7356
rect 5966 7318 5996 7328
rect 5997 7318 6155 7328
rect 6159 7318 6189 7328
rect 6193 7318 6223 7332
rect 6251 7318 6264 7356
rect 6336 7370 6365 7386
rect 6379 7370 6408 7386
rect 6423 7376 6453 7392
rect 6481 7370 6487 7418
rect 6490 7412 6509 7418
rect 6524 7412 6554 7420
rect 6490 7404 6554 7412
rect 6490 7388 6570 7404
rect 6586 7397 6648 7428
rect 6664 7397 6726 7428
rect 6795 7426 6844 7451
rect 6859 7426 6889 7442
rect 6758 7412 6788 7420
rect 6795 7418 6905 7426
rect 6758 7404 6803 7412
rect 6490 7386 6509 7388
rect 6524 7386 6570 7388
rect 6490 7370 6570 7386
rect 6597 7384 6632 7397
rect 6673 7394 6710 7397
rect 6673 7392 6715 7394
rect 6602 7381 6632 7384
rect 6611 7377 6618 7381
rect 6618 7376 6619 7377
rect 6577 7370 6587 7376
rect 6336 7362 6371 7370
rect 6336 7336 6337 7362
rect 6344 7336 6371 7362
rect 6279 7318 6309 7332
rect 6336 7328 6371 7336
rect 6373 7362 6414 7370
rect 6373 7336 6388 7362
rect 6395 7336 6414 7362
rect 6478 7358 6509 7370
rect 6524 7358 6627 7370
rect 6639 7360 6665 7386
rect 6680 7381 6710 7392
rect 6742 7388 6804 7404
rect 6742 7386 6788 7388
rect 6742 7370 6804 7386
rect 6816 7370 6822 7418
rect 6825 7410 6905 7418
rect 6825 7408 6844 7410
rect 6859 7408 6893 7410
rect 6825 7392 6905 7408
rect 6825 7370 6844 7392
rect 6859 7376 6889 7392
rect 6917 7386 6923 7460
rect 6926 7386 6945 7530
rect 6960 7386 6966 7530
rect 6975 7460 6988 7530
rect 7040 7526 7062 7530
rect 7033 7504 7062 7518
rect 7115 7504 7131 7518
rect 7169 7514 7175 7516
rect 7182 7514 7290 7530
rect 7297 7514 7303 7516
rect 7311 7514 7326 7530
rect 7392 7524 7411 7527
rect 7033 7502 7131 7504
rect 7158 7502 7326 7514
rect 7341 7504 7357 7518
rect 7392 7505 7414 7524
rect 7424 7518 7440 7519
rect 7423 7516 7440 7518
rect 7424 7511 7440 7516
rect 7414 7504 7420 7505
rect 7423 7504 7452 7511
rect 7341 7503 7452 7504
rect 7341 7502 7458 7503
rect 7017 7494 7068 7502
rect 7115 7494 7149 7502
rect 7017 7482 7042 7494
rect 7049 7482 7068 7494
rect 7122 7492 7149 7494
rect 7158 7492 7379 7502
rect 7414 7499 7420 7502
rect 7122 7488 7379 7492
rect 7017 7474 7068 7482
rect 7115 7474 7379 7488
rect 7423 7494 7458 7502
rect 6969 7426 6988 7460
rect 7033 7466 7062 7474
rect 7033 7460 7050 7466
rect 7033 7458 7067 7460
rect 7115 7458 7131 7474
rect 7132 7464 7340 7474
rect 7341 7464 7357 7474
rect 7405 7470 7420 7485
rect 7423 7482 7424 7494
rect 7431 7482 7458 7494
rect 7423 7474 7458 7482
rect 7423 7473 7452 7474
rect 7143 7460 7357 7464
rect 7158 7458 7357 7460
rect 7392 7460 7405 7470
rect 7423 7460 7440 7473
rect 7392 7458 7440 7460
rect 7034 7454 7067 7458
rect 7030 7452 7067 7454
rect 7030 7451 7097 7452
rect 7030 7446 7061 7451
rect 7067 7446 7097 7451
rect 7030 7442 7097 7446
rect 7003 7439 7097 7442
rect 7003 7432 7052 7439
rect 7003 7426 7033 7432
rect 7052 7427 7057 7432
rect 6969 7410 7049 7426
rect 7061 7418 7097 7439
rect 7158 7434 7347 7458
rect 7392 7457 7439 7458
rect 7405 7452 7439 7457
rect 7173 7431 7347 7434
rect 7166 7428 7347 7431
rect 7375 7451 7439 7452
rect 6969 7408 6988 7410
rect 7003 7408 7037 7410
rect 6969 7392 7049 7408
rect 6969 7386 6988 7392
rect 6685 7360 6788 7370
rect 6639 7358 6788 7360
rect 6809 7358 6844 7370
rect 6478 7356 6640 7358
rect 6490 7336 6509 7356
rect 6524 7354 6554 7356
rect 6373 7328 6414 7336
rect 6496 7332 6509 7336
rect 6561 7340 6640 7356
rect 6672 7356 6844 7358
rect 6672 7340 6751 7356
rect 6758 7354 6788 7356
rect 6336 7318 6365 7328
rect 6379 7318 6408 7328
rect 6423 7318 6453 7332
rect 6496 7318 6539 7332
rect 6561 7328 6751 7340
rect 6816 7336 6822 7356
rect 6546 7318 6576 7328
rect 6577 7318 6735 7328
rect 6739 7318 6769 7328
rect 6773 7318 6803 7332
rect 6831 7318 6844 7356
rect 6916 7370 6945 7386
rect 6959 7370 6988 7386
rect 7003 7376 7033 7392
rect 7061 7370 7067 7418
rect 7070 7412 7089 7418
rect 7104 7412 7134 7420
rect 7070 7404 7134 7412
rect 7070 7388 7150 7404
rect 7166 7397 7228 7428
rect 7244 7397 7306 7428
rect 7375 7426 7424 7451
rect 7439 7426 7469 7442
rect 7338 7412 7368 7420
rect 7375 7418 7485 7426
rect 7338 7404 7383 7412
rect 7070 7386 7089 7388
rect 7104 7386 7150 7388
rect 7070 7370 7150 7386
rect 7177 7384 7212 7397
rect 7253 7394 7290 7397
rect 7253 7392 7295 7394
rect 7182 7381 7212 7384
rect 7191 7377 7198 7381
rect 7198 7376 7199 7377
rect 7157 7370 7167 7376
rect 6916 7362 6951 7370
rect 6916 7336 6917 7362
rect 6924 7336 6951 7362
rect 6859 7318 6889 7332
rect 6916 7328 6951 7336
rect 6953 7362 6994 7370
rect 6953 7336 6968 7362
rect 6975 7336 6994 7362
rect 7058 7358 7089 7370
rect 7104 7358 7207 7370
rect 7219 7360 7245 7386
rect 7260 7381 7290 7392
rect 7322 7388 7384 7404
rect 7322 7386 7368 7388
rect 7322 7370 7384 7386
rect 7396 7370 7402 7418
rect 7405 7410 7485 7418
rect 7405 7408 7424 7410
rect 7439 7408 7473 7410
rect 7405 7392 7485 7408
rect 7405 7370 7424 7392
rect 7439 7376 7469 7392
rect 7497 7386 7503 7460
rect 7506 7386 7525 7530
rect 7540 7386 7546 7530
rect 7555 7460 7568 7530
rect 7620 7526 7642 7530
rect 7613 7504 7642 7518
rect 7695 7504 7711 7518
rect 7749 7514 7755 7516
rect 7762 7514 7870 7530
rect 7877 7514 7883 7516
rect 7891 7514 7906 7530
rect 7972 7524 7991 7527
rect 7613 7502 7711 7504
rect 7738 7502 7906 7514
rect 7921 7504 7937 7518
rect 7972 7505 7994 7524
rect 8004 7518 8020 7519
rect 8003 7516 8020 7518
rect 8004 7511 8020 7516
rect 7994 7504 8000 7505
rect 8003 7504 8032 7511
rect 7921 7503 8032 7504
rect 7921 7502 8038 7503
rect 7597 7494 7648 7502
rect 7695 7494 7729 7502
rect 7597 7482 7622 7494
rect 7629 7482 7648 7494
rect 7702 7492 7729 7494
rect 7738 7492 7959 7502
rect 7994 7499 8000 7502
rect 7702 7488 7959 7492
rect 7597 7474 7648 7482
rect 7695 7474 7959 7488
rect 8003 7494 8038 7502
rect 7549 7426 7568 7460
rect 7613 7466 7642 7474
rect 7613 7460 7630 7466
rect 7613 7458 7647 7460
rect 7695 7458 7711 7474
rect 7712 7464 7920 7474
rect 7921 7464 7937 7474
rect 7985 7470 8000 7485
rect 8003 7482 8004 7494
rect 8011 7482 8038 7494
rect 8003 7474 8038 7482
rect 8003 7473 8032 7474
rect 7723 7460 7937 7464
rect 7738 7458 7937 7460
rect 7972 7460 7985 7470
rect 8003 7460 8020 7473
rect 7972 7458 8020 7460
rect 7614 7454 7647 7458
rect 7610 7452 7647 7454
rect 7610 7451 7677 7452
rect 7610 7446 7641 7451
rect 7647 7446 7677 7451
rect 7610 7442 7677 7446
rect 7583 7439 7677 7442
rect 7583 7432 7632 7439
rect 7583 7426 7613 7432
rect 7632 7427 7637 7432
rect 7549 7410 7629 7426
rect 7641 7418 7677 7439
rect 7738 7434 7927 7458
rect 7972 7457 8019 7458
rect 7985 7452 8019 7457
rect 7753 7431 7927 7434
rect 7746 7428 7927 7431
rect 7955 7451 8019 7452
rect 7549 7408 7568 7410
rect 7583 7408 7617 7410
rect 7549 7392 7629 7408
rect 7549 7386 7568 7392
rect 7265 7360 7368 7370
rect 7219 7358 7368 7360
rect 7389 7358 7424 7370
rect 7058 7356 7220 7358
rect 7070 7336 7089 7356
rect 7104 7354 7134 7356
rect 6953 7328 6994 7336
rect 7076 7332 7089 7336
rect 7141 7340 7220 7356
rect 7252 7356 7424 7358
rect 7252 7340 7331 7356
rect 7338 7354 7368 7356
rect 6916 7318 6945 7328
rect 6959 7318 6988 7328
rect 7003 7318 7033 7332
rect 7076 7318 7119 7332
rect 7141 7328 7331 7340
rect 7396 7336 7402 7356
rect 7126 7318 7156 7328
rect 7157 7318 7315 7328
rect 7319 7318 7349 7328
rect 7353 7318 7383 7332
rect 7411 7318 7424 7356
rect 7496 7370 7525 7386
rect 7539 7370 7568 7386
rect 7583 7376 7613 7392
rect 7641 7370 7647 7418
rect 7650 7412 7669 7418
rect 7684 7412 7714 7420
rect 7650 7404 7714 7412
rect 7650 7388 7730 7404
rect 7746 7397 7808 7428
rect 7824 7397 7886 7428
rect 7955 7426 8004 7451
rect 8019 7426 8049 7442
rect 7918 7412 7948 7420
rect 7955 7418 8065 7426
rect 7918 7404 7963 7412
rect 7650 7386 7669 7388
rect 7684 7386 7730 7388
rect 7650 7370 7730 7386
rect 7757 7384 7792 7397
rect 7833 7394 7870 7397
rect 7833 7392 7875 7394
rect 7762 7381 7792 7384
rect 7771 7377 7778 7381
rect 7778 7376 7779 7377
rect 7737 7370 7747 7376
rect 7496 7362 7531 7370
rect 7496 7336 7497 7362
rect 7504 7336 7531 7362
rect 7439 7318 7469 7332
rect 7496 7328 7531 7336
rect 7533 7362 7574 7370
rect 7533 7336 7548 7362
rect 7555 7336 7574 7362
rect 7638 7358 7669 7370
rect 7684 7358 7787 7370
rect 7799 7360 7825 7386
rect 7840 7381 7870 7392
rect 7902 7388 7964 7404
rect 7902 7386 7948 7388
rect 7902 7370 7964 7386
rect 7976 7370 7982 7418
rect 7985 7410 8065 7418
rect 7985 7408 8004 7410
rect 8019 7408 8053 7410
rect 7985 7392 8065 7408
rect 7985 7370 8004 7392
rect 8019 7376 8049 7392
rect 8077 7386 8083 7460
rect 8086 7386 8105 7530
rect 8120 7386 8126 7530
rect 8135 7460 8148 7530
rect 8200 7526 8222 7530
rect 8193 7504 8222 7518
rect 8275 7504 8291 7518
rect 8329 7514 8335 7516
rect 8342 7514 8450 7530
rect 8457 7514 8463 7516
rect 8471 7514 8486 7530
rect 8552 7524 8571 7527
rect 8193 7502 8291 7504
rect 8318 7502 8486 7514
rect 8501 7504 8517 7518
rect 8552 7505 8574 7524
rect 8584 7518 8600 7519
rect 8583 7516 8600 7518
rect 8584 7511 8600 7516
rect 8574 7504 8580 7505
rect 8583 7504 8612 7511
rect 8501 7503 8612 7504
rect 8501 7502 8618 7503
rect 8177 7494 8228 7502
rect 8275 7494 8309 7502
rect 8177 7482 8202 7494
rect 8209 7482 8228 7494
rect 8282 7492 8309 7494
rect 8318 7492 8539 7502
rect 8574 7499 8580 7502
rect 8282 7488 8539 7492
rect 8177 7474 8228 7482
rect 8275 7474 8539 7488
rect 8583 7494 8618 7502
rect 8129 7426 8148 7460
rect 8193 7466 8222 7474
rect 8193 7460 8210 7466
rect 8193 7458 8227 7460
rect 8275 7458 8291 7474
rect 8292 7464 8500 7474
rect 8501 7464 8517 7474
rect 8565 7470 8580 7485
rect 8583 7482 8584 7494
rect 8591 7482 8618 7494
rect 8583 7474 8618 7482
rect 8583 7473 8612 7474
rect 8303 7460 8517 7464
rect 8318 7458 8517 7460
rect 8552 7460 8565 7470
rect 8583 7460 8600 7473
rect 8552 7458 8600 7460
rect 8194 7454 8227 7458
rect 8190 7452 8227 7454
rect 8190 7451 8257 7452
rect 8190 7446 8221 7451
rect 8227 7446 8257 7451
rect 8190 7442 8257 7446
rect 8163 7439 8257 7442
rect 8163 7432 8212 7439
rect 8163 7426 8193 7432
rect 8212 7427 8217 7432
rect 8129 7410 8209 7426
rect 8221 7418 8257 7439
rect 8318 7434 8507 7458
rect 8552 7457 8599 7458
rect 8565 7452 8599 7457
rect 8333 7431 8507 7434
rect 8326 7428 8507 7431
rect 8535 7451 8599 7452
rect 8129 7408 8148 7410
rect 8163 7408 8197 7410
rect 8129 7392 8209 7408
rect 8129 7386 8148 7392
rect 7845 7360 7948 7370
rect 7799 7358 7948 7360
rect 7969 7358 8004 7370
rect 7638 7356 7800 7358
rect 7650 7336 7669 7356
rect 7684 7354 7714 7356
rect 7533 7328 7574 7336
rect 7656 7332 7669 7336
rect 7721 7340 7800 7356
rect 7832 7356 8004 7358
rect 7832 7340 7911 7356
rect 7918 7354 7948 7356
rect 7496 7318 7525 7328
rect 7539 7318 7568 7328
rect 7583 7318 7613 7332
rect 7656 7318 7699 7332
rect 7721 7328 7911 7340
rect 7976 7336 7982 7356
rect 7706 7318 7736 7328
rect 7737 7318 7895 7328
rect 7899 7318 7929 7328
rect 7933 7318 7963 7332
rect 7991 7318 8004 7356
rect 8076 7370 8105 7386
rect 8119 7370 8148 7386
rect 8163 7376 8193 7392
rect 8221 7370 8227 7418
rect 8230 7412 8249 7418
rect 8264 7412 8294 7420
rect 8230 7404 8294 7412
rect 8230 7388 8310 7404
rect 8326 7397 8388 7428
rect 8404 7397 8466 7428
rect 8535 7426 8584 7451
rect 8599 7426 8629 7442
rect 8498 7412 8528 7420
rect 8535 7418 8645 7426
rect 8498 7404 8543 7412
rect 8230 7386 8249 7388
rect 8264 7386 8310 7388
rect 8230 7370 8310 7386
rect 8337 7384 8372 7397
rect 8413 7394 8450 7397
rect 8413 7392 8455 7394
rect 8342 7381 8372 7384
rect 8351 7377 8358 7381
rect 8358 7376 8359 7377
rect 8317 7370 8327 7376
rect 8076 7362 8111 7370
rect 8076 7336 8077 7362
rect 8084 7336 8111 7362
rect 8019 7318 8049 7332
rect 8076 7328 8111 7336
rect 8113 7362 8154 7370
rect 8113 7336 8128 7362
rect 8135 7336 8154 7362
rect 8218 7358 8249 7370
rect 8264 7358 8367 7370
rect 8379 7360 8405 7386
rect 8420 7381 8450 7392
rect 8482 7388 8544 7404
rect 8482 7386 8528 7388
rect 8482 7370 8544 7386
rect 8556 7370 8562 7418
rect 8565 7410 8645 7418
rect 8565 7408 8584 7410
rect 8599 7408 8633 7410
rect 8565 7392 8645 7408
rect 8565 7370 8584 7392
rect 8599 7376 8629 7392
rect 8657 7386 8663 7460
rect 8666 7386 8685 7530
rect 8700 7386 8706 7530
rect 8715 7460 8728 7530
rect 8780 7526 8802 7530
rect 8773 7504 8802 7518
rect 8855 7504 8871 7518
rect 8909 7514 8915 7516
rect 8922 7514 9030 7530
rect 9037 7514 9043 7516
rect 9051 7514 9066 7530
rect 9132 7524 9151 7527
rect 8773 7502 8871 7504
rect 8898 7502 9066 7514
rect 9081 7504 9097 7518
rect 9132 7505 9154 7524
rect 9164 7518 9180 7519
rect 9163 7516 9180 7518
rect 9164 7511 9180 7516
rect 9154 7504 9160 7505
rect 9163 7504 9192 7511
rect 9081 7503 9192 7504
rect 9081 7502 9198 7503
rect 8757 7494 8808 7502
rect 8855 7494 8889 7502
rect 8757 7482 8782 7494
rect 8789 7482 8808 7494
rect 8862 7492 8889 7494
rect 8898 7492 9119 7502
rect 9154 7499 9160 7502
rect 8862 7488 9119 7492
rect 8757 7474 8808 7482
rect 8855 7474 9119 7488
rect 9163 7494 9198 7502
rect 8709 7426 8728 7460
rect 8773 7466 8802 7474
rect 8773 7460 8790 7466
rect 8773 7458 8807 7460
rect 8855 7458 8871 7474
rect 8872 7464 9080 7474
rect 9081 7464 9097 7474
rect 9145 7470 9160 7485
rect 9163 7482 9164 7494
rect 9171 7482 9198 7494
rect 9163 7474 9198 7482
rect 9163 7473 9192 7474
rect 8883 7460 9097 7464
rect 8898 7458 9097 7460
rect 9132 7460 9145 7470
rect 9163 7460 9180 7473
rect 9132 7458 9180 7460
rect 8774 7454 8807 7458
rect 8770 7452 8807 7454
rect 8770 7451 8837 7452
rect 8770 7446 8801 7451
rect 8807 7446 8837 7451
rect 8770 7442 8837 7446
rect 8743 7439 8837 7442
rect 8743 7432 8792 7439
rect 8743 7426 8773 7432
rect 8792 7427 8797 7432
rect 8709 7410 8789 7426
rect 8801 7418 8837 7439
rect 8898 7434 9087 7458
rect 9132 7457 9179 7458
rect 9145 7452 9179 7457
rect 8913 7431 9087 7434
rect 8906 7428 9087 7431
rect 9115 7451 9179 7452
rect 8709 7408 8728 7410
rect 8743 7408 8777 7410
rect 8709 7392 8789 7408
rect 8709 7386 8728 7392
rect 8425 7360 8528 7370
rect 8379 7358 8528 7360
rect 8549 7358 8584 7370
rect 8218 7356 8380 7358
rect 8230 7336 8249 7356
rect 8264 7354 8294 7356
rect 8113 7328 8154 7336
rect 8236 7332 8249 7336
rect 8301 7340 8380 7356
rect 8412 7356 8584 7358
rect 8412 7340 8491 7356
rect 8498 7354 8528 7356
rect 8076 7318 8105 7328
rect 8119 7318 8148 7328
rect 8163 7318 8193 7332
rect 8236 7318 8279 7332
rect 8301 7328 8491 7340
rect 8556 7336 8562 7356
rect 8286 7318 8316 7328
rect 8317 7318 8475 7328
rect 8479 7318 8509 7328
rect 8513 7318 8543 7332
rect 8571 7318 8584 7356
rect 8656 7370 8685 7386
rect 8699 7370 8728 7386
rect 8743 7376 8773 7392
rect 8801 7370 8807 7418
rect 8810 7412 8829 7418
rect 8844 7412 8874 7420
rect 8810 7404 8874 7412
rect 8810 7388 8890 7404
rect 8906 7397 8968 7428
rect 8984 7397 9046 7428
rect 9115 7426 9164 7451
rect 9179 7426 9209 7442
rect 9078 7412 9108 7420
rect 9115 7418 9225 7426
rect 9078 7404 9123 7412
rect 8810 7386 8829 7388
rect 8844 7386 8890 7388
rect 8810 7370 8890 7386
rect 8917 7384 8952 7397
rect 8993 7394 9030 7397
rect 8993 7392 9035 7394
rect 8922 7381 8952 7384
rect 8931 7377 8938 7381
rect 8938 7376 8939 7377
rect 8897 7370 8907 7376
rect 8656 7362 8691 7370
rect 8656 7336 8657 7362
rect 8664 7336 8691 7362
rect 8599 7318 8629 7332
rect 8656 7328 8691 7336
rect 8693 7362 8734 7370
rect 8693 7336 8708 7362
rect 8715 7336 8734 7362
rect 8798 7358 8829 7370
rect 8844 7358 8947 7370
rect 8959 7360 8985 7386
rect 9000 7381 9030 7392
rect 9062 7388 9124 7404
rect 9062 7386 9108 7388
rect 9062 7370 9124 7386
rect 9136 7370 9142 7418
rect 9145 7410 9225 7418
rect 9145 7408 9164 7410
rect 9179 7408 9213 7410
rect 9145 7392 9225 7408
rect 9145 7370 9164 7392
rect 9179 7376 9209 7392
rect 9237 7386 9243 7460
rect 9246 7386 9265 7530
rect 9280 7386 9286 7530
rect 9295 7460 9308 7530
rect 9360 7526 9382 7530
rect 9353 7504 9382 7518
rect 9435 7504 9451 7518
rect 9489 7514 9495 7516
rect 9502 7514 9610 7530
rect 9617 7514 9623 7516
rect 9631 7514 9646 7530
rect 9712 7524 9731 7527
rect 9353 7502 9451 7504
rect 9478 7502 9646 7514
rect 9661 7504 9677 7518
rect 9712 7505 9734 7524
rect 9744 7518 9760 7519
rect 9743 7516 9760 7518
rect 9744 7511 9760 7516
rect 9734 7504 9740 7505
rect 9743 7504 9772 7511
rect 9661 7503 9772 7504
rect 9661 7502 9778 7503
rect 9337 7494 9388 7502
rect 9435 7494 9469 7502
rect 9337 7482 9362 7494
rect 9369 7482 9388 7494
rect 9442 7492 9469 7494
rect 9478 7492 9699 7502
rect 9734 7499 9740 7502
rect 9442 7488 9699 7492
rect 9337 7474 9388 7482
rect 9435 7474 9699 7488
rect 9743 7494 9778 7502
rect 9289 7426 9308 7460
rect 9353 7466 9382 7474
rect 9353 7460 9370 7466
rect 9353 7458 9387 7460
rect 9435 7458 9451 7474
rect 9452 7464 9660 7474
rect 9661 7464 9677 7474
rect 9725 7470 9740 7485
rect 9743 7482 9744 7494
rect 9751 7482 9778 7494
rect 9743 7474 9778 7482
rect 9743 7473 9772 7474
rect 9463 7460 9677 7464
rect 9478 7458 9677 7460
rect 9712 7460 9725 7470
rect 9743 7460 9760 7473
rect 9712 7458 9760 7460
rect 9354 7454 9387 7458
rect 9350 7452 9387 7454
rect 9350 7451 9417 7452
rect 9350 7446 9381 7451
rect 9387 7446 9417 7451
rect 9350 7442 9417 7446
rect 9323 7439 9417 7442
rect 9323 7432 9372 7439
rect 9323 7426 9353 7432
rect 9372 7427 9377 7432
rect 9289 7410 9369 7426
rect 9381 7418 9417 7439
rect 9478 7434 9667 7458
rect 9712 7457 9759 7458
rect 9725 7452 9759 7457
rect 9493 7431 9667 7434
rect 9486 7428 9667 7431
rect 9695 7451 9759 7452
rect 9289 7408 9308 7410
rect 9323 7408 9357 7410
rect 9289 7392 9369 7408
rect 9289 7386 9308 7392
rect 9005 7360 9108 7370
rect 8959 7358 9108 7360
rect 9129 7358 9164 7370
rect 8798 7356 8960 7358
rect 8810 7336 8829 7356
rect 8844 7354 8874 7356
rect 8693 7328 8734 7336
rect 8816 7332 8829 7336
rect 8881 7340 8960 7356
rect 8992 7356 9164 7358
rect 8992 7340 9071 7356
rect 9078 7354 9108 7356
rect 8656 7318 8685 7328
rect 8699 7318 8728 7328
rect 8743 7318 8773 7332
rect 8816 7318 8859 7332
rect 8881 7328 9071 7340
rect 9136 7336 9142 7356
rect 8866 7318 8896 7328
rect 8897 7318 9055 7328
rect 9059 7318 9089 7328
rect 9093 7318 9123 7332
rect 9151 7318 9164 7356
rect 9236 7370 9265 7386
rect 9279 7370 9308 7386
rect 9323 7376 9353 7392
rect 9381 7370 9387 7418
rect 9390 7412 9409 7418
rect 9424 7412 9454 7420
rect 9390 7404 9454 7412
rect 9390 7388 9470 7404
rect 9486 7397 9548 7428
rect 9564 7397 9626 7428
rect 9695 7426 9744 7451
rect 9759 7426 9789 7442
rect 9658 7412 9688 7420
rect 9695 7418 9805 7426
rect 9658 7404 9703 7412
rect 9390 7386 9409 7388
rect 9424 7386 9470 7388
rect 9390 7370 9470 7386
rect 9497 7384 9532 7397
rect 9573 7394 9610 7397
rect 9573 7392 9615 7394
rect 9502 7381 9532 7384
rect 9511 7377 9518 7381
rect 9518 7376 9519 7377
rect 9477 7370 9487 7376
rect 9236 7362 9271 7370
rect 9236 7336 9237 7362
rect 9244 7336 9271 7362
rect 9179 7318 9209 7332
rect 9236 7328 9271 7336
rect 9273 7362 9314 7370
rect 9273 7336 9288 7362
rect 9295 7336 9314 7362
rect 9378 7358 9409 7370
rect 9424 7358 9527 7370
rect 9539 7360 9565 7386
rect 9580 7381 9610 7392
rect 9642 7388 9704 7404
rect 9642 7386 9688 7388
rect 9642 7370 9704 7386
rect 9716 7370 9722 7418
rect 9725 7410 9805 7418
rect 9725 7408 9744 7410
rect 9759 7408 9793 7410
rect 9725 7392 9805 7408
rect 9725 7370 9744 7392
rect 9759 7376 9789 7392
rect 9817 7386 9823 7460
rect 9826 7386 9845 7530
rect 9860 7386 9866 7530
rect 9875 7460 9888 7530
rect 9940 7526 9962 7530
rect 9933 7504 9962 7518
rect 10015 7504 10031 7518
rect 10069 7514 10075 7516
rect 10082 7514 10190 7530
rect 10197 7514 10203 7516
rect 10211 7514 10226 7530
rect 10292 7524 10311 7527
rect 9933 7502 10031 7504
rect 10058 7502 10226 7514
rect 10241 7504 10257 7518
rect 10292 7505 10314 7524
rect 10324 7518 10340 7519
rect 10323 7516 10340 7518
rect 10324 7511 10340 7516
rect 10314 7504 10320 7505
rect 10323 7504 10352 7511
rect 10241 7503 10352 7504
rect 10241 7502 10358 7503
rect 9917 7494 9968 7502
rect 10015 7494 10049 7502
rect 9917 7482 9942 7494
rect 9949 7482 9968 7494
rect 10022 7492 10049 7494
rect 10058 7492 10279 7502
rect 10314 7499 10320 7502
rect 10022 7488 10279 7492
rect 9917 7474 9968 7482
rect 10015 7474 10279 7488
rect 10323 7494 10358 7502
rect 9869 7426 9888 7460
rect 9933 7466 9962 7474
rect 9933 7460 9950 7466
rect 9933 7458 9967 7460
rect 10015 7458 10031 7474
rect 10032 7464 10240 7474
rect 10241 7464 10257 7474
rect 10305 7470 10320 7485
rect 10323 7482 10324 7494
rect 10331 7482 10358 7494
rect 10323 7474 10358 7482
rect 10323 7473 10352 7474
rect 10043 7460 10257 7464
rect 10058 7458 10257 7460
rect 10292 7460 10305 7470
rect 10323 7460 10340 7473
rect 10292 7458 10340 7460
rect 9934 7454 9967 7458
rect 9930 7452 9967 7454
rect 9930 7451 9997 7452
rect 9930 7446 9961 7451
rect 9967 7446 9997 7451
rect 9930 7442 9997 7446
rect 9903 7439 9997 7442
rect 9903 7432 9952 7439
rect 9903 7426 9933 7432
rect 9952 7427 9957 7432
rect 9869 7410 9949 7426
rect 9961 7418 9997 7439
rect 10058 7434 10247 7458
rect 10292 7457 10339 7458
rect 10305 7452 10339 7457
rect 10073 7431 10247 7434
rect 10066 7428 10247 7431
rect 10275 7451 10339 7452
rect 9869 7408 9888 7410
rect 9903 7408 9937 7410
rect 9869 7392 9949 7408
rect 9869 7386 9888 7392
rect 9585 7360 9688 7370
rect 9539 7358 9688 7360
rect 9709 7358 9744 7370
rect 9378 7356 9540 7358
rect 9390 7336 9409 7356
rect 9424 7354 9454 7356
rect 9273 7328 9314 7336
rect 9396 7332 9409 7336
rect 9461 7340 9540 7356
rect 9572 7356 9744 7358
rect 9572 7340 9651 7356
rect 9658 7354 9688 7356
rect 9236 7318 9265 7328
rect 9279 7318 9308 7328
rect 9323 7318 9353 7332
rect 9396 7318 9439 7332
rect 9461 7328 9651 7340
rect 9716 7336 9722 7356
rect 9446 7318 9476 7328
rect 9477 7318 9635 7328
rect 9639 7318 9669 7328
rect 9673 7318 9703 7332
rect 9731 7318 9744 7356
rect 9816 7370 9845 7386
rect 9859 7370 9888 7386
rect 9903 7376 9933 7392
rect 9961 7370 9967 7418
rect 9970 7412 9989 7418
rect 10004 7412 10034 7420
rect 9970 7404 10034 7412
rect 9970 7388 10050 7404
rect 10066 7397 10128 7428
rect 10144 7397 10206 7428
rect 10275 7426 10324 7451
rect 10339 7426 10369 7442
rect 10238 7412 10268 7420
rect 10275 7418 10385 7426
rect 10238 7404 10283 7412
rect 9970 7386 9989 7388
rect 10004 7386 10050 7388
rect 9970 7370 10050 7386
rect 10077 7384 10112 7397
rect 10153 7394 10190 7397
rect 10153 7392 10195 7394
rect 10082 7381 10112 7384
rect 10091 7377 10098 7381
rect 10098 7376 10099 7377
rect 10057 7370 10067 7376
rect 9816 7362 9851 7370
rect 9816 7336 9817 7362
rect 9824 7336 9851 7362
rect 9759 7318 9789 7332
rect 9816 7328 9851 7336
rect 9853 7362 9894 7370
rect 9853 7336 9868 7362
rect 9875 7336 9894 7362
rect 9958 7358 9989 7370
rect 10004 7358 10107 7370
rect 10119 7360 10145 7386
rect 10160 7381 10190 7392
rect 10222 7388 10284 7404
rect 10222 7386 10268 7388
rect 10222 7370 10284 7386
rect 10296 7370 10302 7418
rect 10305 7410 10385 7418
rect 10305 7408 10324 7410
rect 10339 7408 10373 7410
rect 10305 7392 10385 7408
rect 10305 7370 10324 7392
rect 10339 7376 10369 7392
rect 10397 7386 10403 7460
rect 10406 7386 10425 7530
rect 10440 7386 10446 7530
rect 10455 7460 10468 7530
rect 10520 7526 10542 7530
rect 10513 7504 10542 7518
rect 10595 7504 10611 7518
rect 10649 7514 10655 7516
rect 10662 7514 10770 7530
rect 10777 7514 10783 7516
rect 10791 7514 10806 7530
rect 10872 7524 10891 7527
rect 10513 7502 10611 7504
rect 10638 7502 10806 7514
rect 10821 7504 10837 7518
rect 10872 7505 10894 7524
rect 10904 7518 10920 7519
rect 10903 7516 10920 7518
rect 10904 7511 10920 7516
rect 10894 7504 10900 7505
rect 10903 7504 10932 7511
rect 10821 7503 10932 7504
rect 10821 7502 10938 7503
rect 10497 7494 10548 7502
rect 10595 7494 10629 7502
rect 10497 7482 10522 7494
rect 10529 7482 10548 7494
rect 10602 7492 10629 7494
rect 10638 7492 10859 7502
rect 10894 7499 10900 7502
rect 10602 7488 10859 7492
rect 10497 7474 10548 7482
rect 10595 7474 10859 7488
rect 10903 7494 10938 7502
rect 10449 7426 10468 7460
rect 10513 7466 10542 7474
rect 10513 7460 10530 7466
rect 10513 7458 10547 7460
rect 10595 7458 10611 7474
rect 10612 7464 10820 7474
rect 10821 7464 10837 7474
rect 10885 7470 10900 7485
rect 10903 7482 10904 7494
rect 10911 7482 10938 7494
rect 10903 7474 10938 7482
rect 10903 7473 10932 7474
rect 10623 7460 10837 7464
rect 10638 7458 10837 7460
rect 10872 7460 10885 7470
rect 10903 7460 10920 7473
rect 10872 7458 10920 7460
rect 10514 7454 10547 7458
rect 10510 7452 10547 7454
rect 10510 7451 10577 7452
rect 10510 7446 10541 7451
rect 10547 7446 10577 7451
rect 10510 7442 10577 7446
rect 10483 7439 10577 7442
rect 10483 7432 10532 7439
rect 10483 7426 10513 7432
rect 10532 7427 10537 7432
rect 10449 7410 10529 7426
rect 10541 7418 10577 7439
rect 10638 7434 10827 7458
rect 10872 7457 10919 7458
rect 10885 7452 10919 7457
rect 10653 7431 10827 7434
rect 10646 7428 10827 7431
rect 10855 7451 10919 7452
rect 10449 7408 10468 7410
rect 10483 7408 10517 7410
rect 10449 7392 10529 7408
rect 10449 7386 10468 7392
rect 10165 7360 10268 7370
rect 10119 7358 10268 7360
rect 10289 7358 10324 7370
rect 9958 7356 10120 7358
rect 9970 7336 9989 7356
rect 10004 7354 10034 7356
rect 9853 7328 9894 7336
rect 9976 7332 9989 7336
rect 10041 7340 10120 7356
rect 10152 7356 10324 7358
rect 10152 7340 10231 7356
rect 10238 7354 10268 7356
rect 9816 7318 9845 7328
rect 9859 7318 9888 7328
rect 9903 7318 9933 7332
rect 9976 7318 10019 7332
rect 10041 7328 10231 7340
rect 10296 7336 10302 7356
rect 10026 7318 10056 7328
rect 10057 7318 10215 7328
rect 10219 7318 10249 7328
rect 10253 7318 10283 7332
rect 10311 7318 10324 7356
rect 10396 7370 10425 7386
rect 10439 7370 10468 7386
rect 10483 7376 10513 7392
rect 10541 7370 10547 7418
rect 10550 7412 10569 7418
rect 10584 7412 10614 7420
rect 10550 7404 10614 7412
rect 10550 7388 10630 7404
rect 10646 7397 10708 7428
rect 10724 7397 10786 7428
rect 10855 7426 10904 7451
rect 10919 7426 10949 7442
rect 10818 7412 10848 7420
rect 10855 7418 10965 7426
rect 10818 7404 10863 7412
rect 10550 7386 10569 7388
rect 10584 7386 10630 7388
rect 10550 7370 10630 7386
rect 10657 7384 10692 7397
rect 10733 7394 10770 7397
rect 10733 7392 10775 7394
rect 10662 7381 10692 7384
rect 10671 7377 10678 7381
rect 10678 7376 10679 7377
rect 10637 7370 10647 7376
rect 10396 7362 10431 7370
rect 10396 7336 10397 7362
rect 10404 7336 10431 7362
rect 10339 7318 10369 7332
rect 10396 7328 10431 7336
rect 10433 7362 10474 7370
rect 10433 7336 10448 7362
rect 10455 7336 10474 7362
rect 10538 7358 10569 7370
rect 10584 7358 10687 7370
rect 10699 7360 10725 7386
rect 10740 7381 10770 7392
rect 10802 7388 10864 7404
rect 10802 7386 10848 7388
rect 10802 7370 10864 7386
rect 10876 7370 10882 7418
rect 10885 7410 10965 7418
rect 10885 7408 10904 7410
rect 10919 7408 10953 7410
rect 10885 7392 10965 7408
rect 10885 7370 10904 7392
rect 10919 7376 10949 7392
rect 10977 7386 10983 7460
rect 10986 7386 11005 7530
rect 11020 7386 11026 7530
rect 11035 7460 11048 7530
rect 11100 7526 11122 7530
rect 11093 7504 11122 7518
rect 11175 7504 11191 7518
rect 11229 7514 11235 7516
rect 11242 7514 11350 7530
rect 11357 7514 11363 7516
rect 11371 7514 11386 7530
rect 11452 7524 11471 7527
rect 11093 7502 11191 7504
rect 11218 7502 11386 7514
rect 11401 7504 11417 7518
rect 11452 7505 11474 7524
rect 11484 7518 11500 7519
rect 11483 7516 11500 7518
rect 11484 7511 11500 7516
rect 11474 7504 11480 7505
rect 11483 7504 11512 7511
rect 11401 7503 11512 7504
rect 11401 7502 11518 7503
rect 11077 7494 11128 7502
rect 11175 7494 11209 7502
rect 11077 7482 11102 7494
rect 11109 7482 11128 7494
rect 11182 7492 11209 7494
rect 11218 7492 11439 7502
rect 11474 7499 11480 7502
rect 11182 7488 11439 7492
rect 11077 7474 11128 7482
rect 11175 7474 11439 7488
rect 11483 7494 11518 7502
rect 11029 7426 11048 7460
rect 11093 7466 11122 7474
rect 11093 7460 11110 7466
rect 11093 7458 11127 7460
rect 11175 7458 11191 7474
rect 11192 7464 11400 7474
rect 11401 7464 11417 7474
rect 11465 7470 11480 7485
rect 11483 7482 11484 7494
rect 11491 7482 11518 7494
rect 11483 7474 11518 7482
rect 11483 7473 11512 7474
rect 11203 7460 11417 7464
rect 11218 7458 11417 7460
rect 11452 7460 11465 7470
rect 11483 7460 11500 7473
rect 11452 7458 11500 7460
rect 11094 7454 11127 7458
rect 11090 7452 11127 7454
rect 11090 7451 11157 7452
rect 11090 7446 11121 7451
rect 11127 7446 11157 7451
rect 11090 7442 11157 7446
rect 11063 7439 11157 7442
rect 11063 7432 11112 7439
rect 11063 7426 11093 7432
rect 11112 7427 11117 7432
rect 11029 7410 11109 7426
rect 11121 7418 11157 7439
rect 11218 7434 11407 7458
rect 11452 7457 11499 7458
rect 11465 7452 11499 7457
rect 11233 7431 11407 7434
rect 11226 7428 11407 7431
rect 11435 7451 11499 7452
rect 11029 7408 11048 7410
rect 11063 7408 11097 7410
rect 11029 7392 11109 7408
rect 11029 7386 11048 7392
rect 10745 7360 10848 7370
rect 10699 7358 10848 7360
rect 10869 7358 10904 7370
rect 10538 7356 10700 7358
rect 10550 7336 10569 7356
rect 10584 7354 10614 7356
rect 10433 7328 10474 7336
rect 10556 7332 10569 7336
rect 10621 7340 10700 7356
rect 10732 7356 10904 7358
rect 10732 7340 10811 7356
rect 10818 7354 10848 7356
rect 10396 7318 10425 7328
rect 10439 7318 10468 7328
rect 10483 7318 10513 7332
rect 10556 7318 10599 7332
rect 10621 7328 10811 7340
rect 10876 7336 10882 7356
rect 10606 7318 10636 7328
rect 10637 7318 10795 7328
rect 10799 7318 10829 7328
rect 10833 7318 10863 7332
rect 10891 7318 10904 7356
rect 10976 7370 11005 7386
rect 11019 7370 11048 7386
rect 11063 7376 11093 7392
rect 11121 7370 11127 7418
rect 11130 7412 11149 7418
rect 11164 7412 11194 7420
rect 11130 7404 11194 7412
rect 11130 7388 11210 7404
rect 11226 7397 11288 7428
rect 11304 7397 11366 7428
rect 11435 7426 11484 7451
rect 11499 7426 11529 7442
rect 11398 7412 11428 7420
rect 11435 7418 11545 7426
rect 11398 7404 11443 7412
rect 11130 7386 11149 7388
rect 11164 7386 11210 7388
rect 11130 7370 11210 7386
rect 11237 7384 11272 7397
rect 11313 7394 11350 7397
rect 11313 7392 11355 7394
rect 11242 7381 11272 7384
rect 11251 7377 11258 7381
rect 11258 7376 11259 7377
rect 11217 7370 11227 7376
rect 10976 7362 11011 7370
rect 10976 7336 10977 7362
rect 10984 7336 11011 7362
rect 10919 7318 10949 7332
rect 10976 7328 11011 7336
rect 11013 7362 11054 7370
rect 11013 7336 11028 7362
rect 11035 7336 11054 7362
rect 11118 7358 11149 7370
rect 11164 7358 11267 7370
rect 11279 7360 11305 7386
rect 11320 7381 11350 7392
rect 11382 7388 11444 7404
rect 11382 7386 11428 7388
rect 11382 7370 11444 7386
rect 11456 7370 11462 7418
rect 11465 7410 11545 7418
rect 11465 7408 11484 7410
rect 11499 7408 11533 7410
rect 11465 7392 11545 7408
rect 11465 7370 11484 7392
rect 11499 7376 11529 7392
rect 11557 7386 11563 7460
rect 11566 7386 11585 7530
rect 11600 7386 11606 7530
rect 11615 7460 11628 7530
rect 11680 7526 11702 7530
rect 11673 7504 11702 7518
rect 11755 7504 11771 7518
rect 11809 7514 11815 7516
rect 11822 7514 11930 7530
rect 11937 7514 11943 7516
rect 11951 7514 11966 7530
rect 12032 7524 12051 7527
rect 11673 7502 11771 7504
rect 11798 7502 11966 7514
rect 11981 7504 11997 7518
rect 12032 7505 12054 7524
rect 12064 7518 12080 7519
rect 12063 7516 12080 7518
rect 12064 7511 12080 7516
rect 12054 7504 12060 7505
rect 12063 7504 12092 7511
rect 11981 7503 12092 7504
rect 11981 7502 12098 7503
rect 11657 7494 11708 7502
rect 11755 7494 11789 7502
rect 11657 7482 11682 7494
rect 11689 7482 11708 7494
rect 11762 7492 11789 7494
rect 11798 7492 12019 7502
rect 12054 7499 12060 7502
rect 11762 7488 12019 7492
rect 11657 7474 11708 7482
rect 11755 7474 12019 7488
rect 12063 7494 12098 7502
rect 11609 7426 11628 7460
rect 11673 7466 11702 7474
rect 11673 7460 11690 7466
rect 11673 7458 11707 7460
rect 11755 7458 11771 7474
rect 11772 7464 11980 7474
rect 11981 7464 11997 7474
rect 12045 7470 12060 7485
rect 12063 7482 12064 7494
rect 12071 7482 12098 7494
rect 12063 7474 12098 7482
rect 12063 7473 12092 7474
rect 11783 7460 11997 7464
rect 11798 7458 11997 7460
rect 12032 7460 12045 7470
rect 12063 7460 12080 7473
rect 12032 7458 12080 7460
rect 11674 7454 11707 7458
rect 11670 7452 11707 7454
rect 11670 7451 11737 7452
rect 11670 7446 11701 7451
rect 11707 7446 11737 7451
rect 11670 7442 11737 7446
rect 11643 7439 11737 7442
rect 11643 7432 11692 7439
rect 11643 7426 11673 7432
rect 11692 7427 11697 7432
rect 11609 7410 11689 7426
rect 11701 7418 11737 7439
rect 11798 7434 11987 7458
rect 12032 7457 12079 7458
rect 12045 7452 12079 7457
rect 11813 7431 11987 7434
rect 11806 7428 11987 7431
rect 12015 7451 12079 7452
rect 11609 7408 11628 7410
rect 11643 7408 11677 7410
rect 11609 7392 11689 7408
rect 11609 7386 11628 7392
rect 11325 7360 11428 7370
rect 11279 7358 11428 7360
rect 11449 7358 11484 7370
rect 11118 7356 11280 7358
rect 11130 7336 11149 7356
rect 11164 7354 11194 7356
rect 11013 7328 11054 7336
rect 11136 7332 11149 7336
rect 11201 7340 11280 7356
rect 11312 7356 11484 7358
rect 11312 7340 11391 7356
rect 11398 7354 11428 7356
rect 10976 7318 11005 7328
rect 11019 7318 11048 7328
rect 11063 7318 11093 7332
rect 11136 7318 11179 7332
rect 11201 7328 11391 7340
rect 11456 7336 11462 7356
rect 11186 7318 11216 7328
rect 11217 7318 11375 7328
rect 11379 7318 11409 7328
rect 11413 7318 11443 7332
rect 11471 7318 11484 7356
rect 11556 7370 11585 7386
rect 11599 7370 11628 7386
rect 11643 7376 11673 7392
rect 11701 7370 11707 7418
rect 11710 7412 11729 7418
rect 11744 7412 11774 7420
rect 11710 7404 11774 7412
rect 11710 7388 11790 7404
rect 11806 7397 11868 7428
rect 11884 7397 11946 7428
rect 12015 7426 12064 7451
rect 12079 7426 12109 7442
rect 11978 7412 12008 7420
rect 12015 7418 12125 7426
rect 11978 7404 12023 7412
rect 11710 7386 11729 7388
rect 11744 7386 11790 7388
rect 11710 7370 11790 7386
rect 11817 7384 11852 7397
rect 11893 7394 11930 7397
rect 11893 7392 11935 7394
rect 11822 7381 11852 7384
rect 11831 7377 11838 7381
rect 11838 7376 11839 7377
rect 11797 7370 11807 7376
rect 11556 7362 11591 7370
rect 11556 7336 11557 7362
rect 11564 7336 11591 7362
rect 11499 7318 11529 7332
rect 11556 7328 11591 7336
rect 11593 7362 11634 7370
rect 11593 7336 11608 7362
rect 11615 7336 11634 7362
rect 11698 7358 11729 7370
rect 11744 7358 11847 7370
rect 11859 7360 11885 7386
rect 11900 7381 11930 7392
rect 11962 7388 12024 7404
rect 11962 7386 12008 7388
rect 11962 7370 12024 7386
rect 12036 7370 12042 7418
rect 12045 7410 12125 7418
rect 12045 7408 12064 7410
rect 12079 7408 12113 7410
rect 12045 7392 12125 7408
rect 12045 7370 12064 7392
rect 12079 7376 12109 7392
rect 12137 7386 12143 7460
rect 12146 7386 12165 7530
rect 12180 7386 12186 7530
rect 12195 7460 12208 7530
rect 12260 7526 12282 7530
rect 12253 7504 12282 7518
rect 12335 7504 12351 7518
rect 12389 7514 12395 7516
rect 12402 7514 12510 7530
rect 12517 7514 12523 7516
rect 12531 7514 12546 7530
rect 12612 7524 12631 7527
rect 12253 7502 12351 7504
rect 12378 7502 12546 7514
rect 12561 7504 12577 7518
rect 12612 7505 12634 7524
rect 12644 7518 12660 7519
rect 12643 7516 12660 7518
rect 12644 7511 12660 7516
rect 12634 7504 12640 7505
rect 12643 7504 12672 7511
rect 12561 7503 12672 7504
rect 12561 7502 12678 7503
rect 12237 7494 12288 7502
rect 12335 7494 12369 7502
rect 12237 7482 12262 7494
rect 12269 7482 12288 7494
rect 12342 7492 12369 7494
rect 12378 7492 12599 7502
rect 12634 7499 12640 7502
rect 12342 7488 12599 7492
rect 12237 7474 12288 7482
rect 12335 7474 12599 7488
rect 12643 7494 12678 7502
rect 12189 7426 12208 7460
rect 12253 7466 12282 7474
rect 12253 7460 12270 7466
rect 12253 7458 12287 7460
rect 12335 7458 12351 7474
rect 12352 7464 12560 7474
rect 12561 7464 12577 7474
rect 12625 7470 12640 7485
rect 12643 7482 12644 7494
rect 12651 7482 12678 7494
rect 12643 7474 12678 7482
rect 12643 7473 12672 7474
rect 12363 7460 12577 7464
rect 12378 7458 12577 7460
rect 12612 7460 12625 7470
rect 12643 7460 12660 7473
rect 12612 7458 12660 7460
rect 12254 7454 12287 7458
rect 12250 7452 12287 7454
rect 12250 7451 12317 7452
rect 12250 7446 12281 7451
rect 12287 7446 12317 7451
rect 12250 7442 12317 7446
rect 12223 7439 12317 7442
rect 12223 7432 12272 7439
rect 12223 7426 12253 7432
rect 12272 7427 12277 7432
rect 12189 7410 12269 7426
rect 12281 7418 12317 7439
rect 12378 7434 12567 7458
rect 12612 7457 12659 7458
rect 12625 7452 12659 7457
rect 12393 7431 12567 7434
rect 12386 7428 12567 7431
rect 12595 7451 12659 7452
rect 12189 7408 12208 7410
rect 12223 7408 12257 7410
rect 12189 7392 12269 7408
rect 12189 7386 12208 7392
rect 11905 7360 12008 7370
rect 11859 7358 12008 7360
rect 12029 7358 12064 7370
rect 11698 7356 11860 7358
rect 11710 7336 11729 7356
rect 11744 7354 11774 7356
rect 11593 7328 11634 7336
rect 11716 7332 11729 7336
rect 11781 7340 11860 7356
rect 11892 7356 12064 7358
rect 11892 7340 11971 7356
rect 11978 7354 12008 7356
rect 11556 7318 11585 7328
rect 11599 7318 11628 7328
rect 11643 7318 11673 7332
rect 11716 7318 11759 7332
rect 11781 7328 11971 7340
rect 12036 7336 12042 7356
rect 11766 7318 11796 7328
rect 11797 7318 11955 7328
rect 11959 7318 11989 7328
rect 11993 7318 12023 7332
rect 12051 7318 12064 7356
rect 12136 7370 12165 7386
rect 12179 7370 12208 7386
rect 12223 7376 12253 7392
rect 12281 7370 12287 7418
rect 12290 7412 12309 7418
rect 12324 7412 12354 7420
rect 12290 7404 12354 7412
rect 12290 7388 12370 7404
rect 12386 7397 12448 7428
rect 12464 7397 12526 7428
rect 12595 7426 12644 7451
rect 12659 7426 12689 7442
rect 12558 7412 12588 7420
rect 12595 7418 12705 7426
rect 12558 7404 12603 7412
rect 12290 7386 12309 7388
rect 12324 7386 12370 7388
rect 12290 7370 12370 7386
rect 12397 7384 12432 7397
rect 12473 7394 12510 7397
rect 12473 7392 12515 7394
rect 12402 7381 12432 7384
rect 12411 7377 12418 7381
rect 12418 7376 12419 7377
rect 12377 7370 12387 7376
rect 12136 7362 12171 7370
rect 12136 7336 12137 7362
rect 12144 7336 12171 7362
rect 12079 7318 12109 7332
rect 12136 7328 12171 7336
rect 12173 7362 12214 7370
rect 12173 7336 12188 7362
rect 12195 7336 12214 7362
rect 12278 7358 12309 7370
rect 12324 7358 12427 7370
rect 12439 7360 12465 7386
rect 12480 7381 12510 7392
rect 12542 7388 12604 7404
rect 12542 7386 12588 7388
rect 12542 7370 12604 7386
rect 12616 7370 12622 7418
rect 12625 7410 12705 7418
rect 12625 7408 12644 7410
rect 12659 7408 12693 7410
rect 12625 7392 12705 7408
rect 12625 7370 12644 7392
rect 12659 7376 12689 7392
rect 12717 7386 12723 7460
rect 12726 7386 12745 7530
rect 12760 7386 12766 7530
rect 12775 7460 12788 7530
rect 12840 7526 12862 7530
rect 12833 7504 12862 7518
rect 12915 7504 12931 7518
rect 12969 7514 12975 7516
rect 12982 7514 13090 7530
rect 13097 7514 13103 7516
rect 13111 7514 13126 7530
rect 13192 7524 13211 7527
rect 12833 7502 12931 7504
rect 12958 7502 13126 7514
rect 13141 7504 13157 7518
rect 13192 7505 13214 7524
rect 13224 7518 13240 7519
rect 13223 7516 13240 7518
rect 13224 7511 13240 7516
rect 13214 7504 13220 7505
rect 13223 7504 13252 7511
rect 13141 7503 13252 7504
rect 13141 7502 13258 7503
rect 12817 7494 12868 7502
rect 12915 7494 12949 7502
rect 12817 7482 12842 7494
rect 12849 7482 12868 7494
rect 12922 7492 12949 7494
rect 12958 7492 13179 7502
rect 13214 7499 13220 7502
rect 12922 7488 13179 7492
rect 12817 7474 12868 7482
rect 12915 7474 13179 7488
rect 13223 7494 13258 7502
rect 12769 7426 12788 7460
rect 12833 7466 12862 7474
rect 12833 7460 12850 7466
rect 12833 7458 12867 7460
rect 12915 7458 12931 7474
rect 12932 7464 13140 7474
rect 13141 7464 13157 7474
rect 13205 7470 13220 7485
rect 13223 7482 13224 7494
rect 13231 7482 13258 7494
rect 13223 7474 13258 7482
rect 13223 7473 13252 7474
rect 12943 7460 13157 7464
rect 12958 7458 13157 7460
rect 13192 7460 13205 7470
rect 13223 7460 13240 7473
rect 13192 7458 13240 7460
rect 12834 7454 12867 7458
rect 12830 7452 12867 7454
rect 12830 7451 12897 7452
rect 12830 7446 12861 7451
rect 12867 7446 12897 7451
rect 12830 7442 12897 7446
rect 12803 7439 12897 7442
rect 12803 7432 12852 7439
rect 12803 7426 12833 7432
rect 12852 7427 12857 7432
rect 12769 7410 12849 7426
rect 12861 7418 12897 7439
rect 12958 7434 13147 7458
rect 13192 7457 13239 7458
rect 13205 7452 13239 7457
rect 12973 7431 13147 7434
rect 12966 7428 13147 7431
rect 13175 7451 13239 7452
rect 12769 7408 12788 7410
rect 12803 7408 12837 7410
rect 12769 7392 12849 7408
rect 12769 7386 12788 7392
rect 12485 7360 12588 7370
rect 12439 7358 12588 7360
rect 12609 7358 12644 7370
rect 12278 7356 12440 7358
rect 12290 7336 12309 7356
rect 12324 7354 12354 7356
rect 12173 7328 12214 7336
rect 12296 7332 12309 7336
rect 12361 7340 12440 7356
rect 12472 7356 12644 7358
rect 12472 7340 12551 7356
rect 12558 7354 12588 7356
rect 12136 7318 12165 7328
rect 12179 7318 12208 7328
rect 12223 7318 12253 7332
rect 12296 7318 12339 7332
rect 12361 7328 12551 7340
rect 12616 7336 12622 7356
rect 12346 7318 12376 7328
rect 12377 7318 12535 7328
rect 12539 7318 12569 7328
rect 12573 7318 12603 7332
rect 12631 7318 12644 7356
rect 12716 7370 12745 7386
rect 12759 7370 12788 7386
rect 12803 7376 12833 7392
rect 12861 7370 12867 7418
rect 12870 7412 12889 7418
rect 12904 7412 12934 7420
rect 12870 7404 12934 7412
rect 12870 7388 12950 7404
rect 12966 7397 13028 7428
rect 13044 7397 13106 7428
rect 13175 7426 13224 7451
rect 13239 7426 13269 7442
rect 13138 7412 13168 7420
rect 13175 7418 13285 7426
rect 13138 7404 13183 7412
rect 12870 7386 12889 7388
rect 12904 7386 12950 7388
rect 12870 7370 12950 7386
rect 12977 7384 13012 7397
rect 13053 7394 13090 7397
rect 13053 7392 13095 7394
rect 12982 7381 13012 7384
rect 12991 7377 12998 7381
rect 12998 7376 12999 7377
rect 12957 7370 12967 7376
rect 12716 7362 12751 7370
rect 12716 7336 12717 7362
rect 12724 7336 12751 7362
rect 12659 7318 12689 7332
rect 12716 7328 12751 7336
rect 12753 7362 12794 7370
rect 12753 7336 12768 7362
rect 12775 7336 12794 7362
rect 12858 7358 12889 7370
rect 12904 7358 13007 7370
rect 13019 7360 13045 7386
rect 13060 7381 13090 7392
rect 13122 7388 13184 7404
rect 13122 7386 13168 7388
rect 13122 7370 13184 7386
rect 13196 7370 13202 7418
rect 13205 7410 13285 7418
rect 13205 7408 13224 7410
rect 13239 7408 13273 7410
rect 13205 7392 13285 7408
rect 13205 7370 13224 7392
rect 13239 7376 13269 7392
rect 13297 7386 13303 7460
rect 13306 7386 13325 7530
rect 13340 7386 13346 7530
rect 13355 7460 13368 7530
rect 13420 7526 13442 7530
rect 13413 7504 13442 7518
rect 13495 7504 13511 7518
rect 13549 7514 13555 7516
rect 13562 7514 13670 7530
rect 13677 7514 13683 7516
rect 13691 7514 13706 7530
rect 13772 7524 13791 7527
rect 13413 7502 13511 7504
rect 13538 7502 13706 7514
rect 13721 7504 13737 7518
rect 13772 7505 13794 7524
rect 13804 7518 13820 7519
rect 13803 7516 13820 7518
rect 13804 7511 13820 7516
rect 13794 7504 13800 7505
rect 13803 7504 13832 7511
rect 13721 7503 13832 7504
rect 13721 7502 13838 7503
rect 13397 7494 13448 7502
rect 13495 7494 13529 7502
rect 13397 7482 13422 7494
rect 13429 7482 13448 7494
rect 13502 7492 13529 7494
rect 13538 7492 13759 7502
rect 13794 7499 13800 7502
rect 13502 7488 13759 7492
rect 13397 7474 13448 7482
rect 13495 7474 13759 7488
rect 13803 7494 13838 7502
rect 13349 7426 13368 7460
rect 13413 7466 13442 7474
rect 13413 7460 13430 7466
rect 13413 7458 13447 7460
rect 13495 7458 13511 7474
rect 13512 7464 13720 7474
rect 13721 7464 13737 7474
rect 13785 7470 13800 7485
rect 13803 7482 13804 7494
rect 13811 7482 13838 7494
rect 13803 7474 13838 7482
rect 13803 7473 13832 7474
rect 13523 7460 13737 7464
rect 13538 7458 13737 7460
rect 13772 7460 13785 7470
rect 13803 7460 13820 7473
rect 13772 7458 13820 7460
rect 13414 7454 13447 7458
rect 13410 7452 13447 7454
rect 13410 7451 13477 7452
rect 13410 7446 13441 7451
rect 13447 7446 13477 7451
rect 13410 7442 13477 7446
rect 13383 7439 13477 7442
rect 13383 7432 13432 7439
rect 13383 7426 13413 7432
rect 13432 7427 13437 7432
rect 13349 7410 13429 7426
rect 13441 7418 13477 7439
rect 13538 7434 13727 7458
rect 13772 7457 13819 7458
rect 13785 7452 13819 7457
rect 13553 7431 13727 7434
rect 13546 7428 13727 7431
rect 13755 7451 13819 7452
rect 13349 7408 13368 7410
rect 13383 7408 13417 7410
rect 13349 7392 13429 7408
rect 13349 7386 13368 7392
rect 13065 7360 13168 7370
rect 13019 7358 13168 7360
rect 13189 7358 13224 7370
rect 12858 7356 13020 7358
rect 12870 7336 12889 7356
rect 12904 7354 12934 7356
rect 12753 7328 12794 7336
rect 12876 7332 12889 7336
rect 12941 7340 13020 7356
rect 13052 7356 13224 7358
rect 13052 7340 13131 7356
rect 13138 7354 13168 7356
rect 12716 7318 12745 7328
rect 12759 7318 12788 7328
rect 12803 7318 12833 7332
rect 12876 7318 12919 7332
rect 12941 7328 13131 7340
rect 13196 7336 13202 7356
rect 12926 7318 12956 7328
rect 12957 7318 13115 7328
rect 13119 7318 13149 7328
rect 13153 7318 13183 7332
rect 13211 7318 13224 7356
rect 13296 7370 13325 7386
rect 13339 7370 13368 7386
rect 13383 7376 13413 7392
rect 13441 7370 13447 7418
rect 13450 7412 13469 7418
rect 13484 7412 13514 7420
rect 13450 7404 13514 7412
rect 13450 7388 13530 7404
rect 13546 7397 13608 7428
rect 13624 7397 13686 7428
rect 13755 7426 13804 7451
rect 13819 7426 13849 7442
rect 13718 7412 13748 7420
rect 13755 7418 13865 7426
rect 13718 7404 13763 7412
rect 13450 7386 13469 7388
rect 13484 7386 13530 7388
rect 13450 7370 13530 7386
rect 13557 7384 13592 7397
rect 13633 7394 13670 7397
rect 13633 7392 13675 7394
rect 13562 7381 13592 7384
rect 13571 7377 13578 7381
rect 13578 7376 13579 7377
rect 13537 7370 13547 7376
rect 13296 7362 13331 7370
rect 13296 7336 13297 7362
rect 13304 7336 13331 7362
rect 13239 7318 13269 7332
rect 13296 7328 13331 7336
rect 13333 7362 13374 7370
rect 13333 7336 13348 7362
rect 13355 7336 13374 7362
rect 13438 7358 13469 7370
rect 13484 7358 13587 7370
rect 13599 7360 13625 7386
rect 13640 7381 13670 7392
rect 13702 7388 13764 7404
rect 13702 7386 13748 7388
rect 13702 7370 13764 7386
rect 13776 7370 13782 7418
rect 13785 7410 13865 7418
rect 13785 7408 13804 7410
rect 13819 7408 13853 7410
rect 13785 7392 13865 7408
rect 13785 7370 13804 7392
rect 13819 7376 13849 7392
rect 13877 7386 13883 7460
rect 13886 7386 13905 7530
rect 13920 7386 13926 7530
rect 13935 7460 13948 7530
rect 14000 7526 14022 7530
rect 13993 7504 14022 7518
rect 14075 7504 14091 7518
rect 14129 7514 14135 7516
rect 14142 7514 14250 7530
rect 14257 7514 14263 7516
rect 14271 7514 14286 7530
rect 14352 7524 14371 7527
rect 13993 7502 14091 7504
rect 14118 7502 14286 7514
rect 14301 7504 14317 7518
rect 14352 7505 14374 7524
rect 14384 7518 14400 7519
rect 14383 7516 14400 7518
rect 14384 7511 14400 7516
rect 14374 7504 14380 7505
rect 14383 7504 14412 7511
rect 14301 7503 14412 7504
rect 14301 7502 14418 7503
rect 13977 7494 14028 7502
rect 14075 7494 14109 7502
rect 13977 7482 14002 7494
rect 14009 7482 14028 7494
rect 14082 7492 14109 7494
rect 14118 7492 14339 7502
rect 14374 7499 14380 7502
rect 14082 7488 14339 7492
rect 13977 7474 14028 7482
rect 14075 7474 14339 7488
rect 14383 7494 14418 7502
rect 13929 7426 13948 7460
rect 13993 7466 14022 7474
rect 13993 7460 14010 7466
rect 13993 7458 14027 7460
rect 14075 7458 14091 7474
rect 14092 7464 14300 7474
rect 14301 7464 14317 7474
rect 14365 7470 14380 7485
rect 14383 7482 14384 7494
rect 14391 7482 14418 7494
rect 14383 7474 14418 7482
rect 14383 7473 14412 7474
rect 14103 7460 14317 7464
rect 14118 7458 14317 7460
rect 14352 7460 14365 7470
rect 14383 7460 14400 7473
rect 14352 7458 14400 7460
rect 13994 7454 14027 7458
rect 13990 7452 14027 7454
rect 13990 7451 14057 7452
rect 13990 7446 14021 7451
rect 14027 7446 14057 7451
rect 13990 7442 14057 7446
rect 13963 7439 14057 7442
rect 13963 7432 14012 7439
rect 13963 7426 13993 7432
rect 14012 7427 14017 7432
rect 13929 7410 14009 7426
rect 14021 7418 14057 7439
rect 14118 7434 14307 7458
rect 14352 7457 14399 7458
rect 14365 7452 14399 7457
rect 14133 7431 14307 7434
rect 14126 7428 14307 7431
rect 14335 7451 14399 7452
rect 13929 7408 13948 7410
rect 13963 7408 13997 7410
rect 13929 7392 14009 7408
rect 13929 7386 13948 7392
rect 13645 7360 13748 7370
rect 13599 7358 13748 7360
rect 13769 7358 13804 7370
rect 13438 7356 13600 7358
rect 13450 7336 13469 7356
rect 13484 7354 13514 7356
rect 13333 7328 13374 7336
rect 13456 7332 13469 7336
rect 13521 7340 13600 7356
rect 13632 7356 13804 7358
rect 13632 7340 13711 7356
rect 13718 7354 13748 7356
rect 13296 7318 13325 7328
rect 13339 7318 13368 7328
rect 13383 7318 13413 7332
rect 13456 7318 13499 7332
rect 13521 7328 13711 7340
rect 13776 7336 13782 7356
rect 13506 7318 13536 7328
rect 13537 7318 13695 7328
rect 13699 7318 13729 7328
rect 13733 7318 13763 7332
rect 13791 7318 13804 7356
rect 13876 7370 13905 7386
rect 13919 7370 13948 7386
rect 13963 7376 13993 7392
rect 14021 7370 14027 7418
rect 14030 7412 14049 7418
rect 14064 7412 14094 7420
rect 14030 7404 14094 7412
rect 14030 7388 14110 7404
rect 14126 7397 14188 7428
rect 14204 7397 14266 7428
rect 14335 7426 14384 7451
rect 14399 7426 14429 7442
rect 14298 7412 14328 7420
rect 14335 7418 14445 7426
rect 14298 7404 14343 7412
rect 14030 7386 14049 7388
rect 14064 7386 14110 7388
rect 14030 7370 14110 7386
rect 14137 7384 14172 7397
rect 14213 7394 14250 7397
rect 14213 7392 14255 7394
rect 14142 7381 14172 7384
rect 14151 7377 14158 7381
rect 14158 7376 14159 7377
rect 14117 7370 14127 7376
rect 13876 7362 13911 7370
rect 13876 7336 13877 7362
rect 13884 7336 13911 7362
rect 13819 7318 13849 7332
rect 13876 7328 13911 7336
rect 13913 7362 13954 7370
rect 13913 7336 13928 7362
rect 13935 7336 13954 7362
rect 14018 7358 14049 7370
rect 14064 7358 14167 7370
rect 14179 7360 14205 7386
rect 14220 7381 14250 7392
rect 14282 7388 14344 7404
rect 14282 7386 14328 7388
rect 14282 7370 14344 7386
rect 14356 7370 14362 7418
rect 14365 7410 14445 7418
rect 14365 7408 14384 7410
rect 14399 7408 14433 7410
rect 14365 7392 14445 7408
rect 14365 7370 14384 7392
rect 14399 7376 14429 7392
rect 14457 7386 14463 7460
rect 14466 7386 14485 7530
rect 14500 7386 14506 7530
rect 14515 7460 14528 7530
rect 14580 7526 14602 7530
rect 14573 7504 14602 7518
rect 14655 7504 14671 7518
rect 14709 7514 14715 7516
rect 14722 7514 14830 7530
rect 14837 7514 14843 7516
rect 14851 7514 14866 7530
rect 14932 7524 14951 7527
rect 14573 7502 14671 7504
rect 14698 7502 14866 7514
rect 14881 7504 14897 7518
rect 14932 7505 14954 7524
rect 14964 7518 14980 7519
rect 14963 7516 14980 7518
rect 14964 7511 14980 7516
rect 14954 7504 14960 7505
rect 14963 7504 14992 7511
rect 14881 7503 14992 7504
rect 14881 7502 14998 7503
rect 14557 7494 14608 7502
rect 14655 7494 14689 7502
rect 14557 7482 14582 7494
rect 14589 7482 14608 7494
rect 14662 7492 14689 7494
rect 14698 7492 14919 7502
rect 14954 7499 14960 7502
rect 14662 7488 14919 7492
rect 14557 7474 14608 7482
rect 14655 7474 14919 7488
rect 14963 7494 14998 7502
rect 14509 7426 14528 7460
rect 14573 7466 14602 7474
rect 14573 7460 14590 7466
rect 14573 7458 14607 7460
rect 14655 7458 14671 7474
rect 14672 7464 14880 7474
rect 14881 7464 14897 7474
rect 14945 7470 14960 7485
rect 14963 7482 14964 7494
rect 14971 7482 14998 7494
rect 14963 7474 14998 7482
rect 14963 7473 14992 7474
rect 14683 7460 14897 7464
rect 14698 7458 14897 7460
rect 14932 7460 14945 7470
rect 14963 7460 14980 7473
rect 14932 7458 14980 7460
rect 14574 7454 14607 7458
rect 14570 7452 14607 7454
rect 14570 7451 14637 7452
rect 14570 7446 14601 7451
rect 14607 7446 14637 7451
rect 14570 7442 14637 7446
rect 14543 7439 14637 7442
rect 14543 7432 14592 7439
rect 14543 7426 14573 7432
rect 14592 7427 14597 7432
rect 14509 7410 14589 7426
rect 14601 7418 14637 7439
rect 14698 7434 14887 7458
rect 14932 7457 14979 7458
rect 14945 7452 14979 7457
rect 14713 7431 14887 7434
rect 14706 7428 14887 7431
rect 14915 7451 14979 7452
rect 14509 7408 14528 7410
rect 14543 7408 14577 7410
rect 14509 7392 14589 7408
rect 14509 7386 14528 7392
rect 14225 7360 14328 7370
rect 14179 7358 14328 7360
rect 14349 7358 14384 7370
rect 14018 7356 14180 7358
rect 14030 7336 14049 7356
rect 14064 7354 14094 7356
rect 13913 7328 13954 7336
rect 14036 7332 14049 7336
rect 14101 7340 14180 7356
rect 14212 7356 14384 7358
rect 14212 7340 14291 7356
rect 14298 7354 14328 7356
rect 13876 7318 13905 7328
rect 13919 7318 13948 7328
rect 13963 7318 13993 7332
rect 14036 7318 14079 7332
rect 14101 7328 14291 7340
rect 14356 7336 14362 7356
rect 14086 7318 14116 7328
rect 14117 7318 14275 7328
rect 14279 7318 14309 7328
rect 14313 7318 14343 7332
rect 14371 7318 14384 7356
rect 14456 7370 14485 7386
rect 14499 7370 14528 7386
rect 14543 7376 14573 7392
rect 14601 7370 14607 7418
rect 14610 7412 14629 7418
rect 14644 7412 14674 7420
rect 14610 7404 14674 7412
rect 14610 7388 14690 7404
rect 14706 7397 14768 7428
rect 14784 7397 14846 7428
rect 14915 7426 14964 7451
rect 14979 7426 15009 7442
rect 14878 7412 14908 7420
rect 14915 7418 15025 7426
rect 14878 7404 14923 7412
rect 14610 7386 14629 7388
rect 14644 7386 14690 7388
rect 14610 7370 14690 7386
rect 14717 7384 14752 7397
rect 14793 7394 14830 7397
rect 14793 7392 14835 7394
rect 14722 7381 14752 7384
rect 14731 7377 14738 7381
rect 14738 7376 14739 7377
rect 14697 7370 14707 7376
rect 14456 7362 14491 7370
rect 14456 7336 14457 7362
rect 14464 7336 14491 7362
rect 14399 7318 14429 7332
rect 14456 7328 14491 7336
rect 14493 7362 14534 7370
rect 14493 7336 14508 7362
rect 14515 7336 14534 7362
rect 14598 7358 14629 7370
rect 14644 7358 14747 7370
rect 14759 7360 14785 7386
rect 14800 7381 14830 7392
rect 14862 7388 14924 7404
rect 14862 7386 14908 7388
rect 14862 7370 14924 7386
rect 14936 7370 14942 7418
rect 14945 7410 15025 7418
rect 14945 7408 14964 7410
rect 14979 7408 15013 7410
rect 14945 7392 15025 7408
rect 14945 7370 14964 7392
rect 14979 7376 15009 7392
rect 15037 7386 15043 7460
rect 15046 7386 15065 7530
rect 15080 7386 15086 7530
rect 15095 7460 15108 7530
rect 15160 7526 15182 7530
rect 15153 7504 15182 7518
rect 15235 7504 15251 7518
rect 15289 7514 15295 7516
rect 15302 7514 15410 7530
rect 15417 7514 15423 7516
rect 15431 7514 15446 7530
rect 15512 7524 15531 7527
rect 15153 7502 15251 7504
rect 15278 7502 15446 7514
rect 15461 7504 15477 7518
rect 15512 7505 15534 7524
rect 15544 7518 15560 7519
rect 15543 7516 15560 7518
rect 15544 7511 15560 7516
rect 15534 7504 15540 7505
rect 15543 7504 15572 7511
rect 15461 7503 15572 7504
rect 15461 7502 15578 7503
rect 15137 7494 15188 7502
rect 15235 7494 15269 7502
rect 15137 7482 15162 7494
rect 15169 7482 15188 7494
rect 15242 7492 15269 7494
rect 15278 7492 15499 7502
rect 15534 7499 15540 7502
rect 15242 7488 15499 7492
rect 15137 7474 15188 7482
rect 15235 7474 15499 7488
rect 15543 7494 15578 7502
rect 15089 7426 15108 7460
rect 15153 7466 15182 7474
rect 15153 7460 15170 7466
rect 15153 7458 15187 7460
rect 15235 7458 15251 7474
rect 15252 7464 15460 7474
rect 15461 7464 15477 7474
rect 15525 7470 15540 7485
rect 15543 7482 15544 7494
rect 15551 7482 15578 7494
rect 15543 7474 15578 7482
rect 15543 7473 15572 7474
rect 15263 7460 15477 7464
rect 15278 7458 15477 7460
rect 15512 7460 15525 7470
rect 15543 7460 15560 7473
rect 15512 7458 15560 7460
rect 15154 7454 15187 7458
rect 15150 7452 15187 7454
rect 15150 7451 15217 7452
rect 15150 7446 15181 7451
rect 15187 7446 15217 7451
rect 15150 7442 15217 7446
rect 15123 7439 15217 7442
rect 15123 7432 15172 7439
rect 15123 7426 15153 7432
rect 15172 7427 15177 7432
rect 15089 7410 15169 7426
rect 15181 7418 15217 7439
rect 15278 7434 15467 7458
rect 15512 7457 15559 7458
rect 15525 7452 15559 7457
rect 15293 7431 15467 7434
rect 15286 7428 15467 7431
rect 15495 7451 15559 7452
rect 15089 7408 15108 7410
rect 15123 7408 15157 7410
rect 15089 7392 15169 7408
rect 15089 7386 15108 7392
rect 14805 7360 14908 7370
rect 14759 7358 14908 7360
rect 14929 7358 14964 7370
rect 14598 7356 14760 7358
rect 14610 7336 14629 7356
rect 14644 7354 14674 7356
rect 14493 7328 14534 7336
rect 14616 7332 14629 7336
rect 14681 7340 14760 7356
rect 14792 7356 14964 7358
rect 14792 7340 14871 7356
rect 14878 7354 14908 7356
rect 14456 7318 14485 7328
rect 14499 7318 14528 7328
rect 14543 7318 14573 7332
rect 14616 7318 14659 7332
rect 14681 7328 14871 7340
rect 14936 7336 14942 7356
rect 14666 7318 14696 7328
rect 14697 7318 14855 7328
rect 14859 7318 14889 7328
rect 14893 7318 14923 7332
rect 14951 7318 14964 7356
rect 15036 7370 15065 7386
rect 15079 7370 15108 7386
rect 15123 7376 15153 7392
rect 15181 7370 15187 7418
rect 15190 7412 15209 7418
rect 15224 7412 15254 7420
rect 15190 7404 15254 7412
rect 15190 7388 15270 7404
rect 15286 7397 15348 7428
rect 15364 7397 15426 7428
rect 15495 7426 15544 7451
rect 15559 7426 15589 7442
rect 15458 7412 15488 7420
rect 15495 7418 15605 7426
rect 15458 7404 15503 7412
rect 15190 7386 15209 7388
rect 15224 7386 15270 7388
rect 15190 7370 15270 7386
rect 15297 7384 15332 7397
rect 15373 7394 15410 7397
rect 15373 7392 15415 7394
rect 15302 7381 15332 7384
rect 15311 7377 15318 7381
rect 15318 7376 15319 7377
rect 15277 7370 15287 7376
rect 15036 7362 15071 7370
rect 15036 7336 15037 7362
rect 15044 7336 15071 7362
rect 14979 7318 15009 7332
rect 15036 7328 15071 7336
rect 15073 7362 15114 7370
rect 15073 7336 15088 7362
rect 15095 7336 15114 7362
rect 15178 7358 15209 7370
rect 15224 7358 15327 7370
rect 15339 7360 15365 7386
rect 15380 7381 15410 7392
rect 15442 7388 15504 7404
rect 15442 7386 15488 7388
rect 15442 7370 15504 7386
rect 15516 7370 15522 7418
rect 15525 7410 15605 7418
rect 15525 7408 15544 7410
rect 15559 7408 15593 7410
rect 15525 7392 15605 7408
rect 15525 7370 15544 7392
rect 15559 7376 15589 7392
rect 15617 7386 15623 7460
rect 15626 7386 15645 7530
rect 15660 7386 15666 7530
rect 15675 7460 15688 7530
rect 15740 7526 15762 7530
rect 15733 7504 15762 7518
rect 15815 7504 15831 7518
rect 15869 7514 15875 7516
rect 15882 7514 15990 7530
rect 15997 7514 16003 7516
rect 16011 7514 16026 7530
rect 16092 7524 16111 7527
rect 15733 7502 15831 7504
rect 15858 7502 16026 7514
rect 16041 7504 16057 7518
rect 16092 7505 16114 7524
rect 16124 7518 16140 7519
rect 16123 7516 16140 7518
rect 16124 7511 16140 7516
rect 16114 7504 16120 7505
rect 16123 7504 16152 7511
rect 16041 7503 16152 7504
rect 16041 7502 16158 7503
rect 15717 7494 15768 7502
rect 15815 7494 15849 7502
rect 15717 7482 15742 7494
rect 15749 7482 15768 7494
rect 15822 7492 15849 7494
rect 15858 7492 16079 7502
rect 16114 7499 16120 7502
rect 15822 7488 16079 7492
rect 15717 7474 15768 7482
rect 15815 7474 16079 7488
rect 16123 7494 16158 7502
rect 15669 7426 15688 7460
rect 15733 7466 15762 7474
rect 15733 7460 15750 7466
rect 15733 7458 15767 7460
rect 15815 7458 15831 7474
rect 15832 7464 16040 7474
rect 16041 7464 16057 7474
rect 16105 7470 16120 7485
rect 16123 7482 16124 7494
rect 16131 7482 16158 7494
rect 16123 7474 16158 7482
rect 16123 7473 16152 7474
rect 15843 7460 16057 7464
rect 15858 7458 16057 7460
rect 16092 7460 16105 7470
rect 16123 7460 16140 7473
rect 16092 7458 16140 7460
rect 15734 7454 15767 7458
rect 15730 7452 15767 7454
rect 15730 7451 15797 7452
rect 15730 7446 15761 7451
rect 15767 7446 15797 7451
rect 15730 7442 15797 7446
rect 15703 7439 15797 7442
rect 15703 7432 15752 7439
rect 15703 7426 15733 7432
rect 15752 7427 15757 7432
rect 15669 7410 15749 7426
rect 15761 7418 15797 7439
rect 15858 7434 16047 7458
rect 16092 7457 16139 7458
rect 16105 7452 16139 7457
rect 15873 7431 16047 7434
rect 15866 7428 16047 7431
rect 16075 7451 16139 7452
rect 15669 7408 15688 7410
rect 15703 7408 15737 7410
rect 15669 7392 15749 7408
rect 15669 7386 15688 7392
rect 15385 7360 15488 7370
rect 15339 7358 15488 7360
rect 15509 7358 15544 7370
rect 15178 7356 15340 7358
rect 15190 7336 15209 7356
rect 15224 7354 15254 7356
rect 15073 7328 15114 7336
rect 15196 7332 15209 7336
rect 15261 7340 15340 7356
rect 15372 7356 15544 7358
rect 15372 7340 15451 7356
rect 15458 7354 15488 7356
rect 15036 7318 15065 7328
rect 15079 7318 15108 7328
rect 15123 7318 15153 7332
rect 15196 7318 15239 7332
rect 15261 7328 15451 7340
rect 15516 7336 15522 7356
rect 15246 7318 15276 7328
rect 15277 7318 15435 7328
rect 15439 7318 15469 7328
rect 15473 7318 15503 7332
rect 15531 7318 15544 7356
rect 15616 7370 15645 7386
rect 15659 7370 15688 7386
rect 15703 7376 15733 7392
rect 15761 7370 15767 7418
rect 15770 7412 15789 7418
rect 15804 7412 15834 7420
rect 15770 7404 15834 7412
rect 15770 7388 15850 7404
rect 15866 7397 15928 7428
rect 15944 7397 16006 7428
rect 16075 7426 16124 7451
rect 16139 7426 16169 7442
rect 16038 7412 16068 7420
rect 16075 7418 16185 7426
rect 16038 7404 16083 7412
rect 15770 7386 15789 7388
rect 15804 7386 15850 7388
rect 15770 7370 15850 7386
rect 15877 7384 15912 7397
rect 15953 7394 15990 7397
rect 15953 7392 15995 7394
rect 15882 7381 15912 7384
rect 15891 7377 15898 7381
rect 15898 7376 15899 7377
rect 15857 7370 15867 7376
rect 15616 7362 15651 7370
rect 15616 7336 15617 7362
rect 15624 7336 15651 7362
rect 15559 7318 15589 7332
rect 15616 7328 15651 7336
rect 15653 7362 15694 7370
rect 15653 7336 15668 7362
rect 15675 7336 15694 7362
rect 15758 7358 15789 7370
rect 15804 7358 15907 7370
rect 15919 7360 15945 7386
rect 15960 7381 15990 7392
rect 16022 7388 16084 7404
rect 16022 7386 16068 7388
rect 16022 7370 16084 7386
rect 16096 7370 16102 7418
rect 16105 7410 16185 7418
rect 16105 7408 16124 7410
rect 16139 7408 16173 7410
rect 16105 7392 16185 7408
rect 16105 7370 16124 7392
rect 16139 7376 16169 7392
rect 16197 7386 16203 7460
rect 16206 7386 16225 7530
rect 16240 7386 16246 7530
rect 16255 7460 16268 7530
rect 16320 7526 16342 7530
rect 16313 7504 16342 7518
rect 16395 7504 16411 7518
rect 16449 7514 16455 7516
rect 16462 7514 16570 7530
rect 16577 7514 16583 7516
rect 16591 7514 16606 7530
rect 16672 7524 16691 7527
rect 16313 7502 16411 7504
rect 16438 7502 16606 7514
rect 16621 7504 16637 7518
rect 16672 7505 16694 7524
rect 16704 7518 16720 7519
rect 16703 7516 16720 7518
rect 16704 7511 16720 7516
rect 16694 7504 16700 7505
rect 16703 7504 16732 7511
rect 16621 7503 16732 7504
rect 16621 7502 16738 7503
rect 16297 7494 16348 7502
rect 16395 7494 16429 7502
rect 16297 7482 16322 7494
rect 16329 7482 16348 7494
rect 16402 7492 16429 7494
rect 16438 7492 16659 7502
rect 16694 7499 16700 7502
rect 16402 7488 16659 7492
rect 16297 7474 16348 7482
rect 16395 7474 16659 7488
rect 16703 7494 16738 7502
rect 16249 7426 16268 7460
rect 16313 7466 16342 7474
rect 16313 7460 16330 7466
rect 16313 7458 16347 7460
rect 16395 7458 16411 7474
rect 16412 7464 16620 7474
rect 16621 7464 16637 7474
rect 16685 7470 16700 7485
rect 16703 7482 16704 7494
rect 16711 7482 16738 7494
rect 16703 7474 16738 7482
rect 16703 7473 16732 7474
rect 16423 7460 16637 7464
rect 16438 7458 16637 7460
rect 16672 7460 16685 7470
rect 16703 7460 16720 7473
rect 16672 7458 16720 7460
rect 16314 7454 16347 7458
rect 16310 7452 16347 7454
rect 16310 7451 16377 7452
rect 16310 7446 16341 7451
rect 16347 7446 16377 7451
rect 16310 7442 16377 7446
rect 16283 7439 16377 7442
rect 16283 7432 16332 7439
rect 16283 7426 16313 7432
rect 16332 7427 16337 7432
rect 16249 7410 16329 7426
rect 16341 7418 16377 7439
rect 16438 7434 16627 7458
rect 16672 7457 16719 7458
rect 16685 7452 16719 7457
rect 16453 7431 16627 7434
rect 16446 7428 16627 7431
rect 16655 7451 16719 7452
rect 16249 7408 16268 7410
rect 16283 7408 16317 7410
rect 16249 7392 16329 7408
rect 16249 7386 16268 7392
rect 15965 7360 16068 7370
rect 15919 7358 16068 7360
rect 16089 7358 16124 7370
rect 15758 7356 15920 7358
rect 15770 7336 15789 7356
rect 15804 7354 15834 7356
rect 15653 7328 15694 7336
rect 15776 7332 15789 7336
rect 15841 7340 15920 7356
rect 15952 7356 16124 7358
rect 15952 7340 16031 7356
rect 16038 7354 16068 7356
rect 15616 7318 15645 7328
rect 15659 7318 15688 7328
rect 15703 7318 15733 7332
rect 15776 7318 15819 7332
rect 15841 7328 16031 7340
rect 16096 7336 16102 7356
rect 15826 7318 15856 7328
rect 15857 7318 16015 7328
rect 16019 7318 16049 7328
rect 16053 7318 16083 7332
rect 16111 7318 16124 7356
rect 16196 7370 16225 7386
rect 16239 7370 16268 7386
rect 16283 7376 16313 7392
rect 16341 7370 16347 7418
rect 16350 7412 16369 7418
rect 16384 7412 16414 7420
rect 16350 7404 16414 7412
rect 16350 7388 16430 7404
rect 16446 7397 16508 7428
rect 16524 7397 16586 7428
rect 16655 7426 16704 7451
rect 16719 7426 16749 7442
rect 16618 7412 16648 7420
rect 16655 7418 16765 7426
rect 16618 7404 16663 7412
rect 16350 7386 16369 7388
rect 16384 7386 16430 7388
rect 16350 7370 16430 7386
rect 16457 7384 16492 7397
rect 16533 7394 16570 7397
rect 16533 7392 16575 7394
rect 16462 7381 16492 7384
rect 16471 7377 16478 7381
rect 16478 7376 16479 7377
rect 16437 7370 16447 7376
rect 16196 7362 16231 7370
rect 16196 7336 16197 7362
rect 16204 7336 16231 7362
rect 16139 7318 16169 7332
rect 16196 7328 16231 7336
rect 16233 7362 16274 7370
rect 16233 7336 16248 7362
rect 16255 7336 16274 7362
rect 16338 7358 16369 7370
rect 16384 7358 16487 7370
rect 16499 7360 16525 7386
rect 16540 7381 16570 7392
rect 16602 7388 16664 7404
rect 16602 7386 16648 7388
rect 16602 7370 16664 7386
rect 16676 7370 16682 7418
rect 16685 7410 16765 7418
rect 16685 7408 16704 7410
rect 16719 7408 16753 7410
rect 16685 7392 16765 7408
rect 16685 7370 16704 7392
rect 16719 7376 16749 7392
rect 16777 7386 16783 7460
rect 16786 7386 16805 7530
rect 16820 7386 16826 7530
rect 16835 7460 16848 7530
rect 16900 7526 16922 7530
rect 16893 7504 16922 7518
rect 16975 7504 16991 7518
rect 17029 7514 17035 7516
rect 17042 7514 17150 7530
rect 17157 7514 17163 7516
rect 17171 7514 17186 7530
rect 17252 7524 17271 7527
rect 16893 7502 16991 7504
rect 17018 7502 17186 7514
rect 17201 7504 17217 7518
rect 17252 7505 17274 7524
rect 17284 7518 17300 7519
rect 17283 7516 17300 7518
rect 17284 7511 17300 7516
rect 17274 7504 17280 7505
rect 17283 7504 17312 7511
rect 17201 7503 17312 7504
rect 17201 7502 17318 7503
rect 16877 7494 16928 7502
rect 16975 7494 17009 7502
rect 16877 7482 16902 7494
rect 16909 7482 16928 7494
rect 16982 7492 17009 7494
rect 17018 7492 17239 7502
rect 17274 7499 17280 7502
rect 16982 7488 17239 7492
rect 16877 7474 16928 7482
rect 16975 7474 17239 7488
rect 17283 7494 17318 7502
rect 16829 7426 16848 7460
rect 16893 7466 16922 7474
rect 16893 7460 16910 7466
rect 16893 7458 16927 7460
rect 16975 7458 16991 7474
rect 16992 7464 17200 7474
rect 17201 7464 17217 7474
rect 17265 7470 17280 7485
rect 17283 7482 17284 7494
rect 17291 7482 17318 7494
rect 17283 7474 17318 7482
rect 17283 7473 17312 7474
rect 17003 7460 17217 7464
rect 17018 7458 17217 7460
rect 17252 7460 17265 7470
rect 17283 7460 17300 7473
rect 17252 7458 17300 7460
rect 16894 7454 16927 7458
rect 16890 7452 16927 7454
rect 16890 7451 16957 7452
rect 16890 7446 16921 7451
rect 16927 7446 16957 7451
rect 16890 7442 16957 7446
rect 16863 7439 16957 7442
rect 16863 7432 16912 7439
rect 16863 7426 16893 7432
rect 16912 7427 16917 7432
rect 16829 7410 16909 7426
rect 16921 7418 16957 7439
rect 17018 7434 17207 7458
rect 17252 7457 17299 7458
rect 17265 7452 17299 7457
rect 17033 7431 17207 7434
rect 17026 7428 17207 7431
rect 17235 7451 17299 7452
rect 16829 7408 16848 7410
rect 16863 7408 16897 7410
rect 16829 7392 16909 7408
rect 16829 7386 16848 7392
rect 16545 7360 16648 7370
rect 16499 7358 16648 7360
rect 16669 7358 16704 7370
rect 16338 7356 16500 7358
rect 16350 7336 16369 7356
rect 16384 7354 16414 7356
rect 16233 7328 16274 7336
rect 16356 7332 16369 7336
rect 16421 7340 16500 7356
rect 16532 7356 16704 7358
rect 16532 7340 16611 7356
rect 16618 7354 16648 7356
rect 16196 7318 16225 7328
rect 16239 7318 16268 7328
rect 16283 7318 16313 7332
rect 16356 7318 16399 7332
rect 16421 7328 16611 7340
rect 16676 7336 16682 7356
rect 16406 7318 16436 7328
rect 16437 7318 16595 7328
rect 16599 7318 16629 7328
rect 16633 7318 16663 7332
rect 16691 7318 16704 7356
rect 16776 7370 16805 7386
rect 16819 7370 16848 7386
rect 16863 7376 16893 7392
rect 16921 7370 16927 7418
rect 16930 7412 16949 7418
rect 16964 7412 16994 7420
rect 16930 7404 16994 7412
rect 16930 7388 17010 7404
rect 17026 7397 17088 7428
rect 17104 7397 17166 7428
rect 17235 7426 17284 7451
rect 17299 7426 17329 7442
rect 17198 7412 17228 7420
rect 17235 7418 17345 7426
rect 17198 7404 17243 7412
rect 16930 7386 16949 7388
rect 16964 7386 17010 7388
rect 16930 7370 17010 7386
rect 17037 7384 17072 7397
rect 17113 7394 17150 7397
rect 17113 7392 17155 7394
rect 17042 7381 17072 7384
rect 17051 7377 17058 7381
rect 17058 7376 17059 7377
rect 17017 7370 17027 7376
rect 16776 7362 16811 7370
rect 16776 7336 16777 7362
rect 16784 7336 16811 7362
rect 16719 7318 16749 7332
rect 16776 7328 16811 7336
rect 16813 7362 16854 7370
rect 16813 7336 16828 7362
rect 16835 7336 16854 7362
rect 16918 7358 16949 7370
rect 16964 7358 17067 7370
rect 17079 7360 17105 7386
rect 17120 7381 17150 7392
rect 17182 7388 17244 7404
rect 17182 7386 17228 7388
rect 17182 7370 17244 7386
rect 17256 7370 17262 7418
rect 17265 7410 17345 7418
rect 17265 7408 17284 7410
rect 17299 7408 17333 7410
rect 17265 7392 17345 7408
rect 17265 7370 17284 7392
rect 17299 7376 17329 7392
rect 17357 7386 17363 7460
rect 17366 7386 17385 7530
rect 17400 7386 17406 7530
rect 17415 7460 17428 7530
rect 17480 7526 17502 7530
rect 17473 7504 17502 7518
rect 17555 7504 17571 7518
rect 17609 7514 17615 7516
rect 17622 7514 17730 7530
rect 17737 7514 17743 7516
rect 17751 7514 17766 7530
rect 17832 7524 17851 7527
rect 17473 7502 17571 7504
rect 17598 7502 17766 7514
rect 17781 7504 17797 7518
rect 17832 7505 17854 7524
rect 17864 7518 17880 7519
rect 17863 7516 17880 7518
rect 17864 7511 17880 7516
rect 17854 7504 17860 7505
rect 17863 7504 17892 7511
rect 17781 7503 17892 7504
rect 17781 7502 17898 7503
rect 17457 7494 17508 7502
rect 17555 7494 17589 7502
rect 17457 7482 17482 7494
rect 17489 7482 17508 7494
rect 17562 7492 17589 7494
rect 17598 7492 17819 7502
rect 17854 7499 17860 7502
rect 17562 7488 17819 7492
rect 17457 7474 17508 7482
rect 17555 7474 17819 7488
rect 17863 7494 17898 7502
rect 17409 7426 17428 7460
rect 17473 7466 17502 7474
rect 17473 7460 17490 7466
rect 17473 7458 17507 7460
rect 17555 7458 17571 7474
rect 17572 7464 17780 7474
rect 17781 7464 17797 7474
rect 17845 7470 17860 7485
rect 17863 7482 17864 7494
rect 17871 7482 17898 7494
rect 17863 7474 17898 7482
rect 17863 7473 17892 7474
rect 17583 7460 17797 7464
rect 17598 7458 17797 7460
rect 17832 7460 17845 7470
rect 17863 7460 17880 7473
rect 17832 7458 17880 7460
rect 17474 7454 17507 7458
rect 17470 7452 17507 7454
rect 17470 7451 17537 7452
rect 17470 7446 17501 7451
rect 17507 7446 17537 7451
rect 17470 7442 17537 7446
rect 17443 7439 17537 7442
rect 17443 7432 17492 7439
rect 17443 7426 17473 7432
rect 17492 7427 17497 7432
rect 17409 7410 17489 7426
rect 17501 7418 17537 7439
rect 17598 7434 17787 7458
rect 17832 7457 17879 7458
rect 17845 7452 17879 7457
rect 17613 7431 17787 7434
rect 17606 7428 17787 7431
rect 17815 7451 17879 7452
rect 17409 7408 17428 7410
rect 17443 7408 17477 7410
rect 17409 7392 17489 7408
rect 17409 7386 17428 7392
rect 17125 7360 17228 7370
rect 17079 7358 17228 7360
rect 17249 7358 17284 7370
rect 16918 7356 17080 7358
rect 16930 7336 16949 7356
rect 16964 7354 16994 7356
rect 16813 7328 16854 7336
rect 16936 7332 16949 7336
rect 17001 7340 17080 7356
rect 17112 7356 17284 7358
rect 17112 7340 17191 7356
rect 17198 7354 17228 7356
rect 16776 7318 16805 7328
rect 16819 7318 16848 7328
rect 16863 7318 16893 7332
rect 16936 7318 16979 7332
rect 17001 7328 17191 7340
rect 17256 7336 17262 7356
rect 16986 7318 17016 7328
rect 17017 7318 17175 7328
rect 17179 7318 17209 7328
rect 17213 7318 17243 7332
rect 17271 7318 17284 7356
rect 17356 7370 17385 7386
rect 17399 7370 17428 7386
rect 17443 7376 17473 7392
rect 17501 7370 17507 7418
rect 17510 7412 17529 7418
rect 17544 7412 17574 7420
rect 17510 7404 17574 7412
rect 17510 7388 17590 7404
rect 17606 7397 17668 7428
rect 17684 7397 17746 7428
rect 17815 7426 17864 7451
rect 17879 7426 17909 7442
rect 17778 7412 17808 7420
rect 17815 7418 17925 7426
rect 17778 7404 17823 7412
rect 17510 7386 17529 7388
rect 17544 7386 17590 7388
rect 17510 7370 17590 7386
rect 17617 7384 17652 7397
rect 17693 7394 17730 7397
rect 17693 7392 17735 7394
rect 17622 7381 17652 7384
rect 17631 7377 17638 7381
rect 17638 7376 17639 7377
rect 17597 7370 17607 7376
rect 17356 7362 17391 7370
rect 17356 7336 17357 7362
rect 17364 7336 17391 7362
rect 17299 7318 17329 7332
rect 17356 7328 17391 7336
rect 17393 7362 17434 7370
rect 17393 7336 17408 7362
rect 17415 7336 17434 7362
rect 17498 7358 17529 7370
rect 17544 7358 17647 7370
rect 17659 7360 17685 7386
rect 17700 7381 17730 7392
rect 17762 7388 17824 7404
rect 17762 7386 17808 7388
rect 17762 7370 17824 7386
rect 17836 7370 17842 7418
rect 17845 7410 17925 7418
rect 17845 7408 17864 7410
rect 17879 7408 17913 7410
rect 17845 7392 17925 7408
rect 17845 7370 17864 7392
rect 17879 7376 17909 7392
rect 17937 7386 17943 7460
rect 17946 7386 17965 7530
rect 17980 7386 17986 7530
rect 17995 7460 18008 7530
rect 18060 7526 18082 7530
rect 18053 7504 18082 7518
rect 18135 7504 18151 7518
rect 18189 7514 18195 7516
rect 18202 7514 18310 7530
rect 18317 7514 18323 7516
rect 18331 7514 18346 7530
rect 18412 7524 18431 7527
rect 18053 7502 18151 7504
rect 18178 7502 18346 7514
rect 18361 7504 18377 7518
rect 18412 7505 18434 7524
rect 18444 7518 18460 7519
rect 18443 7516 18460 7518
rect 18444 7511 18460 7516
rect 18434 7504 18440 7505
rect 18443 7504 18472 7511
rect 18361 7503 18472 7504
rect 18361 7502 18478 7503
rect 18037 7494 18088 7502
rect 18135 7494 18169 7502
rect 18037 7482 18062 7494
rect 18069 7482 18088 7494
rect 18142 7492 18169 7494
rect 18178 7492 18399 7502
rect 18434 7499 18440 7502
rect 18142 7488 18399 7492
rect 18037 7474 18088 7482
rect 18135 7474 18399 7488
rect 18443 7494 18478 7502
rect 17989 7426 18008 7460
rect 18053 7466 18082 7474
rect 18053 7460 18070 7466
rect 18053 7458 18087 7460
rect 18135 7458 18151 7474
rect 18152 7464 18360 7474
rect 18361 7464 18377 7474
rect 18425 7470 18440 7485
rect 18443 7482 18444 7494
rect 18451 7482 18478 7494
rect 18443 7474 18478 7482
rect 18443 7473 18472 7474
rect 18163 7460 18377 7464
rect 18178 7458 18377 7460
rect 18412 7460 18425 7470
rect 18443 7460 18460 7473
rect 18412 7458 18460 7460
rect 18054 7454 18087 7458
rect 18050 7452 18087 7454
rect 18050 7451 18117 7452
rect 18050 7446 18081 7451
rect 18087 7446 18117 7451
rect 18050 7442 18117 7446
rect 18023 7439 18117 7442
rect 18023 7432 18072 7439
rect 18023 7426 18053 7432
rect 18072 7427 18077 7432
rect 17989 7410 18069 7426
rect 18081 7418 18117 7439
rect 18178 7434 18367 7458
rect 18412 7457 18459 7458
rect 18425 7452 18459 7457
rect 18193 7431 18367 7434
rect 18186 7428 18367 7431
rect 18395 7451 18459 7452
rect 17989 7408 18008 7410
rect 18023 7408 18057 7410
rect 17989 7392 18069 7408
rect 17989 7386 18008 7392
rect 17705 7360 17808 7370
rect 17659 7358 17808 7360
rect 17829 7358 17864 7370
rect 17498 7356 17660 7358
rect 17510 7336 17529 7356
rect 17544 7354 17574 7356
rect 17393 7328 17434 7336
rect 17516 7332 17529 7336
rect 17581 7340 17660 7356
rect 17692 7356 17864 7358
rect 17692 7340 17771 7356
rect 17778 7354 17808 7356
rect 17356 7318 17385 7328
rect 17399 7318 17428 7328
rect 17443 7318 17473 7332
rect 17516 7318 17559 7332
rect 17581 7328 17771 7340
rect 17836 7336 17842 7356
rect 17566 7318 17596 7328
rect 17597 7318 17755 7328
rect 17759 7318 17789 7328
rect 17793 7318 17823 7332
rect 17851 7318 17864 7356
rect 17936 7370 17965 7386
rect 17979 7370 18008 7386
rect 18023 7376 18053 7392
rect 18081 7370 18087 7418
rect 18090 7412 18109 7418
rect 18124 7412 18154 7420
rect 18090 7404 18154 7412
rect 18090 7388 18170 7404
rect 18186 7397 18248 7428
rect 18264 7397 18326 7428
rect 18395 7426 18444 7451
rect 18459 7426 18489 7442
rect 18358 7412 18388 7420
rect 18395 7418 18505 7426
rect 18358 7404 18403 7412
rect 18090 7386 18109 7388
rect 18124 7386 18170 7388
rect 18090 7370 18170 7386
rect 18197 7384 18232 7397
rect 18273 7394 18310 7397
rect 18273 7392 18315 7394
rect 18202 7381 18232 7384
rect 18211 7377 18218 7381
rect 18218 7376 18219 7377
rect 18177 7370 18187 7376
rect 17936 7362 17971 7370
rect 17936 7336 17937 7362
rect 17944 7336 17971 7362
rect 17879 7318 17909 7332
rect 17936 7328 17971 7336
rect 17973 7362 18014 7370
rect 17973 7336 17988 7362
rect 17995 7336 18014 7362
rect 18078 7358 18109 7370
rect 18124 7358 18227 7370
rect 18239 7360 18265 7386
rect 18280 7381 18310 7392
rect 18342 7388 18404 7404
rect 18342 7386 18388 7388
rect 18342 7370 18404 7386
rect 18416 7370 18422 7418
rect 18425 7410 18505 7418
rect 18425 7408 18444 7410
rect 18459 7408 18493 7410
rect 18425 7392 18505 7408
rect 18425 7370 18444 7392
rect 18459 7376 18489 7392
rect 18517 7386 18523 7460
rect 18532 7386 18545 7530
rect 18285 7360 18388 7370
rect 18239 7358 18388 7360
rect 18409 7358 18444 7370
rect 18078 7356 18240 7358
rect 18090 7336 18109 7356
rect 18124 7354 18154 7356
rect 17973 7328 18014 7336
rect 18096 7332 18109 7336
rect 18161 7340 18240 7356
rect 18272 7356 18444 7358
rect 18272 7340 18351 7356
rect 18358 7354 18388 7356
rect 17936 7318 17965 7328
rect 17979 7318 18008 7328
rect 18023 7318 18053 7332
rect 18096 7318 18139 7332
rect 18161 7328 18351 7340
rect 18416 7336 18422 7356
rect 18146 7318 18176 7328
rect 18177 7318 18335 7328
rect 18339 7318 18369 7328
rect 18373 7318 18403 7332
rect 18431 7318 18444 7356
rect 18516 7370 18545 7386
rect 18516 7362 18551 7370
rect 18516 7336 18517 7362
rect 18524 7336 18551 7362
rect 18459 7318 18489 7332
rect 18516 7328 18551 7336
rect 18516 7318 18545 7328
rect -1 7312 18545 7318
rect 0 7304 18545 7312
rect 15 7274 28 7304
rect 43 7290 73 7304
rect 116 7290 159 7304
rect 166 7290 386 7304
rect 393 7290 423 7304
rect 83 7276 98 7288
rect 117 7276 130 7290
rect 198 7286 351 7290
rect 80 7274 102 7276
rect 180 7274 372 7286
rect 451 7274 464 7304
rect 479 7290 509 7304
rect 546 7274 565 7304
rect 580 7274 586 7304
rect 595 7274 608 7304
rect 623 7290 653 7304
rect 696 7290 739 7304
rect 746 7290 966 7304
rect 973 7290 1003 7304
rect 663 7276 678 7288
rect 697 7276 710 7290
rect 778 7286 931 7290
rect 660 7274 682 7276
rect 760 7274 952 7286
rect 1031 7274 1044 7304
rect 1059 7290 1089 7304
rect 1126 7274 1145 7304
rect 1160 7274 1166 7304
rect 1175 7274 1188 7304
rect 1203 7290 1233 7304
rect 1276 7290 1319 7304
rect 1326 7290 1546 7304
rect 1553 7290 1583 7304
rect 1243 7276 1258 7288
rect 1277 7276 1290 7290
rect 1358 7286 1511 7290
rect 1240 7274 1262 7276
rect 1340 7274 1532 7286
rect 1611 7274 1624 7304
rect 1639 7290 1669 7304
rect 1706 7274 1725 7304
rect 1740 7274 1746 7304
rect 1755 7274 1768 7304
rect 1783 7290 1813 7304
rect 1856 7290 1899 7304
rect 1906 7290 2126 7304
rect 2133 7290 2163 7304
rect 1823 7276 1838 7288
rect 1857 7276 1870 7290
rect 1938 7286 2091 7290
rect 1820 7274 1842 7276
rect 1920 7274 2112 7286
rect 2191 7274 2204 7304
rect 2219 7290 2249 7304
rect 2286 7274 2305 7304
rect 2320 7274 2326 7304
rect 2335 7274 2348 7304
rect 2363 7290 2393 7304
rect 2436 7290 2479 7304
rect 2486 7290 2706 7304
rect 2713 7290 2743 7304
rect 2403 7276 2418 7288
rect 2437 7276 2450 7290
rect 2518 7286 2671 7290
rect 2400 7274 2422 7276
rect 2500 7274 2692 7286
rect 2771 7274 2784 7304
rect 2799 7290 2829 7304
rect 2866 7274 2885 7304
rect 2900 7274 2906 7304
rect 2915 7274 2928 7304
rect 2943 7290 2973 7304
rect 3016 7290 3059 7304
rect 3066 7290 3286 7304
rect 3293 7290 3323 7304
rect 2983 7276 2998 7288
rect 3017 7276 3030 7290
rect 3098 7286 3251 7290
rect 2980 7274 3002 7276
rect 3080 7274 3272 7286
rect 3351 7274 3364 7304
rect 3379 7290 3409 7304
rect 3446 7274 3465 7304
rect 3480 7274 3486 7304
rect 3495 7274 3508 7304
rect 3523 7290 3553 7304
rect 3596 7290 3639 7304
rect 3646 7290 3866 7304
rect 3873 7290 3903 7304
rect 3563 7276 3578 7288
rect 3597 7276 3610 7290
rect 3678 7286 3831 7290
rect 3560 7274 3582 7276
rect 3660 7274 3852 7286
rect 3931 7274 3944 7304
rect 3959 7290 3989 7304
rect 4026 7274 4045 7304
rect 4060 7274 4066 7304
rect 4075 7274 4088 7304
rect 4103 7290 4133 7304
rect 4176 7290 4219 7304
rect 4226 7290 4446 7304
rect 4453 7290 4483 7304
rect 4143 7276 4158 7288
rect 4177 7276 4190 7290
rect 4258 7286 4411 7290
rect 4140 7274 4162 7276
rect 4240 7274 4432 7286
rect 4511 7274 4524 7304
rect 4539 7290 4569 7304
rect 4606 7274 4625 7304
rect 4640 7274 4646 7304
rect 4655 7274 4668 7304
rect 4683 7290 4713 7304
rect 4756 7290 4799 7304
rect 4806 7290 5026 7304
rect 5033 7290 5063 7304
rect 4723 7276 4738 7288
rect 4757 7276 4770 7290
rect 4838 7286 4991 7290
rect 4720 7274 4742 7276
rect 4820 7274 5012 7286
rect 5091 7274 5104 7304
rect 5119 7290 5149 7304
rect 5186 7274 5205 7304
rect 5220 7274 5226 7304
rect 5235 7274 5248 7304
rect 5263 7290 5293 7304
rect 5336 7290 5379 7304
rect 5386 7290 5606 7304
rect 5613 7290 5643 7304
rect 5303 7276 5318 7288
rect 5337 7276 5350 7290
rect 5418 7286 5571 7290
rect 5300 7274 5322 7276
rect 5400 7274 5592 7286
rect 5671 7274 5684 7304
rect 5699 7290 5729 7304
rect 5766 7274 5785 7304
rect 5800 7274 5806 7304
rect 5815 7274 5828 7304
rect 5843 7290 5873 7304
rect 5916 7290 5959 7304
rect 5966 7290 6186 7304
rect 6193 7290 6223 7304
rect 5883 7276 5898 7288
rect 5917 7276 5930 7290
rect 5998 7286 6151 7290
rect 5880 7274 5902 7276
rect 5980 7274 6172 7286
rect 6251 7274 6264 7304
rect 6279 7290 6309 7304
rect 6346 7274 6365 7304
rect 6380 7274 6386 7304
rect 6395 7274 6408 7304
rect 6423 7290 6453 7304
rect 6496 7290 6539 7304
rect 6546 7290 6766 7304
rect 6773 7290 6803 7304
rect 6463 7276 6478 7288
rect 6497 7276 6510 7290
rect 6578 7286 6731 7290
rect 6460 7274 6482 7276
rect 6560 7274 6752 7286
rect 6831 7274 6844 7304
rect 6859 7290 6889 7304
rect 6926 7274 6945 7304
rect 6960 7274 6966 7304
rect 6975 7274 6988 7304
rect 7003 7290 7033 7304
rect 7076 7290 7119 7304
rect 7126 7290 7346 7304
rect 7353 7290 7383 7304
rect 7043 7276 7058 7288
rect 7077 7276 7090 7290
rect 7158 7286 7311 7290
rect 7040 7274 7062 7276
rect 7140 7274 7332 7286
rect 7411 7274 7424 7304
rect 7439 7290 7469 7304
rect 7506 7274 7525 7304
rect 7540 7274 7546 7304
rect 7555 7274 7568 7304
rect 7583 7290 7613 7304
rect 7656 7290 7699 7304
rect 7706 7290 7926 7304
rect 7933 7290 7963 7304
rect 7623 7276 7638 7288
rect 7657 7276 7670 7290
rect 7738 7286 7891 7290
rect 7620 7274 7642 7276
rect 7720 7274 7912 7286
rect 7991 7274 8004 7304
rect 8019 7290 8049 7304
rect 8086 7274 8105 7304
rect 8120 7274 8126 7304
rect 8135 7274 8148 7304
rect 8163 7290 8193 7304
rect 8236 7290 8279 7304
rect 8286 7290 8506 7304
rect 8513 7290 8543 7304
rect 8203 7276 8218 7288
rect 8237 7276 8250 7290
rect 8318 7286 8471 7290
rect 8200 7274 8222 7276
rect 8300 7274 8492 7286
rect 8571 7274 8584 7304
rect 8599 7290 8629 7304
rect 8666 7274 8685 7304
rect 8700 7274 8706 7304
rect 8715 7274 8728 7304
rect 8743 7290 8773 7304
rect 8816 7290 8859 7304
rect 8866 7290 9086 7304
rect 9093 7290 9123 7304
rect 8783 7276 8798 7288
rect 8817 7276 8830 7290
rect 8898 7286 9051 7290
rect 8780 7274 8802 7276
rect 8880 7274 9072 7286
rect 9151 7274 9164 7304
rect 9179 7290 9209 7304
rect 9246 7274 9265 7304
rect 9280 7274 9286 7304
rect 9295 7274 9308 7304
rect 9323 7290 9353 7304
rect 9396 7290 9439 7304
rect 9446 7290 9666 7304
rect 9673 7290 9703 7304
rect 9363 7276 9378 7288
rect 9397 7276 9410 7290
rect 9478 7286 9631 7290
rect 9360 7274 9382 7276
rect 9460 7274 9652 7286
rect 9731 7274 9744 7304
rect 9759 7290 9789 7304
rect 9826 7274 9845 7304
rect 9860 7274 9866 7304
rect 9875 7274 9888 7304
rect 9903 7290 9933 7304
rect 9976 7290 10019 7304
rect 10026 7290 10246 7304
rect 10253 7290 10283 7304
rect 9943 7276 9958 7288
rect 9977 7276 9990 7290
rect 10058 7286 10211 7290
rect 9940 7274 9962 7276
rect 10040 7274 10232 7286
rect 10311 7274 10324 7304
rect 10339 7290 10369 7304
rect 10406 7274 10425 7304
rect 10440 7274 10446 7304
rect 10455 7274 10468 7304
rect 10483 7290 10513 7304
rect 10556 7290 10599 7304
rect 10606 7290 10826 7304
rect 10833 7290 10863 7304
rect 10523 7276 10538 7288
rect 10557 7276 10570 7290
rect 10638 7286 10791 7290
rect 10520 7274 10542 7276
rect 10620 7274 10812 7286
rect 10891 7274 10904 7304
rect 10919 7290 10949 7304
rect 10986 7274 11005 7304
rect 11020 7274 11026 7304
rect 11035 7274 11048 7304
rect 11063 7290 11093 7304
rect 11136 7290 11179 7304
rect 11186 7290 11406 7304
rect 11413 7290 11443 7304
rect 11103 7276 11118 7288
rect 11137 7276 11150 7290
rect 11218 7286 11371 7290
rect 11100 7274 11122 7276
rect 11200 7274 11392 7286
rect 11471 7274 11484 7304
rect 11499 7290 11529 7304
rect 11566 7274 11585 7304
rect 11600 7274 11606 7304
rect 11615 7274 11628 7304
rect 11643 7290 11673 7304
rect 11716 7290 11759 7304
rect 11766 7290 11986 7304
rect 11993 7290 12023 7304
rect 11683 7276 11698 7288
rect 11717 7276 11730 7290
rect 11798 7286 11951 7290
rect 11680 7274 11702 7276
rect 11780 7274 11972 7286
rect 12051 7274 12064 7304
rect 12079 7290 12109 7304
rect 12146 7274 12165 7304
rect 12180 7274 12186 7304
rect 12195 7274 12208 7304
rect 12223 7290 12253 7304
rect 12296 7290 12339 7304
rect 12346 7290 12566 7304
rect 12573 7290 12603 7304
rect 12263 7276 12278 7288
rect 12297 7276 12310 7290
rect 12378 7286 12531 7290
rect 12260 7274 12282 7276
rect 12360 7274 12552 7286
rect 12631 7274 12644 7304
rect 12659 7290 12689 7304
rect 12726 7274 12745 7304
rect 12760 7274 12766 7304
rect 12775 7274 12788 7304
rect 12803 7290 12833 7304
rect 12876 7290 12919 7304
rect 12926 7290 13146 7304
rect 13153 7290 13183 7304
rect 12843 7276 12858 7288
rect 12877 7276 12890 7290
rect 12958 7286 13111 7290
rect 12840 7274 12862 7276
rect 12940 7274 13132 7286
rect 13211 7274 13224 7304
rect 13239 7290 13269 7304
rect 13306 7274 13325 7304
rect 13340 7274 13346 7304
rect 13355 7274 13368 7304
rect 13383 7290 13413 7304
rect 13456 7290 13499 7304
rect 13506 7290 13726 7304
rect 13733 7290 13763 7304
rect 13423 7276 13438 7288
rect 13457 7276 13470 7290
rect 13538 7286 13691 7290
rect 13420 7274 13442 7276
rect 13520 7274 13712 7286
rect 13791 7274 13804 7304
rect 13819 7290 13849 7304
rect 13886 7274 13905 7304
rect 13920 7274 13926 7304
rect 13935 7274 13948 7304
rect 13963 7290 13993 7304
rect 14036 7290 14079 7304
rect 14086 7290 14306 7304
rect 14313 7290 14343 7304
rect 14003 7276 14018 7288
rect 14037 7276 14050 7290
rect 14118 7286 14271 7290
rect 14000 7274 14022 7276
rect 14100 7274 14292 7286
rect 14371 7274 14384 7304
rect 14399 7290 14429 7304
rect 14466 7274 14485 7304
rect 14500 7274 14506 7304
rect 14515 7274 14528 7304
rect 14543 7290 14573 7304
rect 14616 7290 14659 7304
rect 14666 7290 14886 7304
rect 14893 7290 14923 7304
rect 14583 7276 14598 7288
rect 14617 7276 14630 7290
rect 14698 7286 14851 7290
rect 14580 7274 14602 7276
rect 14680 7274 14872 7286
rect 14951 7274 14964 7304
rect 14979 7290 15009 7304
rect 15046 7274 15065 7304
rect 15080 7274 15086 7304
rect 15095 7274 15108 7304
rect 15123 7290 15153 7304
rect 15196 7290 15239 7304
rect 15246 7290 15466 7304
rect 15473 7290 15503 7304
rect 15163 7276 15178 7288
rect 15197 7276 15210 7290
rect 15278 7286 15431 7290
rect 15160 7274 15182 7276
rect 15260 7274 15452 7286
rect 15531 7274 15544 7304
rect 15559 7290 15589 7304
rect 15626 7274 15645 7304
rect 15660 7274 15666 7304
rect 15675 7274 15688 7304
rect 15703 7290 15733 7304
rect 15776 7290 15819 7304
rect 15826 7290 16046 7304
rect 16053 7290 16083 7304
rect 15743 7276 15758 7288
rect 15777 7276 15790 7290
rect 15858 7286 16011 7290
rect 15740 7274 15762 7276
rect 15840 7274 16032 7286
rect 16111 7274 16124 7304
rect 16139 7290 16169 7304
rect 16206 7274 16225 7304
rect 16240 7274 16246 7304
rect 16255 7274 16268 7304
rect 16283 7290 16313 7304
rect 16356 7290 16399 7304
rect 16406 7290 16626 7304
rect 16633 7290 16663 7304
rect 16323 7276 16338 7288
rect 16357 7276 16370 7290
rect 16438 7286 16591 7290
rect 16320 7274 16342 7276
rect 16420 7274 16612 7286
rect 16691 7274 16704 7304
rect 16719 7290 16749 7304
rect 16786 7274 16805 7304
rect 16820 7274 16826 7304
rect 16835 7274 16848 7304
rect 16863 7290 16893 7304
rect 16936 7290 16979 7304
rect 16986 7290 17206 7304
rect 17213 7290 17243 7304
rect 16903 7276 16918 7288
rect 16937 7276 16950 7290
rect 17018 7286 17171 7290
rect 16900 7274 16922 7276
rect 17000 7274 17192 7286
rect 17271 7274 17284 7304
rect 17299 7290 17329 7304
rect 17366 7274 17385 7304
rect 17400 7274 17406 7304
rect 17415 7274 17428 7304
rect 17443 7290 17473 7304
rect 17516 7290 17559 7304
rect 17566 7290 17786 7304
rect 17793 7290 17823 7304
rect 17483 7276 17498 7288
rect 17517 7276 17530 7290
rect 17598 7286 17751 7290
rect 17480 7274 17502 7276
rect 17580 7274 17772 7286
rect 17851 7274 17864 7304
rect 17879 7290 17909 7304
rect 17946 7274 17965 7304
rect 17980 7274 17986 7304
rect 17995 7274 18008 7304
rect 18023 7290 18053 7304
rect 18096 7290 18139 7304
rect 18146 7290 18366 7304
rect 18373 7290 18403 7304
rect 18063 7276 18078 7288
rect 18097 7276 18110 7290
rect 18178 7286 18331 7290
rect 18060 7274 18082 7276
rect 18160 7274 18352 7286
rect 18431 7274 18444 7304
rect 18459 7290 18489 7304
rect 18532 7274 18545 7304
rect 0 7260 18545 7274
rect 15 7190 28 7260
rect 80 7256 102 7260
rect 73 7234 102 7248
rect 155 7234 171 7248
rect 209 7244 215 7246
rect 222 7244 330 7260
rect 337 7244 343 7246
rect 351 7244 366 7260
rect 432 7254 451 7257
rect 73 7232 171 7234
rect 198 7232 366 7244
rect 381 7234 397 7248
rect 432 7235 454 7254
rect 464 7248 480 7249
rect 463 7246 480 7248
rect 464 7241 480 7246
rect 454 7234 460 7235
rect 463 7234 492 7241
rect 381 7233 492 7234
rect 381 7232 498 7233
rect 57 7224 108 7232
rect 155 7224 189 7232
rect 57 7212 82 7224
rect 89 7212 108 7224
rect 162 7222 189 7224
rect 198 7222 419 7232
rect 454 7229 460 7232
rect 162 7218 419 7222
rect 57 7204 108 7212
rect 155 7204 419 7218
rect 463 7224 498 7232
rect 9 7156 28 7190
rect 73 7196 102 7204
rect 73 7190 90 7196
rect 73 7188 107 7190
rect 155 7188 171 7204
rect 172 7194 380 7204
rect 381 7194 397 7204
rect 445 7200 460 7215
rect 463 7212 464 7224
rect 471 7212 498 7224
rect 463 7204 498 7212
rect 463 7203 492 7204
rect 183 7190 397 7194
rect 198 7188 397 7190
rect 432 7190 445 7200
rect 463 7190 480 7203
rect 432 7188 480 7190
rect 74 7184 107 7188
rect 70 7182 107 7184
rect 70 7181 137 7182
rect 70 7176 101 7181
rect 107 7176 137 7181
rect 70 7172 137 7176
rect 43 7169 137 7172
rect 43 7162 92 7169
rect 43 7156 73 7162
rect 92 7157 97 7162
rect 9 7140 89 7156
rect 101 7148 137 7169
rect 198 7164 387 7188
rect 432 7187 479 7188
rect 445 7182 479 7187
rect 213 7161 387 7164
rect 206 7158 387 7161
rect 415 7181 479 7182
rect 9 7138 28 7140
rect 43 7138 77 7140
rect 9 7122 89 7138
rect 9 7116 28 7122
rect -1 7100 28 7116
rect 43 7106 73 7122
rect 101 7100 107 7148
rect 110 7142 129 7148
rect 144 7142 174 7150
rect 110 7134 174 7142
rect 110 7118 190 7134
rect 206 7127 268 7158
rect 284 7127 346 7158
rect 415 7156 464 7181
rect 479 7156 509 7172
rect 378 7142 408 7150
rect 415 7148 525 7156
rect 378 7134 423 7142
rect 110 7116 129 7118
rect 144 7116 190 7118
rect 110 7100 190 7116
rect 217 7114 252 7127
rect 293 7124 330 7127
rect 293 7122 335 7124
rect 222 7111 252 7114
rect 231 7107 238 7111
rect 238 7106 239 7107
rect 197 7100 207 7106
rect -7 7092 34 7100
rect -7 7066 8 7092
rect 15 7066 34 7092
rect 98 7088 129 7100
rect 144 7088 247 7100
rect 259 7090 285 7116
rect 300 7111 330 7122
rect 362 7118 424 7134
rect 362 7116 408 7118
rect 362 7100 424 7116
rect 436 7100 442 7148
rect 445 7140 525 7148
rect 445 7138 464 7140
rect 479 7138 513 7140
rect 445 7122 525 7138
rect 445 7100 464 7122
rect 479 7106 509 7122
rect 537 7116 543 7190
rect 546 7116 565 7260
rect 580 7116 586 7260
rect 595 7190 608 7260
rect 660 7256 682 7260
rect 653 7234 682 7248
rect 735 7234 751 7248
rect 789 7244 795 7246
rect 802 7244 910 7260
rect 917 7244 923 7246
rect 931 7244 946 7260
rect 1012 7254 1031 7257
rect 653 7232 751 7234
rect 778 7232 946 7244
rect 961 7234 977 7248
rect 1012 7235 1034 7254
rect 1044 7248 1060 7249
rect 1043 7246 1060 7248
rect 1044 7241 1060 7246
rect 1034 7234 1040 7235
rect 1043 7234 1072 7241
rect 961 7233 1072 7234
rect 961 7232 1078 7233
rect 637 7224 688 7232
rect 735 7224 769 7232
rect 637 7212 662 7224
rect 669 7212 688 7224
rect 742 7222 769 7224
rect 778 7222 999 7232
rect 1034 7229 1040 7232
rect 742 7218 999 7222
rect 637 7204 688 7212
rect 735 7204 999 7218
rect 1043 7224 1078 7232
rect 589 7156 608 7190
rect 653 7196 682 7204
rect 653 7190 670 7196
rect 653 7188 687 7190
rect 735 7188 751 7204
rect 752 7194 960 7204
rect 961 7194 977 7204
rect 1025 7200 1040 7215
rect 1043 7212 1044 7224
rect 1051 7212 1078 7224
rect 1043 7204 1078 7212
rect 1043 7203 1072 7204
rect 763 7190 977 7194
rect 778 7188 977 7190
rect 1012 7190 1025 7200
rect 1043 7190 1060 7203
rect 1012 7188 1060 7190
rect 654 7184 687 7188
rect 650 7182 687 7184
rect 650 7181 717 7182
rect 650 7176 681 7181
rect 687 7176 717 7181
rect 650 7172 717 7176
rect 623 7169 717 7172
rect 623 7162 672 7169
rect 623 7156 653 7162
rect 672 7157 677 7162
rect 589 7140 669 7156
rect 681 7148 717 7169
rect 778 7164 967 7188
rect 1012 7187 1059 7188
rect 1025 7182 1059 7187
rect 793 7161 967 7164
rect 786 7158 967 7161
rect 995 7181 1059 7182
rect 589 7138 608 7140
rect 623 7138 657 7140
rect 589 7122 669 7138
rect 589 7116 608 7122
rect 305 7090 408 7100
rect 259 7088 408 7090
rect 429 7088 464 7100
rect 98 7086 260 7088
rect 110 7066 129 7086
rect 144 7084 174 7086
rect -7 7058 34 7066
rect 116 7062 129 7066
rect 181 7070 260 7086
rect 292 7086 464 7088
rect 292 7070 371 7086
rect 378 7084 408 7086
rect -1 7048 28 7058
rect 43 7048 73 7062
rect 116 7048 159 7062
rect 181 7058 371 7070
rect 436 7066 442 7086
rect 166 7048 196 7058
rect 197 7048 355 7058
rect 359 7048 389 7058
rect 393 7048 423 7062
rect 451 7048 464 7086
rect 536 7100 565 7116
rect 579 7100 608 7116
rect 623 7106 653 7122
rect 681 7100 687 7148
rect 690 7142 709 7148
rect 724 7142 754 7150
rect 690 7134 754 7142
rect 690 7118 770 7134
rect 786 7127 848 7158
rect 864 7127 926 7158
rect 995 7156 1044 7181
rect 1059 7156 1089 7172
rect 958 7142 988 7150
rect 995 7148 1105 7156
rect 958 7134 1003 7142
rect 690 7116 709 7118
rect 724 7116 770 7118
rect 690 7100 770 7116
rect 797 7114 832 7127
rect 873 7124 910 7127
rect 873 7122 915 7124
rect 802 7111 832 7114
rect 811 7107 818 7111
rect 818 7106 819 7107
rect 777 7100 787 7106
rect 536 7092 571 7100
rect 536 7066 537 7092
rect 544 7066 571 7092
rect 479 7048 509 7062
rect 536 7058 571 7066
rect 573 7092 614 7100
rect 573 7066 588 7092
rect 595 7066 614 7092
rect 678 7088 709 7100
rect 724 7088 827 7100
rect 839 7090 865 7116
rect 880 7111 910 7122
rect 942 7118 1004 7134
rect 942 7116 988 7118
rect 942 7100 1004 7116
rect 1016 7100 1022 7148
rect 1025 7140 1105 7148
rect 1025 7138 1044 7140
rect 1059 7138 1093 7140
rect 1025 7122 1105 7138
rect 1025 7100 1044 7122
rect 1059 7106 1089 7122
rect 1117 7116 1123 7190
rect 1126 7116 1145 7260
rect 1160 7116 1166 7260
rect 1175 7190 1188 7260
rect 1240 7256 1262 7260
rect 1233 7234 1262 7248
rect 1315 7234 1331 7248
rect 1369 7244 1375 7246
rect 1382 7244 1490 7260
rect 1497 7244 1503 7246
rect 1511 7244 1526 7260
rect 1592 7254 1611 7257
rect 1233 7232 1331 7234
rect 1358 7232 1526 7244
rect 1541 7234 1557 7248
rect 1592 7235 1614 7254
rect 1624 7248 1640 7249
rect 1623 7246 1640 7248
rect 1624 7241 1640 7246
rect 1614 7234 1620 7235
rect 1623 7234 1652 7241
rect 1541 7233 1652 7234
rect 1541 7232 1658 7233
rect 1217 7224 1268 7232
rect 1315 7224 1349 7232
rect 1217 7212 1242 7224
rect 1249 7212 1268 7224
rect 1322 7222 1349 7224
rect 1358 7222 1579 7232
rect 1614 7229 1620 7232
rect 1322 7218 1579 7222
rect 1217 7204 1268 7212
rect 1315 7204 1579 7218
rect 1623 7224 1658 7232
rect 1169 7156 1188 7190
rect 1233 7196 1262 7204
rect 1233 7190 1250 7196
rect 1233 7188 1267 7190
rect 1315 7188 1331 7204
rect 1332 7194 1540 7204
rect 1541 7194 1557 7204
rect 1605 7200 1620 7215
rect 1623 7212 1624 7224
rect 1631 7212 1658 7224
rect 1623 7204 1658 7212
rect 1623 7203 1652 7204
rect 1343 7190 1557 7194
rect 1358 7188 1557 7190
rect 1592 7190 1605 7200
rect 1623 7190 1640 7203
rect 1592 7188 1640 7190
rect 1234 7184 1267 7188
rect 1230 7182 1267 7184
rect 1230 7181 1297 7182
rect 1230 7176 1261 7181
rect 1267 7176 1297 7181
rect 1230 7172 1297 7176
rect 1203 7169 1297 7172
rect 1203 7162 1252 7169
rect 1203 7156 1233 7162
rect 1252 7157 1257 7162
rect 1169 7140 1249 7156
rect 1261 7148 1297 7169
rect 1358 7164 1547 7188
rect 1592 7187 1639 7188
rect 1605 7182 1639 7187
rect 1373 7161 1547 7164
rect 1366 7158 1547 7161
rect 1575 7181 1639 7182
rect 1169 7138 1188 7140
rect 1203 7138 1237 7140
rect 1169 7122 1249 7138
rect 1169 7116 1188 7122
rect 885 7090 988 7100
rect 839 7088 988 7090
rect 1009 7088 1044 7100
rect 678 7086 840 7088
rect 690 7066 709 7086
rect 724 7084 754 7086
rect 573 7058 614 7066
rect 696 7062 709 7066
rect 761 7070 840 7086
rect 872 7086 1044 7088
rect 872 7070 951 7086
rect 958 7084 988 7086
rect 536 7048 565 7058
rect 579 7048 608 7058
rect 623 7048 653 7062
rect 696 7048 739 7062
rect 761 7058 951 7070
rect 1016 7066 1022 7086
rect 746 7048 776 7058
rect 777 7048 935 7058
rect 939 7048 969 7058
rect 973 7048 1003 7062
rect 1031 7048 1044 7086
rect 1116 7100 1145 7116
rect 1159 7100 1188 7116
rect 1203 7106 1233 7122
rect 1261 7100 1267 7148
rect 1270 7142 1289 7148
rect 1304 7142 1334 7150
rect 1270 7134 1334 7142
rect 1270 7118 1350 7134
rect 1366 7127 1428 7158
rect 1444 7127 1506 7158
rect 1575 7156 1624 7181
rect 1639 7156 1669 7172
rect 1538 7142 1568 7150
rect 1575 7148 1685 7156
rect 1538 7134 1583 7142
rect 1270 7116 1289 7118
rect 1304 7116 1350 7118
rect 1270 7100 1350 7116
rect 1377 7114 1412 7127
rect 1453 7124 1490 7127
rect 1453 7122 1495 7124
rect 1382 7111 1412 7114
rect 1391 7107 1398 7111
rect 1398 7106 1399 7107
rect 1357 7100 1367 7106
rect 1116 7092 1151 7100
rect 1116 7066 1117 7092
rect 1124 7066 1151 7092
rect 1059 7048 1089 7062
rect 1116 7058 1151 7066
rect 1153 7092 1194 7100
rect 1153 7066 1168 7092
rect 1175 7066 1194 7092
rect 1258 7088 1289 7100
rect 1304 7088 1407 7100
rect 1419 7090 1445 7116
rect 1460 7111 1490 7122
rect 1522 7118 1584 7134
rect 1522 7116 1568 7118
rect 1522 7100 1584 7116
rect 1596 7100 1602 7148
rect 1605 7140 1685 7148
rect 1605 7138 1624 7140
rect 1639 7138 1673 7140
rect 1605 7122 1685 7138
rect 1605 7100 1624 7122
rect 1639 7106 1669 7122
rect 1697 7116 1703 7190
rect 1706 7116 1725 7260
rect 1740 7116 1746 7260
rect 1755 7190 1768 7260
rect 1820 7256 1842 7260
rect 1813 7234 1842 7248
rect 1895 7234 1911 7248
rect 1949 7244 1955 7246
rect 1962 7244 2070 7260
rect 2077 7244 2083 7246
rect 2091 7244 2106 7260
rect 2172 7254 2191 7257
rect 1813 7232 1911 7234
rect 1938 7232 2106 7244
rect 2121 7234 2137 7248
rect 2172 7235 2194 7254
rect 2204 7248 2220 7249
rect 2203 7246 2220 7248
rect 2204 7241 2220 7246
rect 2194 7234 2200 7235
rect 2203 7234 2232 7241
rect 2121 7233 2232 7234
rect 2121 7232 2238 7233
rect 1797 7224 1848 7232
rect 1895 7224 1929 7232
rect 1797 7212 1822 7224
rect 1829 7212 1848 7224
rect 1902 7222 1929 7224
rect 1938 7222 2159 7232
rect 2194 7229 2200 7232
rect 1902 7218 2159 7222
rect 1797 7204 1848 7212
rect 1895 7204 2159 7218
rect 2203 7224 2238 7232
rect 1749 7156 1768 7190
rect 1813 7196 1842 7204
rect 1813 7190 1830 7196
rect 1813 7188 1847 7190
rect 1895 7188 1911 7204
rect 1912 7194 2120 7204
rect 2121 7194 2137 7204
rect 2185 7200 2200 7215
rect 2203 7212 2204 7224
rect 2211 7212 2238 7224
rect 2203 7204 2238 7212
rect 2203 7203 2232 7204
rect 1923 7190 2137 7194
rect 1938 7188 2137 7190
rect 2172 7190 2185 7200
rect 2203 7190 2220 7203
rect 2172 7188 2220 7190
rect 1814 7184 1847 7188
rect 1810 7182 1847 7184
rect 1810 7181 1877 7182
rect 1810 7176 1841 7181
rect 1847 7176 1877 7181
rect 1810 7172 1877 7176
rect 1783 7169 1877 7172
rect 1783 7162 1832 7169
rect 1783 7156 1813 7162
rect 1832 7157 1837 7162
rect 1749 7140 1829 7156
rect 1841 7148 1877 7169
rect 1938 7164 2127 7188
rect 2172 7187 2219 7188
rect 2185 7182 2219 7187
rect 1953 7161 2127 7164
rect 1946 7158 2127 7161
rect 2155 7181 2219 7182
rect 1749 7138 1768 7140
rect 1783 7138 1817 7140
rect 1749 7122 1829 7138
rect 1749 7116 1768 7122
rect 1465 7090 1568 7100
rect 1419 7088 1568 7090
rect 1589 7088 1624 7100
rect 1258 7086 1420 7088
rect 1270 7066 1289 7086
rect 1304 7084 1334 7086
rect 1153 7058 1194 7066
rect 1276 7062 1289 7066
rect 1341 7070 1420 7086
rect 1452 7086 1624 7088
rect 1452 7070 1531 7086
rect 1538 7084 1568 7086
rect 1116 7048 1145 7058
rect 1159 7048 1188 7058
rect 1203 7048 1233 7062
rect 1276 7048 1319 7062
rect 1341 7058 1531 7070
rect 1596 7066 1602 7086
rect 1326 7048 1356 7058
rect 1357 7048 1515 7058
rect 1519 7048 1549 7058
rect 1553 7048 1583 7062
rect 1611 7048 1624 7086
rect 1696 7100 1725 7116
rect 1739 7100 1768 7116
rect 1783 7106 1813 7122
rect 1841 7100 1847 7148
rect 1850 7142 1869 7148
rect 1884 7142 1914 7150
rect 1850 7134 1914 7142
rect 1850 7118 1930 7134
rect 1946 7127 2008 7158
rect 2024 7127 2086 7158
rect 2155 7156 2204 7181
rect 2219 7156 2249 7172
rect 2118 7142 2148 7150
rect 2155 7148 2265 7156
rect 2118 7134 2163 7142
rect 1850 7116 1869 7118
rect 1884 7116 1930 7118
rect 1850 7100 1930 7116
rect 1957 7114 1992 7127
rect 2033 7124 2070 7127
rect 2033 7122 2075 7124
rect 1962 7111 1992 7114
rect 1971 7107 1978 7111
rect 1978 7106 1979 7107
rect 1937 7100 1947 7106
rect 1696 7092 1731 7100
rect 1696 7066 1697 7092
rect 1704 7066 1731 7092
rect 1639 7048 1669 7062
rect 1696 7058 1731 7066
rect 1733 7092 1774 7100
rect 1733 7066 1748 7092
rect 1755 7066 1774 7092
rect 1838 7088 1869 7100
rect 1884 7088 1987 7100
rect 1999 7090 2025 7116
rect 2040 7111 2070 7122
rect 2102 7118 2164 7134
rect 2102 7116 2148 7118
rect 2102 7100 2164 7116
rect 2176 7100 2182 7148
rect 2185 7140 2265 7148
rect 2185 7138 2204 7140
rect 2219 7138 2253 7140
rect 2185 7122 2265 7138
rect 2185 7100 2204 7122
rect 2219 7106 2249 7122
rect 2277 7116 2283 7190
rect 2286 7116 2305 7260
rect 2320 7116 2326 7260
rect 2335 7190 2348 7260
rect 2400 7256 2422 7260
rect 2393 7234 2422 7248
rect 2475 7234 2491 7248
rect 2529 7244 2535 7246
rect 2542 7244 2650 7260
rect 2657 7244 2663 7246
rect 2671 7244 2686 7260
rect 2752 7254 2771 7257
rect 2393 7232 2491 7234
rect 2518 7232 2686 7244
rect 2701 7234 2717 7248
rect 2752 7235 2774 7254
rect 2784 7248 2800 7249
rect 2783 7246 2800 7248
rect 2784 7241 2800 7246
rect 2774 7234 2780 7235
rect 2783 7234 2812 7241
rect 2701 7233 2812 7234
rect 2701 7232 2818 7233
rect 2377 7224 2428 7232
rect 2475 7224 2509 7232
rect 2377 7212 2402 7224
rect 2409 7212 2428 7224
rect 2482 7222 2509 7224
rect 2518 7222 2739 7232
rect 2774 7229 2780 7232
rect 2482 7218 2739 7222
rect 2377 7204 2428 7212
rect 2475 7204 2739 7218
rect 2783 7224 2818 7232
rect 2329 7156 2348 7190
rect 2393 7196 2422 7204
rect 2393 7190 2410 7196
rect 2393 7188 2427 7190
rect 2475 7188 2491 7204
rect 2492 7194 2700 7204
rect 2701 7194 2717 7204
rect 2765 7200 2780 7215
rect 2783 7212 2784 7224
rect 2791 7212 2818 7224
rect 2783 7204 2818 7212
rect 2783 7203 2812 7204
rect 2503 7190 2717 7194
rect 2518 7188 2717 7190
rect 2752 7190 2765 7200
rect 2783 7190 2800 7203
rect 2752 7188 2800 7190
rect 2394 7184 2427 7188
rect 2390 7182 2427 7184
rect 2390 7181 2457 7182
rect 2390 7176 2421 7181
rect 2427 7176 2457 7181
rect 2390 7172 2457 7176
rect 2363 7169 2457 7172
rect 2363 7162 2412 7169
rect 2363 7156 2393 7162
rect 2412 7157 2417 7162
rect 2329 7140 2409 7156
rect 2421 7148 2457 7169
rect 2518 7164 2707 7188
rect 2752 7187 2799 7188
rect 2765 7182 2799 7187
rect 2533 7161 2707 7164
rect 2526 7158 2707 7161
rect 2735 7181 2799 7182
rect 2329 7138 2348 7140
rect 2363 7138 2397 7140
rect 2329 7122 2409 7138
rect 2329 7116 2348 7122
rect 2045 7090 2148 7100
rect 1999 7088 2148 7090
rect 2169 7088 2204 7100
rect 1838 7086 2000 7088
rect 1850 7066 1869 7086
rect 1884 7084 1914 7086
rect 1733 7058 1774 7066
rect 1856 7062 1869 7066
rect 1921 7070 2000 7086
rect 2032 7086 2204 7088
rect 2032 7070 2111 7086
rect 2118 7084 2148 7086
rect 1696 7048 1725 7058
rect 1739 7048 1768 7058
rect 1783 7048 1813 7062
rect 1856 7048 1899 7062
rect 1921 7058 2111 7070
rect 2176 7066 2182 7086
rect 1906 7048 1936 7058
rect 1937 7048 2095 7058
rect 2099 7048 2129 7058
rect 2133 7048 2163 7062
rect 2191 7048 2204 7086
rect 2276 7100 2305 7116
rect 2319 7100 2348 7116
rect 2363 7106 2393 7122
rect 2421 7100 2427 7148
rect 2430 7142 2449 7148
rect 2464 7142 2494 7150
rect 2430 7134 2494 7142
rect 2430 7118 2510 7134
rect 2526 7127 2588 7158
rect 2604 7127 2666 7158
rect 2735 7156 2784 7181
rect 2799 7156 2829 7172
rect 2698 7142 2728 7150
rect 2735 7148 2845 7156
rect 2698 7134 2743 7142
rect 2430 7116 2449 7118
rect 2464 7116 2510 7118
rect 2430 7100 2510 7116
rect 2537 7114 2572 7127
rect 2613 7124 2650 7127
rect 2613 7122 2655 7124
rect 2542 7111 2572 7114
rect 2551 7107 2558 7111
rect 2558 7106 2559 7107
rect 2517 7100 2527 7106
rect 2276 7092 2311 7100
rect 2276 7066 2277 7092
rect 2284 7066 2311 7092
rect 2219 7048 2249 7062
rect 2276 7058 2311 7066
rect 2313 7092 2354 7100
rect 2313 7066 2328 7092
rect 2335 7066 2354 7092
rect 2418 7088 2449 7100
rect 2464 7088 2567 7100
rect 2579 7090 2605 7116
rect 2620 7111 2650 7122
rect 2682 7118 2744 7134
rect 2682 7116 2728 7118
rect 2682 7100 2744 7116
rect 2756 7100 2762 7148
rect 2765 7140 2845 7148
rect 2765 7138 2784 7140
rect 2799 7138 2833 7140
rect 2765 7122 2845 7138
rect 2765 7100 2784 7122
rect 2799 7106 2829 7122
rect 2857 7116 2863 7190
rect 2866 7116 2885 7260
rect 2900 7116 2906 7260
rect 2915 7190 2928 7260
rect 2980 7256 3002 7260
rect 2973 7234 3002 7248
rect 3055 7234 3071 7248
rect 3109 7244 3115 7246
rect 3122 7244 3230 7260
rect 3237 7244 3243 7246
rect 3251 7244 3266 7260
rect 3332 7254 3351 7257
rect 2973 7232 3071 7234
rect 3098 7232 3266 7244
rect 3281 7234 3297 7248
rect 3332 7235 3354 7254
rect 3364 7248 3380 7249
rect 3363 7246 3380 7248
rect 3364 7241 3380 7246
rect 3354 7234 3360 7235
rect 3363 7234 3392 7241
rect 3281 7233 3392 7234
rect 3281 7232 3398 7233
rect 2957 7224 3008 7232
rect 3055 7224 3089 7232
rect 2957 7212 2982 7224
rect 2989 7212 3008 7224
rect 3062 7222 3089 7224
rect 3098 7222 3319 7232
rect 3354 7229 3360 7232
rect 3062 7218 3319 7222
rect 2957 7204 3008 7212
rect 3055 7204 3319 7218
rect 3363 7224 3398 7232
rect 2909 7156 2928 7190
rect 2973 7196 3002 7204
rect 2973 7190 2990 7196
rect 2973 7188 3007 7190
rect 3055 7188 3071 7204
rect 3072 7194 3280 7204
rect 3281 7194 3297 7204
rect 3345 7200 3360 7215
rect 3363 7212 3364 7224
rect 3371 7212 3398 7224
rect 3363 7204 3398 7212
rect 3363 7203 3392 7204
rect 3083 7190 3297 7194
rect 3098 7188 3297 7190
rect 3332 7190 3345 7200
rect 3363 7190 3380 7203
rect 3332 7188 3380 7190
rect 2974 7184 3007 7188
rect 2970 7182 3007 7184
rect 2970 7181 3037 7182
rect 2970 7176 3001 7181
rect 3007 7176 3037 7181
rect 2970 7172 3037 7176
rect 2943 7169 3037 7172
rect 2943 7162 2992 7169
rect 2943 7156 2973 7162
rect 2992 7157 2997 7162
rect 2909 7140 2989 7156
rect 3001 7148 3037 7169
rect 3098 7164 3287 7188
rect 3332 7187 3379 7188
rect 3345 7182 3379 7187
rect 3113 7161 3287 7164
rect 3106 7158 3287 7161
rect 3315 7181 3379 7182
rect 2909 7138 2928 7140
rect 2943 7138 2977 7140
rect 2909 7122 2989 7138
rect 2909 7116 2928 7122
rect 2625 7090 2728 7100
rect 2579 7088 2728 7090
rect 2749 7088 2784 7100
rect 2418 7086 2580 7088
rect 2430 7066 2449 7086
rect 2464 7084 2494 7086
rect 2313 7058 2354 7066
rect 2436 7062 2449 7066
rect 2501 7070 2580 7086
rect 2612 7086 2784 7088
rect 2612 7070 2691 7086
rect 2698 7084 2728 7086
rect 2276 7048 2305 7058
rect 2319 7048 2348 7058
rect 2363 7048 2393 7062
rect 2436 7048 2479 7062
rect 2501 7058 2691 7070
rect 2756 7066 2762 7086
rect 2486 7048 2516 7058
rect 2517 7048 2675 7058
rect 2679 7048 2709 7058
rect 2713 7048 2743 7062
rect 2771 7048 2784 7086
rect 2856 7100 2885 7116
rect 2899 7100 2928 7116
rect 2943 7106 2973 7122
rect 3001 7100 3007 7148
rect 3010 7142 3029 7148
rect 3044 7142 3074 7150
rect 3010 7134 3074 7142
rect 3010 7118 3090 7134
rect 3106 7127 3168 7158
rect 3184 7127 3246 7158
rect 3315 7156 3364 7181
rect 3379 7156 3409 7172
rect 3278 7142 3308 7150
rect 3315 7148 3425 7156
rect 3278 7134 3323 7142
rect 3010 7116 3029 7118
rect 3044 7116 3090 7118
rect 3010 7100 3090 7116
rect 3117 7114 3152 7127
rect 3193 7124 3230 7127
rect 3193 7122 3235 7124
rect 3122 7111 3152 7114
rect 3131 7107 3138 7111
rect 3138 7106 3139 7107
rect 3097 7100 3107 7106
rect 2856 7092 2891 7100
rect 2856 7066 2857 7092
rect 2864 7066 2891 7092
rect 2799 7048 2829 7062
rect 2856 7058 2891 7066
rect 2893 7092 2934 7100
rect 2893 7066 2908 7092
rect 2915 7066 2934 7092
rect 2998 7088 3029 7100
rect 3044 7088 3147 7100
rect 3159 7090 3185 7116
rect 3200 7111 3230 7122
rect 3262 7118 3324 7134
rect 3262 7116 3308 7118
rect 3262 7100 3324 7116
rect 3336 7100 3342 7148
rect 3345 7140 3425 7148
rect 3345 7138 3364 7140
rect 3379 7138 3413 7140
rect 3345 7122 3425 7138
rect 3345 7100 3364 7122
rect 3379 7106 3409 7122
rect 3437 7116 3443 7190
rect 3446 7116 3465 7260
rect 3480 7116 3486 7260
rect 3495 7190 3508 7260
rect 3560 7256 3582 7260
rect 3553 7234 3582 7248
rect 3635 7234 3651 7248
rect 3689 7244 3695 7246
rect 3702 7244 3810 7260
rect 3817 7244 3823 7246
rect 3831 7244 3846 7260
rect 3912 7254 3931 7257
rect 3553 7232 3651 7234
rect 3678 7232 3846 7244
rect 3861 7234 3877 7248
rect 3912 7235 3934 7254
rect 3944 7248 3960 7249
rect 3943 7246 3960 7248
rect 3944 7241 3960 7246
rect 3934 7234 3940 7235
rect 3943 7234 3972 7241
rect 3861 7233 3972 7234
rect 3861 7232 3978 7233
rect 3537 7224 3588 7232
rect 3635 7224 3669 7232
rect 3537 7212 3562 7224
rect 3569 7212 3588 7224
rect 3642 7222 3669 7224
rect 3678 7222 3899 7232
rect 3934 7229 3940 7232
rect 3642 7218 3899 7222
rect 3537 7204 3588 7212
rect 3635 7204 3899 7218
rect 3943 7224 3978 7232
rect 3489 7156 3508 7190
rect 3553 7196 3582 7204
rect 3553 7190 3570 7196
rect 3553 7188 3587 7190
rect 3635 7188 3651 7204
rect 3652 7194 3860 7204
rect 3861 7194 3877 7204
rect 3925 7200 3940 7215
rect 3943 7212 3944 7224
rect 3951 7212 3978 7224
rect 3943 7204 3978 7212
rect 3943 7203 3972 7204
rect 3663 7190 3877 7194
rect 3678 7188 3877 7190
rect 3912 7190 3925 7200
rect 3943 7190 3960 7203
rect 3912 7188 3960 7190
rect 3554 7184 3587 7188
rect 3550 7182 3587 7184
rect 3550 7181 3617 7182
rect 3550 7176 3581 7181
rect 3587 7176 3617 7181
rect 3550 7172 3617 7176
rect 3523 7169 3617 7172
rect 3523 7162 3572 7169
rect 3523 7156 3553 7162
rect 3572 7157 3577 7162
rect 3489 7140 3569 7156
rect 3581 7148 3617 7169
rect 3678 7164 3867 7188
rect 3912 7187 3959 7188
rect 3925 7182 3959 7187
rect 3693 7161 3867 7164
rect 3686 7158 3867 7161
rect 3895 7181 3959 7182
rect 3489 7138 3508 7140
rect 3523 7138 3557 7140
rect 3489 7122 3569 7138
rect 3489 7116 3508 7122
rect 3205 7090 3308 7100
rect 3159 7088 3308 7090
rect 3329 7088 3364 7100
rect 2998 7086 3160 7088
rect 3010 7066 3029 7086
rect 3044 7084 3074 7086
rect 2893 7058 2934 7066
rect 3016 7062 3029 7066
rect 3081 7070 3160 7086
rect 3192 7086 3364 7088
rect 3192 7070 3271 7086
rect 3278 7084 3308 7086
rect 2856 7048 2885 7058
rect 2899 7048 2928 7058
rect 2943 7048 2973 7062
rect 3016 7048 3059 7062
rect 3081 7058 3271 7070
rect 3336 7066 3342 7086
rect 3066 7048 3096 7058
rect 3097 7048 3255 7058
rect 3259 7048 3289 7058
rect 3293 7048 3323 7062
rect 3351 7048 3364 7086
rect 3436 7100 3465 7116
rect 3479 7100 3508 7116
rect 3523 7106 3553 7122
rect 3581 7100 3587 7148
rect 3590 7142 3609 7148
rect 3624 7142 3654 7150
rect 3590 7134 3654 7142
rect 3590 7118 3670 7134
rect 3686 7127 3748 7158
rect 3764 7127 3826 7158
rect 3895 7156 3944 7181
rect 3959 7156 3989 7172
rect 3858 7142 3888 7150
rect 3895 7148 4005 7156
rect 3858 7134 3903 7142
rect 3590 7116 3609 7118
rect 3624 7116 3670 7118
rect 3590 7100 3670 7116
rect 3697 7114 3732 7127
rect 3773 7124 3810 7127
rect 3773 7122 3815 7124
rect 3702 7111 3732 7114
rect 3711 7107 3718 7111
rect 3718 7106 3719 7107
rect 3677 7100 3687 7106
rect 3436 7092 3471 7100
rect 3436 7066 3437 7092
rect 3444 7066 3471 7092
rect 3379 7048 3409 7062
rect 3436 7058 3471 7066
rect 3473 7092 3514 7100
rect 3473 7066 3488 7092
rect 3495 7066 3514 7092
rect 3578 7088 3609 7100
rect 3624 7088 3727 7100
rect 3739 7090 3765 7116
rect 3780 7111 3810 7122
rect 3842 7118 3904 7134
rect 3842 7116 3888 7118
rect 3842 7100 3904 7116
rect 3916 7100 3922 7148
rect 3925 7140 4005 7148
rect 3925 7138 3944 7140
rect 3959 7138 3993 7140
rect 3925 7122 4005 7138
rect 3925 7100 3944 7122
rect 3959 7106 3989 7122
rect 4017 7116 4023 7190
rect 4026 7116 4045 7260
rect 4060 7116 4066 7260
rect 4075 7190 4088 7260
rect 4140 7256 4162 7260
rect 4133 7234 4162 7248
rect 4215 7234 4231 7248
rect 4269 7244 4275 7246
rect 4282 7244 4390 7260
rect 4397 7244 4403 7246
rect 4411 7244 4426 7260
rect 4492 7254 4511 7257
rect 4133 7232 4231 7234
rect 4258 7232 4426 7244
rect 4441 7234 4457 7248
rect 4492 7235 4514 7254
rect 4524 7248 4540 7249
rect 4523 7246 4540 7248
rect 4524 7241 4540 7246
rect 4514 7234 4520 7235
rect 4523 7234 4552 7241
rect 4441 7233 4552 7234
rect 4441 7232 4558 7233
rect 4117 7224 4168 7232
rect 4215 7224 4249 7232
rect 4117 7212 4142 7224
rect 4149 7212 4168 7224
rect 4222 7222 4249 7224
rect 4258 7222 4479 7232
rect 4514 7229 4520 7232
rect 4222 7218 4479 7222
rect 4117 7204 4168 7212
rect 4215 7204 4479 7218
rect 4523 7224 4558 7232
rect 4069 7156 4088 7190
rect 4133 7196 4162 7204
rect 4133 7190 4150 7196
rect 4133 7188 4167 7190
rect 4215 7188 4231 7204
rect 4232 7194 4440 7204
rect 4441 7194 4457 7204
rect 4505 7200 4520 7215
rect 4523 7212 4524 7224
rect 4531 7212 4558 7224
rect 4523 7204 4558 7212
rect 4523 7203 4552 7204
rect 4243 7190 4457 7194
rect 4258 7188 4457 7190
rect 4492 7190 4505 7200
rect 4523 7190 4540 7203
rect 4492 7188 4540 7190
rect 4134 7184 4167 7188
rect 4130 7182 4167 7184
rect 4130 7181 4197 7182
rect 4130 7176 4161 7181
rect 4167 7176 4197 7181
rect 4130 7172 4197 7176
rect 4103 7169 4197 7172
rect 4103 7162 4152 7169
rect 4103 7156 4133 7162
rect 4152 7157 4157 7162
rect 4069 7140 4149 7156
rect 4161 7148 4197 7169
rect 4258 7164 4447 7188
rect 4492 7187 4539 7188
rect 4505 7182 4539 7187
rect 4273 7161 4447 7164
rect 4266 7158 4447 7161
rect 4475 7181 4539 7182
rect 4069 7138 4088 7140
rect 4103 7138 4137 7140
rect 4069 7122 4149 7138
rect 4069 7116 4088 7122
rect 3785 7090 3888 7100
rect 3739 7088 3888 7090
rect 3909 7088 3944 7100
rect 3578 7086 3740 7088
rect 3590 7066 3609 7086
rect 3624 7084 3654 7086
rect 3473 7058 3514 7066
rect 3596 7062 3609 7066
rect 3661 7070 3740 7086
rect 3772 7086 3944 7088
rect 3772 7070 3851 7086
rect 3858 7084 3888 7086
rect 3436 7048 3465 7058
rect 3479 7048 3508 7058
rect 3523 7048 3553 7062
rect 3596 7048 3639 7062
rect 3661 7058 3851 7070
rect 3916 7066 3922 7086
rect 3646 7048 3676 7058
rect 3677 7048 3835 7058
rect 3839 7048 3869 7058
rect 3873 7048 3903 7062
rect 3931 7048 3944 7086
rect 4016 7100 4045 7116
rect 4059 7100 4088 7116
rect 4103 7106 4133 7122
rect 4161 7100 4167 7148
rect 4170 7142 4189 7148
rect 4204 7142 4234 7150
rect 4170 7134 4234 7142
rect 4170 7118 4250 7134
rect 4266 7127 4328 7158
rect 4344 7127 4406 7158
rect 4475 7156 4524 7181
rect 4539 7156 4569 7172
rect 4438 7142 4468 7150
rect 4475 7148 4585 7156
rect 4438 7134 4483 7142
rect 4170 7116 4189 7118
rect 4204 7116 4250 7118
rect 4170 7100 4250 7116
rect 4277 7114 4312 7127
rect 4353 7124 4390 7127
rect 4353 7122 4395 7124
rect 4282 7111 4312 7114
rect 4291 7107 4298 7111
rect 4298 7106 4299 7107
rect 4257 7100 4267 7106
rect 4016 7092 4051 7100
rect 4016 7066 4017 7092
rect 4024 7066 4051 7092
rect 3959 7048 3989 7062
rect 4016 7058 4051 7066
rect 4053 7092 4094 7100
rect 4053 7066 4068 7092
rect 4075 7066 4094 7092
rect 4158 7088 4189 7100
rect 4204 7088 4307 7100
rect 4319 7090 4345 7116
rect 4360 7111 4390 7122
rect 4422 7118 4484 7134
rect 4422 7116 4468 7118
rect 4422 7100 4484 7116
rect 4496 7100 4502 7148
rect 4505 7140 4585 7148
rect 4505 7138 4524 7140
rect 4539 7138 4573 7140
rect 4505 7122 4585 7138
rect 4505 7100 4524 7122
rect 4539 7106 4569 7122
rect 4597 7116 4603 7190
rect 4606 7116 4625 7260
rect 4640 7116 4646 7260
rect 4655 7190 4668 7260
rect 4720 7256 4742 7260
rect 4713 7234 4742 7248
rect 4795 7234 4811 7248
rect 4849 7244 4855 7246
rect 4862 7244 4970 7260
rect 4977 7244 4983 7246
rect 4991 7244 5006 7260
rect 5072 7254 5091 7257
rect 4713 7232 4811 7234
rect 4838 7232 5006 7244
rect 5021 7234 5037 7248
rect 5072 7235 5094 7254
rect 5104 7248 5120 7249
rect 5103 7246 5120 7248
rect 5104 7241 5120 7246
rect 5094 7234 5100 7235
rect 5103 7234 5132 7241
rect 5021 7233 5132 7234
rect 5021 7232 5138 7233
rect 4697 7224 4748 7232
rect 4795 7224 4829 7232
rect 4697 7212 4722 7224
rect 4729 7212 4748 7224
rect 4802 7222 4829 7224
rect 4838 7222 5059 7232
rect 5094 7229 5100 7232
rect 4802 7218 5059 7222
rect 4697 7204 4748 7212
rect 4795 7204 5059 7218
rect 5103 7224 5138 7232
rect 4649 7156 4668 7190
rect 4713 7196 4742 7204
rect 4713 7190 4730 7196
rect 4713 7188 4747 7190
rect 4795 7188 4811 7204
rect 4812 7194 5020 7204
rect 5021 7194 5037 7204
rect 5085 7200 5100 7215
rect 5103 7212 5104 7224
rect 5111 7212 5138 7224
rect 5103 7204 5138 7212
rect 5103 7203 5132 7204
rect 4823 7190 5037 7194
rect 4838 7188 5037 7190
rect 5072 7190 5085 7200
rect 5103 7190 5120 7203
rect 5072 7188 5120 7190
rect 4714 7184 4747 7188
rect 4710 7182 4747 7184
rect 4710 7181 4777 7182
rect 4710 7176 4741 7181
rect 4747 7176 4777 7181
rect 4710 7172 4777 7176
rect 4683 7169 4777 7172
rect 4683 7162 4732 7169
rect 4683 7156 4713 7162
rect 4732 7157 4737 7162
rect 4649 7140 4729 7156
rect 4741 7148 4777 7169
rect 4838 7164 5027 7188
rect 5072 7187 5119 7188
rect 5085 7182 5119 7187
rect 4853 7161 5027 7164
rect 4846 7158 5027 7161
rect 5055 7181 5119 7182
rect 4649 7138 4668 7140
rect 4683 7138 4717 7140
rect 4649 7122 4729 7138
rect 4649 7116 4668 7122
rect 4365 7090 4468 7100
rect 4319 7088 4468 7090
rect 4489 7088 4524 7100
rect 4158 7086 4320 7088
rect 4170 7066 4189 7086
rect 4204 7084 4234 7086
rect 4053 7058 4094 7066
rect 4176 7062 4189 7066
rect 4241 7070 4320 7086
rect 4352 7086 4524 7088
rect 4352 7070 4431 7086
rect 4438 7084 4468 7086
rect 4016 7048 4045 7058
rect 4059 7048 4088 7058
rect 4103 7048 4133 7062
rect 4176 7048 4219 7062
rect 4241 7058 4431 7070
rect 4496 7066 4502 7086
rect 4226 7048 4256 7058
rect 4257 7048 4415 7058
rect 4419 7048 4449 7058
rect 4453 7048 4483 7062
rect 4511 7048 4524 7086
rect 4596 7100 4625 7116
rect 4639 7100 4668 7116
rect 4683 7106 4713 7122
rect 4741 7100 4747 7148
rect 4750 7142 4769 7148
rect 4784 7142 4814 7150
rect 4750 7134 4814 7142
rect 4750 7118 4830 7134
rect 4846 7127 4908 7158
rect 4924 7127 4986 7158
rect 5055 7156 5104 7181
rect 5119 7156 5149 7172
rect 5018 7142 5048 7150
rect 5055 7148 5165 7156
rect 5018 7134 5063 7142
rect 4750 7116 4769 7118
rect 4784 7116 4830 7118
rect 4750 7100 4830 7116
rect 4857 7114 4892 7127
rect 4933 7124 4970 7127
rect 4933 7122 4975 7124
rect 4862 7111 4892 7114
rect 4871 7107 4878 7111
rect 4878 7106 4879 7107
rect 4837 7100 4847 7106
rect 4596 7092 4631 7100
rect 4596 7066 4597 7092
rect 4604 7066 4631 7092
rect 4539 7048 4569 7062
rect 4596 7058 4631 7066
rect 4633 7092 4674 7100
rect 4633 7066 4648 7092
rect 4655 7066 4674 7092
rect 4738 7088 4769 7100
rect 4784 7088 4887 7100
rect 4899 7090 4925 7116
rect 4940 7111 4970 7122
rect 5002 7118 5064 7134
rect 5002 7116 5048 7118
rect 5002 7100 5064 7116
rect 5076 7100 5082 7148
rect 5085 7140 5165 7148
rect 5085 7138 5104 7140
rect 5119 7138 5153 7140
rect 5085 7122 5165 7138
rect 5085 7100 5104 7122
rect 5119 7106 5149 7122
rect 5177 7116 5183 7190
rect 5186 7116 5205 7260
rect 5220 7116 5226 7260
rect 5235 7190 5248 7260
rect 5300 7256 5322 7260
rect 5293 7234 5322 7248
rect 5375 7234 5391 7248
rect 5429 7244 5435 7246
rect 5442 7244 5550 7260
rect 5557 7244 5563 7246
rect 5571 7244 5586 7260
rect 5652 7254 5671 7257
rect 5293 7232 5391 7234
rect 5418 7232 5586 7244
rect 5601 7234 5617 7248
rect 5652 7235 5674 7254
rect 5684 7248 5700 7249
rect 5683 7246 5700 7248
rect 5684 7241 5700 7246
rect 5674 7234 5680 7235
rect 5683 7234 5712 7241
rect 5601 7233 5712 7234
rect 5601 7232 5718 7233
rect 5277 7224 5328 7232
rect 5375 7224 5409 7232
rect 5277 7212 5302 7224
rect 5309 7212 5328 7224
rect 5382 7222 5409 7224
rect 5418 7222 5639 7232
rect 5674 7229 5680 7232
rect 5382 7218 5639 7222
rect 5277 7204 5328 7212
rect 5375 7204 5639 7218
rect 5683 7224 5718 7232
rect 5229 7156 5248 7190
rect 5293 7196 5322 7204
rect 5293 7190 5310 7196
rect 5293 7188 5327 7190
rect 5375 7188 5391 7204
rect 5392 7194 5600 7204
rect 5601 7194 5617 7204
rect 5665 7200 5680 7215
rect 5683 7212 5684 7224
rect 5691 7212 5718 7224
rect 5683 7204 5718 7212
rect 5683 7203 5712 7204
rect 5403 7190 5617 7194
rect 5418 7188 5617 7190
rect 5652 7190 5665 7200
rect 5683 7190 5700 7203
rect 5652 7188 5700 7190
rect 5294 7184 5327 7188
rect 5290 7182 5327 7184
rect 5290 7181 5357 7182
rect 5290 7176 5321 7181
rect 5327 7176 5357 7181
rect 5290 7172 5357 7176
rect 5263 7169 5357 7172
rect 5263 7162 5312 7169
rect 5263 7156 5293 7162
rect 5312 7157 5317 7162
rect 5229 7140 5309 7156
rect 5321 7148 5357 7169
rect 5418 7164 5607 7188
rect 5652 7187 5699 7188
rect 5665 7182 5699 7187
rect 5433 7161 5607 7164
rect 5426 7158 5607 7161
rect 5635 7181 5699 7182
rect 5229 7138 5248 7140
rect 5263 7138 5297 7140
rect 5229 7122 5309 7138
rect 5229 7116 5248 7122
rect 4945 7090 5048 7100
rect 4899 7088 5048 7090
rect 5069 7088 5104 7100
rect 4738 7086 4900 7088
rect 4750 7066 4769 7086
rect 4784 7084 4814 7086
rect 4633 7058 4674 7066
rect 4756 7062 4769 7066
rect 4821 7070 4900 7086
rect 4932 7086 5104 7088
rect 4932 7070 5011 7086
rect 5018 7084 5048 7086
rect 4596 7048 4625 7058
rect 4639 7048 4668 7058
rect 4683 7048 4713 7062
rect 4756 7048 4799 7062
rect 4821 7058 5011 7070
rect 5076 7066 5082 7086
rect 4806 7048 4836 7058
rect 4837 7048 4995 7058
rect 4999 7048 5029 7058
rect 5033 7048 5063 7062
rect 5091 7048 5104 7086
rect 5176 7100 5205 7116
rect 5219 7100 5248 7116
rect 5263 7106 5293 7122
rect 5321 7100 5327 7148
rect 5330 7142 5349 7148
rect 5364 7142 5394 7150
rect 5330 7134 5394 7142
rect 5330 7118 5410 7134
rect 5426 7127 5488 7158
rect 5504 7127 5566 7158
rect 5635 7156 5684 7181
rect 5699 7156 5729 7172
rect 5598 7142 5628 7150
rect 5635 7148 5745 7156
rect 5598 7134 5643 7142
rect 5330 7116 5349 7118
rect 5364 7116 5410 7118
rect 5330 7100 5410 7116
rect 5437 7114 5472 7127
rect 5513 7124 5550 7127
rect 5513 7122 5555 7124
rect 5442 7111 5472 7114
rect 5451 7107 5458 7111
rect 5458 7106 5459 7107
rect 5417 7100 5427 7106
rect 5176 7092 5211 7100
rect 5176 7066 5177 7092
rect 5184 7066 5211 7092
rect 5119 7048 5149 7062
rect 5176 7058 5211 7066
rect 5213 7092 5254 7100
rect 5213 7066 5228 7092
rect 5235 7066 5254 7092
rect 5318 7088 5349 7100
rect 5364 7088 5467 7100
rect 5479 7090 5505 7116
rect 5520 7111 5550 7122
rect 5582 7118 5644 7134
rect 5582 7116 5628 7118
rect 5582 7100 5644 7116
rect 5656 7100 5662 7148
rect 5665 7140 5745 7148
rect 5665 7138 5684 7140
rect 5699 7138 5733 7140
rect 5665 7122 5745 7138
rect 5665 7100 5684 7122
rect 5699 7106 5729 7122
rect 5757 7116 5763 7190
rect 5766 7116 5785 7260
rect 5800 7116 5806 7260
rect 5815 7190 5828 7260
rect 5880 7256 5902 7260
rect 5873 7234 5902 7248
rect 5955 7234 5971 7248
rect 6009 7244 6015 7246
rect 6022 7244 6130 7260
rect 6137 7244 6143 7246
rect 6151 7244 6166 7260
rect 6232 7254 6251 7257
rect 5873 7232 5971 7234
rect 5998 7232 6166 7244
rect 6181 7234 6197 7248
rect 6232 7235 6254 7254
rect 6264 7248 6280 7249
rect 6263 7246 6280 7248
rect 6264 7241 6280 7246
rect 6254 7234 6260 7235
rect 6263 7234 6292 7241
rect 6181 7233 6292 7234
rect 6181 7232 6298 7233
rect 5857 7224 5908 7232
rect 5955 7224 5989 7232
rect 5857 7212 5882 7224
rect 5889 7212 5908 7224
rect 5962 7222 5989 7224
rect 5998 7222 6219 7232
rect 6254 7229 6260 7232
rect 5962 7218 6219 7222
rect 5857 7204 5908 7212
rect 5955 7204 6219 7218
rect 6263 7224 6298 7232
rect 5809 7156 5828 7190
rect 5873 7196 5902 7204
rect 5873 7190 5890 7196
rect 5873 7188 5907 7190
rect 5955 7188 5971 7204
rect 5972 7194 6180 7204
rect 6181 7194 6197 7204
rect 6245 7200 6260 7215
rect 6263 7212 6264 7224
rect 6271 7212 6298 7224
rect 6263 7204 6298 7212
rect 6263 7203 6292 7204
rect 5983 7190 6197 7194
rect 5998 7188 6197 7190
rect 6232 7190 6245 7200
rect 6263 7190 6280 7203
rect 6232 7188 6280 7190
rect 5874 7184 5907 7188
rect 5870 7182 5907 7184
rect 5870 7181 5937 7182
rect 5870 7176 5901 7181
rect 5907 7176 5937 7181
rect 5870 7172 5937 7176
rect 5843 7169 5937 7172
rect 5843 7162 5892 7169
rect 5843 7156 5873 7162
rect 5892 7157 5897 7162
rect 5809 7140 5889 7156
rect 5901 7148 5937 7169
rect 5998 7164 6187 7188
rect 6232 7187 6279 7188
rect 6245 7182 6279 7187
rect 6013 7161 6187 7164
rect 6006 7158 6187 7161
rect 6215 7181 6279 7182
rect 5809 7138 5828 7140
rect 5843 7138 5877 7140
rect 5809 7122 5889 7138
rect 5809 7116 5828 7122
rect 5525 7090 5628 7100
rect 5479 7088 5628 7090
rect 5649 7088 5684 7100
rect 5318 7086 5480 7088
rect 5330 7066 5349 7086
rect 5364 7084 5394 7086
rect 5213 7058 5254 7066
rect 5336 7062 5349 7066
rect 5401 7070 5480 7086
rect 5512 7086 5684 7088
rect 5512 7070 5591 7086
rect 5598 7084 5628 7086
rect 5176 7048 5205 7058
rect 5219 7048 5248 7058
rect 5263 7048 5293 7062
rect 5336 7048 5379 7062
rect 5401 7058 5591 7070
rect 5656 7066 5662 7086
rect 5386 7048 5416 7058
rect 5417 7048 5575 7058
rect 5579 7048 5609 7058
rect 5613 7048 5643 7062
rect 5671 7048 5684 7086
rect 5756 7100 5785 7116
rect 5799 7100 5828 7116
rect 5843 7106 5873 7122
rect 5901 7100 5907 7148
rect 5910 7142 5929 7148
rect 5944 7142 5974 7150
rect 5910 7134 5974 7142
rect 5910 7118 5990 7134
rect 6006 7127 6068 7158
rect 6084 7127 6146 7158
rect 6215 7156 6264 7181
rect 6279 7156 6309 7172
rect 6178 7142 6208 7150
rect 6215 7148 6325 7156
rect 6178 7134 6223 7142
rect 5910 7116 5929 7118
rect 5944 7116 5990 7118
rect 5910 7100 5990 7116
rect 6017 7114 6052 7127
rect 6093 7124 6130 7127
rect 6093 7122 6135 7124
rect 6022 7111 6052 7114
rect 6031 7107 6038 7111
rect 6038 7106 6039 7107
rect 5997 7100 6007 7106
rect 5756 7092 5791 7100
rect 5756 7066 5757 7092
rect 5764 7066 5791 7092
rect 5699 7048 5729 7062
rect 5756 7058 5791 7066
rect 5793 7092 5834 7100
rect 5793 7066 5808 7092
rect 5815 7066 5834 7092
rect 5898 7088 5929 7100
rect 5944 7088 6047 7100
rect 6059 7090 6085 7116
rect 6100 7111 6130 7122
rect 6162 7118 6224 7134
rect 6162 7116 6208 7118
rect 6162 7100 6224 7116
rect 6236 7100 6242 7148
rect 6245 7140 6325 7148
rect 6245 7138 6264 7140
rect 6279 7138 6313 7140
rect 6245 7122 6325 7138
rect 6245 7100 6264 7122
rect 6279 7106 6309 7122
rect 6337 7116 6343 7190
rect 6346 7116 6365 7260
rect 6380 7116 6386 7260
rect 6395 7190 6408 7260
rect 6460 7256 6482 7260
rect 6453 7234 6482 7248
rect 6535 7234 6551 7248
rect 6589 7244 6595 7246
rect 6602 7244 6710 7260
rect 6717 7244 6723 7246
rect 6731 7244 6746 7260
rect 6812 7254 6831 7257
rect 6453 7232 6551 7234
rect 6578 7232 6746 7244
rect 6761 7234 6777 7248
rect 6812 7235 6834 7254
rect 6844 7248 6860 7249
rect 6843 7246 6860 7248
rect 6844 7241 6860 7246
rect 6834 7234 6840 7235
rect 6843 7234 6872 7241
rect 6761 7233 6872 7234
rect 6761 7232 6878 7233
rect 6437 7224 6488 7232
rect 6535 7224 6569 7232
rect 6437 7212 6462 7224
rect 6469 7212 6488 7224
rect 6542 7222 6569 7224
rect 6578 7222 6799 7232
rect 6834 7229 6840 7232
rect 6542 7218 6799 7222
rect 6437 7204 6488 7212
rect 6535 7204 6799 7218
rect 6843 7224 6878 7232
rect 6389 7156 6408 7190
rect 6453 7196 6482 7204
rect 6453 7190 6470 7196
rect 6453 7188 6487 7190
rect 6535 7188 6551 7204
rect 6552 7194 6760 7204
rect 6761 7194 6777 7204
rect 6825 7200 6840 7215
rect 6843 7212 6844 7224
rect 6851 7212 6878 7224
rect 6843 7204 6878 7212
rect 6843 7203 6872 7204
rect 6563 7190 6777 7194
rect 6578 7188 6777 7190
rect 6812 7190 6825 7200
rect 6843 7190 6860 7203
rect 6812 7188 6860 7190
rect 6454 7184 6487 7188
rect 6450 7182 6487 7184
rect 6450 7181 6517 7182
rect 6450 7176 6481 7181
rect 6487 7176 6517 7181
rect 6450 7172 6517 7176
rect 6423 7169 6517 7172
rect 6423 7162 6472 7169
rect 6423 7156 6453 7162
rect 6472 7157 6477 7162
rect 6389 7140 6469 7156
rect 6481 7148 6517 7169
rect 6578 7164 6767 7188
rect 6812 7187 6859 7188
rect 6825 7182 6859 7187
rect 6593 7161 6767 7164
rect 6586 7158 6767 7161
rect 6795 7181 6859 7182
rect 6389 7138 6408 7140
rect 6423 7138 6457 7140
rect 6389 7122 6469 7138
rect 6389 7116 6408 7122
rect 6105 7090 6208 7100
rect 6059 7088 6208 7090
rect 6229 7088 6264 7100
rect 5898 7086 6060 7088
rect 5910 7066 5929 7086
rect 5944 7084 5974 7086
rect 5793 7058 5834 7066
rect 5916 7062 5929 7066
rect 5981 7070 6060 7086
rect 6092 7086 6264 7088
rect 6092 7070 6171 7086
rect 6178 7084 6208 7086
rect 5756 7048 5785 7058
rect 5799 7048 5828 7058
rect 5843 7048 5873 7062
rect 5916 7048 5959 7062
rect 5981 7058 6171 7070
rect 6236 7066 6242 7086
rect 5966 7048 5996 7058
rect 5997 7048 6155 7058
rect 6159 7048 6189 7058
rect 6193 7048 6223 7062
rect 6251 7048 6264 7086
rect 6336 7100 6365 7116
rect 6379 7100 6408 7116
rect 6423 7106 6453 7122
rect 6481 7100 6487 7148
rect 6490 7142 6509 7148
rect 6524 7142 6554 7150
rect 6490 7134 6554 7142
rect 6490 7118 6570 7134
rect 6586 7127 6648 7158
rect 6664 7127 6726 7158
rect 6795 7156 6844 7181
rect 6859 7156 6889 7172
rect 6758 7142 6788 7150
rect 6795 7148 6905 7156
rect 6758 7134 6803 7142
rect 6490 7116 6509 7118
rect 6524 7116 6570 7118
rect 6490 7100 6570 7116
rect 6597 7114 6632 7127
rect 6673 7124 6710 7127
rect 6673 7122 6715 7124
rect 6602 7111 6632 7114
rect 6611 7107 6618 7111
rect 6618 7106 6619 7107
rect 6577 7100 6587 7106
rect 6336 7092 6371 7100
rect 6336 7066 6337 7092
rect 6344 7066 6371 7092
rect 6279 7048 6309 7062
rect 6336 7058 6371 7066
rect 6373 7092 6414 7100
rect 6373 7066 6388 7092
rect 6395 7066 6414 7092
rect 6478 7088 6509 7100
rect 6524 7088 6627 7100
rect 6639 7090 6665 7116
rect 6680 7111 6710 7122
rect 6742 7118 6804 7134
rect 6742 7116 6788 7118
rect 6742 7100 6804 7116
rect 6816 7100 6822 7148
rect 6825 7140 6905 7148
rect 6825 7138 6844 7140
rect 6859 7138 6893 7140
rect 6825 7122 6905 7138
rect 6825 7100 6844 7122
rect 6859 7106 6889 7122
rect 6917 7116 6923 7190
rect 6926 7116 6945 7260
rect 6960 7116 6966 7260
rect 6975 7190 6988 7260
rect 7040 7256 7062 7260
rect 7033 7234 7062 7248
rect 7115 7234 7131 7248
rect 7169 7244 7175 7246
rect 7182 7244 7290 7260
rect 7297 7244 7303 7246
rect 7311 7244 7326 7260
rect 7392 7254 7411 7257
rect 7033 7232 7131 7234
rect 7158 7232 7326 7244
rect 7341 7234 7357 7248
rect 7392 7235 7414 7254
rect 7424 7248 7440 7249
rect 7423 7246 7440 7248
rect 7424 7241 7440 7246
rect 7414 7234 7420 7235
rect 7423 7234 7452 7241
rect 7341 7233 7452 7234
rect 7341 7232 7458 7233
rect 7017 7224 7068 7232
rect 7115 7224 7149 7232
rect 7017 7212 7042 7224
rect 7049 7212 7068 7224
rect 7122 7222 7149 7224
rect 7158 7222 7379 7232
rect 7414 7229 7420 7232
rect 7122 7218 7379 7222
rect 7017 7204 7068 7212
rect 7115 7204 7379 7218
rect 7423 7224 7458 7232
rect 6969 7156 6988 7190
rect 7033 7196 7062 7204
rect 7033 7190 7050 7196
rect 7033 7188 7067 7190
rect 7115 7188 7131 7204
rect 7132 7194 7340 7204
rect 7341 7194 7357 7204
rect 7405 7200 7420 7215
rect 7423 7212 7424 7224
rect 7431 7212 7458 7224
rect 7423 7204 7458 7212
rect 7423 7203 7452 7204
rect 7143 7190 7357 7194
rect 7158 7188 7357 7190
rect 7392 7190 7405 7200
rect 7423 7190 7440 7203
rect 7392 7188 7440 7190
rect 7034 7184 7067 7188
rect 7030 7182 7067 7184
rect 7030 7181 7097 7182
rect 7030 7176 7061 7181
rect 7067 7176 7097 7181
rect 7030 7172 7097 7176
rect 7003 7169 7097 7172
rect 7003 7162 7052 7169
rect 7003 7156 7033 7162
rect 7052 7157 7057 7162
rect 6969 7140 7049 7156
rect 7061 7148 7097 7169
rect 7158 7164 7347 7188
rect 7392 7187 7439 7188
rect 7405 7182 7439 7187
rect 7173 7161 7347 7164
rect 7166 7158 7347 7161
rect 7375 7181 7439 7182
rect 6969 7138 6988 7140
rect 7003 7138 7037 7140
rect 6969 7122 7049 7138
rect 6969 7116 6988 7122
rect 6685 7090 6788 7100
rect 6639 7088 6788 7090
rect 6809 7088 6844 7100
rect 6478 7086 6640 7088
rect 6490 7066 6509 7086
rect 6524 7084 6554 7086
rect 6373 7058 6414 7066
rect 6496 7062 6509 7066
rect 6561 7070 6640 7086
rect 6672 7086 6844 7088
rect 6672 7070 6751 7086
rect 6758 7084 6788 7086
rect 6336 7048 6365 7058
rect 6379 7048 6408 7058
rect 6423 7048 6453 7062
rect 6496 7048 6539 7062
rect 6561 7058 6751 7070
rect 6816 7066 6822 7086
rect 6546 7048 6576 7058
rect 6577 7048 6735 7058
rect 6739 7048 6769 7058
rect 6773 7048 6803 7062
rect 6831 7048 6844 7086
rect 6916 7100 6945 7116
rect 6959 7100 6988 7116
rect 7003 7106 7033 7122
rect 7061 7100 7067 7148
rect 7070 7142 7089 7148
rect 7104 7142 7134 7150
rect 7070 7134 7134 7142
rect 7070 7118 7150 7134
rect 7166 7127 7228 7158
rect 7244 7127 7306 7158
rect 7375 7156 7424 7181
rect 7439 7156 7469 7172
rect 7338 7142 7368 7150
rect 7375 7148 7485 7156
rect 7338 7134 7383 7142
rect 7070 7116 7089 7118
rect 7104 7116 7150 7118
rect 7070 7100 7150 7116
rect 7177 7114 7212 7127
rect 7253 7124 7290 7127
rect 7253 7122 7295 7124
rect 7182 7111 7212 7114
rect 7191 7107 7198 7111
rect 7198 7106 7199 7107
rect 7157 7100 7167 7106
rect 6916 7092 6951 7100
rect 6916 7066 6917 7092
rect 6924 7066 6951 7092
rect 6859 7048 6889 7062
rect 6916 7058 6951 7066
rect 6953 7092 6994 7100
rect 6953 7066 6968 7092
rect 6975 7066 6994 7092
rect 7058 7088 7089 7100
rect 7104 7088 7207 7100
rect 7219 7090 7245 7116
rect 7260 7111 7290 7122
rect 7322 7118 7384 7134
rect 7322 7116 7368 7118
rect 7322 7100 7384 7116
rect 7396 7100 7402 7148
rect 7405 7140 7485 7148
rect 7405 7138 7424 7140
rect 7439 7138 7473 7140
rect 7405 7122 7485 7138
rect 7405 7100 7424 7122
rect 7439 7106 7469 7122
rect 7497 7116 7503 7190
rect 7506 7116 7525 7260
rect 7540 7116 7546 7260
rect 7555 7190 7568 7260
rect 7620 7256 7642 7260
rect 7613 7234 7642 7248
rect 7695 7234 7711 7248
rect 7749 7244 7755 7246
rect 7762 7244 7870 7260
rect 7877 7244 7883 7246
rect 7891 7244 7906 7260
rect 7972 7254 7991 7257
rect 7613 7232 7711 7234
rect 7738 7232 7906 7244
rect 7921 7234 7937 7248
rect 7972 7235 7994 7254
rect 8004 7248 8020 7249
rect 8003 7246 8020 7248
rect 8004 7241 8020 7246
rect 7994 7234 8000 7235
rect 8003 7234 8032 7241
rect 7921 7233 8032 7234
rect 7921 7232 8038 7233
rect 7597 7224 7648 7232
rect 7695 7224 7729 7232
rect 7597 7212 7622 7224
rect 7629 7212 7648 7224
rect 7702 7222 7729 7224
rect 7738 7222 7959 7232
rect 7994 7229 8000 7232
rect 7702 7218 7959 7222
rect 7597 7204 7648 7212
rect 7695 7204 7959 7218
rect 8003 7224 8038 7232
rect 7549 7156 7568 7190
rect 7613 7196 7642 7204
rect 7613 7190 7630 7196
rect 7613 7188 7647 7190
rect 7695 7188 7711 7204
rect 7712 7194 7920 7204
rect 7921 7194 7937 7204
rect 7985 7200 8000 7215
rect 8003 7212 8004 7224
rect 8011 7212 8038 7224
rect 8003 7204 8038 7212
rect 8003 7203 8032 7204
rect 7723 7190 7937 7194
rect 7738 7188 7937 7190
rect 7972 7190 7985 7200
rect 8003 7190 8020 7203
rect 7972 7188 8020 7190
rect 7614 7184 7647 7188
rect 7610 7182 7647 7184
rect 7610 7181 7677 7182
rect 7610 7176 7641 7181
rect 7647 7176 7677 7181
rect 7610 7172 7677 7176
rect 7583 7169 7677 7172
rect 7583 7162 7632 7169
rect 7583 7156 7613 7162
rect 7632 7157 7637 7162
rect 7549 7140 7629 7156
rect 7641 7148 7677 7169
rect 7738 7164 7927 7188
rect 7972 7187 8019 7188
rect 7985 7182 8019 7187
rect 7753 7161 7927 7164
rect 7746 7158 7927 7161
rect 7955 7181 8019 7182
rect 7549 7138 7568 7140
rect 7583 7138 7617 7140
rect 7549 7122 7629 7138
rect 7549 7116 7568 7122
rect 7265 7090 7368 7100
rect 7219 7088 7368 7090
rect 7389 7088 7424 7100
rect 7058 7086 7220 7088
rect 7070 7066 7089 7086
rect 7104 7084 7134 7086
rect 6953 7058 6994 7066
rect 7076 7062 7089 7066
rect 7141 7070 7220 7086
rect 7252 7086 7424 7088
rect 7252 7070 7331 7086
rect 7338 7084 7368 7086
rect 6916 7048 6945 7058
rect 6959 7048 6988 7058
rect 7003 7048 7033 7062
rect 7076 7048 7119 7062
rect 7141 7058 7331 7070
rect 7396 7066 7402 7086
rect 7126 7048 7156 7058
rect 7157 7048 7315 7058
rect 7319 7048 7349 7058
rect 7353 7048 7383 7062
rect 7411 7048 7424 7086
rect 7496 7100 7525 7116
rect 7539 7100 7568 7116
rect 7583 7106 7613 7122
rect 7641 7100 7647 7148
rect 7650 7142 7669 7148
rect 7684 7142 7714 7150
rect 7650 7134 7714 7142
rect 7650 7118 7730 7134
rect 7746 7127 7808 7158
rect 7824 7127 7886 7158
rect 7955 7156 8004 7181
rect 8019 7156 8049 7172
rect 7918 7142 7948 7150
rect 7955 7148 8065 7156
rect 7918 7134 7963 7142
rect 7650 7116 7669 7118
rect 7684 7116 7730 7118
rect 7650 7100 7730 7116
rect 7757 7114 7792 7127
rect 7833 7124 7870 7127
rect 7833 7122 7875 7124
rect 7762 7111 7792 7114
rect 7771 7107 7778 7111
rect 7778 7106 7779 7107
rect 7737 7100 7747 7106
rect 7496 7092 7531 7100
rect 7496 7066 7497 7092
rect 7504 7066 7531 7092
rect 7439 7048 7469 7062
rect 7496 7058 7531 7066
rect 7533 7092 7574 7100
rect 7533 7066 7548 7092
rect 7555 7066 7574 7092
rect 7638 7088 7669 7100
rect 7684 7088 7787 7100
rect 7799 7090 7825 7116
rect 7840 7111 7870 7122
rect 7902 7118 7964 7134
rect 7902 7116 7948 7118
rect 7902 7100 7964 7116
rect 7976 7100 7982 7148
rect 7985 7140 8065 7148
rect 7985 7138 8004 7140
rect 8019 7138 8053 7140
rect 7985 7122 8065 7138
rect 7985 7100 8004 7122
rect 8019 7106 8049 7122
rect 8077 7116 8083 7190
rect 8086 7116 8105 7260
rect 8120 7116 8126 7260
rect 8135 7190 8148 7260
rect 8200 7256 8222 7260
rect 8193 7234 8222 7248
rect 8275 7234 8291 7248
rect 8329 7244 8335 7246
rect 8342 7244 8450 7260
rect 8457 7244 8463 7246
rect 8471 7244 8486 7260
rect 8552 7254 8571 7257
rect 8193 7232 8291 7234
rect 8318 7232 8486 7244
rect 8501 7234 8517 7248
rect 8552 7235 8574 7254
rect 8584 7248 8600 7249
rect 8583 7246 8600 7248
rect 8584 7241 8600 7246
rect 8574 7234 8580 7235
rect 8583 7234 8612 7241
rect 8501 7233 8612 7234
rect 8501 7232 8618 7233
rect 8177 7224 8228 7232
rect 8275 7224 8309 7232
rect 8177 7212 8202 7224
rect 8209 7212 8228 7224
rect 8282 7222 8309 7224
rect 8318 7222 8539 7232
rect 8574 7229 8580 7232
rect 8282 7218 8539 7222
rect 8177 7204 8228 7212
rect 8275 7204 8539 7218
rect 8583 7224 8618 7232
rect 8129 7156 8148 7190
rect 8193 7196 8222 7204
rect 8193 7190 8210 7196
rect 8193 7188 8227 7190
rect 8275 7188 8291 7204
rect 8292 7194 8500 7204
rect 8501 7194 8517 7204
rect 8565 7200 8580 7215
rect 8583 7212 8584 7224
rect 8591 7212 8618 7224
rect 8583 7204 8618 7212
rect 8583 7203 8612 7204
rect 8303 7190 8517 7194
rect 8318 7188 8517 7190
rect 8552 7190 8565 7200
rect 8583 7190 8600 7203
rect 8552 7188 8600 7190
rect 8194 7184 8227 7188
rect 8190 7182 8227 7184
rect 8190 7181 8257 7182
rect 8190 7176 8221 7181
rect 8227 7176 8257 7181
rect 8190 7172 8257 7176
rect 8163 7169 8257 7172
rect 8163 7162 8212 7169
rect 8163 7156 8193 7162
rect 8212 7157 8217 7162
rect 8129 7140 8209 7156
rect 8221 7148 8257 7169
rect 8318 7164 8507 7188
rect 8552 7187 8599 7188
rect 8565 7182 8599 7187
rect 8333 7161 8507 7164
rect 8326 7158 8507 7161
rect 8535 7181 8599 7182
rect 8129 7138 8148 7140
rect 8163 7138 8197 7140
rect 8129 7122 8209 7138
rect 8129 7116 8148 7122
rect 7845 7090 7948 7100
rect 7799 7088 7948 7090
rect 7969 7088 8004 7100
rect 7638 7086 7800 7088
rect 7650 7066 7669 7086
rect 7684 7084 7714 7086
rect 7533 7058 7574 7066
rect 7656 7062 7669 7066
rect 7721 7070 7800 7086
rect 7832 7086 8004 7088
rect 7832 7070 7911 7086
rect 7918 7084 7948 7086
rect 7496 7048 7525 7058
rect 7539 7048 7568 7058
rect 7583 7048 7613 7062
rect 7656 7048 7699 7062
rect 7721 7058 7911 7070
rect 7976 7066 7982 7086
rect 7706 7048 7736 7058
rect 7737 7048 7895 7058
rect 7899 7048 7929 7058
rect 7933 7048 7963 7062
rect 7991 7048 8004 7086
rect 8076 7100 8105 7116
rect 8119 7100 8148 7116
rect 8163 7106 8193 7122
rect 8221 7100 8227 7148
rect 8230 7142 8249 7148
rect 8264 7142 8294 7150
rect 8230 7134 8294 7142
rect 8230 7118 8310 7134
rect 8326 7127 8388 7158
rect 8404 7127 8466 7158
rect 8535 7156 8584 7181
rect 8599 7156 8629 7172
rect 8498 7142 8528 7150
rect 8535 7148 8645 7156
rect 8498 7134 8543 7142
rect 8230 7116 8249 7118
rect 8264 7116 8310 7118
rect 8230 7100 8310 7116
rect 8337 7114 8372 7127
rect 8413 7124 8450 7127
rect 8413 7122 8455 7124
rect 8342 7111 8372 7114
rect 8351 7107 8358 7111
rect 8358 7106 8359 7107
rect 8317 7100 8327 7106
rect 8076 7092 8111 7100
rect 8076 7066 8077 7092
rect 8084 7066 8111 7092
rect 8019 7048 8049 7062
rect 8076 7058 8111 7066
rect 8113 7092 8154 7100
rect 8113 7066 8128 7092
rect 8135 7066 8154 7092
rect 8218 7088 8249 7100
rect 8264 7088 8367 7100
rect 8379 7090 8405 7116
rect 8420 7111 8450 7122
rect 8482 7118 8544 7134
rect 8482 7116 8528 7118
rect 8482 7100 8544 7116
rect 8556 7100 8562 7148
rect 8565 7140 8645 7148
rect 8565 7138 8584 7140
rect 8599 7138 8633 7140
rect 8565 7122 8645 7138
rect 8565 7100 8584 7122
rect 8599 7106 8629 7122
rect 8657 7116 8663 7190
rect 8666 7116 8685 7260
rect 8700 7116 8706 7260
rect 8715 7190 8728 7260
rect 8780 7256 8802 7260
rect 8773 7234 8802 7248
rect 8855 7234 8871 7248
rect 8909 7244 8915 7246
rect 8922 7244 9030 7260
rect 9037 7244 9043 7246
rect 9051 7244 9066 7260
rect 9132 7254 9151 7257
rect 8773 7232 8871 7234
rect 8898 7232 9066 7244
rect 9081 7234 9097 7248
rect 9132 7235 9154 7254
rect 9164 7248 9180 7249
rect 9163 7246 9180 7248
rect 9164 7241 9180 7246
rect 9154 7234 9160 7235
rect 9163 7234 9192 7241
rect 9081 7233 9192 7234
rect 9081 7232 9198 7233
rect 8757 7224 8808 7232
rect 8855 7224 8889 7232
rect 8757 7212 8782 7224
rect 8789 7212 8808 7224
rect 8862 7222 8889 7224
rect 8898 7222 9119 7232
rect 9154 7229 9160 7232
rect 8862 7218 9119 7222
rect 8757 7204 8808 7212
rect 8855 7204 9119 7218
rect 9163 7224 9198 7232
rect 8709 7156 8728 7190
rect 8773 7196 8802 7204
rect 8773 7190 8790 7196
rect 8773 7188 8807 7190
rect 8855 7188 8871 7204
rect 8872 7194 9080 7204
rect 9081 7194 9097 7204
rect 9145 7200 9160 7215
rect 9163 7212 9164 7224
rect 9171 7212 9198 7224
rect 9163 7204 9198 7212
rect 9163 7203 9192 7204
rect 8883 7190 9097 7194
rect 8898 7188 9097 7190
rect 9132 7190 9145 7200
rect 9163 7190 9180 7203
rect 9132 7188 9180 7190
rect 8774 7184 8807 7188
rect 8770 7182 8807 7184
rect 8770 7181 8837 7182
rect 8770 7176 8801 7181
rect 8807 7176 8837 7181
rect 8770 7172 8837 7176
rect 8743 7169 8837 7172
rect 8743 7162 8792 7169
rect 8743 7156 8773 7162
rect 8792 7157 8797 7162
rect 8709 7140 8789 7156
rect 8801 7148 8837 7169
rect 8898 7164 9087 7188
rect 9132 7187 9179 7188
rect 9145 7182 9179 7187
rect 8913 7161 9087 7164
rect 8906 7158 9087 7161
rect 9115 7181 9179 7182
rect 8709 7138 8728 7140
rect 8743 7138 8777 7140
rect 8709 7122 8789 7138
rect 8709 7116 8728 7122
rect 8425 7090 8528 7100
rect 8379 7088 8528 7090
rect 8549 7088 8584 7100
rect 8218 7086 8380 7088
rect 8230 7066 8249 7086
rect 8264 7084 8294 7086
rect 8113 7058 8154 7066
rect 8236 7062 8249 7066
rect 8301 7070 8380 7086
rect 8412 7086 8584 7088
rect 8412 7070 8491 7086
rect 8498 7084 8528 7086
rect 8076 7048 8105 7058
rect 8119 7048 8148 7058
rect 8163 7048 8193 7062
rect 8236 7048 8279 7062
rect 8301 7058 8491 7070
rect 8556 7066 8562 7086
rect 8286 7048 8316 7058
rect 8317 7048 8475 7058
rect 8479 7048 8509 7058
rect 8513 7048 8543 7062
rect 8571 7048 8584 7086
rect 8656 7100 8685 7116
rect 8699 7100 8728 7116
rect 8743 7106 8773 7122
rect 8801 7100 8807 7148
rect 8810 7142 8829 7148
rect 8844 7142 8874 7150
rect 8810 7134 8874 7142
rect 8810 7118 8890 7134
rect 8906 7127 8968 7158
rect 8984 7127 9046 7158
rect 9115 7156 9164 7181
rect 9179 7156 9209 7172
rect 9078 7142 9108 7150
rect 9115 7148 9225 7156
rect 9078 7134 9123 7142
rect 8810 7116 8829 7118
rect 8844 7116 8890 7118
rect 8810 7100 8890 7116
rect 8917 7114 8952 7127
rect 8993 7124 9030 7127
rect 8993 7122 9035 7124
rect 8922 7111 8952 7114
rect 8931 7107 8938 7111
rect 8938 7106 8939 7107
rect 8897 7100 8907 7106
rect 8656 7092 8691 7100
rect 8656 7066 8657 7092
rect 8664 7066 8691 7092
rect 8599 7048 8629 7062
rect 8656 7058 8691 7066
rect 8693 7092 8734 7100
rect 8693 7066 8708 7092
rect 8715 7066 8734 7092
rect 8798 7088 8829 7100
rect 8844 7088 8947 7100
rect 8959 7090 8985 7116
rect 9000 7111 9030 7122
rect 9062 7118 9124 7134
rect 9062 7116 9108 7118
rect 9062 7100 9124 7116
rect 9136 7100 9142 7148
rect 9145 7140 9225 7148
rect 9145 7138 9164 7140
rect 9179 7138 9213 7140
rect 9145 7122 9225 7138
rect 9145 7100 9164 7122
rect 9179 7106 9209 7122
rect 9237 7116 9243 7190
rect 9246 7116 9265 7260
rect 9280 7116 9286 7260
rect 9295 7190 9308 7260
rect 9360 7256 9382 7260
rect 9353 7234 9382 7248
rect 9435 7234 9451 7248
rect 9489 7244 9495 7246
rect 9502 7244 9610 7260
rect 9617 7244 9623 7246
rect 9631 7244 9646 7260
rect 9712 7254 9731 7257
rect 9353 7232 9451 7234
rect 9478 7232 9646 7244
rect 9661 7234 9677 7248
rect 9712 7235 9734 7254
rect 9744 7248 9760 7249
rect 9743 7246 9760 7248
rect 9744 7241 9760 7246
rect 9734 7234 9740 7235
rect 9743 7234 9772 7241
rect 9661 7233 9772 7234
rect 9661 7232 9778 7233
rect 9337 7224 9388 7232
rect 9435 7224 9469 7232
rect 9337 7212 9362 7224
rect 9369 7212 9388 7224
rect 9442 7222 9469 7224
rect 9478 7222 9699 7232
rect 9734 7229 9740 7232
rect 9442 7218 9699 7222
rect 9337 7204 9388 7212
rect 9435 7204 9699 7218
rect 9743 7224 9778 7232
rect 9289 7156 9308 7190
rect 9353 7196 9382 7204
rect 9353 7190 9370 7196
rect 9353 7188 9387 7190
rect 9435 7188 9451 7204
rect 9452 7194 9660 7204
rect 9661 7194 9677 7204
rect 9725 7200 9740 7215
rect 9743 7212 9744 7224
rect 9751 7212 9778 7224
rect 9743 7204 9778 7212
rect 9743 7203 9772 7204
rect 9463 7190 9677 7194
rect 9478 7188 9677 7190
rect 9712 7190 9725 7200
rect 9743 7190 9760 7203
rect 9712 7188 9760 7190
rect 9354 7184 9387 7188
rect 9350 7182 9387 7184
rect 9350 7181 9417 7182
rect 9350 7176 9381 7181
rect 9387 7176 9417 7181
rect 9350 7172 9417 7176
rect 9323 7169 9417 7172
rect 9323 7162 9372 7169
rect 9323 7156 9353 7162
rect 9372 7157 9377 7162
rect 9289 7140 9369 7156
rect 9381 7148 9417 7169
rect 9478 7164 9667 7188
rect 9712 7187 9759 7188
rect 9725 7182 9759 7187
rect 9493 7161 9667 7164
rect 9486 7158 9667 7161
rect 9695 7181 9759 7182
rect 9289 7138 9308 7140
rect 9323 7138 9357 7140
rect 9289 7122 9369 7138
rect 9289 7116 9308 7122
rect 9005 7090 9108 7100
rect 8959 7088 9108 7090
rect 9129 7088 9164 7100
rect 8798 7086 8960 7088
rect 8810 7066 8829 7086
rect 8844 7084 8874 7086
rect 8693 7058 8734 7066
rect 8816 7062 8829 7066
rect 8881 7070 8960 7086
rect 8992 7086 9164 7088
rect 8992 7070 9071 7086
rect 9078 7084 9108 7086
rect 8656 7048 8685 7058
rect 8699 7048 8728 7058
rect 8743 7048 8773 7062
rect 8816 7048 8859 7062
rect 8881 7058 9071 7070
rect 9136 7066 9142 7086
rect 8866 7048 8896 7058
rect 8897 7048 9055 7058
rect 9059 7048 9089 7058
rect 9093 7048 9123 7062
rect 9151 7048 9164 7086
rect 9236 7100 9265 7116
rect 9279 7100 9308 7116
rect 9323 7106 9353 7122
rect 9381 7100 9387 7148
rect 9390 7142 9409 7148
rect 9424 7142 9454 7150
rect 9390 7134 9454 7142
rect 9390 7118 9470 7134
rect 9486 7127 9548 7158
rect 9564 7127 9626 7158
rect 9695 7156 9744 7181
rect 9759 7156 9789 7172
rect 9658 7142 9688 7150
rect 9695 7148 9805 7156
rect 9658 7134 9703 7142
rect 9390 7116 9409 7118
rect 9424 7116 9470 7118
rect 9390 7100 9470 7116
rect 9497 7114 9532 7127
rect 9573 7124 9610 7127
rect 9573 7122 9615 7124
rect 9502 7111 9532 7114
rect 9511 7107 9518 7111
rect 9518 7106 9519 7107
rect 9477 7100 9487 7106
rect 9236 7092 9271 7100
rect 9236 7066 9237 7092
rect 9244 7066 9271 7092
rect 9179 7048 9209 7062
rect 9236 7058 9271 7066
rect 9273 7092 9314 7100
rect 9273 7066 9288 7092
rect 9295 7066 9314 7092
rect 9378 7088 9409 7100
rect 9424 7088 9527 7100
rect 9539 7090 9565 7116
rect 9580 7111 9610 7122
rect 9642 7118 9704 7134
rect 9642 7116 9688 7118
rect 9642 7100 9704 7116
rect 9716 7100 9722 7148
rect 9725 7140 9805 7148
rect 9725 7138 9744 7140
rect 9759 7138 9793 7140
rect 9725 7122 9805 7138
rect 9725 7100 9744 7122
rect 9759 7106 9789 7122
rect 9817 7116 9823 7190
rect 9826 7116 9845 7260
rect 9860 7116 9866 7260
rect 9875 7190 9888 7260
rect 9940 7256 9962 7260
rect 9933 7234 9962 7248
rect 10015 7234 10031 7248
rect 10069 7244 10075 7246
rect 10082 7244 10190 7260
rect 10197 7244 10203 7246
rect 10211 7244 10226 7260
rect 10292 7254 10311 7257
rect 9933 7232 10031 7234
rect 10058 7232 10226 7244
rect 10241 7234 10257 7248
rect 10292 7235 10314 7254
rect 10324 7248 10340 7249
rect 10323 7246 10340 7248
rect 10324 7241 10340 7246
rect 10314 7234 10320 7235
rect 10323 7234 10352 7241
rect 10241 7233 10352 7234
rect 10241 7232 10358 7233
rect 9917 7224 9968 7232
rect 10015 7224 10049 7232
rect 9917 7212 9942 7224
rect 9949 7212 9968 7224
rect 10022 7222 10049 7224
rect 10058 7222 10279 7232
rect 10314 7229 10320 7232
rect 10022 7218 10279 7222
rect 9917 7204 9968 7212
rect 10015 7204 10279 7218
rect 10323 7224 10358 7232
rect 9869 7156 9888 7190
rect 9933 7196 9962 7204
rect 9933 7190 9950 7196
rect 9933 7188 9967 7190
rect 10015 7188 10031 7204
rect 10032 7194 10240 7204
rect 10241 7194 10257 7204
rect 10305 7200 10320 7215
rect 10323 7212 10324 7224
rect 10331 7212 10358 7224
rect 10323 7204 10358 7212
rect 10323 7203 10352 7204
rect 10043 7190 10257 7194
rect 10058 7188 10257 7190
rect 10292 7190 10305 7200
rect 10323 7190 10340 7203
rect 10292 7188 10340 7190
rect 9934 7184 9967 7188
rect 9930 7182 9967 7184
rect 9930 7181 9997 7182
rect 9930 7176 9961 7181
rect 9967 7176 9997 7181
rect 9930 7172 9997 7176
rect 9903 7169 9997 7172
rect 9903 7162 9952 7169
rect 9903 7156 9933 7162
rect 9952 7157 9957 7162
rect 9869 7140 9949 7156
rect 9961 7148 9997 7169
rect 10058 7164 10247 7188
rect 10292 7187 10339 7188
rect 10305 7182 10339 7187
rect 10073 7161 10247 7164
rect 10066 7158 10247 7161
rect 10275 7181 10339 7182
rect 9869 7138 9888 7140
rect 9903 7138 9937 7140
rect 9869 7122 9949 7138
rect 9869 7116 9888 7122
rect 9585 7090 9688 7100
rect 9539 7088 9688 7090
rect 9709 7088 9744 7100
rect 9378 7086 9540 7088
rect 9390 7066 9409 7086
rect 9424 7084 9454 7086
rect 9273 7058 9314 7066
rect 9396 7062 9409 7066
rect 9461 7070 9540 7086
rect 9572 7086 9744 7088
rect 9572 7070 9651 7086
rect 9658 7084 9688 7086
rect 9236 7048 9265 7058
rect 9279 7048 9308 7058
rect 9323 7048 9353 7062
rect 9396 7048 9439 7062
rect 9461 7058 9651 7070
rect 9716 7066 9722 7086
rect 9446 7048 9476 7058
rect 9477 7048 9635 7058
rect 9639 7048 9669 7058
rect 9673 7048 9703 7062
rect 9731 7048 9744 7086
rect 9816 7100 9845 7116
rect 9859 7100 9888 7116
rect 9903 7106 9933 7122
rect 9961 7100 9967 7148
rect 9970 7142 9989 7148
rect 10004 7142 10034 7150
rect 9970 7134 10034 7142
rect 9970 7118 10050 7134
rect 10066 7127 10128 7158
rect 10144 7127 10206 7158
rect 10275 7156 10324 7181
rect 10339 7156 10369 7172
rect 10238 7142 10268 7150
rect 10275 7148 10385 7156
rect 10238 7134 10283 7142
rect 9970 7116 9989 7118
rect 10004 7116 10050 7118
rect 9970 7100 10050 7116
rect 10077 7114 10112 7127
rect 10153 7124 10190 7127
rect 10153 7122 10195 7124
rect 10082 7111 10112 7114
rect 10091 7107 10098 7111
rect 10098 7106 10099 7107
rect 10057 7100 10067 7106
rect 9816 7092 9851 7100
rect 9816 7066 9817 7092
rect 9824 7066 9851 7092
rect 9759 7048 9789 7062
rect 9816 7058 9851 7066
rect 9853 7092 9894 7100
rect 9853 7066 9868 7092
rect 9875 7066 9894 7092
rect 9958 7088 9989 7100
rect 10004 7088 10107 7100
rect 10119 7090 10145 7116
rect 10160 7111 10190 7122
rect 10222 7118 10284 7134
rect 10222 7116 10268 7118
rect 10222 7100 10284 7116
rect 10296 7100 10302 7148
rect 10305 7140 10385 7148
rect 10305 7138 10324 7140
rect 10339 7138 10373 7140
rect 10305 7122 10385 7138
rect 10305 7100 10324 7122
rect 10339 7106 10369 7122
rect 10397 7116 10403 7190
rect 10406 7116 10425 7260
rect 10440 7116 10446 7260
rect 10455 7190 10468 7260
rect 10520 7256 10542 7260
rect 10513 7234 10542 7248
rect 10595 7234 10611 7248
rect 10649 7244 10655 7246
rect 10662 7244 10770 7260
rect 10777 7244 10783 7246
rect 10791 7244 10806 7260
rect 10872 7254 10891 7257
rect 10513 7232 10611 7234
rect 10638 7232 10806 7244
rect 10821 7234 10837 7248
rect 10872 7235 10894 7254
rect 10904 7248 10920 7249
rect 10903 7246 10920 7248
rect 10904 7241 10920 7246
rect 10894 7234 10900 7235
rect 10903 7234 10932 7241
rect 10821 7233 10932 7234
rect 10821 7232 10938 7233
rect 10497 7224 10548 7232
rect 10595 7224 10629 7232
rect 10497 7212 10522 7224
rect 10529 7212 10548 7224
rect 10602 7222 10629 7224
rect 10638 7222 10859 7232
rect 10894 7229 10900 7232
rect 10602 7218 10859 7222
rect 10497 7204 10548 7212
rect 10595 7204 10859 7218
rect 10903 7224 10938 7232
rect 10449 7156 10468 7190
rect 10513 7196 10542 7204
rect 10513 7190 10530 7196
rect 10513 7188 10547 7190
rect 10595 7188 10611 7204
rect 10612 7194 10820 7204
rect 10821 7194 10837 7204
rect 10885 7200 10900 7215
rect 10903 7212 10904 7224
rect 10911 7212 10938 7224
rect 10903 7204 10938 7212
rect 10903 7203 10932 7204
rect 10623 7190 10837 7194
rect 10638 7188 10837 7190
rect 10872 7190 10885 7200
rect 10903 7190 10920 7203
rect 10872 7188 10920 7190
rect 10514 7184 10547 7188
rect 10510 7182 10547 7184
rect 10510 7181 10577 7182
rect 10510 7176 10541 7181
rect 10547 7176 10577 7181
rect 10510 7172 10577 7176
rect 10483 7169 10577 7172
rect 10483 7162 10532 7169
rect 10483 7156 10513 7162
rect 10532 7157 10537 7162
rect 10449 7140 10529 7156
rect 10541 7148 10577 7169
rect 10638 7164 10827 7188
rect 10872 7187 10919 7188
rect 10885 7182 10919 7187
rect 10653 7161 10827 7164
rect 10646 7158 10827 7161
rect 10855 7181 10919 7182
rect 10449 7138 10468 7140
rect 10483 7138 10517 7140
rect 10449 7122 10529 7138
rect 10449 7116 10468 7122
rect 10165 7090 10268 7100
rect 10119 7088 10268 7090
rect 10289 7088 10324 7100
rect 9958 7086 10120 7088
rect 9970 7066 9989 7086
rect 10004 7084 10034 7086
rect 9853 7058 9894 7066
rect 9976 7062 9989 7066
rect 10041 7070 10120 7086
rect 10152 7086 10324 7088
rect 10152 7070 10231 7086
rect 10238 7084 10268 7086
rect 9816 7048 9845 7058
rect 9859 7048 9888 7058
rect 9903 7048 9933 7062
rect 9976 7048 10019 7062
rect 10041 7058 10231 7070
rect 10296 7066 10302 7086
rect 10026 7048 10056 7058
rect 10057 7048 10215 7058
rect 10219 7048 10249 7058
rect 10253 7048 10283 7062
rect 10311 7048 10324 7086
rect 10396 7100 10425 7116
rect 10439 7100 10468 7116
rect 10483 7106 10513 7122
rect 10541 7100 10547 7148
rect 10550 7142 10569 7148
rect 10584 7142 10614 7150
rect 10550 7134 10614 7142
rect 10550 7118 10630 7134
rect 10646 7127 10708 7158
rect 10724 7127 10786 7158
rect 10855 7156 10904 7181
rect 10919 7156 10949 7172
rect 10818 7142 10848 7150
rect 10855 7148 10965 7156
rect 10818 7134 10863 7142
rect 10550 7116 10569 7118
rect 10584 7116 10630 7118
rect 10550 7100 10630 7116
rect 10657 7114 10692 7127
rect 10733 7124 10770 7127
rect 10733 7122 10775 7124
rect 10662 7111 10692 7114
rect 10671 7107 10678 7111
rect 10678 7106 10679 7107
rect 10637 7100 10647 7106
rect 10396 7092 10431 7100
rect 10396 7066 10397 7092
rect 10404 7066 10431 7092
rect 10339 7048 10369 7062
rect 10396 7058 10431 7066
rect 10433 7092 10474 7100
rect 10433 7066 10448 7092
rect 10455 7066 10474 7092
rect 10538 7088 10569 7100
rect 10584 7088 10687 7100
rect 10699 7090 10725 7116
rect 10740 7111 10770 7122
rect 10802 7118 10864 7134
rect 10802 7116 10848 7118
rect 10802 7100 10864 7116
rect 10876 7100 10882 7148
rect 10885 7140 10965 7148
rect 10885 7138 10904 7140
rect 10919 7138 10953 7140
rect 10885 7122 10965 7138
rect 10885 7100 10904 7122
rect 10919 7106 10949 7122
rect 10977 7116 10983 7190
rect 10986 7116 11005 7260
rect 11020 7116 11026 7260
rect 11035 7190 11048 7260
rect 11100 7256 11122 7260
rect 11093 7234 11122 7248
rect 11175 7234 11191 7248
rect 11229 7244 11235 7246
rect 11242 7244 11350 7260
rect 11357 7244 11363 7246
rect 11371 7244 11386 7260
rect 11452 7254 11471 7257
rect 11093 7232 11191 7234
rect 11218 7232 11386 7244
rect 11401 7234 11417 7248
rect 11452 7235 11474 7254
rect 11484 7248 11500 7249
rect 11483 7246 11500 7248
rect 11484 7241 11500 7246
rect 11474 7234 11480 7235
rect 11483 7234 11512 7241
rect 11401 7233 11512 7234
rect 11401 7232 11518 7233
rect 11077 7224 11128 7232
rect 11175 7224 11209 7232
rect 11077 7212 11102 7224
rect 11109 7212 11128 7224
rect 11182 7222 11209 7224
rect 11218 7222 11439 7232
rect 11474 7229 11480 7232
rect 11182 7218 11439 7222
rect 11077 7204 11128 7212
rect 11175 7204 11439 7218
rect 11483 7224 11518 7232
rect 11029 7156 11048 7190
rect 11093 7196 11122 7204
rect 11093 7190 11110 7196
rect 11093 7188 11127 7190
rect 11175 7188 11191 7204
rect 11192 7194 11400 7204
rect 11401 7194 11417 7204
rect 11465 7200 11480 7215
rect 11483 7212 11484 7224
rect 11491 7212 11518 7224
rect 11483 7204 11518 7212
rect 11483 7203 11512 7204
rect 11203 7190 11417 7194
rect 11218 7188 11417 7190
rect 11452 7190 11465 7200
rect 11483 7190 11500 7203
rect 11452 7188 11500 7190
rect 11094 7184 11127 7188
rect 11090 7182 11127 7184
rect 11090 7181 11157 7182
rect 11090 7176 11121 7181
rect 11127 7176 11157 7181
rect 11090 7172 11157 7176
rect 11063 7169 11157 7172
rect 11063 7162 11112 7169
rect 11063 7156 11093 7162
rect 11112 7157 11117 7162
rect 11029 7140 11109 7156
rect 11121 7148 11157 7169
rect 11218 7164 11407 7188
rect 11452 7187 11499 7188
rect 11465 7182 11499 7187
rect 11233 7161 11407 7164
rect 11226 7158 11407 7161
rect 11435 7181 11499 7182
rect 11029 7138 11048 7140
rect 11063 7138 11097 7140
rect 11029 7122 11109 7138
rect 11029 7116 11048 7122
rect 10745 7090 10848 7100
rect 10699 7088 10848 7090
rect 10869 7088 10904 7100
rect 10538 7086 10700 7088
rect 10550 7066 10569 7086
rect 10584 7084 10614 7086
rect 10433 7058 10474 7066
rect 10556 7062 10569 7066
rect 10621 7070 10700 7086
rect 10732 7086 10904 7088
rect 10732 7070 10811 7086
rect 10818 7084 10848 7086
rect 10396 7048 10425 7058
rect 10439 7048 10468 7058
rect 10483 7048 10513 7062
rect 10556 7048 10599 7062
rect 10621 7058 10811 7070
rect 10876 7066 10882 7086
rect 10606 7048 10636 7058
rect 10637 7048 10795 7058
rect 10799 7048 10829 7058
rect 10833 7048 10863 7062
rect 10891 7048 10904 7086
rect 10976 7100 11005 7116
rect 11019 7100 11048 7116
rect 11063 7106 11093 7122
rect 11121 7100 11127 7148
rect 11130 7142 11149 7148
rect 11164 7142 11194 7150
rect 11130 7134 11194 7142
rect 11130 7118 11210 7134
rect 11226 7127 11288 7158
rect 11304 7127 11366 7158
rect 11435 7156 11484 7181
rect 11499 7156 11529 7172
rect 11398 7142 11428 7150
rect 11435 7148 11545 7156
rect 11398 7134 11443 7142
rect 11130 7116 11149 7118
rect 11164 7116 11210 7118
rect 11130 7100 11210 7116
rect 11237 7114 11272 7127
rect 11313 7124 11350 7127
rect 11313 7122 11355 7124
rect 11242 7111 11272 7114
rect 11251 7107 11258 7111
rect 11258 7106 11259 7107
rect 11217 7100 11227 7106
rect 10976 7092 11011 7100
rect 10976 7066 10977 7092
rect 10984 7066 11011 7092
rect 10919 7048 10949 7062
rect 10976 7058 11011 7066
rect 11013 7092 11054 7100
rect 11013 7066 11028 7092
rect 11035 7066 11054 7092
rect 11118 7088 11149 7100
rect 11164 7088 11267 7100
rect 11279 7090 11305 7116
rect 11320 7111 11350 7122
rect 11382 7118 11444 7134
rect 11382 7116 11428 7118
rect 11382 7100 11444 7116
rect 11456 7100 11462 7148
rect 11465 7140 11545 7148
rect 11465 7138 11484 7140
rect 11499 7138 11533 7140
rect 11465 7122 11545 7138
rect 11465 7100 11484 7122
rect 11499 7106 11529 7122
rect 11557 7116 11563 7190
rect 11566 7116 11585 7260
rect 11600 7116 11606 7260
rect 11615 7190 11628 7260
rect 11680 7256 11702 7260
rect 11673 7234 11702 7248
rect 11755 7234 11771 7248
rect 11809 7244 11815 7246
rect 11822 7244 11930 7260
rect 11937 7244 11943 7246
rect 11951 7244 11966 7260
rect 12032 7254 12051 7257
rect 11673 7232 11771 7234
rect 11798 7232 11966 7244
rect 11981 7234 11997 7248
rect 12032 7235 12054 7254
rect 12064 7248 12080 7249
rect 12063 7246 12080 7248
rect 12064 7241 12080 7246
rect 12054 7234 12060 7235
rect 12063 7234 12092 7241
rect 11981 7233 12092 7234
rect 11981 7232 12098 7233
rect 11657 7224 11708 7232
rect 11755 7224 11789 7232
rect 11657 7212 11682 7224
rect 11689 7212 11708 7224
rect 11762 7222 11789 7224
rect 11798 7222 12019 7232
rect 12054 7229 12060 7232
rect 11762 7218 12019 7222
rect 11657 7204 11708 7212
rect 11755 7204 12019 7218
rect 12063 7224 12098 7232
rect 11609 7156 11628 7190
rect 11673 7196 11702 7204
rect 11673 7190 11690 7196
rect 11673 7188 11707 7190
rect 11755 7188 11771 7204
rect 11772 7194 11980 7204
rect 11981 7194 11997 7204
rect 12045 7200 12060 7215
rect 12063 7212 12064 7224
rect 12071 7212 12098 7224
rect 12063 7204 12098 7212
rect 12063 7203 12092 7204
rect 11783 7190 11997 7194
rect 11798 7188 11997 7190
rect 12032 7190 12045 7200
rect 12063 7190 12080 7203
rect 12032 7188 12080 7190
rect 11674 7184 11707 7188
rect 11670 7182 11707 7184
rect 11670 7181 11737 7182
rect 11670 7176 11701 7181
rect 11707 7176 11737 7181
rect 11670 7172 11737 7176
rect 11643 7169 11737 7172
rect 11643 7162 11692 7169
rect 11643 7156 11673 7162
rect 11692 7157 11697 7162
rect 11609 7140 11689 7156
rect 11701 7148 11737 7169
rect 11798 7164 11987 7188
rect 12032 7187 12079 7188
rect 12045 7182 12079 7187
rect 11813 7161 11987 7164
rect 11806 7158 11987 7161
rect 12015 7181 12079 7182
rect 11609 7138 11628 7140
rect 11643 7138 11677 7140
rect 11609 7122 11689 7138
rect 11609 7116 11628 7122
rect 11325 7090 11428 7100
rect 11279 7088 11428 7090
rect 11449 7088 11484 7100
rect 11118 7086 11280 7088
rect 11130 7066 11149 7086
rect 11164 7084 11194 7086
rect 11013 7058 11054 7066
rect 11136 7062 11149 7066
rect 11201 7070 11280 7086
rect 11312 7086 11484 7088
rect 11312 7070 11391 7086
rect 11398 7084 11428 7086
rect 10976 7048 11005 7058
rect 11019 7048 11048 7058
rect 11063 7048 11093 7062
rect 11136 7048 11179 7062
rect 11201 7058 11391 7070
rect 11456 7066 11462 7086
rect 11186 7048 11216 7058
rect 11217 7048 11375 7058
rect 11379 7048 11409 7058
rect 11413 7048 11443 7062
rect 11471 7048 11484 7086
rect 11556 7100 11585 7116
rect 11599 7100 11628 7116
rect 11643 7106 11673 7122
rect 11701 7100 11707 7148
rect 11710 7142 11729 7148
rect 11744 7142 11774 7150
rect 11710 7134 11774 7142
rect 11710 7118 11790 7134
rect 11806 7127 11868 7158
rect 11884 7127 11946 7158
rect 12015 7156 12064 7181
rect 12079 7156 12109 7172
rect 11978 7142 12008 7150
rect 12015 7148 12125 7156
rect 11978 7134 12023 7142
rect 11710 7116 11729 7118
rect 11744 7116 11790 7118
rect 11710 7100 11790 7116
rect 11817 7114 11852 7127
rect 11893 7124 11930 7127
rect 11893 7122 11935 7124
rect 11822 7111 11852 7114
rect 11831 7107 11838 7111
rect 11838 7106 11839 7107
rect 11797 7100 11807 7106
rect 11556 7092 11591 7100
rect 11556 7066 11557 7092
rect 11564 7066 11591 7092
rect 11499 7048 11529 7062
rect 11556 7058 11591 7066
rect 11593 7092 11634 7100
rect 11593 7066 11608 7092
rect 11615 7066 11634 7092
rect 11698 7088 11729 7100
rect 11744 7088 11847 7100
rect 11859 7090 11885 7116
rect 11900 7111 11930 7122
rect 11962 7118 12024 7134
rect 11962 7116 12008 7118
rect 11962 7100 12024 7116
rect 12036 7100 12042 7148
rect 12045 7140 12125 7148
rect 12045 7138 12064 7140
rect 12079 7138 12113 7140
rect 12045 7122 12125 7138
rect 12045 7100 12064 7122
rect 12079 7106 12109 7122
rect 12137 7116 12143 7190
rect 12146 7116 12165 7260
rect 12180 7116 12186 7260
rect 12195 7190 12208 7260
rect 12260 7256 12282 7260
rect 12253 7234 12282 7248
rect 12335 7234 12351 7248
rect 12389 7244 12395 7246
rect 12402 7244 12510 7260
rect 12517 7244 12523 7246
rect 12531 7244 12546 7260
rect 12612 7254 12631 7257
rect 12253 7232 12351 7234
rect 12378 7232 12546 7244
rect 12561 7234 12577 7248
rect 12612 7235 12634 7254
rect 12644 7248 12660 7249
rect 12643 7246 12660 7248
rect 12644 7241 12660 7246
rect 12634 7234 12640 7235
rect 12643 7234 12672 7241
rect 12561 7233 12672 7234
rect 12561 7232 12678 7233
rect 12237 7224 12288 7232
rect 12335 7224 12369 7232
rect 12237 7212 12262 7224
rect 12269 7212 12288 7224
rect 12342 7222 12369 7224
rect 12378 7222 12599 7232
rect 12634 7229 12640 7232
rect 12342 7218 12599 7222
rect 12237 7204 12288 7212
rect 12335 7204 12599 7218
rect 12643 7224 12678 7232
rect 12189 7156 12208 7190
rect 12253 7196 12282 7204
rect 12253 7190 12270 7196
rect 12253 7188 12287 7190
rect 12335 7188 12351 7204
rect 12352 7194 12560 7204
rect 12561 7194 12577 7204
rect 12625 7200 12640 7215
rect 12643 7212 12644 7224
rect 12651 7212 12678 7224
rect 12643 7204 12678 7212
rect 12643 7203 12672 7204
rect 12363 7190 12577 7194
rect 12378 7188 12577 7190
rect 12612 7190 12625 7200
rect 12643 7190 12660 7203
rect 12612 7188 12660 7190
rect 12254 7184 12287 7188
rect 12250 7182 12287 7184
rect 12250 7181 12317 7182
rect 12250 7176 12281 7181
rect 12287 7176 12317 7181
rect 12250 7172 12317 7176
rect 12223 7169 12317 7172
rect 12223 7162 12272 7169
rect 12223 7156 12253 7162
rect 12272 7157 12277 7162
rect 12189 7140 12269 7156
rect 12281 7148 12317 7169
rect 12378 7164 12567 7188
rect 12612 7187 12659 7188
rect 12625 7182 12659 7187
rect 12393 7161 12567 7164
rect 12386 7158 12567 7161
rect 12595 7181 12659 7182
rect 12189 7138 12208 7140
rect 12223 7138 12257 7140
rect 12189 7122 12269 7138
rect 12189 7116 12208 7122
rect 11905 7090 12008 7100
rect 11859 7088 12008 7090
rect 12029 7088 12064 7100
rect 11698 7086 11860 7088
rect 11710 7066 11729 7086
rect 11744 7084 11774 7086
rect 11593 7058 11634 7066
rect 11716 7062 11729 7066
rect 11781 7070 11860 7086
rect 11892 7086 12064 7088
rect 11892 7070 11971 7086
rect 11978 7084 12008 7086
rect 11556 7048 11585 7058
rect 11599 7048 11628 7058
rect 11643 7048 11673 7062
rect 11716 7048 11759 7062
rect 11781 7058 11971 7070
rect 12036 7066 12042 7086
rect 11766 7048 11796 7058
rect 11797 7048 11955 7058
rect 11959 7048 11989 7058
rect 11993 7048 12023 7062
rect 12051 7048 12064 7086
rect 12136 7100 12165 7116
rect 12179 7100 12208 7116
rect 12223 7106 12253 7122
rect 12281 7100 12287 7148
rect 12290 7142 12309 7148
rect 12324 7142 12354 7150
rect 12290 7134 12354 7142
rect 12290 7118 12370 7134
rect 12386 7127 12448 7158
rect 12464 7127 12526 7158
rect 12595 7156 12644 7181
rect 12659 7156 12689 7172
rect 12558 7142 12588 7150
rect 12595 7148 12705 7156
rect 12558 7134 12603 7142
rect 12290 7116 12309 7118
rect 12324 7116 12370 7118
rect 12290 7100 12370 7116
rect 12397 7114 12432 7127
rect 12473 7124 12510 7127
rect 12473 7122 12515 7124
rect 12402 7111 12432 7114
rect 12411 7107 12418 7111
rect 12418 7106 12419 7107
rect 12377 7100 12387 7106
rect 12136 7092 12171 7100
rect 12136 7066 12137 7092
rect 12144 7066 12171 7092
rect 12079 7048 12109 7062
rect 12136 7058 12171 7066
rect 12173 7092 12214 7100
rect 12173 7066 12188 7092
rect 12195 7066 12214 7092
rect 12278 7088 12309 7100
rect 12324 7088 12427 7100
rect 12439 7090 12465 7116
rect 12480 7111 12510 7122
rect 12542 7118 12604 7134
rect 12542 7116 12588 7118
rect 12542 7100 12604 7116
rect 12616 7100 12622 7148
rect 12625 7140 12705 7148
rect 12625 7138 12644 7140
rect 12659 7138 12693 7140
rect 12625 7122 12705 7138
rect 12625 7100 12644 7122
rect 12659 7106 12689 7122
rect 12717 7116 12723 7190
rect 12726 7116 12745 7260
rect 12760 7116 12766 7260
rect 12775 7190 12788 7260
rect 12840 7256 12862 7260
rect 12833 7234 12862 7248
rect 12915 7234 12931 7248
rect 12969 7244 12975 7246
rect 12982 7244 13090 7260
rect 13097 7244 13103 7246
rect 13111 7244 13126 7260
rect 13192 7254 13211 7257
rect 12833 7232 12931 7234
rect 12958 7232 13126 7244
rect 13141 7234 13157 7248
rect 13192 7235 13214 7254
rect 13224 7248 13240 7249
rect 13223 7246 13240 7248
rect 13224 7241 13240 7246
rect 13214 7234 13220 7235
rect 13223 7234 13252 7241
rect 13141 7233 13252 7234
rect 13141 7232 13258 7233
rect 12817 7224 12868 7232
rect 12915 7224 12949 7232
rect 12817 7212 12842 7224
rect 12849 7212 12868 7224
rect 12922 7222 12949 7224
rect 12958 7222 13179 7232
rect 13214 7229 13220 7232
rect 12922 7218 13179 7222
rect 12817 7204 12868 7212
rect 12915 7204 13179 7218
rect 13223 7224 13258 7232
rect 12769 7156 12788 7190
rect 12833 7196 12862 7204
rect 12833 7190 12850 7196
rect 12833 7188 12867 7190
rect 12915 7188 12931 7204
rect 12932 7194 13140 7204
rect 13141 7194 13157 7204
rect 13205 7200 13220 7215
rect 13223 7212 13224 7224
rect 13231 7212 13258 7224
rect 13223 7204 13258 7212
rect 13223 7203 13252 7204
rect 12943 7190 13157 7194
rect 12958 7188 13157 7190
rect 13192 7190 13205 7200
rect 13223 7190 13240 7203
rect 13192 7188 13240 7190
rect 12834 7184 12867 7188
rect 12830 7182 12867 7184
rect 12830 7181 12897 7182
rect 12830 7176 12861 7181
rect 12867 7176 12897 7181
rect 12830 7172 12897 7176
rect 12803 7169 12897 7172
rect 12803 7162 12852 7169
rect 12803 7156 12833 7162
rect 12852 7157 12857 7162
rect 12769 7140 12849 7156
rect 12861 7148 12897 7169
rect 12958 7164 13147 7188
rect 13192 7187 13239 7188
rect 13205 7182 13239 7187
rect 12973 7161 13147 7164
rect 12966 7158 13147 7161
rect 13175 7181 13239 7182
rect 12769 7138 12788 7140
rect 12803 7138 12837 7140
rect 12769 7122 12849 7138
rect 12769 7116 12788 7122
rect 12485 7090 12588 7100
rect 12439 7088 12588 7090
rect 12609 7088 12644 7100
rect 12278 7086 12440 7088
rect 12290 7066 12309 7086
rect 12324 7084 12354 7086
rect 12173 7058 12214 7066
rect 12296 7062 12309 7066
rect 12361 7070 12440 7086
rect 12472 7086 12644 7088
rect 12472 7070 12551 7086
rect 12558 7084 12588 7086
rect 12136 7048 12165 7058
rect 12179 7048 12208 7058
rect 12223 7048 12253 7062
rect 12296 7048 12339 7062
rect 12361 7058 12551 7070
rect 12616 7066 12622 7086
rect 12346 7048 12376 7058
rect 12377 7048 12535 7058
rect 12539 7048 12569 7058
rect 12573 7048 12603 7062
rect 12631 7048 12644 7086
rect 12716 7100 12745 7116
rect 12759 7100 12788 7116
rect 12803 7106 12833 7122
rect 12861 7100 12867 7148
rect 12870 7142 12889 7148
rect 12904 7142 12934 7150
rect 12870 7134 12934 7142
rect 12870 7118 12950 7134
rect 12966 7127 13028 7158
rect 13044 7127 13106 7158
rect 13175 7156 13224 7181
rect 13239 7156 13269 7172
rect 13138 7142 13168 7150
rect 13175 7148 13285 7156
rect 13138 7134 13183 7142
rect 12870 7116 12889 7118
rect 12904 7116 12950 7118
rect 12870 7100 12950 7116
rect 12977 7114 13012 7127
rect 13053 7124 13090 7127
rect 13053 7122 13095 7124
rect 12982 7111 13012 7114
rect 12991 7107 12998 7111
rect 12998 7106 12999 7107
rect 12957 7100 12967 7106
rect 12716 7092 12751 7100
rect 12716 7066 12717 7092
rect 12724 7066 12751 7092
rect 12659 7048 12689 7062
rect 12716 7058 12751 7066
rect 12753 7092 12794 7100
rect 12753 7066 12768 7092
rect 12775 7066 12794 7092
rect 12858 7088 12889 7100
rect 12904 7088 13007 7100
rect 13019 7090 13045 7116
rect 13060 7111 13090 7122
rect 13122 7118 13184 7134
rect 13122 7116 13168 7118
rect 13122 7100 13184 7116
rect 13196 7100 13202 7148
rect 13205 7140 13285 7148
rect 13205 7138 13224 7140
rect 13239 7138 13273 7140
rect 13205 7122 13285 7138
rect 13205 7100 13224 7122
rect 13239 7106 13269 7122
rect 13297 7116 13303 7190
rect 13306 7116 13325 7260
rect 13340 7116 13346 7260
rect 13355 7190 13368 7260
rect 13420 7256 13442 7260
rect 13413 7234 13442 7248
rect 13495 7234 13511 7248
rect 13549 7244 13555 7246
rect 13562 7244 13670 7260
rect 13677 7244 13683 7246
rect 13691 7244 13706 7260
rect 13772 7254 13791 7257
rect 13413 7232 13511 7234
rect 13538 7232 13706 7244
rect 13721 7234 13737 7248
rect 13772 7235 13794 7254
rect 13804 7248 13820 7249
rect 13803 7246 13820 7248
rect 13804 7241 13820 7246
rect 13794 7234 13800 7235
rect 13803 7234 13832 7241
rect 13721 7233 13832 7234
rect 13721 7232 13838 7233
rect 13397 7224 13448 7232
rect 13495 7224 13529 7232
rect 13397 7212 13422 7224
rect 13429 7212 13448 7224
rect 13502 7222 13529 7224
rect 13538 7222 13759 7232
rect 13794 7229 13800 7232
rect 13502 7218 13759 7222
rect 13397 7204 13448 7212
rect 13495 7204 13759 7218
rect 13803 7224 13838 7232
rect 13349 7156 13368 7190
rect 13413 7196 13442 7204
rect 13413 7190 13430 7196
rect 13413 7188 13447 7190
rect 13495 7188 13511 7204
rect 13512 7194 13720 7204
rect 13721 7194 13737 7204
rect 13785 7200 13800 7215
rect 13803 7212 13804 7224
rect 13811 7212 13838 7224
rect 13803 7204 13838 7212
rect 13803 7203 13832 7204
rect 13523 7190 13737 7194
rect 13538 7188 13737 7190
rect 13772 7190 13785 7200
rect 13803 7190 13820 7203
rect 13772 7188 13820 7190
rect 13414 7184 13447 7188
rect 13410 7182 13447 7184
rect 13410 7181 13477 7182
rect 13410 7176 13441 7181
rect 13447 7176 13477 7181
rect 13410 7172 13477 7176
rect 13383 7169 13477 7172
rect 13383 7162 13432 7169
rect 13383 7156 13413 7162
rect 13432 7157 13437 7162
rect 13349 7140 13429 7156
rect 13441 7148 13477 7169
rect 13538 7164 13727 7188
rect 13772 7187 13819 7188
rect 13785 7182 13819 7187
rect 13553 7161 13727 7164
rect 13546 7158 13727 7161
rect 13755 7181 13819 7182
rect 13349 7138 13368 7140
rect 13383 7138 13417 7140
rect 13349 7122 13429 7138
rect 13349 7116 13368 7122
rect 13065 7090 13168 7100
rect 13019 7088 13168 7090
rect 13189 7088 13224 7100
rect 12858 7086 13020 7088
rect 12870 7066 12889 7086
rect 12904 7084 12934 7086
rect 12753 7058 12794 7066
rect 12876 7062 12889 7066
rect 12941 7070 13020 7086
rect 13052 7086 13224 7088
rect 13052 7070 13131 7086
rect 13138 7084 13168 7086
rect 12716 7048 12745 7058
rect 12759 7048 12788 7058
rect 12803 7048 12833 7062
rect 12876 7048 12919 7062
rect 12941 7058 13131 7070
rect 13196 7066 13202 7086
rect 12926 7048 12956 7058
rect 12957 7048 13115 7058
rect 13119 7048 13149 7058
rect 13153 7048 13183 7062
rect 13211 7048 13224 7086
rect 13296 7100 13325 7116
rect 13339 7100 13368 7116
rect 13383 7106 13413 7122
rect 13441 7100 13447 7148
rect 13450 7142 13469 7148
rect 13484 7142 13514 7150
rect 13450 7134 13514 7142
rect 13450 7118 13530 7134
rect 13546 7127 13608 7158
rect 13624 7127 13686 7158
rect 13755 7156 13804 7181
rect 13819 7156 13849 7172
rect 13718 7142 13748 7150
rect 13755 7148 13865 7156
rect 13718 7134 13763 7142
rect 13450 7116 13469 7118
rect 13484 7116 13530 7118
rect 13450 7100 13530 7116
rect 13557 7114 13592 7127
rect 13633 7124 13670 7127
rect 13633 7122 13675 7124
rect 13562 7111 13592 7114
rect 13571 7107 13578 7111
rect 13578 7106 13579 7107
rect 13537 7100 13547 7106
rect 13296 7092 13331 7100
rect 13296 7066 13297 7092
rect 13304 7066 13331 7092
rect 13239 7048 13269 7062
rect 13296 7058 13331 7066
rect 13333 7092 13374 7100
rect 13333 7066 13348 7092
rect 13355 7066 13374 7092
rect 13438 7088 13469 7100
rect 13484 7088 13587 7100
rect 13599 7090 13625 7116
rect 13640 7111 13670 7122
rect 13702 7118 13764 7134
rect 13702 7116 13748 7118
rect 13702 7100 13764 7116
rect 13776 7100 13782 7148
rect 13785 7140 13865 7148
rect 13785 7138 13804 7140
rect 13819 7138 13853 7140
rect 13785 7122 13865 7138
rect 13785 7100 13804 7122
rect 13819 7106 13849 7122
rect 13877 7116 13883 7190
rect 13886 7116 13905 7260
rect 13920 7116 13926 7260
rect 13935 7190 13948 7260
rect 14000 7256 14022 7260
rect 13993 7234 14022 7248
rect 14075 7234 14091 7248
rect 14129 7244 14135 7246
rect 14142 7244 14250 7260
rect 14257 7244 14263 7246
rect 14271 7244 14286 7260
rect 14352 7254 14371 7257
rect 13993 7232 14091 7234
rect 14118 7232 14286 7244
rect 14301 7234 14317 7248
rect 14352 7235 14374 7254
rect 14384 7248 14400 7249
rect 14383 7246 14400 7248
rect 14384 7241 14400 7246
rect 14374 7234 14380 7235
rect 14383 7234 14412 7241
rect 14301 7233 14412 7234
rect 14301 7232 14418 7233
rect 13977 7224 14028 7232
rect 14075 7224 14109 7232
rect 13977 7212 14002 7224
rect 14009 7212 14028 7224
rect 14082 7222 14109 7224
rect 14118 7222 14339 7232
rect 14374 7229 14380 7232
rect 14082 7218 14339 7222
rect 13977 7204 14028 7212
rect 14075 7204 14339 7218
rect 14383 7224 14418 7232
rect 13929 7156 13948 7190
rect 13993 7196 14022 7204
rect 13993 7190 14010 7196
rect 13993 7188 14027 7190
rect 14075 7188 14091 7204
rect 14092 7194 14300 7204
rect 14301 7194 14317 7204
rect 14365 7200 14380 7215
rect 14383 7212 14384 7224
rect 14391 7212 14418 7224
rect 14383 7204 14418 7212
rect 14383 7203 14412 7204
rect 14103 7190 14317 7194
rect 14118 7188 14317 7190
rect 14352 7190 14365 7200
rect 14383 7190 14400 7203
rect 14352 7188 14400 7190
rect 13994 7184 14027 7188
rect 13990 7182 14027 7184
rect 13990 7181 14057 7182
rect 13990 7176 14021 7181
rect 14027 7176 14057 7181
rect 13990 7172 14057 7176
rect 13963 7169 14057 7172
rect 13963 7162 14012 7169
rect 13963 7156 13993 7162
rect 14012 7157 14017 7162
rect 13929 7140 14009 7156
rect 14021 7148 14057 7169
rect 14118 7164 14307 7188
rect 14352 7187 14399 7188
rect 14365 7182 14399 7187
rect 14133 7161 14307 7164
rect 14126 7158 14307 7161
rect 14335 7181 14399 7182
rect 13929 7138 13948 7140
rect 13963 7138 13997 7140
rect 13929 7122 14009 7138
rect 13929 7116 13948 7122
rect 13645 7090 13748 7100
rect 13599 7088 13748 7090
rect 13769 7088 13804 7100
rect 13438 7086 13600 7088
rect 13450 7066 13469 7086
rect 13484 7084 13514 7086
rect 13333 7058 13374 7066
rect 13456 7062 13469 7066
rect 13521 7070 13600 7086
rect 13632 7086 13804 7088
rect 13632 7070 13711 7086
rect 13718 7084 13748 7086
rect 13296 7048 13325 7058
rect 13339 7048 13368 7058
rect 13383 7048 13413 7062
rect 13456 7048 13499 7062
rect 13521 7058 13711 7070
rect 13776 7066 13782 7086
rect 13506 7048 13536 7058
rect 13537 7048 13695 7058
rect 13699 7048 13729 7058
rect 13733 7048 13763 7062
rect 13791 7048 13804 7086
rect 13876 7100 13905 7116
rect 13919 7100 13948 7116
rect 13963 7106 13993 7122
rect 14021 7100 14027 7148
rect 14030 7142 14049 7148
rect 14064 7142 14094 7150
rect 14030 7134 14094 7142
rect 14030 7118 14110 7134
rect 14126 7127 14188 7158
rect 14204 7127 14266 7158
rect 14335 7156 14384 7181
rect 14399 7156 14429 7172
rect 14298 7142 14328 7150
rect 14335 7148 14445 7156
rect 14298 7134 14343 7142
rect 14030 7116 14049 7118
rect 14064 7116 14110 7118
rect 14030 7100 14110 7116
rect 14137 7114 14172 7127
rect 14213 7124 14250 7127
rect 14213 7122 14255 7124
rect 14142 7111 14172 7114
rect 14151 7107 14158 7111
rect 14158 7106 14159 7107
rect 14117 7100 14127 7106
rect 13876 7092 13911 7100
rect 13876 7066 13877 7092
rect 13884 7066 13911 7092
rect 13819 7048 13849 7062
rect 13876 7058 13911 7066
rect 13913 7092 13954 7100
rect 13913 7066 13928 7092
rect 13935 7066 13954 7092
rect 14018 7088 14049 7100
rect 14064 7088 14167 7100
rect 14179 7090 14205 7116
rect 14220 7111 14250 7122
rect 14282 7118 14344 7134
rect 14282 7116 14328 7118
rect 14282 7100 14344 7116
rect 14356 7100 14362 7148
rect 14365 7140 14445 7148
rect 14365 7138 14384 7140
rect 14399 7138 14433 7140
rect 14365 7122 14445 7138
rect 14365 7100 14384 7122
rect 14399 7106 14429 7122
rect 14457 7116 14463 7190
rect 14466 7116 14485 7260
rect 14500 7116 14506 7260
rect 14515 7190 14528 7260
rect 14580 7256 14602 7260
rect 14573 7234 14602 7248
rect 14655 7234 14671 7248
rect 14709 7244 14715 7246
rect 14722 7244 14830 7260
rect 14837 7244 14843 7246
rect 14851 7244 14866 7260
rect 14932 7254 14951 7257
rect 14573 7232 14671 7234
rect 14698 7232 14866 7244
rect 14881 7234 14897 7248
rect 14932 7235 14954 7254
rect 14964 7248 14980 7249
rect 14963 7246 14980 7248
rect 14964 7241 14980 7246
rect 14954 7234 14960 7235
rect 14963 7234 14992 7241
rect 14881 7233 14992 7234
rect 14881 7232 14998 7233
rect 14557 7224 14608 7232
rect 14655 7224 14689 7232
rect 14557 7212 14582 7224
rect 14589 7212 14608 7224
rect 14662 7222 14689 7224
rect 14698 7222 14919 7232
rect 14954 7229 14960 7232
rect 14662 7218 14919 7222
rect 14557 7204 14608 7212
rect 14655 7204 14919 7218
rect 14963 7224 14998 7232
rect 14509 7156 14528 7190
rect 14573 7196 14602 7204
rect 14573 7190 14590 7196
rect 14573 7188 14607 7190
rect 14655 7188 14671 7204
rect 14672 7194 14880 7204
rect 14881 7194 14897 7204
rect 14945 7200 14960 7215
rect 14963 7212 14964 7224
rect 14971 7212 14998 7224
rect 14963 7204 14998 7212
rect 14963 7203 14992 7204
rect 14683 7190 14897 7194
rect 14698 7188 14897 7190
rect 14932 7190 14945 7200
rect 14963 7190 14980 7203
rect 14932 7188 14980 7190
rect 14574 7184 14607 7188
rect 14570 7182 14607 7184
rect 14570 7181 14637 7182
rect 14570 7176 14601 7181
rect 14607 7176 14637 7181
rect 14570 7172 14637 7176
rect 14543 7169 14637 7172
rect 14543 7162 14592 7169
rect 14543 7156 14573 7162
rect 14592 7157 14597 7162
rect 14509 7140 14589 7156
rect 14601 7148 14637 7169
rect 14698 7164 14887 7188
rect 14932 7187 14979 7188
rect 14945 7182 14979 7187
rect 14713 7161 14887 7164
rect 14706 7158 14887 7161
rect 14915 7181 14979 7182
rect 14509 7138 14528 7140
rect 14543 7138 14577 7140
rect 14509 7122 14589 7138
rect 14509 7116 14528 7122
rect 14225 7090 14328 7100
rect 14179 7088 14328 7090
rect 14349 7088 14384 7100
rect 14018 7086 14180 7088
rect 14030 7066 14049 7086
rect 14064 7084 14094 7086
rect 13913 7058 13954 7066
rect 14036 7062 14049 7066
rect 14101 7070 14180 7086
rect 14212 7086 14384 7088
rect 14212 7070 14291 7086
rect 14298 7084 14328 7086
rect 13876 7048 13905 7058
rect 13919 7048 13948 7058
rect 13963 7048 13993 7062
rect 14036 7048 14079 7062
rect 14101 7058 14291 7070
rect 14356 7066 14362 7086
rect 14086 7048 14116 7058
rect 14117 7048 14275 7058
rect 14279 7048 14309 7058
rect 14313 7048 14343 7062
rect 14371 7048 14384 7086
rect 14456 7100 14485 7116
rect 14499 7100 14528 7116
rect 14543 7106 14573 7122
rect 14601 7100 14607 7148
rect 14610 7142 14629 7148
rect 14644 7142 14674 7150
rect 14610 7134 14674 7142
rect 14610 7118 14690 7134
rect 14706 7127 14768 7158
rect 14784 7127 14846 7158
rect 14915 7156 14964 7181
rect 14979 7156 15009 7172
rect 14878 7142 14908 7150
rect 14915 7148 15025 7156
rect 14878 7134 14923 7142
rect 14610 7116 14629 7118
rect 14644 7116 14690 7118
rect 14610 7100 14690 7116
rect 14717 7114 14752 7127
rect 14793 7124 14830 7127
rect 14793 7122 14835 7124
rect 14722 7111 14752 7114
rect 14731 7107 14738 7111
rect 14738 7106 14739 7107
rect 14697 7100 14707 7106
rect 14456 7092 14491 7100
rect 14456 7066 14457 7092
rect 14464 7066 14491 7092
rect 14399 7048 14429 7062
rect 14456 7058 14491 7066
rect 14493 7092 14534 7100
rect 14493 7066 14508 7092
rect 14515 7066 14534 7092
rect 14598 7088 14629 7100
rect 14644 7088 14747 7100
rect 14759 7090 14785 7116
rect 14800 7111 14830 7122
rect 14862 7118 14924 7134
rect 14862 7116 14908 7118
rect 14862 7100 14924 7116
rect 14936 7100 14942 7148
rect 14945 7140 15025 7148
rect 14945 7138 14964 7140
rect 14979 7138 15013 7140
rect 14945 7122 15025 7138
rect 14945 7100 14964 7122
rect 14979 7106 15009 7122
rect 15037 7116 15043 7190
rect 15046 7116 15065 7260
rect 15080 7116 15086 7260
rect 15095 7190 15108 7260
rect 15160 7256 15182 7260
rect 15153 7234 15182 7248
rect 15235 7234 15251 7248
rect 15289 7244 15295 7246
rect 15302 7244 15410 7260
rect 15417 7244 15423 7246
rect 15431 7244 15446 7260
rect 15512 7254 15531 7257
rect 15153 7232 15251 7234
rect 15278 7232 15446 7244
rect 15461 7234 15477 7248
rect 15512 7235 15534 7254
rect 15544 7248 15560 7249
rect 15543 7246 15560 7248
rect 15544 7241 15560 7246
rect 15534 7234 15540 7235
rect 15543 7234 15572 7241
rect 15461 7233 15572 7234
rect 15461 7232 15578 7233
rect 15137 7224 15188 7232
rect 15235 7224 15269 7232
rect 15137 7212 15162 7224
rect 15169 7212 15188 7224
rect 15242 7222 15269 7224
rect 15278 7222 15499 7232
rect 15534 7229 15540 7232
rect 15242 7218 15499 7222
rect 15137 7204 15188 7212
rect 15235 7204 15499 7218
rect 15543 7224 15578 7232
rect 15089 7156 15108 7190
rect 15153 7196 15182 7204
rect 15153 7190 15170 7196
rect 15153 7188 15187 7190
rect 15235 7188 15251 7204
rect 15252 7194 15460 7204
rect 15461 7194 15477 7204
rect 15525 7200 15540 7215
rect 15543 7212 15544 7224
rect 15551 7212 15578 7224
rect 15543 7204 15578 7212
rect 15543 7203 15572 7204
rect 15263 7190 15477 7194
rect 15278 7188 15477 7190
rect 15512 7190 15525 7200
rect 15543 7190 15560 7203
rect 15512 7188 15560 7190
rect 15154 7184 15187 7188
rect 15150 7182 15187 7184
rect 15150 7181 15217 7182
rect 15150 7176 15181 7181
rect 15187 7176 15217 7181
rect 15150 7172 15217 7176
rect 15123 7169 15217 7172
rect 15123 7162 15172 7169
rect 15123 7156 15153 7162
rect 15172 7157 15177 7162
rect 15089 7140 15169 7156
rect 15181 7148 15217 7169
rect 15278 7164 15467 7188
rect 15512 7187 15559 7188
rect 15525 7182 15559 7187
rect 15293 7161 15467 7164
rect 15286 7158 15467 7161
rect 15495 7181 15559 7182
rect 15089 7138 15108 7140
rect 15123 7138 15157 7140
rect 15089 7122 15169 7138
rect 15089 7116 15108 7122
rect 14805 7090 14908 7100
rect 14759 7088 14908 7090
rect 14929 7088 14964 7100
rect 14598 7086 14760 7088
rect 14610 7066 14629 7086
rect 14644 7084 14674 7086
rect 14493 7058 14534 7066
rect 14616 7062 14629 7066
rect 14681 7070 14760 7086
rect 14792 7086 14964 7088
rect 14792 7070 14871 7086
rect 14878 7084 14908 7086
rect 14456 7048 14485 7058
rect 14499 7048 14528 7058
rect 14543 7048 14573 7062
rect 14616 7048 14659 7062
rect 14681 7058 14871 7070
rect 14936 7066 14942 7086
rect 14666 7048 14696 7058
rect 14697 7048 14855 7058
rect 14859 7048 14889 7058
rect 14893 7048 14923 7062
rect 14951 7048 14964 7086
rect 15036 7100 15065 7116
rect 15079 7100 15108 7116
rect 15123 7106 15153 7122
rect 15181 7100 15187 7148
rect 15190 7142 15209 7148
rect 15224 7142 15254 7150
rect 15190 7134 15254 7142
rect 15190 7118 15270 7134
rect 15286 7127 15348 7158
rect 15364 7127 15426 7158
rect 15495 7156 15544 7181
rect 15559 7156 15589 7172
rect 15458 7142 15488 7150
rect 15495 7148 15605 7156
rect 15458 7134 15503 7142
rect 15190 7116 15209 7118
rect 15224 7116 15270 7118
rect 15190 7100 15270 7116
rect 15297 7114 15332 7127
rect 15373 7124 15410 7127
rect 15373 7122 15415 7124
rect 15302 7111 15332 7114
rect 15311 7107 15318 7111
rect 15318 7106 15319 7107
rect 15277 7100 15287 7106
rect 15036 7092 15071 7100
rect 15036 7066 15037 7092
rect 15044 7066 15071 7092
rect 14979 7048 15009 7062
rect 15036 7058 15071 7066
rect 15073 7092 15114 7100
rect 15073 7066 15088 7092
rect 15095 7066 15114 7092
rect 15178 7088 15209 7100
rect 15224 7088 15327 7100
rect 15339 7090 15365 7116
rect 15380 7111 15410 7122
rect 15442 7118 15504 7134
rect 15442 7116 15488 7118
rect 15442 7100 15504 7116
rect 15516 7100 15522 7148
rect 15525 7140 15605 7148
rect 15525 7138 15544 7140
rect 15559 7138 15593 7140
rect 15525 7122 15605 7138
rect 15525 7100 15544 7122
rect 15559 7106 15589 7122
rect 15617 7116 15623 7190
rect 15626 7116 15645 7260
rect 15660 7116 15666 7260
rect 15675 7190 15688 7260
rect 15740 7256 15762 7260
rect 15733 7234 15762 7248
rect 15815 7234 15831 7248
rect 15869 7244 15875 7246
rect 15882 7244 15990 7260
rect 15997 7244 16003 7246
rect 16011 7244 16026 7260
rect 16092 7254 16111 7257
rect 15733 7232 15831 7234
rect 15858 7232 16026 7244
rect 16041 7234 16057 7248
rect 16092 7235 16114 7254
rect 16124 7248 16140 7249
rect 16123 7246 16140 7248
rect 16124 7241 16140 7246
rect 16114 7234 16120 7235
rect 16123 7234 16152 7241
rect 16041 7233 16152 7234
rect 16041 7232 16158 7233
rect 15717 7224 15768 7232
rect 15815 7224 15849 7232
rect 15717 7212 15742 7224
rect 15749 7212 15768 7224
rect 15822 7222 15849 7224
rect 15858 7222 16079 7232
rect 16114 7229 16120 7232
rect 15822 7218 16079 7222
rect 15717 7204 15768 7212
rect 15815 7204 16079 7218
rect 16123 7224 16158 7232
rect 15669 7156 15688 7190
rect 15733 7196 15762 7204
rect 15733 7190 15750 7196
rect 15733 7188 15767 7190
rect 15815 7188 15831 7204
rect 15832 7194 16040 7204
rect 16041 7194 16057 7204
rect 16105 7200 16120 7215
rect 16123 7212 16124 7224
rect 16131 7212 16158 7224
rect 16123 7204 16158 7212
rect 16123 7203 16152 7204
rect 15843 7190 16057 7194
rect 15858 7188 16057 7190
rect 16092 7190 16105 7200
rect 16123 7190 16140 7203
rect 16092 7188 16140 7190
rect 15734 7184 15767 7188
rect 15730 7182 15767 7184
rect 15730 7181 15797 7182
rect 15730 7176 15761 7181
rect 15767 7176 15797 7181
rect 15730 7172 15797 7176
rect 15703 7169 15797 7172
rect 15703 7162 15752 7169
rect 15703 7156 15733 7162
rect 15752 7157 15757 7162
rect 15669 7140 15749 7156
rect 15761 7148 15797 7169
rect 15858 7164 16047 7188
rect 16092 7187 16139 7188
rect 16105 7182 16139 7187
rect 15873 7161 16047 7164
rect 15866 7158 16047 7161
rect 16075 7181 16139 7182
rect 15669 7138 15688 7140
rect 15703 7138 15737 7140
rect 15669 7122 15749 7138
rect 15669 7116 15688 7122
rect 15385 7090 15488 7100
rect 15339 7088 15488 7090
rect 15509 7088 15544 7100
rect 15178 7086 15340 7088
rect 15190 7066 15209 7086
rect 15224 7084 15254 7086
rect 15073 7058 15114 7066
rect 15196 7062 15209 7066
rect 15261 7070 15340 7086
rect 15372 7086 15544 7088
rect 15372 7070 15451 7086
rect 15458 7084 15488 7086
rect 15036 7048 15065 7058
rect 15079 7048 15108 7058
rect 15123 7048 15153 7062
rect 15196 7048 15239 7062
rect 15261 7058 15451 7070
rect 15516 7066 15522 7086
rect 15246 7048 15276 7058
rect 15277 7048 15435 7058
rect 15439 7048 15469 7058
rect 15473 7048 15503 7062
rect 15531 7048 15544 7086
rect 15616 7100 15645 7116
rect 15659 7100 15688 7116
rect 15703 7106 15733 7122
rect 15761 7100 15767 7148
rect 15770 7142 15789 7148
rect 15804 7142 15834 7150
rect 15770 7134 15834 7142
rect 15770 7118 15850 7134
rect 15866 7127 15928 7158
rect 15944 7127 16006 7158
rect 16075 7156 16124 7181
rect 16139 7156 16169 7172
rect 16038 7142 16068 7150
rect 16075 7148 16185 7156
rect 16038 7134 16083 7142
rect 15770 7116 15789 7118
rect 15804 7116 15850 7118
rect 15770 7100 15850 7116
rect 15877 7114 15912 7127
rect 15953 7124 15990 7127
rect 15953 7122 15995 7124
rect 15882 7111 15912 7114
rect 15891 7107 15898 7111
rect 15898 7106 15899 7107
rect 15857 7100 15867 7106
rect 15616 7092 15651 7100
rect 15616 7066 15617 7092
rect 15624 7066 15651 7092
rect 15559 7048 15589 7062
rect 15616 7058 15651 7066
rect 15653 7092 15694 7100
rect 15653 7066 15668 7092
rect 15675 7066 15694 7092
rect 15758 7088 15789 7100
rect 15804 7088 15907 7100
rect 15919 7090 15945 7116
rect 15960 7111 15990 7122
rect 16022 7118 16084 7134
rect 16022 7116 16068 7118
rect 16022 7100 16084 7116
rect 16096 7100 16102 7148
rect 16105 7140 16185 7148
rect 16105 7138 16124 7140
rect 16139 7138 16173 7140
rect 16105 7122 16185 7138
rect 16105 7100 16124 7122
rect 16139 7106 16169 7122
rect 16197 7116 16203 7190
rect 16206 7116 16225 7260
rect 16240 7116 16246 7260
rect 16255 7190 16268 7260
rect 16320 7256 16342 7260
rect 16313 7234 16342 7248
rect 16395 7234 16411 7248
rect 16449 7244 16455 7246
rect 16462 7244 16570 7260
rect 16577 7244 16583 7246
rect 16591 7244 16606 7260
rect 16672 7254 16691 7257
rect 16313 7232 16411 7234
rect 16438 7232 16606 7244
rect 16621 7234 16637 7248
rect 16672 7235 16694 7254
rect 16704 7248 16720 7249
rect 16703 7246 16720 7248
rect 16704 7241 16720 7246
rect 16694 7234 16700 7235
rect 16703 7234 16732 7241
rect 16621 7233 16732 7234
rect 16621 7232 16738 7233
rect 16297 7224 16348 7232
rect 16395 7224 16429 7232
rect 16297 7212 16322 7224
rect 16329 7212 16348 7224
rect 16402 7222 16429 7224
rect 16438 7222 16659 7232
rect 16694 7229 16700 7232
rect 16402 7218 16659 7222
rect 16297 7204 16348 7212
rect 16395 7204 16659 7218
rect 16703 7224 16738 7232
rect 16249 7156 16268 7190
rect 16313 7196 16342 7204
rect 16313 7190 16330 7196
rect 16313 7188 16347 7190
rect 16395 7188 16411 7204
rect 16412 7194 16620 7204
rect 16621 7194 16637 7204
rect 16685 7200 16700 7215
rect 16703 7212 16704 7224
rect 16711 7212 16738 7224
rect 16703 7204 16738 7212
rect 16703 7203 16732 7204
rect 16423 7190 16637 7194
rect 16438 7188 16637 7190
rect 16672 7190 16685 7200
rect 16703 7190 16720 7203
rect 16672 7188 16720 7190
rect 16314 7184 16347 7188
rect 16310 7182 16347 7184
rect 16310 7181 16377 7182
rect 16310 7176 16341 7181
rect 16347 7176 16377 7181
rect 16310 7172 16377 7176
rect 16283 7169 16377 7172
rect 16283 7162 16332 7169
rect 16283 7156 16313 7162
rect 16332 7157 16337 7162
rect 16249 7140 16329 7156
rect 16341 7148 16377 7169
rect 16438 7164 16627 7188
rect 16672 7187 16719 7188
rect 16685 7182 16719 7187
rect 16453 7161 16627 7164
rect 16446 7158 16627 7161
rect 16655 7181 16719 7182
rect 16249 7138 16268 7140
rect 16283 7138 16317 7140
rect 16249 7122 16329 7138
rect 16249 7116 16268 7122
rect 15965 7090 16068 7100
rect 15919 7088 16068 7090
rect 16089 7088 16124 7100
rect 15758 7086 15920 7088
rect 15770 7066 15789 7086
rect 15804 7084 15834 7086
rect 15653 7058 15694 7066
rect 15776 7062 15789 7066
rect 15841 7070 15920 7086
rect 15952 7086 16124 7088
rect 15952 7070 16031 7086
rect 16038 7084 16068 7086
rect 15616 7048 15645 7058
rect 15659 7048 15688 7058
rect 15703 7048 15733 7062
rect 15776 7048 15819 7062
rect 15841 7058 16031 7070
rect 16096 7066 16102 7086
rect 15826 7048 15856 7058
rect 15857 7048 16015 7058
rect 16019 7048 16049 7058
rect 16053 7048 16083 7062
rect 16111 7048 16124 7086
rect 16196 7100 16225 7116
rect 16239 7100 16268 7116
rect 16283 7106 16313 7122
rect 16341 7100 16347 7148
rect 16350 7142 16369 7148
rect 16384 7142 16414 7150
rect 16350 7134 16414 7142
rect 16350 7118 16430 7134
rect 16446 7127 16508 7158
rect 16524 7127 16586 7158
rect 16655 7156 16704 7181
rect 16719 7156 16749 7172
rect 16618 7142 16648 7150
rect 16655 7148 16765 7156
rect 16618 7134 16663 7142
rect 16350 7116 16369 7118
rect 16384 7116 16430 7118
rect 16350 7100 16430 7116
rect 16457 7114 16492 7127
rect 16533 7124 16570 7127
rect 16533 7122 16575 7124
rect 16462 7111 16492 7114
rect 16471 7107 16478 7111
rect 16478 7106 16479 7107
rect 16437 7100 16447 7106
rect 16196 7092 16231 7100
rect 16196 7066 16197 7092
rect 16204 7066 16231 7092
rect 16139 7048 16169 7062
rect 16196 7058 16231 7066
rect 16233 7092 16274 7100
rect 16233 7066 16248 7092
rect 16255 7066 16274 7092
rect 16338 7088 16369 7100
rect 16384 7088 16487 7100
rect 16499 7090 16525 7116
rect 16540 7111 16570 7122
rect 16602 7118 16664 7134
rect 16602 7116 16648 7118
rect 16602 7100 16664 7116
rect 16676 7100 16682 7148
rect 16685 7140 16765 7148
rect 16685 7138 16704 7140
rect 16719 7138 16753 7140
rect 16685 7122 16765 7138
rect 16685 7100 16704 7122
rect 16719 7106 16749 7122
rect 16777 7116 16783 7190
rect 16786 7116 16805 7260
rect 16820 7116 16826 7260
rect 16835 7190 16848 7260
rect 16900 7256 16922 7260
rect 16893 7234 16922 7248
rect 16975 7234 16991 7248
rect 17029 7244 17035 7246
rect 17042 7244 17150 7260
rect 17157 7244 17163 7246
rect 17171 7244 17186 7260
rect 17252 7254 17271 7257
rect 16893 7232 16991 7234
rect 17018 7232 17186 7244
rect 17201 7234 17217 7248
rect 17252 7235 17274 7254
rect 17284 7248 17300 7249
rect 17283 7246 17300 7248
rect 17284 7241 17300 7246
rect 17274 7234 17280 7235
rect 17283 7234 17312 7241
rect 17201 7233 17312 7234
rect 17201 7232 17318 7233
rect 16877 7224 16928 7232
rect 16975 7224 17009 7232
rect 16877 7212 16902 7224
rect 16909 7212 16928 7224
rect 16982 7222 17009 7224
rect 17018 7222 17239 7232
rect 17274 7229 17280 7232
rect 16982 7218 17239 7222
rect 16877 7204 16928 7212
rect 16975 7204 17239 7218
rect 17283 7224 17318 7232
rect 16829 7156 16848 7190
rect 16893 7196 16922 7204
rect 16893 7190 16910 7196
rect 16893 7188 16927 7190
rect 16975 7188 16991 7204
rect 16992 7194 17200 7204
rect 17201 7194 17217 7204
rect 17265 7200 17280 7215
rect 17283 7212 17284 7224
rect 17291 7212 17318 7224
rect 17283 7204 17318 7212
rect 17283 7203 17312 7204
rect 17003 7190 17217 7194
rect 17018 7188 17217 7190
rect 17252 7190 17265 7200
rect 17283 7190 17300 7203
rect 17252 7188 17300 7190
rect 16894 7184 16927 7188
rect 16890 7182 16927 7184
rect 16890 7181 16957 7182
rect 16890 7176 16921 7181
rect 16927 7176 16957 7181
rect 16890 7172 16957 7176
rect 16863 7169 16957 7172
rect 16863 7162 16912 7169
rect 16863 7156 16893 7162
rect 16912 7157 16917 7162
rect 16829 7140 16909 7156
rect 16921 7148 16957 7169
rect 17018 7164 17207 7188
rect 17252 7187 17299 7188
rect 17265 7182 17299 7187
rect 17033 7161 17207 7164
rect 17026 7158 17207 7161
rect 17235 7181 17299 7182
rect 16829 7138 16848 7140
rect 16863 7138 16897 7140
rect 16829 7122 16909 7138
rect 16829 7116 16848 7122
rect 16545 7090 16648 7100
rect 16499 7088 16648 7090
rect 16669 7088 16704 7100
rect 16338 7086 16500 7088
rect 16350 7066 16369 7086
rect 16384 7084 16414 7086
rect 16233 7058 16274 7066
rect 16356 7062 16369 7066
rect 16421 7070 16500 7086
rect 16532 7086 16704 7088
rect 16532 7070 16611 7086
rect 16618 7084 16648 7086
rect 16196 7048 16225 7058
rect 16239 7048 16268 7058
rect 16283 7048 16313 7062
rect 16356 7048 16399 7062
rect 16421 7058 16611 7070
rect 16676 7066 16682 7086
rect 16406 7048 16436 7058
rect 16437 7048 16595 7058
rect 16599 7048 16629 7058
rect 16633 7048 16663 7062
rect 16691 7048 16704 7086
rect 16776 7100 16805 7116
rect 16819 7100 16848 7116
rect 16863 7106 16893 7122
rect 16921 7100 16927 7148
rect 16930 7142 16949 7148
rect 16964 7142 16994 7150
rect 16930 7134 16994 7142
rect 16930 7118 17010 7134
rect 17026 7127 17088 7158
rect 17104 7127 17166 7158
rect 17235 7156 17284 7181
rect 17299 7156 17329 7172
rect 17198 7142 17228 7150
rect 17235 7148 17345 7156
rect 17198 7134 17243 7142
rect 16930 7116 16949 7118
rect 16964 7116 17010 7118
rect 16930 7100 17010 7116
rect 17037 7114 17072 7127
rect 17113 7124 17150 7127
rect 17113 7122 17155 7124
rect 17042 7111 17072 7114
rect 17051 7107 17058 7111
rect 17058 7106 17059 7107
rect 17017 7100 17027 7106
rect 16776 7092 16811 7100
rect 16776 7066 16777 7092
rect 16784 7066 16811 7092
rect 16719 7048 16749 7062
rect 16776 7058 16811 7066
rect 16813 7092 16854 7100
rect 16813 7066 16828 7092
rect 16835 7066 16854 7092
rect 16918 7088 16949 7100
rect 16964 7088 17067 7100
rect 17079 7090 17105 7116
rect 17120 7111 17150 7122
rect 17182 7118 17244 7134
rect 17182 7116 17228 7118
rect 17182 7100 17244 7116
rect 17256 7100 17262 7148
rect 17265 7140 17345 7148
rect 17265 7138 17284 7140
rect 17299 7138 17333 7140
rect 17265 7122 17345 7138
rect 17265 7100 17284 7122
rect 17299 7106 17329 7122
rect 17357 7116 17363 7190
rect 17366 7116 17385 7260
rect 17400 7116 17406 7260
rect 17415 7190 17428 7260
rect 17480 7256 17502 7260
rect 17473 7234 17502 7248
rect 17555 7234 17571 7248
rect 17609 7244 17615 7246
rect 17622 7244 17730 7260
rect 17737 7244 17743 7246
rect 17751 7244 17766 7260
rect 17832 7254 17851 7257
rect 17473 7232 17571 7234
rect 17598 7232 17766 7244
rect 17781 7234 17797 7248
rect 17832 7235 17854 7254
rect 17864 7248 17880 7249
rect 17863 7246 17880 7248
rect 17864 7241 17880 7246
rect 17854 7234 17860 7235
rect 17863 7234 17892 7241
rect 17781 7233 17892 7234
rect 17781 7232 17898 7233
rect 17457 7224 17508 7232
rect 17555 7224 17589 7232
rect 17457 7212 17482 7224
rect 17489 7212 17508 7224
rect 17562 7222 17589 7224
rect 17598 7222 17819 7232
rect 17854 7229 17860 7232
rect 17562 7218 17819 7222
rect 17457 7204 17508 7212
rect 17555 7204 17819 7218
rect 17863 7224 17898 7232
rect 17409 7156 17428 7190
rect 17473 7196 17502 7204
rect 17473 7190 17490 7196
rect 17473 7188 17507 7190
rect 17555 7188 17571 7204
rect 17572 7194 17780 7204
rect 17781 7194 17797 7204
rect 17845 7200 17860 7215
rect 17863 7212 17864 7224
rect 17871 7212 17898 7224
rect 17863 7204 17898 7212
rect 17863 7203 17892 7204
rect 17583 7190 17797 7194
rect 17598 7188 17797 7190
rect 17832 7190 17845 7200
rect 17863 7190 17880 7203
rect 17832 7188 17880 7190
rect 17474 7184 17507 7188
rect 17470 7182 17507 7184
rect 17470 7181 17537 7182
rect 17470 7176 17501 7181
rect 17507 7176 17537 7181
rect 17470 7172 17537 7176
rect 17443 7169 17537 7172
rect 17443 7162 17492 7169
rect 17443 7156 17473 7162
rect 17492 7157 17497 7162
rect 17409 7140 17489 7156
rect 17501 7148 17537 7169
rect 17598 7164 17787 7188
rect 17832 7187 17879 7188
rect 17845 7182 17879 7187
rect 17613 7161 17787 7164
rect 17606 7158 17787 7161
rect 17815 7181 17879 7182
rect 17409 7138 17428 7140
rect 17443 7138 17477 7140
rect 17409 7122 17489 7138
rect 17409 7116 17428 7122
rect 17125 7090 17228 7100
rect 17079 7088 17228 7090
rect 17249 7088 17284 7100
rect 16918 7086 17080 7088
rect 16930 7066 16949 7086
rect 16964 7084 16994 7086
rect 16813 7058 16854 7066
rect 16936 7062 16949 7066
rect 17001 7070 17080 7086
rect 17112 7086 17284 7088
rect 17112 7070 17191 7086
rect 17198 7084 17228 7086
rect 16776 7048 16805 7058
rect 16819 7048 16848 7058
rect 16863 7048 16893 7062
rect 16936 7048 16979 7062
rect 17001 7058 17191 7070
rect 17256 7066 17262 7086
rect 16986 7048 17016 7058
rect 17017 7048 17175 7058
rect 17179 7048 17209 7058
rect 17213 7048 17243 7062
rect 17271 7048 17284 7086
rect 17356 7100 17385 7116
rect 17399 7100 17428 7116
rect 17443 7106 17473 7122
rect 17501 7100 17507 7148
rect 17510 7142 17529 7148
rect 17544 7142 17574 7150
rect 17510 7134 17574 7142
rect 17510 7118 17590 7134
rect 17606 7127 17668 7158
rect 17684 7127 17746 7158
rect 17815 7156 17864 7181
rect 17879 7156 17909 7172
rect 17778 7142 17808 7150
rect 17815 7148 17925 7156
rect 17778 7134 17823 7142
rect 17510 7116 17529 7118
rect 17544 7116 17590 7118
rect 17510 7100 17590 7116
rect 17617 7114 17652 7127
rect 17693 7124 17730 7127
rect 17693 7122 17735 7124
rect 17622 7111 17652 7114
rect 17631 7107 17638 7111
rect 17638 7106 17639 7107
rect 17597 7100 17607 7106
rect 17356 7092 17391 7100
rect 17356 7066 17357 7092
rect 17364 7066 17391 7092
rect 17299 7048 17329 7062
rect 17356 7058 17391 7066
rect 17393 7092 17434 7100
rect 17393 7066 17408 7092
rect 17415 7066 17434 7092
rect 17498 7088 17529 7100
rect 17544 7088 17647 7100
rect 17659 7090 17685 7116
rect 17700 7111 17730 7122
rect 17762 7118 17824 7134
rect 17762 7116 17808 7118
rect 17762 7100 17824 7116
rect 17836 7100 17842 7148
rect 17845 7140 17925 7148
rect 17845 7138 17864 7140
rect 17879 7138 17913 7140
rect 17845 7122 17925 7138
rect 17845 7100 17864 7122
rect 17879 7106 17909 7122
rect 17937 7116 17943 7190
rect 17946 7116 17965 7260
rect 17980 7116 17986 7260
rect 17995 7190 18008 7260
rect 18060 7256 18082 7260
rect 18053 7234 18082 7248
rect 18135 7234 18151 7248
rect 18189 7244 18195 7246
rect 18202 7244 18310 7260
rect 18317 7244 18323 7246
rect 18331 7244 18346 7260
rect 18412 7254 18431 7257
rect 18053 7232 18151 7234
rect 18178 7232 18346 7244
rect 18361 7234 18377 7248
rect 18412 7235 18434 7254
rect 18444 7248 18460 7249
rect 18443 7246 18460 7248
rect 18444 7241 18460 7246
rect 18434 7234 18440 7235
rect 18443 7234 18472 7241
rect 18361 7233 18472 7234
rect 18361 7232 18478 7233
rect 18037 7224 18088 7232
rect 18135 7224 18169 7232
rect 18037 7212 18062 7224
rect 18069 7212 18088 7224
rect 18142 7222 18169 7224
rect 18178 7222 18399 7232
rect 18434 7229 18440 7232
rect 18142 7218 18399 7222
rect 18037 7204 18088 7212
rect 18135 7204 18399 7218
rect 18443 7224 18478 7232
rect 17989 7156 18008 7190
rect 18053 7196 18082 7204
rect 18053 7190 18070 7196
rect 18053 7188 18087 7190
rect 18135 7188 18151 7204
rect 18152 7194 18360 7204
rect 18361 7194 18377 7204
rect 18425 7200 18440 7215
rect 18443 7212 18444 7224
rect 18451 7212 18478 7224
rect 18443 7204 18478 7212
rect 18443 7203 18472 7204
rect 18163 7190 18377 7194
rect 18178 7188 18377 7190
rect 18412 7190 18425 7200
rect 18443 7190 18460 7203
rect 18412 7188 18460 7190
rect 18054 7184 18087 7188
rect 18050 7182 18087 7184
rect 18050 7181 18117 7182
rect 18050 7176 18081 7181
rect 18087 7176 18117 7181
rect 18050 7172 18117 7176
rect 18023 7169 18117 7172
rect 18023 7162 18072 7169
rect 18023 7156 18053 7162
rect 18072 7157 18077 7162
rect 17989 7140 18069 7156
rect 18081 7148 18117 7169
rect 18178 7164 18367 7188
rect 18412 7187 18459 7188
rect 18425 7182 18459 7187
rect 18193 7161 18367 7164
rect 18186 7158 18367 7161
rect 18395 7181 18459 7182
rect 17989 7138 18008 7140
rect 18023 7138 18057 7140
rect 17989 7122 18069 7138
rect 17989 7116 18008 7122
rect 17705 7090 17808 7100
rect 17659 7088 17808 7090
rect 17829 7088 17864 7100
rect 17498 7086 17660 7088
rect 17510 7066 17529 7086
rect 17544 7084 17574 7086
rect 17393 7058 17434 7066
rect 17516 7062 17529 7066
rect 17581 7070 17660 7086
rect 17692 7086 17864 7088
rect 17692 7070 17771 7086
rect 17778 7084 17808 7086
rect 17356 7048 17385 7058
rect 17399 7048 17428 7058
rect 17443 7048 17473 7062
rect 17516 7048 17559 7062
rect 17581 7058 17771 7070
rect 17836 7066 17842 7086
rect 17566 7048 17596 7058
rect 17597 7048 17755 7058
rect 17759 7048 17789 7058
rect 17793 7048 17823 7062
rect 17851 7048 17864 7086
rect 17936 7100 17965 7116
rect 17979 7100 18008 7116
rect 18023 7106 18053 7122
rect 18081 7100 18087 7148
rect 18090 7142 18109 7148
rect 18124 7142 18154 7150
rect 18090 7134 18154 7142
rect 18090 7118 18170 7134
rect 18186 7127 18248 7158
rect 18264 7127 18326 7158
rect 18395 7156 18444 7181
rect 18459 7156 18489 7172
rect 18358 7142 18388 7150
rect 18395 7148 18505 7156
rect 18358 7134 18403 7142
rect 18090 7116 18109 7118
rect 18124 7116 18170 7118
rect 18090 7100 18170 7116
rect 18197 7114 18232 7127
rect 18273 7124 18310 7127
rect 18273 7122 18315 7124
rect 18202 7111 18232 7114
rect 18211 7107 18218 7111
rect 18218 7106 18219 7107
rect 18177 7100 18187 7106
rect 17936 7092 17971 7100
rect 17936 7066 17937 7092
rect 17944 7066 17971 7092
rect 17879 7048 17909 7062
rect 17936 7058 17971 7066
rect 17973 7092 18014 7100
rect 17973 7066 17988 7092
rect 17995 7066 18014 7092
rect 18078 7088 18109 7100
rect 18124 7088 18227 7100
rect 18239 7090 18265 7116
rect 18280 7111 18310 7122
rect 18342 7118 18404 7134
rect 18342 7116 18388 7118
rect 18342 7100 18404 7116
rect 18416 7100 18422 7148
rect 18425 7140 18505 7148
rect 18425 7138 18444 7140
rect 18459 7138 18493 7140
rect 18425 7122 18505 7138
rect 18425 7100 18444 7122
rect 18459 7106 18489 7122
rect 18517 7116 18523 7190
rect 18532 7116 18545 7260
rect 18285 7090 18388 7100
rect 18239 7088 18388 7090
rect 18409 7088 18444 7100
rect 18078 7086 18240 7088
rect 18090 7066 18109 7086
rect 18124 7084 18154 7086
rect 17973 7058 18014 7066
rect 18096 7062 18109 7066
rect 18161 7070 18240 7086
rect 18272 7086 18444 7088
rect 18272 7070 18351 7086
rect 18358 7084 18388 7086
rect 17936 7048 17965 7058
rect 17979 7048 18008 7058
rect 18023 7048 18053 7062
rect 18096 7048 18139 7062
rect 18161 7058 18351 7070
rect 18416 7066 18422 7086
rect 18146 7048 18176 7058
rect 18177 7048 18335 7058
rect 18339 7048 18369 7058
rect 18373 7048 18403 7062
rect 18431 7048 18444 7086
rect 18516 7100 18545 7116
rect 18516 7092 18551 7100
rect 18516 7066 18517 7092
rect 18524 7066 18551 7092
rect 18459 7048 18489 7062
rect 18516 7058 18551 7066
rect 18516 7048 18545 7058
rect -1 7042 18545 7048
rect 0 7034 18545 7042
rect 15 7004 28 7034
rect 43 7020 73 7034
rect 116 7020 159 7034
rect 166 7020 386 7034
rect 393 7020 423 7034
rect 83 7006 98 7018
rect 117 7006 130 7020
rect 198 7016 351 7020
rect 80 7004 102 7006
rect 180 7004 372 7016
rect 451 7004 464 7034
rect 479 7020 509 7034
rect 546 7004 565 7034
rect 580 7004 586 7034
rect 595 7004 608 7034
rect 623 7020 653 7034
rect 696 7020 739 7034
rect 746 7020 966 7034
rect 973 7020 1003 7034
rect 663 7006 678 7018
rect 697 7006 710 7020
rect 778 7016 931 7020
rect 660 7004 682 7006
rect 760 7004 952 7016
rect 1031 7004 1044 7034
rect 1059 7020 1089 7034
rect 1126 7004 1145 7034
rect 1160 7004 1166 7034
rect 1175 7004 1188 7034
rect 1203 7020 1233 7034
rect 1276 7020 1319 7034
rect 1326 7020 1546 7034
rect 1553 7020 1583 7034
rect 1243 7006 1258 7018
rect 1277 7006 1290 7020
rect 1358 7016 1511 7020
rect 1240 7004 1262 7006
rect 1340 7004 1532 7016
rect 1611 7004 1624 7034
rect 1639 7020 1669 7034
rect 1706 7004 1725 7034
rect 1740 7004 1746 7034
rect 1755 7004 1768 7034
rect 1783 7020 1813 7034
rect 1856 7020 1899 7034
rect 1906 7020 2126 7034
rect 2133 7020 2163 7034
rect 1823 7006 1838 7018
rect 1857 7006 1870 7020
rect 1938 7016 2091 7020
rect 1820 7004 1842 7006
rect 1920 7004 2112 7016
rect 2191 7004 2204 7034
rect 2219 7020 2249 7034
rect 2286 7004 2305 7034
rect 2320 7004 2326 7034
rect 2335 7004 2348 7034
rect 2363 7020 2393 7034
rect 2436 7020 2479 7034
rect 2486 7020 2706 7034
rect 2713 7020 2743 7034
rect 2403 7006 2418 7018
rect 2437 7006 2450 7020
rect 2518 7016 2671 7020
rect 2400 7004 2422 7006
rect 2500 7004 2692 7016
rect 2771 7004 2784 7034
rect 2799 7020 2829 7034
rect 2866 7004 2885 7034
rect 2900 7004 2906 7034
rect 2915 7004 2928 7034
rect 2943 7020 2973 7034
rect 3016 7020 3059 7034
rect 3066 7020 3286 7034
rect 3293 7020 3323 7034
rect 2983 7006 2998 7018
rect 3017 7006 3030 7020
rect 3098 7016 3251 7020
rect 2980 7004 3002 7006
rect 3080 7004 3272 7016
rect 3351 7004 3364 7034
rect 3379 7020 3409 7034
rect 3446 7004 3465 7034
rect 3480 7004 3486 7034
rect 3495 7004 3508 7034
rect 3523 7020 3553 7034
rect 3596 7020 3639 7034
rect 3646 7020 3866 7034
rect 3873 7020 3903 7034
rect 3563 7006 3578 7018
rect 3597 7006 3610 7020
rect 3678 7016 3831 7020
rect 3560 7004 3582 7006
rect 3660 7004 3852 7016
rect 3931 7004 3944 7034
rect 3959 7020 3989 7034
rect 4026 7004 4045 7034
rect 4060 7004 4066 7034
rect 4075 7004 4088 7034
rect 4103 7020 4133 7034
rect 4176 7020 4219 7034
rect 4226 7020 4446 7034
rect 4453 7020 4483 7034
rect 4143 7006 4158 7018
rect 4177 7006 4190 7020
rect 4258 7016 4411 7020
rect 4140 7004 4162 7006
rect 4240 7004 4432 7016
rect 4511 7004 4524 7034
rect 4539 7020 4569 7034
rect 4606 7004 4625 7034
rect 4640 7004 4646 7034
rect 4655 7004 4668 7034
rect 4683 7020 4713 7034
rect 4756 7020 4799 7034
rect 4806 7020 5026 7034
rect 5033 7020 5063 7034
rect 4723 7006 4738 7018
rect 4757 7006 4770 7020
rect 4838 7016 4991 7020
rect 4720 7004 4742 7006
rect 4820 7004 5012 7016
rect 5091 7004 5104 7034
rect 5119 7020 5149 7034
rect 5186 7004 5205 7034
rect 5220 7004 5226 7034
rect 5235 7004 5248 7034
rect 5263 7020 5293 7034
rect 5336 7020 5379 7034
rect 5386 7020 5606 7034
rect 5613 7020 5643 7034
rect 5303 7006 5318 7018
rect 5337 7006 5350 7020
rect 5418 7016 5571 7020
rect 5300 7004 5322 7006
rect 5400 7004 5592 7016
rect 5671 7004 5684 7034
rect 5699 7020 5729 7034
rect 5766 7004 5785 7034
rect 5800 7004 5806 7034
rect 5815 7004 5828 7034
rect 5843 7020 5873 7034
rect 5916 7020 5959 7034
rect 5966 7020 6186 7034
rect 6193 7020 6223 7034
rect 5883 7006 5898 7018
rect 5917 7006 5930 7020
rect 5998 7016 6151 7020
rect 5880 7004 5902 7006
rect 5980 7004 6172 7016
rect 6251 7004 6264 7034
rect 6279 7020 6309 7034
rect 6346 7004 6365 7034
rect 6380 7004 6386 7034
rect 6395 7004 6408 7034
rect 6423 7020 6453 7034
rect 6496 7020 6539 7034
rect 6546 7020 6766 7034
rect 6773 7020 6803 7034
rect 6463 7006 6478 7018
rect 6497 7006 6510 7020
rect 6578 7016 6731 7020
rect 6460 7004 6482 7006
rect 6560 7004 6752 7016
rect 6831 7004 6844 7034
rect 6859 7020 6889 7034
rect 6926 7004 6945 7034
rect 6960 7004 6966 7034
rect 6975 7004 6988 7034
rect 7003 7020 7033 7034
rect 7076 7020 7119 7034
rect 7126 7020 7346 7034
rect 7353 7020 7383 7034
rect 7043 7006 7058 7018
rect 7077 7006 7090 7020
rect 7158 7016 7311 7020
rect 7040 7004 7062 7006
rect 7140 7004 7332 7016
rect 7411 7004 7424 7034
rect 7439 7020 7469 7034
rect 7506 7004 7525 7034
rect 7540 7004 7546 7034
rect 7555 7004 7568 7034
rect 7583 7020 7613 7034
rect 7656 7020 7699 7034
rect 7706 7020 7926 7034
rect 7933 7020 7963 7034
rect 7623 7006 7638 7018
rect 7657 7006 7670 7020
rect 7738 7016 7891 7020
rect 7620 7004 7642 7006
rect 7720 7004 7912 7016
rect 7991 7004 8004 7034
rect 8019 7020 8049 7034
rect 8086 7004 8105 7034
rect 8120 7004 8126 7034
rect 8135 7004 8148 7034
rect 8163 7020 8193 7034
rect 8236 7020 8279 7034
rect 8286 7020 8506 7034
rect 8513 7020 8543 7034
rect 8203 7006 8218 7018
rect 8237 7006 8250 7020
rect 8318 7016 8471 7020
rect 8200 7004 8222 7006
rect 8300 7004 8492 7016
rect 8571 7004 8584 7034
rect 8599 7020 8629 7034
rect 8666 7004 8685 7034
rect 8700 7004 8706 7034
rect 8715 7004 8728 7034
rect 8743 7020 8773 7034
rect 8816 7020 8859 7034
rect 8866 7020 9086 7034
rect 9093 7020 9123 7034
rect 8783 7006 8798 7018
rect 8817 7006 8830 7020
rect 8898 7016 9051 7020
rect 8780 7004 8802 7006
rect 8880 7004 9072 7016
rect 9151 7004 9164 7034
rect 9179 7020 9209 7034
rect 9246 7004 9265 7034
rect 9280 7004 9286 7034
rect 9295 7004 9308 7034
rect 9323 7020 9353 7034
rect 9396 7020 9439 7034
rect 9446 7020 9666 7034
rect 9673 7020 9703 7034
rect 9363 7006 9378 7018
rect 9397 7006 9410 7020
rect 9478 7016 9631 7020
rect 9360 7004 9382 7006
rect 9460 7004 9652 7016
rect 9731 7004 9744 7034
rect 9759 7020 9789 7034
rect 9826 7004 9845 7034
rect 9860 7004 9866 7034
rect 9875 7004 9888 7034
rect 9903 7020 9933 7034
rect 9976 7020 10019 7034
rect 10026 7020 10246 7034
rect 10253 7020 10283 7034
rect 9943 7006 9958 7018
rect 9977 7006 9990 7020
rect 10058 7016 10211 7020
rect 9940 7004 9962 7006
rect 10040 7004 10232 7016
rect 10311 7004 10324 7034
rect 10339 7020 10369 7034
rect 10406 7004 10425 7034
rect 10440 7004 10446 7034
rect 10455 7004 10468 7034
rect 10483 7020 10513 7034
rect 10556 7020 10599 7034
rect 10606 7020 10826 7034
rect 10833 7020 10863 7034
rect 10523 7006 10538 7018
rect 10557 7006 10570 7020
rect 10638 7016 10791 7020
rect 10520 7004 10542 7006
rect 10620 7004 10812 7016
rect 10891 7004 10904 7034
rect 10919 7020 10949 7034
rect 10986 7004 11005 7034
rect 11020 7004 11026 7034
rect 11035 7004 11048 7034
rect 11063 7020 11093 7034
rect 11136 7020 11179 7034
rect 11186 7020 11406 7034
rect 11413 7020 11443 7034
rect 11103 7006 11118 7018
rect 11137 7006 11150 7020
rect 11218 7016 11371 7020
rect 11100 7004 11122 7006
rect 11200 7004 11392 7016
rect 11471 7004 11484 7034
rect 11499 7020 11529 7034
rect 11566 7004 11585 7034
rect 11600 7004 11606 7034
rect 11615 7004 11628 7034
rect 11643 7020 11673 7034
rect 11716 7020 11759 7034
rect 11766 7020 11986 7034
rect 11993 7020 12023 7034
rect 11683 7006 11698 7018
rect 11717 7006 11730 7020
rect 11798 7016 11951 7020
rect 11680 7004 11702 7006
rect 11780 7004 11972 7016
rect 12051 7004 12064 7034
rect 12079 7020 12109 7034
rect 12146 7004 12165 7034
rect 12180 7004 12186 7034
rect 12195 7004 12208 7034
rect 12223 7020 12253 7034
rect 12296 7020 12339 7034
rect 12346 7020 12566 7034
rect 12573 7020 12603 7034
rect 12263 7006 12278 7018
rect 12297 7006 12310 7020
rect 12378 7016 12531 7020
rect 12260 7004 12282 7006
rect 12360 7004 12552 7016
rect 12631 7004 12644 7034
rect 12659 7020 12689 7034
rect 12726 7004 12745 7034
rect 12760 7004 12766 7034
rect 12775 7004 12788 7034
rect 12803 7020 12833 7034
rect 12876 7020 12919 7034
rect 12926 7020 13146 7034
rect 13153 7020 13183 7034
rect 12843 7006 12858 7018
rect 12877 7006 12890 7020
rect 12958 7016 13111 7020
rect 12840 7004 12862 7006
rect 12940 7004 13132 7016
rect 13211 7004 13224 7034
rect 13239 7020 13269 7034
rect 13306 7004 13325 7034
rect 13340 7004 13346 7034
rect 13355 7004 13368 7034
rect 13383 7020 13413 7034
rect 13456 7020 13499 7034
rect 13506 7020 13726 7034
rect 13733 7020 13763 7034
rect 13423 7006 13438 7018
rect 13457 7006 13470 7020
rect 13538 7016 13691 7020
rect 13420 7004 13442 7006
rect 13520 7004 13712 7016
rect 13791 7004 13804 7034
rect 13819 7020 13849 7034
rect 13886 7004 13905 7034
rect 13920 7004 13926 7034
rect 13935 7004 13948 7034
rect 13963 7020 13993 7034
rect 14036 7020 14079 7034
rect 14086 7020 14306 7034
rect 14313 7020 14343 7034
rect 14003 7006 14018 7018
rect 14037 7006 14050 7020
rect 14118 7016 14271 7020
rect 14000 7004 14022 7006
rect 14100 7004 14292 7016
rect 14371 7004 14384 7034
rect 14399 7020 14429 7034
rect 14466 7004 14485 7034
rect 14500 7004 14506 7034
rect 14515 7004 14528 7034
rect 14543 7020 14573 7034
rect 14616 7020 14659 7034
rect 14666 7020 14886 7034
rect 14893 7020 14923 7034
rect 14583 7006 14598 7018
rect 14617 7006 14630 7020
rect 14698 7016 14851 7020
rect 14580 7004 14602 7006
rect 14680 7004 14872 7016
rect 14951 7004 14964 7034
rect 14979 7020 15009 7034
rect 15046 7004 15065 7034
rect 15080 7004 15086 7034
rect 15095 7004 15108 7034
rect 15123 7020 15153 7034
rect 15196 7020 15239 7034
rect 15246 7020 15466 7034
rect 15473 7020 15503 7034
rect 15163 7006 15178 7018
rect 15197 7006 15210 7020
rect 15278 7016 15431 7020
rect 15160 7004 15182 7006
rect 15260 7004 15452 7016
rect 15531 7004 15544 7034
rect 15559 7020 15589 7034
rect 15626 7004 15645 7034
rect 15660 7004 15666 7034
rect 15675 7004 15688 7034
rect 15703 7020 15733 7034
rect 15776 7020 15819 7034
rect 15826 7020 16046 7034
rect 16053 7020 16083 7034
rect 15743 7006 15758 7018
rect 15777 7006 15790 7020
rect 15858 7016 16011 7020
rect 15740 7004 15762 7006
rect 15840 7004 16032 7016
rect 16111 7004 16124 7034
rect 16139 7020 16169 7034
rect 16206 7004 16225 7034
rect 16240 7004 16246 7034
rect 16255 7004 16268 7034
rect 16283 7020 16313 7034
rect 16356 7020 16399 7034
rect 16406 7020 16626 7034
rect 16633 7020 16663 7034
rect 16323 7006 16338 7018
rect 16357 7006 16370 7020
rect 16438 7016 16591 7020
rect 16320 7004 16342 7006
rect 16420 7004 16612 7016
rect 16691 7004 16704 7034
rect 16719 7020 16749 7034
rect 16786 7004 16805 7034
rect 16820 7004 16826 7034
rect 16835 7004 16848 7034
rect 16863 7020 16893 7034
rect 16936 7020 16979 7034
rect 16986 7020 17206 7034
rect 17213 7020 17243 7034
rect 16903 7006 16918 7018
rect 16937 7006 16950 7020
rect 17018 7016 17171 7020
rect 16900 7004 16922 7006
rect 17000 7004 17192 7016
rect 17271 7004 17284 7034
rect 17299 7020 17329 7034
rect 17366 7004 17385 7034
rect 17400 7004 17406 7034
rect 17415 7004 17428 7034
rect 17443 7020 17473 7034
rect 17516 7020 17559 7034
rect 17566 7020 17786 7034
rect 17793 7020 17823 7034
rect 17483 7006 17498 7018
rect 17517 7006 17530 7020
rect 17598 7016 17751 7020
rect 17480 7004 17502 7006
rect 17580 7004 17772 7016
rect 17851 7004 17864 7034
rect 17879 7020 17909 7034
rect 17946 7004 17965 7034
rect 17980 7004 17986 7034
rect 17995 7004 18008 7034
rect 18023 7020 18053 7034
rect 18096 7020 18139 7034
rect 18146 7020 18366 7034
rect 18373 7020 18403 7034
rect 18063 7006 18078 7018
rect 18097 7006 18110 7020
rect 18178 7016 18331 7020
rect 18060 7004 18082 7006
rect 18160 7004 18352 7016
rect 18431 7004 18444 7034
rect 18459 7020 18489 7034
rect 18532 7004 18545 7034
rect 0 6990 18545 7004
rect 15 6920 28 6990
rect 80 6986 102 6990
rect 73 6964 102 6978
rect 155 6964 171 6978
rect 209 6974 215 6976
rect 222 6974 330 6990
rect 337 6974 343 6976
rect 351 6974 366 6990
rect 432 6984 451 6987
rect 73 6962 171 6964
rect 198 6962 366 6974
rect 381 6964 397 6978
rect 432 6965 454 6984
rect 464 6978 480 6979
rect 463 6976 480 6978
rect 464 6971 480 6976
rect 454 6964 460 6965
rect 463 6964 492 6971
rect 381 6963 492 6964
rect 381 6962 498 6963
rect 57 6954 108 6962
rect 155 6954 189 6962
rect 57 6942 82 6954
rect 89 6942 108 6954
rect 162 6952 189 6954
rect 198 6952 419 6962
rect 454 6959 460 6962
rect 162 6948 419 6952
rect 57 6934 108 6942
rect 155 6934 419 6948
rect 463 6954 498 6962
rect 9 6886 28 6920
rect 73 6926 102 6934
rect 73 6920 90 6926
rect 73 6918 107 6920
rect 155 6918 171 6934
rect 172 6924 380 6934
rect 381 6924 397 6934
rect 445 6930 460 6945
rect 463 6942 464 6954
rect 471 6942 498 6954
rect 463 6934 498 6942
rect 463 6933 492 6934
rect 183 6920 397 6924
rect 198 6918 397 6920
rect 432 6920 445 6930
rect 463 6920 480 6933
rect 432 6918 480 6920
rect 74 6914 107 6918
rect 70 6912 107 6914
rect 70 6911 137 6912
rect 70 6906 101 6911
rect 107 6906 137 6911
rect 70 6902 137 6906
rect 43 6899 137 6902
rect 43 6892 92 6899
rect 43 6886 73 6892
rect 92 6887 97 6892
rect 9 6870 89 6886
rect 101 6878 137 6899
rect 198 6894 387 6918
rect 432 6917 479 6918
rect 445 6912 479 6917
rect 213 6891 387 6894
rect 206 6888 387 6891
rect 415 6911 479 6912
rect 9 6868 28 6870
rect 43 6868 77 6870
rect 9 6852 89 6868
rect 9 6846 28 6852
rect -1 6830 28 6846
rect 43 6836 73 6852
rect 101 6830 107 6878
rect 110 6872 129 6878
rect 144 6872 174 6880
rect 110 6864 174 6872
rect 110 6848 190 6864
rect 206 6857 268 6888
rect 284 6857 346 6888
rect 415 6886 464 6911
rect 479 6886 509 6902
rect 378 6872 408 6880
rect 415 6878 525 6886
rect 378 6864 423 6872
rect 110 6846 129 6848
rect 144 6846 190 6848
rect 110 6830 190 6846
rect 217 6844 252 6857
rect 293 6854 330 6857
rect 293 6852 335 6854
rect 222 6841 252 6844
rect 231 6837 238 6841
rect 238 6836 239 6837
rect 197 6830 207 6836
rect -7 6822 34 6830
rect -7 6796 8 6822
rect 15 6796 34 6822
rect 98 6818 129 6830
rect 144 6818 247 6830
rect 259 6820 285 6846
rect 300 6841 330 6852
rect 362 6848 424 6864
rect 362 6846 408 6848
rect 362 6830 424 6846
rect 436 6830 442 6878
rect 445 6870 525 6878
rect 445 6868 464 6870
rect 479 6868 513 6870
rect 445 6852 525 6868
rect 445 6830 464 6852
rect 479 6836 509 6852
rect 537 6846 543 6920
rect 546 6846 565 6990
rect 580 6846 586 6990
rect 595 6920 608 6990
rect 660 6986 682 6990
rect 653 6964 682 6978
rect 735 6964 751 6978
rect 789 6974 795 6976
rect 802 6974 910 6990
rect 917 6974 923 6976
rect 931 6974 946 6990
rect 1012 6984 1031 6987
rect 653 6962 751 6964
rect 778 6962 946 6974
rect 961 6964 977 6978
rect 1012 6965 1034 6984
rect 1044 6978 1060 6979
rect 1043 6976 1060 6978
rect 1044 6971 1060 6976
rect 1034 6964 1040 6965
rect 1043 6964 1072 6971
rect 961 6963 1072 6964
rect 961 6962 1078 6963
rect 637 6954 688 6962
rect 735 6954 769 6962
rect 637 6942 662 6954
rect 669 6942 688 6954
rect 742 6952 769 6954
rect 778 6952 999 6962
rect 1034 6959 1040 6962
rect 742 6948 999 6952
rect 637 6934 688 6942
rect 735 6934 999 6948
rect 1043 6954 1078 6962
rect 589 6886 608 6920
rect 653 6926 682 6934
rect 653 6920 670 6926
rect 653 6918 687 6920
rect 735 6918 751 6934
rect 752 6924 960 6934
rect 961 6924 977 6934
rect 1025 6930 1040 6945
rect 1043 6942 1044 6954
rect 1051 6942 1078 6954
rect 1043 6934 1078 6942
rect 1043 6933 1072 6934
rect 763 6920 977 6924
rect 778 6918 977 6920
rect 1012 6920 1025 6930
rect 1043 6920 1060 6933
rect 1012 6918 1060 6920
rect 654 6914 687 6918
rect 650 6912 687 6914
rect 650 6911 717 6912
rect 650 6906 681 6911
rect 687 6906 717 6911
rect 650 6902 717 6906
rect 623 6899 717 6902
rect 623 6892 672 6899
rect 623 6886 653 6892
rect 672 6887 677 6892
rect 589 6870 669 6886
rect 681 6878 717 6899
rect 778 6894 967 6918
rect 1012 6917 1059 6918
rect 1025 6912 1059 6917
rect 793 6891 967 6894
rect 786 6888 967 6891
rect 995 6911 1059 6912
rect 589 6868 608 6870
rect 623 6868 657 6870
rect 589 6852 669 6868
rect 589 6846 608 6852
rect 305 6820 408 6830
rect 259 6818 408 6820
rect 429 6818 464 6830
rect 98 6816 260 6818
rect 110 6796 129 6816
rect 144 6814 174 6816
rect -7 6788 34 6796
rect 116 6792 129 6796
rect 181 6800 260 6816
rect 292 6816 464 6818
rect 292 6800 371 6816
rect 378 6814 408 6816
rect -1 6778 28 6788
rect 43 6778 73 6792
rect 116 6778 159 6792
rect 181 6788 371 6800
rect 436 6796 442 6816
rect 166 6778 196 6788
rect 197 6778 355 6788
rect 359 6778 389 6788
rect 393 6778 423 6792
rect 451 6778 464 6816
rect 536 6830 565 6846
rect 579 6830 608 6846
rect 623 6836 653 6852
rect 681 6830 687 6878
rect 690 6872 709 6878
rect 724 6872 754 6880
rect 690 6864 754 6872
rect 690 6848 770 6864
rect 786 6857 848 6888
rect 864 6857 926 6888
rect 995 6886 1044 6911
rect 1059 6886 1089 6902
rect 958 6872 988 6880
rect 995 6878 1105 6886
rect 958 6864 1003 6872
rect 690 6846 709 6848
rect 724 6846 770 6848
rect 690 6830 770 6846
rect 797 6844 832 6857
rect 873 6854 910 6857
rect 873 6852 915 6854
rect 802 6841 832 6844
rect 811 6837 818 6841
rect 818 6836 819 6837
rect 777 6830 787 6836
rect 536 6822 571 6830
rect 536 6796 537 6822
rect 544 6796 571 6822
rect 479 6778 509 6792
rect 536 6788 571 6796
rect 573 6822 614 6830
rect 573 6796 588 6822
rect 595 6796 614 6822
rect 678 6818 709 6830
rect 724 6818 827 6830
rect 839 6820 865 6846
rect 880 6841 910 6852
rect 942 6848 1004 6864
rect 942 6846 988 6848
rect 942 6830 1004 6846
rect 1016 6830 1022 6878
rect 1025 6870 1105 6878
rect 1025 6868 1044 6870
rect 1059 6868 1093 6870
rect 1025 6852 1105 6868
rect 1025 6830 1044 6852
rect 1059 6836 1089 6852
rect 1117 6846 1123 6920
rect 1126 6846 1145 6990
rect 1160 6846 1166 6990
rect 1175 6920 1188 6990
rect 1240 6986 1262 6990
rect 1233 6964 1262 6978
rect 1315 6964 1331 6978
rect 1369 6974 1375 6976
rect 1382 6974 1490 6990
rect 1497 6974 1503 6976
rect 1511 6974 1526 6990
rect 1592 6984 1611 6987
rect 1233 6962 1331 6964
rect 1358 6962 1526 6974
rect 1541 6964 1557 6978
rect 1592 6965 1614 6984
rect 1624 6978 1640 6979
rect 1623 6976 1640 6978
rect 1624 6971 1640 6976
rect 1614 6964 1620 6965
rect 1623 6964 1652 6971
rect 1541 6963 1652 6964
rect 1541 6962 1658 6963
rect 1217 6954 1268 6962
rect 1315 6954 1349 6962
rect 1217 6942 1242 6954
rect 1249 6942 1268 6954
rect 1322 6952 1349 6954
rect 1358 6952 1579 6962
rect 1614 6959 1620 6962
rect 1322 6948 1579 6952
rect 1217 6934 1268 6942
rect 1315 6934 1579 6948
rect 1623 6954 1658 6962
rect 1169 6886 1188 6920
rect 1233 6926 1262 6934
rect 1233 6920 1250 6926
rect 1233 6918 1267 6920
rect 1315 6918 1331 6934
rect 1332 6924 1540 6934
rect 1541 6924 1557 6934
rect 1605 6930 1620 6945
rect 1623 6942 1624 6954
rect 1631 6942 1658 6954
rect 1623 6934 1658 6942
rect 1623 6933 1652 6934
rect 1343 6920 1557 6924
rect 1358 6918 1557 6920
rect 1592 6920 1605 6930
rect 1623 6920 1640 6933
rect 1592 6918 1640 6920
rect 1234 6914 1267 6918
rect 1230 6912 1267 6914
rect 1230 6911 1297 6912
rect 1230 6906 1261 6911
rect 1267 6906 1297 6911
rect 1230 6902 1297 6906
rect 1203 6899 1297 6902
rect 1203 6892 1252 6899
rect 1203 6886 1233 6892
rect 1252 6887 1257 6892
rect 1169 6870 1249 6886
rect 1261 6878 1297 6899
rect 1358 6894 1547 6918
rect 1592 6917 1639 6918
rect 1605 6912 1639 6917
rect 1373 6891 1547 6894
rect 1366 6888 1547 6891
rect 1575 6911 1639 6912
rect 1169 6868 1188 6870
rect 1203 6868 1237 6870
rect 1169 6852 1249 6868
rect 1169 6846 1188 6852
rect 885 6820 988 6830
rect 839 6818 988 6820
rect 1009 6818 1044 6830
rect 678 6816 840 6818
rect 690 6796 709 6816
rect 724 6814 754 6816
rect 573 6788 614 6796
rect 696 6792 709 6796
rect 761 6800 840 6816
rect 872 6816 1044 6818
rect 872 6800 951 6816
rect 958 6814 988 6816
rect 536 6778 565 6788
rect 579 6778 608 6788
rect 623 6778 653 6792
rect 696 6778 739 6792
rect 761 6788 951 6800
rect 1016 6796 1022 6816
rect 746 6778 776 6788
rect 777 6778 935 6788
rect 939 6778 969 6788
rect 973 6778 1003 6792
rect 1031 6778 1044 6816
rect 1116 6830 1145 6846
rect 1159 6830 1188 6846
rect 1203 6836 1233 6852
rect 1261 6830 1267 6878
rect 1270 6872 1289 6878
rect 1304 6872 1334 6880
rect 1270 6864 1334 6872
rect 1270 6848 1350 6864
rect 1366 6857 1428 6888
rect 1444 6857 1506 6888
rect 1575 6886 1624 6911
rect 1639 6886 1669 6902
rect 1538 6872 1568 6880
rect 1575 6878 1685 6886
rect 1538 6864 1583 6872
rect 1270 6846 1289 6848
rect 1304 6846 1350 6848
rect 1270 6830 1350 6846
rect 1377 6844 1412 6857
rect 1453 6854 1490 6857
rect 1453 6852 1495 6854
rect 1382 6841 1412 6844
rect 1391 6837 1398 6841
rect 1398 6836 1399 6837
rect 1357 6830 1367 6836
rect 1116 6822 1151 6830
rect 1116 6796 1117 6822
rect 1124 6796 1151 6822
rect 1059 6778 1089 6792
rect 1116 6788 1151 6796
rect 1153 6822 1194 6830
rect 1153 6796 1168 6822
rect 1175 6796 1194 6822
rect 1258 6818 1289 6830
rect 1304 6818 1407 6830
rect 1419 6820 1445 6846
rect 1460 6841 1490 6852
rect 1522 6848 1584 6864
rect 1522 6846 1568 6848
rect 1522 6830 1584 6846
rect 1596 6830 1602 6878
rect 1605 6870 1685 6878
rect 1605 6868 1624 6870
rect 1639 6868 1673 6870
rect 1605 6852 1685 6868
rect 1605 6830 1624 6852
rect 1639 6836 1669 6852
rect 1697 6846 1703 6920
rect 1706 6846 1725 6990
rect 1740 6846 1746 6990
rect 1755 6920 1768 6990
rect 1820 6986 1842 6990
rect 1813 6964 1842 6978
rect 1895 6964 1911 6978
rect 1949 6974 1955 6976
rect 1962 6974 2070 6990
rect 2077 6974 2083 6976
rect 2091 6974 2106 6990
rect 2172 6984 2191 6987
rect 1813 6962 1911 6964
rect 1938 6962 2106 6974
rect 2121 6964 2137 6978
rect 2172 6965 2194 6984
rect 2204 6978 2220 6979
rect 2203 6976 2220 6978
rect 2204 6971 2220 6976
rect 2194 6964 2200 6965
rect 2203 6964 2232 6971
rect 2121 6963 2232 6964
rect 2121 6962 2238 6963
rect 1797 6954 1848 6962
rect 1895 6954 1929 6962
rect 1797 6942 1822 6954
rect 1829 6942 1848 6954
rect 1902 6952 1929 6954
rect 1938 6952 2159 6962
rect 2194 6959 2200 6962
rect 1902 6948 2159 6952
rect 1797 6934 1848 6942
rect 1895 6934 2159 6948
rect 2203 6954 2238 6962
rect 1749 6886 1768 6920
rect 1813 6926 1842 6934
rect 1813 6920 1830 6926
rect 1813 6918 1847 6920
rect 1895 6918 1911 6934
rect 1912 6924 2120 6934
rect 2121 6924 2137 6934
rect 2185 6930 2200 6945
rect 2203 6942 2204 6954
rect 2211 6942 2238 6954
rect 2203 6934 2238 6942
rect 2203 6933 2232 6934
rect 1923 6920 2137 6924
rect 1938 6918 2137 6920
rect 2172 6920 2185 6930
rect 2203 6920 2220 6933
rect 2172 6918 2220 6920
rect 1814 6914 1847 6918
rect 1810 6912 1847 6914
rect 1810 6911 1877 6912
rect 1810 6906 1841 6911
rect 1847 6906 1877 6911
rect 1810 6902 1877 6906
rect 1783 6899 1877 6902
rect 1783 6892 1832 6899
rect 1783 6886 1813 6892
rect 1832 6887 1837 6892
rect 1749 6870 1829 6886
rect 1841 6878 1877 6899
rect 1938 6894 2127 6918
rect 2172 6917 2219 6918
rect 2185 6912 2219 6917
rect 1953 6891 2127 6894
rect 1946 6888 2127 6891
rect 2155 6911 2219 6912
rect 1749 6868 1768 6870
rect 1783 6868 1817 6870
rect 1749 6852 1829 6868
rect 1749 6846 1768 6852
rect 1465 6820 1568 6830
rect 1419 6818 1568 6820
rect 1589 6818 1624 6830
rect 1258 6816 1420 6818
rect 1270 6796 1289 6816
rect 1304 6814 1334 6816
rect 1153 6788 1194 6796
rect 1276 6792 1289 6796
rect 1341 6800 1420 6816
rect 1452 6816 1624 6818
rect 1452 6800 1531 6816
rect 1538 6814 1568 6816
rect 1116 6778 1145 6788
rect 1159 6778 1188 6788
rect 1203 6778 1233 6792
rect 1276 6778 1319 6792
rect 1341 6788 1531 6800
rect 1596 6796 1602 6816
rect 1326 6778 1356 6788
rect 1357 6778 1515 6788
rect 1519 6778 1549 6788
rect 1553 6778 1583 6792
rect 1611 6778 1624 6816
rect 1696 6830 1725 6846
rect 1739 6830 1768 6846
rect 1783 6836 1813 6852
rect 1841 6830 1847 6878
rect 1850 6872 1869 6878
rect 1884 6872 1914 6880
rect 1850 6864 1914 6872
rect 1850 6848 1930 6864
rect 1946 6857 2008 6888
rect 2024 6857 2086 6888
rect 2155 6886 2204 6911
rect 2219 6886 2249 6902
rect 2118 6872 2148 6880
rect 2155 6878 2265 6886
rect 2118 6864 2163 6872
rect 1850 6846 1869 6848
rect 1884 6846 1930 6848
rect 1850 6830 1930 6846
rect 1957 6844 1992 6857
rect 2033 6854 2070 6857
rect 2033 6852 2075 6854
rect 1962 6841 1992 6844
rect 1971 6837 1978 6841
rect 1978 6836 1979 6837
rect 1937 6830 1947 6836
rect 1696 6822 1731 6830
rect 1696 6796 1697 6822
rect 1704 6796 1731 6822
rect 1639 6778 1669 6792
rect 1696 6788 1731 6796
rect 1733 6822 1774 6830
rect 1733 6796 1748 6822
rect 1755 6796 1774 6822
rect 1838 6818 1869 6830
rect 1884 6818 1987 6830
rect 1999 6820 2025 6846
rect 2040 6841 2070 6852
rect 2102 6848 2164 6864
rect 2102 6846 2148 6848
rect 2102 6830 2164 6846
rect 2176 6830 2182 6878
rect 2185 6870 2265 6878
rect 2185 6868 2204 6870
rect 2219 6868 2253 6870
rect 2185 6852 2265 6868
rect 2185 6830 2204 6852
rect 2219 6836 2249 6852
rect 2277 6846 2283 6920
rect 2286 6846 2305 6990
rect 2320 6846 2326 6990
rect 2335 6920 2348 6990
rect 2400 6986 2422 6990
rect 2393 6964 2422 6978
rect 2475 6964 2491 6978
rect 2529 6974 2535 6976
rect 2542 6974 2650 6990
rect 2657 6974 2663 6976
rect 2671 6974 2686 6990
rect 2752 6984 2771 6987
rect 2393 6962 2491 6964
rect 2518 6962 2686 6974
rect 2701 6964 2717 6978
rect 2752 6965 2774 6984
rect 2784 6978 2800 6979
rect 2783 6976 2800 6978
rect 2784 6971 2800 6976
rect 2774 6964 2780 6965
rect 2783 6964 2812 6971
rect 2701 6963 2812 6964
rect 2701 6962 2818 6963
rect 2377 6954 2428 6962
rect 2475 6954 2509 6962
rect 2377 6942 2402 6954
rect 2409 6942 2428 6954
rect 2482 6952 2509 6954
rect 2518 6952 2739 6962
rect 2774 6959 2780 6962
rect 2482 6948 2739 6952
rect 2377 6934 2428 6942
rect 2475 6934 2739 6948
rect 2783 6954 2818 6962
rect 2329 6886 2348 6920
rect 2393 6926 2422 6934
rect 2393 6920 2410 6926
rect 2393 6918 2427 6920
rect 2475 6918 2491 6934
rect 2492 6924 2700 6934
rect 2701 6924 2717 6934
rect 2765 6930 2780 6945
rect 2783 6942 2784 6954
rect 2791 6942 2818 6954
rect 2783 6934 2818 6942
rect 2783 6933 2812 6934
rect 2503 6920 2717 6924
rect 2518 6918 2717 6920
rect 2752 6920 2765 6930
rect 2783 6920 2800 6933
rect 2752 6918 2800 6920
rect 2394 6914 2427 6918
rect 2390 6912 2427 6914
rect 2390 6911 2457 6912
rect 2390 6906 2421 6911
rect 2427 6906 2457 6911
rect 2390 6902 2457 6906
rect 2363 6899 2457 6902
rect 2363 6892 2412 6899
rect 2363 6886 2393 6892
rect 2412 6887 2417 6892
rect 2329 6870 2409 6886
rect 2421 6878 2457 6899
rect 2518 6894 2707 6918
rect 2752 6917 2799 6918
rect 2765 6912 2799 6917
rect 2533 6891 2707 6894
rect 2526 6888 2707 6891
rect 2735 6911 2799 6912
rect 2329 6868 2348 6870
rect 2363 6868 2397 6870
rect 2329 6852 2409 6868
rect 2329 6846 2348 6852
rect 2045 6820 2148 6830
rect 1999 6818 2148 6820
rect 2169 6818 2204 6830
rect 1838 6816 2000 6818
rect 1850 6796 1869 6816
rect 1884 6814 1914 6816
rect 1733 6788 1774 6796
rect 1856 6792 1869 6796
rect 1921 6800 2000 6816
rect 2032 6816 2204 6818
rect 2032 6800 2111 6816
rect 2118 6814 2148 6816
rect 1696 6778 1725 6788
rect 1739 6778 1768 6788
rect 1783 6778 1813 6792
rect 1856 6778 1899 6792
rect 1921 6788 2111 6800
rect 2176 6796 2182 6816
rect 1906 6778 1936 6788
rect 1937 6778 2095 6788
rect 2099 6778 2129 6788
rect 2133 6778 2163 6792
rect 2191 6778 2204 6816
rect 2276 6830 2305 6846
rect 2319 6830 2348 6846
rect 2363 6836 2393 6852
rect 2421 6830 2427 6878
rect 2430 6872 2449 6878
rect 2464 6872 2494 6880
rect 2430 6864 2494 6872
rect 2430 6848 2510 6864
rect 2526 6857 2588 6888
rect 2604 6857 2666 6888
rect 2735 6886 2784 6911
rect 2799 6886 2829 6902
rect 2698 6872 2728 6880
rect 2735 6878 2845 6886
rect 2698 6864 2743 6872
rect 2430 6846 2449 6848
rect 2464 6846 2510 6848
rect 2430 6830 2510 6846
rect 2537 6844 2572 6857
rect 2613 6854 2650 6857
rect 2613 6852 2655 6854
rect 2542 6841 2572 6844
rect 2551 6837 2558 6841
rect 2558 6836 2559 6837
rect 2517 6830 2527 6836
rect 2276 6822 2311 6830
rect 2276 6796 2277 6822
rect 2284 6796 2311 6822
rect 2219 6778 2249 6792
rect 2276 6788 2311 6796
rect 2313 6822 2354 6830
rect 2313 6796 2328 6822
rect 2335 6796 2354 6822
rect 2418 6818 2449 6830
rect 2464 6818 2567 6830
rect 2579 6820 2605 6846
rect 2620 6841 2650 6852
rect 2682 6848 2744 6864
rect 2682 6846 2728 6848
rect 2682 6830 2744 6846
rect 2756 6830 2762 6878
rect 2765 6870 2845 6878
rect 2765 6868 2784 6870
rect 2799 6868 2833 6870
rect 2765 6852 2845 6868
rect 2765 6830 2784 6852
rect 2799 6836 2829 6852
rect 2857 6846 2863 6920
rect 2866 6846 2885 6990
rect 2900 6846 2906 6990
rect 2915 6920 2928 6990
rect 2980 6986 3002 6990
rect 2973 6964 3002 6978
rect 3055 6964 3071 6978
rect 3109 6974 3115 6976
rect 3122 6974 3230 6990
rect 3237 6974 3243 6976
rect 3251 6974 3266 6990
rect 3332 6984 3351 6987
rect 2973 6962 3071 6964
rect 3098 6962 3266 6974
rect 3281 6964 3297 6978
rect 3332 6965 3354 6984
rect 3364 6978 3380 6979
rect 3363 6976 3380 6978
rect 3364 6971 3380 6976
rect 3354 6964 3360 6965
rect 3363 6964 3392 6971
rect 3281 6963 3392 6964
rect 3281 6962 3398 6963
rect 2957 6954 3008 6962
rect 3055 6954 3089 6962
rect 2957 6942 2982 6954
rect 2989 6942 3008 6954
rect 3062 6952 3089 6954
rect 3098 6952 3319 6962
rect 3354 6959 3360 6962
rect 3062 6948 3319 6952
rect 2957 6934 3008 6942
rect 3055 6934 3319 6948
rect 3363 6954 3398 6962
rect 2909 6886 2928 6920
rect 2973 6926 3002 6934
rect 2973 6920 2990 6926
rect 2973 6918 3007 6920
rect 3055 6918 3071 6934
rect 3072 6924 3280 6934
rect 3281 6924 3297 6934
rect 3345 6930 3360 6945
rect 3363 6942 3364 6954
rect 3371 6942 3398 6954
rect 3363 6934 3398 6942
rect 3363 6933 3392 6934
rect 3083 6920 3297 6924
rect 3098 6918 3297 6920
rect 3332 6920 3345 6930
rect 3363 6920 3380 6933
rect 3332 6918 3380 6920
rect 2974 6914 3007 6918
rect 2970 6912 3007 6914
rect 2970 6911 3037 6912
rect 2970 6906 3001 6911
rect 3007 6906 3037 6911
rect 2970 6902 3037 6906
rect 2943 6899 3037 6902
rect 2943 6892 2992 6899
rect 2943 6886 2973 6892
rect 2992 6887 2997 6892
rect 2909 6870 2989 6886
rect 3001 6878 3037 6899
rect 3098 6894 3287 6918
rect 3332 6917 3379 6918
rect 3345 6912 3379 6917
rect 3113 6891 3287 6894
rect 3106 6888 3287 6891
rect 3315 6911 3379 6912
rect 2909 6868 2928 6870
rect 2943 6868 2977 6870
rect 2909 6852 2989 6868
rect 2909 6846 2928 6852
rect 2625 6820 2728 6830
rect 2579 6818 2728 6820
rect 2749 6818 2784 6830
rect 2418 6816 2580 6818
rect 2430 6796 2449 6816
rect 2464 6814 2494 6816
rect 2313 6788 2354 6796
rect 2436 6792 2449 6796
rect 2501 6800 2580 6816
rect 2612 6816 2784 6818
rect 2612 6800 2691 6816
rect 2698 6814 2728 6816
rect 2276 6778 2305 6788
rect 2319 6778 2348 6788
rect 2363 6778 2393 6792
rect 2436 6778 2479 6792
rect 2501 6788 2691 6800
rect 2756 6796 2762 6816
rect 2486 6778 2516 6788
rect 2517 6778 2675 6788
rect 2679 6778 2709 6788
rect 2713 6778 2743 6792
rect 2771 6778 2784 6816
rect 2856 6830 2885 6846
rect 2899 6830 2928 6846
rect 2943 6836 2973 6852
rect 3001 6830 3007 6878
rect 3010 6872 3029 6878
rect 3044 6872 3074 6880
rect 3010 6864 3074 6872
rect 3010 6848 3090 6864
rect 3106 6857 3168 6888
rect 3184 6857 3246 6888
rect 3315 6886 3364 6911
rect 3379 6886 3409 6902
rect 3278 6872 3308 6880
rect 3315 6878 3425 6886
rect 3278 6864 3323 6872
rect 3010 6846 3029 6848
rect 3044 6846 3090 6848
rect 3010 6830 3090 6846
rect 3117 6844 3152 6857
rect 3193 6854 3230 6857
rect 3193 6852 3235 6854
rect 3122 6841 3152 6844
rect 3131 6837 3138 6841
rect 3138 6836 3139 6837
rect 3097 6830 3107 6836
rect 2856 6822 2891 6830
rect 2856 6796 2857 6822
rect 2864 6796 2891 6822
rect 2799 6778 2829 6792
rect 2856 6788 2891 6796
rect 2893 6822 2934 6830
rect 2893 6796 2908 6822
rect 2915 6796 2934 6822
rect 2998 6818 3029 6830
rect 3044 6818 3147 6830
rect 3159 6820 3185 6846
rect 3200 6841 3230 6852
rect 3262 6848 3324 6864
rect 3262 6846 3308 6848
rect 3262 6830 3324 6846
rect 3336 6830 3342 6878
rect 3345 6870 3425 6878
rect 3345 6868 3364 6870
rect 3379 6868 3413 6870
rect 3345 6852 3425 6868
rect 3345 6830 3364 6852
rect 3379 6836 3409 6852
rect 3437 6846 3443 6920
rect 3446 6846 3465 6990
rect 3480 6846 3486 6990
rect 3495 6920 3508 6990
rect 3560 6986 3582 6990
rect 3553 6964 3582 6978
rect 3635 6964 3651 6978
rect 3689 6974 3695 6976
rect 3702 6974 3810 6990
rect 3817 6974 3823 6976
rect 3831 6974 3846 6990
rect 3912 6984 3931 6987
rect 3553 6962 3651 6964
rect 3678 6962 3846 6974
rect 3861 6964 3877 6978
rect 3912 6965 3934 6984
rect 3944 6978 3960 6979
rect 3943 6976 3960 6978
rect 3944 6971 3960 6976
rect 3934 6964 3940 6965
rect 3943 6964 3972 6971
rect 3861 6963 3972 6964
rect 3861 6962 3978 6963
rect 3537 6954 3588 6962
rect 3635 6954 3669 6962
rect 3537 6942 3562 6954
rect 3569 6942 3588 6954
rect 3642 6952 3669 6954
rect 3678 6952 3899 6962
rect 3934 6959 3940 6962
rect 3642 6948 3899 6952
rect 3537 6934 3588 6942
rect 3635 6934 3899 6948
rect 3943 6954 3978 6962
rect 3489 6886 3508 6920
rect 3553 6926 3582 6934
rect 3553 6920 3570 6926
rect 3553 6918 3587 6920
rect 3635 6918 3651 6934
rect 3652 6924 3860 6934
rect 3861 6924 3877 6934
rect 3925 6930 3940 6945
rect 3943 6942 3944 6954
rect 3951 6942 3978 6954
rect 3943 6934 3978 6942
rect 3943 6933 3972 6934
rect 3663 6920 3877 6924
rect 3678 6918 3877 6920
rect 3912 6920 3925 6930
rect 3943 6920 3960 6933
rect 3912 6918 3960 6920
rect 3554 6914 3587 6918
rect 3550 6912 3587 6914
rect 3550 6911 3617 6912
rect 3550 6906 3581 6911
rect 3587 6906 3617 6911
rect 3550 6902 3617 6906
rect 3523 6899 3617 6902
rect 3523 6892 3572 6899
rect 3523 6886 3553 6892
rect 3572 6887 3577 6892
rect 3489 6870 3569 6886
rect 3581 6878 3617 6899
rect 3678 6894 3867 6918
rect 3912 6917 3959 6918
rect 3925 6912 3959 6917
rect 3693 6891 3867 6894
rect 3686 6888 3867 6891
rect 3895 6911 3959 6912
rect 3489 6868 3508 6870
rect 3523 6868 3557 6870
rect 3489 6852 3569 6868
rect 3489 6846 3508 6852
rect 3205 6820 3308 6830
rect 3159 6818 3308 6820
rect 3329 6818 3364 6830
rect 2998 6816 3160 6818
rect 3010 6796 3029 6816
rect 3044 6814 3074 6816
rect 2893 6788 2934 6796
rect 3016 6792 3029 6796
rect 3081 6800 3160 6816
rect 3192 6816 3364 6818
rect 3192 6800 3271 6816
rect 3278 6814 3308 6816
rect 2856 6778 2885 6788
rect 2899 6778 2928 6788
rect 2943 6778 2973 6792
rect 3016 6778 3059 6792
rect 3081 6788 3271 6800
rect 3336 6796 3342 6816
rect 3066 6778 3096 6788
rect 3097 6778 3255 6788
rect 3259 6778 3289 6788
rect 3293 6778 3323 6792
rect 3351 6778 3364 6816
rect 3436 6830 3465 6846
rect 3479 6830 3508 6846
rect 3523 6836 3553 6852
rect 3581 6830 3587 6878
rect 3590 6872 3609 6878
rect 3624 6872 3654 6880
rect 3590 6864 3654 6872
rect 3590 6848 3670 6864
rect 3686 6857 3748 6888
rect 3764 6857 3826 6888
rect 3895 6886 3944 6911
rect 3959 6886 3989 6902
rect 3858 6872 3888 6880
rect 3895 6878 4005 6886
rect 3858 6864 3903 6872
rect 3590 6846 3609 6848
rect 3624 6846 3670 6848
rect 3590 6830 3670 6846
rect 3697 6844 3732 6857
rect 3773 6854 3810 6857
rect 3773 6852 3815 6854
rect 3702 6841 3732 6844
rect 3711 6837 3718 6841
rect 3718 6836 3719 6837
rect 3677 6830 3687 6836
rect 3436 6822 3471 6830
rect 3436 6796 3437 6822
rect 3444 6796 3471 6822
rect 3379 6778 3409 6792
rect 3436 6788 3471 6796
rect 3473 6822 3514 6830
rect 3473 6796 3488 6822
rect 3495 6796 3514 6822
rect 3578 6818 3609 6830
rect 3624 6818 3727 6830
rect 3739 6820 3765 6846
rect 3780 6841 3810 6852
rect 3842 6848 3904 6864
rect 3842 6846 3888 6848
rect 3842 6830 3904 6846
rect 3916 6830 3922 6878
rect 3925 6870 4005 6878
rect 3925 6868 3944 6870
rect 3959 6868 3993 6870
rect 3925 6852 4005 6868
rect 3925 6830 3944 6852
rect 3959 6836 3989 6852
rect 4017 6846 4023 6920
rect 4026 6846 4045 6990
rect 4060 6846 4066 6990
rect 4075 6920 4088 6990
rect 4140 6986 4162 6990
rect 4133 6964 4162 6978
rect 4215 6964 4231 6978
rect 4269 6974 4275 6976
rect 4282 6974 4390 6990
rect 4397 6974 4403 6976
rect 4411 6974 4426 6990
rect 4492 6984 4511 6987
rect 4133 6962 4231 6964
rect 4258 6962 4426 6974
rect 4441 6964 4457 6978
rect 4492 6965 4514 6984
rect 4524 6978 4540 6979
rect 4523 6976 4540 6978
rect 4524 6971 4540 6976
rect 4514 6964 4520 6965
rect 4523 6964 4552 6971
rect 4441 6963 4552 6964
rect 4441 6962 4558 6963
rect 4117 6954 4168 6962
rect 4215 6954 4249 6962
rect 4117 6942 4142 6954
rect 4149 6942 4168 6954
rect 4222 6952 4249 6954
rect 4258 6952 4479 6962
rect 4514 6959 4520 6962
rect 4222 6948 4479 6952
rect 4117 6934 4168 6942
rect 4215 6934 4479 6948
rect 4523 6954 4558 6962
rect 4069 6886 4088 6920
rect 4133 6926 4162 6934
rect 4133 6920 4150 6926
rect 4133 6918 4167 6920
rect 4215 6918 4231 6934
rect 4232 6924 4440 6934
rect 4441 6924 4457 6934
rect 4505 6930 4520 6945
rect 4523 6942 4524 6954
rect 4531 6942 4558 6954
rect 4523 6934 4558 6942
rect 4523 6933 4552 6934
rect 4243 6920 4457 6924
rect 4258 6918 4457 6920
rect 4492 6920 4505 6930
rect 4523 6920 4540 6933
rect 4492 6918 4540 6920
rect 4134 6914 4167 6918
rect 4130 6912 4167 6914
rect 4130 6911 4197 6912
rect 4130 6906 4161 6911
rect 4167 6906 4197 6911
rect 4130 6902 4197 6906
rect 4103 6899 4197 6902
rect 4103 6892 4152 6899
rect 4103 6886 4133 6892
rect 4152 6887 4157 6892
rect 4069 6870 4149 6886
rect 4161 6878 4197 6899
rect 4258 6894 4447 6918
rect 4492 6917 4539 6918
rect 4505 6912 4539 6917
rect 4273 6891 4447 6894
rect 4266 6888 4447 6891
rect 4475 6911 4539 6912
rect 4069 6868 4088 6870
rect 4103 6868 4137 6870
rect 4069 6852 4149 6868
rect 4069 6846 4088 6852
rect 3785 6820 3888 6830
rect 3739 6818 3888 6820
rect 3909 6818 3944 6830
rect 3578 6816 3740 6818
rect 3590 6796 3609 6816
rect 3624 6814 3654 6816
rect 3473 6788 3514 6796
rect 3596 6792 3609 6796
rect 3661 6800 3740 6816
rect 3772 6816 3944 6818
rect 3772 6800 3851 6816
rect 3858 6814 3888 6816
rect 3436 6778 3465 6788
rect 3479 6778 3508 6788
rect 3523 6778 3553 6792
rect 3596 6778 3639 6792
rect 3661 6788 3851 6800
rect 3916 6796 3922 6816
rect 3646 6778 3676 6788
rect 3677 6778 3835 6788
rect 3839 6778 3869 6788
rect 3873 6778 3903 6792
rect 3931 6778 3944 6816
rect 4016 6830 4045 6846
rect 4059 6830 4088 6846
rect 4103 6836 4133 6852
rect 4161 6830 4167 6878
rect 4170 6872 4189 6878
rect 4204 6872 4234 6880
rect 4170 6864 4234 6872
rect 4170 6848 4250 6864
rect 4266 6857 4328 6888
rect 4344 6857 4406 6888
rect 4475 6886 4524 6911
rect 4539 6886 4569 6902
rect 4438 6872 4468 6880
rect 4475 6878 4585 6886
rect 4438 6864 4483 6872
rect 4170 6846 4189 6848
rect 4204 6846 4250 6848
rect 4170 6830 4250 6846
rect 4277 6844 4312 6857
rect 4353 6854 4390 6857
rect 4353 6852 4395 6854
rect 4282 6841 4312 6844
rect 4291 6837 4298 6841
rect 4298 6836 4299 6837
rect 4257 6830 4267 6836
rect 4016 6822 4051 6830
rect 4016 6796 4017 6822
rect 4024 6796 4051 6822
rect 3959 6778 3989 6792
rect 4016 6788 4051 6796
rect 4053 6822 4094 6830
rect 4053 6796 4068 6822
rect 4075 6796 4094 6822
rect 4158 6818 4189 6830
rect 4204 6818 4307 6830
rect 4319 6820 4345 6846
rect 4360 6841 4390 6852
rect 4422 6848 4484 6864
rect 4422 6846 4468 6848
rect 4422 6830 4484 6846
rect 4496 6830 4502 6878
rect 4505 6870 4585 6878
rect 4505 6868 4524 6870
rect 4539 6868 4573 6870
rect 4505 6852 4585 6868
rect 4505 6830 4524 6852
rect 4539 6836 4569 6852
rect 4597 6846 4603 6920
rect 4606 6846 4625 6990
rect 4640 6846 4646 6990
rect 4655 6920 4668 6990
rect 4720 6986 4742 6990
rect 4713 6964 4742 6978
rect 4795 6964 4811 6978
rect 4849 6974 4855 6976
rect 4862 6974 4970 6990
rect 4977 6974 4983 6976
rect 4991 6974 5006 6990
rect 5072 6984 5091 6987
rect 4713 6962 4811 6964
rect 4838 6962 5006 6974
rect 5021 6964 5037 6978
rect 5072 6965 5094 6984
rect 5104 6978 5120 6979
rect 5103 6976 5120 6978
rect 5104 6971 5120 6976
rect 5094 6964 5100 6965
rect 5103 6964 5132 6971
rect 5021 6963 5132 6964
rect 5021 6962 5138 6963
rect 4697 6954 4748 6962
rect 4795 6954 4829 6962
rect 4697 6942 4722 6954
rect 4729 6942 4748 6954
rect 4802 6952 4829 6954
rect 4838 6952 5059 6962
rect 5094 6959 5100 6962
rect 4802 6948 5059 6952
rect 4697 6934 4748 6942
rect 4795 6934 5059 6948
rect 5103 6954 5138 6962
rect 4649 6886 4668 6920
rect 4713 6926 4742 6934
rect 4713 6920 4730 6926
rect 4713 6918 4747 6920
rect 4795 6918 4811 6934
rect 4812 6924 5020 6934
rect 5021 6924 5037 6934
rect 5085 6930 5100 6945
rect 5103 6942 5104 6954
rect 5111 6942 5138 6954
rect 5103 6934 5138 6942
rect 5103 6933 5132 6934
rect 4823 6920 5037 6924
rect 4838 6918 5037 6920
rect 5072 6920 5085 6930
rect 5103 6920 5120 6933
rect 5072 6918 5120 6920
rect 4714 6914 4747 6918
rect 4710 6912 4747 6914
rect 4710 6911 4777 6912
rect 4710 6906 4741 6911
rect 4747 6906 4777 6911
rect 4710 6902 4777 6906
rect 4683 6899 4777 6902
rect 4683 6892 4732 6899
rect 4683 6886 4713 6892
rect 4732 6887 4737 6892
rect 4649 6870 4729 6886
rect 4741 6878 4777 6899
rect 4838 6894 5027 6918
rect 5072 6917 5119 6918
rect 5085 6912 5119 6917
rect 4853 6891 5027 6894
rect 4846 6888 5027 6891
rect 5055 6911 5119 6912
rect 4649 6868 4668 6870
rect 4683 6868 4717 6870
rect 4649 6852 4729 6868
rect 4649 6846 4668 6852
rect 4365 6820 4468 6830
rect 4319 6818 4468 6820
rect 4489 6818 4524 6830
rect 4158 6816 4320 6818
rect 4170 6796 4189 6816
rect 4204 6814 4234 6816
rect 4053 6788 4094 6796
rect 4176 6792 4189 6796
rect 4241 6800 4320 6816
rect 4352 6816 4524 6818
rect 4352 6800 4431 6816
rect 4438 6814 4468 6816
rect 4016 6778 4045 6788
rect 4059 6778 4088 6788
rect 4103 6778 4133 6792
rect 4176 6778 4219 6792
rect 4241 6788 4431 6800
rect 4496 6796 4502 6816
rect 4226 6778 4256 6788
rect 4257 6778 4415 6788
rect 4419 6778 4449 6788
rect 4453 6778 4483 6792
rect 4511 6778 4524 6816
rect 4596 6830 4625 6846
rect 4639 6830 4668 6846
rect 4683 6836 4713 6852
rect 4741 6830 4747 6878
rect 4750 6872 4769 6878
rect 4784 6872 4814 6880
rect 4750 6864 4814 6872
rect 4750 6848 4830 6864
rect 4846 6857 4908 6888
rect 4924 6857 4986 6888
rect 5055 6886 5104 6911
rect 5119 6886 5149 6902
rect 5018 6872 5048 6880
rect 5055 6878 5165 6886
rect 5018 6864 5063 6872
rect 4750 6846 4769 6848
rect 4784 6846 4830 6848
rect 4750 6830 4830 6846
rect 4857 6844 4892 6857
rect 4933 6854 4970 6857
rect 4933 6852 4975 6854
rect 4862 6841 4892 6844
rect 4871 6837 4878 6841
rect 4878 6836 4879 6837
rect 4837 6830 4847 6836
rect 4596 6822 4631 6830
rect 4596 6796 4597 6822
rect 4604 6796 4631 6822
rect 4539 6778 4569 6792
rect 4596 6788 4631 6796
rect 4633 6822 4674 6830
rect 4633 6796 4648 6822
rect 4655 6796 4674 6822
rect 4738 6818 4769 6830
rect 4784 6818 4887 6830
rect 4899 6820 4925 6846
rect 4940 6841 4970 6852
rect 5002 6848 5064 6864
rect 5002 6846 5048 6848
rect 5002 6830 5064 6846
rect 5076 6830 5082 6878
rect 5085 6870 5165 6878
rect 5085 6868 5104 6870
rect 5119 6868 5153 6870
rect 5085 6852 5165 6868
rect 5085 6830 5104 6852
rect 5119 6836 5149 6852
rect 5177 6846 5183 6920
rect 5186 6846 5205 6990
rect 5220 6846 5226 6990
rect 5235 6920 5248 6990
rect 5300 6986 5322 6990
rect 5293 6964 5322 6978
rect 5375 6964 5391 6978
rect 5429 6974 5435 6976
rect 5442 6974 5550 6990
rect 5557 6974 5563 6976
rect 5571 6974 5586 6990
rect 5652 6984 5671 6987
rect 5293 6962 5391 6964
rect 5418 6962 5586 6974
rect 5601 6964 5617 6978
rect 5652 6965 5674 6984
rect 5684 6978 5700 6979
rect 5683 6976 5700 6978
rect 5684 6971 5700 6976
rect 5674 6964 5680 6965
rect 5683 6964 5712 6971
rect 5601 6963 5712 6964
rect 5601 6962 5718 6963
rect 5277 6954 5328 6962
rect 5375 6954 5409 6962
rect 5277 6942 5302 6954
rect 5309 6942 5328 6954
rect 5382 6952 5409 6954
rect 5418 6952 5639 6962
rect 5674 6959 5680 6962
rect 5382 6948 5639 6952
rect 5277 6934 5328 6942
rect 5375 6934 5639 6948
rect 5683 6954 5718 6962
rect 5229 6886 5248 6920
rect 5293 6926 5322 6934
rect 5293 6920 5310 6926
rect 5293 6918 5327 6920
rect 5375 6918 5391 6934
rect 5392 6924 5600 6934
rect 5601 6924 5617 6934
rect 5665 6930 5680 6945
rect 5683 6942 5684 6954
rect 5691 6942 5718 6954
rect 5683 6934 5718 6942
rect 5683 6933 5712 6934
rect 5403 6920 5617 6924
rect 5418 6918 5617 6920
rect 5652 6920 5665 6930
rect 5683 6920 5700 6933
rect 5652 6918 5700 6920
rect 5294 6914 5327 6918
rect 5290 6912 5327 6914
rect 5290 6911 5357 6912
rect 5290 6906 5321 6911
rect 5327 6906 5357 6911
rect 5290 6902 5357 6906
rect 5263 6899 5357 6902
rect 5263 6892 5312 6899
rect 5263 6886 5293 6892
rect 5312 6887 5317 6892
rect 5229 6870 5309 6886
rect 5321 6878 5357 6899
rect 5418 6894 5607 6918
rect 5652 6917 5699 6918
rect 5665 6912 5699 6917
rect 5433 6891 5607 6894
rect 5426 6888 5607 6891
rect 5635 6911 5699 6912
rect 5229 6868 5248 6870
rect 5263 6868 5297 6870
rect 5229 6852 5309 6868
rect 5229 6846 5248 6852
rect 4945 6820 5048 6830
rect 4899 6818 5048 6820
rect 5069 6818 5104 6830
rect 4738 6816 4900 6818
rect 4750 6796 4769 6816
rect 4784 6814 4814 6816
rect 4633 6788 4674 6796
rect 4756 6792 4769 6796
rect 4821 6800 4900 6816
rect 4932 6816 5104 6818
rect 4932 6800 5011 6816
rect 5018 6814 5048 6816
rect 4596 6778 4625 6788
rect 4639 6778 4668 6788
rect 4683 6778 4713 6792
rect 4756 6778 4799 6792
rect 4821 6788 5011 6800
rect 5076 6796 5082 6816
rect 4806 6778 4836 6788
rect 4837 6778 4995 6788
rect 4999 6778 5029 6788
rect 5033 6778 5063 6792
rect 5091 6778 5104 6816
rect 5176 6830 5205 6846
rect 5219 6830 5248 6846
rect 5263 6836 5293 6852
rect 5321 6830 5327 6878
rect 5330 6872 5349 6878
rect 5364 6872 5394 6880
rect 5330 6864 5394 6872
rect 5330 6848 5410 6864
rect 5426 6857 5488 6888
rect 5504 6857 5566 6888
rect 5635 6886 5684 6911
rect 5699 6886 5729 6902
rect 5598 6872 5628 6880
rect 5635 6878 5745 6886
rect 5598 6864 5643 6872
rect 5330 6846 5349 6848
rect 5364 6846 5410 6848
rect 5330 6830 5410 6846
rect 5437 6844 5472 6857
rect 5513 6854 5550 6857
rect 5513 6852 5555 6854
rect 5442 6841 5472 6844
rect 5451 6837 5458 6841
rect 5458 6836 5459 6837
rect 5417 6830 5427 6836
rect 5176 6822 5211 6830
rect 5176 6796 5177 6822
rect 5184 6796 5211 6822
rect 5119 6778 5149 6792
rect 5176 6788 5211 6796
rect 5213 6822 5254 6830
rect 5213 6796 5228 6822
rect 5235 6796 5254 6822
rect 5318 6818 5349 6830
rect 5364 6818 5467 6830
rect 5479 6820 5505 6846
rect 5520 6841 5550 6852
rect 5582 6848 5644 6864
rect 5582 6846 5628 6848
rect 5582 6830 5644 6846
rect 5656 6830 5662 6878
rect 5665 6870 5745 6878
rect 5665 6868 5684 6870
rect 5699 6868 5733 6870
rect 5665 6852 5745 6868
rect 5665 6830 5684 6852
rect 5699 6836 5729 6852
rect 5757 6846 5763 6920
rect 5766 6846 5785 6990
rect 5800 6846 5806 6990
rect 5815 6920 5828 6990
rect 5880 6986 5902 6990
rect 5873 6964 5902 6978
rect 5955 6964 5971 6978
rect 6009 6974 6015 6976
rect 6022 6974 6130 6990
rect 6137 6974 6143 6976
rect 6151 6974 6166 6990
rect 6232 6984 6251 6987
rect 5873 6962 5971 6964
rect 5998 6962 6166 6974
rect 6181 6964 6197 6978
rect 6232 6965 6254 6984
rect 6264 6978 6280 6979
rect 6263 6976 6280 6978
rect 6264 6971 6280 6976
rect 6254 6964 6260 6965
rect 6263 6964 6292 6971
rect 6181 6963 6292 6964
rect 6181 6962 6298 6963
rect 5857 6954 5908 6962
rect 5955 6954 5989 6962
rect 5857 6942 5882 6954
rect 5889 6942 5908 6954
rect 5962 6952 5989 6954
rect 5998 6952 6219 6962
rect 6254 6959 6260 6962
rect 5962 6948 6219 6952
rect 5857 6934 5908 6942
rect 5955 6934 6219 6948
rect 6263 6954 6298 6962
rect 5809 6886 5828 6920
rect 5873 6926 5902 6934
rect 5873 6920 5890 6926
rect 5873 6918 5907 6920
rect 5955 6918 5971 6934
rect 5972 6924 6180 6934
rect 6181 6924 6197 6934
rect 6245 6930 6260 6945
rect 6263 6942 6264 6954
rect 6271 6942 6298 6954
rect 6263 6934 6298 6942
rect 6263 6933 6292 6934
rect 5983 6920 6197 6924
rect 5998 6918 6197 6920
rect 6232 6920 6245 6930
rect 6263 6920 6280 6933
rect 6232 6918 6280 6920
rect 5874 6914 5907 6918
rect 5870 6912 5907 6914
rect 5870 6911 5937 6912
rect 5870 6906 5901 6911
rect 5907 6906 5937 6911
rect 5870 6902 5937 6906
rect 5843 6899 5937 6902
rect 5843 6892 5892 6899
rect 5843 6886 5873 6892
rect 5892 6887 5897 6892
rect 5809 6870 5889 6886
rect 5901 6878 5937 6899
rect 5998 6894 6187 6918
rect 6232 6917 6279 6918
rect 6245 6912 6279 6917
rect 6013 6891 6187 6894
rect 6006 6888 6187 6891
rect 6215 6911 6279 6912
rect 5809 6868 5828 6870
rect 5843 6868 5877 6870
rect 5809 6852 5889 6868
rect 5809 6846 5828 6852
rect 5525 6820 5628 6830
rect 5479 6818 5628 6820
rect 5649 6818 5684 6830
rect 5318 6816 5480 6818
rect 5330 6796 5349 6816
rect 5364 6814 5394 6816
rect 5213 6788 5254 6796
rect 5336 6792 5349 6796
rect 5401 6800 5480 6816
rect 5512 6816 5684 6818
rect 5512 6800 5591 6816
rect 5598 6814 5628 6816
rect 5176 6778 5205 6788
rect 5219 6778 5248 6788
rect 5263 6778 5293 6792
rect 5336 6778 5379 6792
rect 5401 6788 5591 6800
rect 5656 6796 5662 6816
rect 5386 6778 5416 6788
rect 5417 6778 5575 6788
rect 5579 6778 5609 6788
rect 5613 6778 5643 6792
rect 5671 6778 5684 6816
rect 5756 6830 5785 6846
rect 5799 6830 5828 6846
rect 5843 6836 5873 6852
rect 5901 6830 5907 6878
rect 5910 6872 5929 6878
rect 5944 6872 5974 6880
rect 5910 6864 5974 6872
rect 5910 6848 5990 6864
rect 6006 6857 6068 6888
rect 6084 6857 6146 6888
rect 6215 6886 6264 6911
rect 6279 6886 6309 6902
rect 6178 6872 6208 6880
rect 6215 6878 6325 6886
rect 6178 6864 6223 6872
rect 5910 6846 5929 6848
rect 5944 6846 5990 6848
rect 5910 6830 5990 6846
rect 6017 6844 6052 6857
rect 6093 6854 6130 6857
rect 6093 6852 6135 6854
rect 6022 6841 6052 6844
rect 6031 6837 6038 6841
rect 6038 6836 6039 6837
rect 5997 6830 6007 6836
rect 5756 6822 5791 6830
rect 5756 6796 5757 6822
rect 5764 6796 5791 6822
rect 5699 6778 5729 6792
rect 5756 6788 5791 6796
rect 5793 6822 5834 6830
rect 5793 6796 5808 6822
rect 5815 6796 5834 6822
rect 5898 6818 5929 6830
rect 5944 6818 6047 6830
rect 6059 6820 6085 6846
rect 6100 6841 6130 6852
rect 6162 6848 6224 6864
rect 6162 6846 6208 6848
rect 6162 6830 6224 6846
rect 6236 6830 6242 6878
rect 6245 6870 6325 6878
rect 6245 6868 6264 6870
rect 6279 6868 6313 6870
rect 6245 6852 6325 6868
rect 6245 6830 6264 6852
rect 6279 6836 6309 6852
rect 6337 6846 6343 6920
rect 6346 6846 6365 6990
rect 6380 6846 6386 6990
rect 6395 6920 6408 6990
rect 6460 6986 6482 6990
rect 6453 6964 6482 6978
rect 6535 6964 6551 6978
rect 6589 6974 6595 6976
rect 6602 6974 6710 6990
rect 6717 6974 6723 6976
rect 6731 6974 6746 6990
rect 6812 6984 6831 6987
rect 6453 6962 6551 6964
rect 6578 6962 6746 6974
rect 6761 6964 6777 6978
rect 6812 6965 6834 6984
rect 6844 6978 6860 6979
rect 6843 6976 6860 6978
rect 6844 6971 6860 6976
rect 6834 6964 6840 6965
rect 6843 6964 6872 6971
rect 6761 6963 6872 6964
rect 6761 6962 6878 6963
rect 6437 6954 6488 6962
rect 6535 6954 6569 6962
rect 6437 6942 6462 6954
rect 6469 6942 6488 6954
rect 6542 6952 6569 6954
rect 6578 6952 6799 6962
rect 6834 6959 6840 6962
rect 6542 6948 6799 6952
rect 6437 6934 6488 6942
rect 6535 6934 6799 6948
rect 6843 6954 6878 6962
rect 6389 6886 6408 6920
rect 6453 6926 6482 6934
rect 6453 6920 6470 6926
rect 6453 6918 6487 6920
rect 6535 6918 6551 6934
rect 6552 6924 6760 6934
rect 6761 6924 6777 6934
rect 6825 6930 6840 6945
rect 6843 6942 6844 6954
rect 6851 6942 6878 6954
rect 6843 6934 6878 6942
rect 6843 6933 6872 6934
rect 6563 6920 6777 6924
rect 6578 6918 6777 6920
rect 6812 6920 6825 6930
rect 6843 6920 6860 6933
rect 6812 6918 6860 6920
rect 6454 6914 6487 6918
rect 6450 6912 6487 6914
rect 6450 6911 6517 6912
rect 6450 6906 6481 6911
rect 6487 6906 6517 6911
rect 6450 6902 6517 6906
rect 6423 6899 6517 6902
rect 6423 6892 6472 6899
rect 6423 6886 6453 6892
rect 6472 6887 6477 6892
rect 6389 6870 6469 6886
rect 6481 6878 6517 6899
rect 6578 6894 6767 6918
rect 6812 6917 6859 6918
rect 6825 6912 6859 6917
rect 6593 6891 6767 6894
rect 6586 6888 6767 6891
rect 6795 6911 6859 6912
rect 6389 6868 6408 6870
rect 6423 6868 6457 6870
rect 6389 6852 6469 6868
rect 6389 6846 6408 6852
rect 6105 6820 6208 6830
rect 6059 6818 6208 6820
rect 6229 6818 6264 6830
rect 5898 6816 6060 6818
rect 5910 6796 5929 6816
rect 5944 6814 5974 6816
rect 5793 6788 5834 6796
rect 5916 6792 5929 6796
rect 5981 6800 6060 6816
rect 6092 6816 6264 6818
rect 6092 6800 6171 6816
rect 6178 6814 6208 6816
rect 5756 6778 5785 6788
rect 5799 6778 5828 6788
rect 5843 6778 5873 6792
rect 5916 6778 5959 6792
rect 5981 6788 6171 6800
rect 6236 6796 6242 6816
rect 5966 6778 5996 6788
rect 5997 6778 6155 6788
rect 6159 6778 6189 6788
rect 6193 6778 6223 6792
rect 6251 6778 6264 6816
rect 6336 6830 6365 6846
rect 6379 6830 6408 6846
rect 6423 6836 6453 6852
rect 6481 6830 6487 6878
rect 6490 6872 6509 6878
rect 6524 6872 6554 6880
rect 6490 6864 6554 6872
rect 6490 6848 6570 6864
rect 6586 6857 6648 6888
rect 6664 6857 6726 6888
rect 6795 6886 6844 6911
rect 6859 6886 6889 6902
rect 6758 6872 6788 6880
rect 6795 6878 6905 6886
rect 6758 6864 6803 6872
rect 6490 6846 6509 6848
rect 6524 6846 6570 6848
rect 6490 6830 6570 6846
rect 6597 6844 6632 6857
rect 6673 6854 6710 6857
rect 6673 6852 6715 6854
rect 6602 6841 6632 6844
rect 6611 6837 6618 6841
rect 6618 6836 6619 6837
rect 6577 6830 6587 6836
rect 6336 6822 6371 6830
rect 6336 6796 6337 6822
rect 6344 6796 6371 6822
rect 6279 6778 6309 6792
rect 6336 6788 6371 6796
rect 6373 6822 6414 6830
rect 6373 6796 6388 6822
rect 6395 6796 6414 6822
rect 6478 6818 6509 6830
rect 6524 6818 6627 6830
rect 6639 6820 6665 6846
rect 6680 6841 6710 6852
rect 6742 6848 6804 6864
rect 6742 6846 6788 6848
rect 6742 6830 6804 6846
rect 6816 6830 6822 6878
rect 6825 6870 6905 6878
rect 6825 6868 6844 6870
rect 6859 6868 6893 6870
rect 6825 6852 6905 6868
rect 6825 6830 6844 6852
rect 6859 6836 6889 6852
rect 6917 6846 6923 6920
rect 6926 6846 6945 6990
rect 6960 6846 6966 6990
rect 6975 6920 6988 6990
rect 7040 6986 7062 6990
rect 7033 6964 7062 6978
rect 7115 6964 7131 6978
rect 7169 6974 7175 6976
rect 7182 6974 7290 6990
rect 7297 6974 7303 6976
rect 7311 6974 7326 6990
rect 7392 6984 7411 6987
rect 7033 6962 7131 6964
rect 7158 6962 7326 6974
rect 7341 6964 7357 6978
rect 7392 6965 7414 6984
rect 7424 6978 7440 6979
rect 7423 6976 7440 6978
rect 7424 6971 7440 6976
rect 7414 6964 7420 6965
rect 7423 6964 7452 6971
rect 7341 6963 7452 6964
rect 7341 6962 7458 6963
rect 7017 6954 7068 6962
rect 7115 6954 7149 6962
rect 7017 6942 7042 6954
rect 7049 6942 7068 6954
rect 7122 6952 7149 6954
rect 7158 6952 7379 6962
rect 7414 6959 7420 6962
rect 7122 6948 7379 6952
rect 7017 6934 7068 6942
rect 7115 6934 7379 6948
rect 7423 6954 7458 6962
rect 6969 6886 6988 6920
rect 7033 6926 7062 6934
rect 7033 6920 7050 6926
rect 7033 6918 7067 6920
rect 7115 6918 7131 6934
rect 7132 6924 7340 6934
rect 7341 6924 7357 6934
rect 7405 6930 7420 6945
rect 7423 6942 7424 6954
rect 7431 6942 7458 6954
rect 7423 6934 7458 6942
rect 7423 6933 7452 6934
rect 7143 6920 7357 6924
rect 7158 6918 7357 6920
rect 7392 6920 7405 6930
rect 7423 6920 7440 6933
rect 7392 6918 7440 6920
rect 7034 6914 7067 6918
rect 7030 6912 7067 6914
rect 7030 6911 7097 6912
rect 7030 6906 7061 6911
rect 7067 6906 7097 6911
rect 7030 6902 7097 6906
rect 7003 6899 7097 6902
rect 7003 6892 7052 6899
rect 7003 6886 7033 6892
rect 7052 6887 7057 6892
rect 6969 6870 7049 6886
rect 7061 6878 7097 6899
rect 7158 6894 7347 6918
rect 7392 6917 7439 6918
rect 7405 6912 7439 6917
rect 7173 6891 7347 6894
rect 7166 6888 7347 6891
rect 7375 6911 7439 6912
rect 6969 6868 6988 6870
rect 7003 6868 7037 6870
rect 6969 6852 7049 6868
rect 6969 6846 6988 6852
rect 6685 6820 6788 6830
rect 6639 6818 6788 6820
rect 6809 6818 6844 6830
rect 6478 6816 6640 6818
rect 6490 6796 6509 6816
rect 6524 6814 6554 6816
rect 6373 6788 6414 6796
rect 6496 6792 6509 6796
rect 6561 6800 6640 6816
rect 6672 6816 6844 6818
rect 6672 6800 6751 6816
rect 6758 6814 6788 6816
rect 6336 6778 6365 6788
rect 6379 6778 6408 6788
rect 6423 6778 6453 6792
rect 6496 6778 6539 6792
rect 6561 6788 6751 6800
rect 6816 6796 6822 6816
rect 6546 6778 6576 6788
rect 6577 6778 6735 6788
rect 6739 6778 6769 6788
rect 6773 6778 6803 6792
rect 6831 6778 6844 6816
rect 6916 6830 6945 6846
rect 6959 6830 6988 6846
rect 7003 6836 7033 6852
rect 7061 6830 7067 6878
rect 7070 6872 7089 6878
rect 7104 6872 7134 6880
rect 7070 6864 7134 6872
rect 7070 6848 7150 6864
rect 7166 6857 7228 6888
rect 7244 6857 7306 6888
rect 7375 6886 7424 6911
rect 7439 6886 7469 6902
rect 7338 6872 7368 6880
rect 7375 6878 7485 6886
rect 7338 6864 7383 6872
rect 7070 6846 7089 6848
rect 7104 6846 7150 6848
rect 7070 6830 7150 6846
rect 7177 6844 7212 6857
rect 7253 6854 7290 6857
rect 7253 6852 7295 6854
rect 7182 6841 7212 6844
rect 7191 6837 7198 6841
rect 7198 6836 7199 6837
rect 7157 6830 7167 6836
rect 6916 6822 6951 6830
rect 6916 6796 6917 6822
rect 6924 6796 6951 6822
rect 6859 6778 6889 6792
rect 6916 6788 6951 6796
rect 6953 6822 6994 6830
rect 6953 6796 6968 6822
rect 6975 6796 6994 6822
rect 7058 6818 7089 6830
rect 7104 6818 7207 6830
rect 7219 6820 7245 6846
rect 7260 6841 7290 6852
rect 7322 6848 7384 6864
rect 7322 6846 7368 6848
rect 7322 6830 7384 6846
rect 7396 6830 7402 6878
rect 7405 6870 7485 6878
rect 7405 6868 7424 6870
rect 7439 6868 7473 6870
rect 7405 6852 7485 6868
rect 7405 6830 7424 6852
rect 7439 6836 7469 6852
rect 7497 6846 7503 6920
rect 7506 6846 7525 6990
rect 7540 6846 7546 6990
rect 7555 6920 7568 6990
rect 7620 6986 7642 6990
rect 7613 6964 7642 6978
rect 7695 6964 7711 6978
rect 7749 6974 7755 6976
rect 7762 6974 7870 6990
rect 7877 6974 7883 6976
rect 7891 6974 7906 6990
rect 7972 6984 7991 6987
rect 7613 6962 7711 6964
rect 7738 6962 7906 6974
rect 7921 6964 7937 6978
rect 7972 6965 7994 6984
rect 8004 6978 8020 6979
rect 8003 6976 8020 6978
rect 8004 6971 8020 6976
rect 7994 6964 8000 6965
rect 8003 6964 8032 6971
rect 7921 6963 8032 6964
rect 7921 6962 8038 6963
rect 7597 6954 7648 6962
rect 7695 6954 7729 6962
rect 7597 6942 7622 6954
rect 7629 6942 7648 6954
rect 7702 6952 7729 6954
rect 7738 6952 7959 6962
rect 7994 6959 8000 6962
rect 7702 6948 7959 6952
rect 7597 6934 7648 6942
rect 7695 6934 7959 6948
rect 8003 6954 8038 6962
rect 7549 6886 7568 6920
rect 7613 6926 7642 6934
rect 7613 6920 7630 6926
rect 7613 6918 7647 6920
rect 7695 6918 7711 6934
rect 7712 6924 7920 6934
rect 7921 6924 7937 6934
rect 7985 6930 8000 6945
rect 8003 6942 8004 6954
rect 8011 6942 8038 6954
rect 8003 6934 8038 6942
rect 8003 6933 8032 6934
rect 7723 6920 7937 6924
rect 7738 6918 7937 6920
rect 7972 6920 7985 6930
rect 8003 6920 8020 6933
rect 7972 6918 8020 6920
rect 7614 6914 7647 6918
rect 7610 6912 7647 6914
rect 7610 6911 7677 6912
rect 7610 6906 7641 6911
rect 7647 6906 7677 6911
rect 7610 6902 7677 6906
rect 7583 6899 7677 6902
rect 7583 6892 7632 6899
rect 7583 6886 7613 6892
rect 7632 6887 7637 6892
rect 7549 6870 7629 6886
rect 7641 6878 7677 6899
rect 7738 6894 7927 6918
rect 7972 6917 8019 6918
rect 7985 6912 8019 6917
rect 7753 6891 7927 6894
rect 7746 6888 7927 6891
rect 7955 6911 8019 6912
rect 7549 6868 7568 6870
rect 7583 6868 7617 6870
rect 7549 6852 7629 6868
rect 7549 6846 7568 6852
rect 7265 6820 7368 6830
rect 7219 6818 7368 6820
rect 7389 6818 7424 6830
rect 7058 6816 7220 6818
rect 7070 6796 7089 6816
rect 7104 6814 7134 6816
rect 6953 6788 6994 6796
rect 7076 6792 7089 6796
rect 7141 6800 7220 6816
rect 7252 6816 7424 6818
rect 7252 6800 7331 6816
rect 7338 6814 7368 6816
rect 6916 6778 6945 6788
rect 6959 6778 6988 6788
rect 7003 6778 7033 6792
rect 7076 6778 7119 6792
rect 7141 6788 7331 6800
rect 7396 6796 7402 6816
rect 7126 6778 7156 6788
rect 7157 6778 7315 6788
rect 7319 6778 7349 6788
rect 7353 6778 7383 6792
rect 7411 6778 7424 6816
rect 7496 6830 7525 6846
rect 7539 6830 7568 6846
rect 7583 6836 7613 6852
rect 7641 6830 7647 6878
rect 7650 6872 7669 6878
rect 7684 6872 7714 6880
rect 7650 6864 7714 6872
rect 7650 6848 7730 6864
rect 7746 6857 7808 6888
rect 7824 6857 7886 6888
rect 7955 6886 8004 6911
rect 8019 6886 8049 6902
rect 7918 6872 7948 6880
rect 7955 6878 8065 6886
rect 7918 6864 7963 6872
rect 7650 6846 7669 6848
rect 7684 6846 7730 6848
rect 7650 6830 7730 6846
rect 7757 6844 7792 6857
rect 7833 6854 7870 6857
rect 7833 6852 7875 6854
rect 7762 6841 7792 6844
rect 7771 6837 7778 6841
rect 7778 6836 7779 6837
rect 7737 6830 7747 6836
rect 7496 6822 7531 6830
rect 7496 6796 7497 6822
rect 7504 6796 7531 6822
rect 7439 6778 7469 6792
rect 7496 6788 7531 6796
rect 7533 6822 7574 6830
rect 7533 6796 7548 6822
rect 7555 6796 7574 6822
rect 7638 6818 7669 6830
rect 7684 6818 7787 6830
rect 7799 6820 7825 6846
rect 7840 6841 7870 6852
rect 7902 6848 7964 6864
rect 7902 6846 7948 6848
rect 7902 6830 7964 6846
rect 7976 6830 7982 6878
rect 7985 6870 8065 6878
rect 7985 6868 8004 6870
rect 8019 6868 8053 6870
rect 7985 6852 8065 6868
rect 7985 6830 8004 6852
rect 8019 6836 8049 6852
rect 8077 6846 8083 6920
rect 8086 6846 8105 6990
rect 8120 6846 8126 6990
rect 8135 6920 8148 6990
rect 8200 6986 8222 6990
rect 8193 6964 8222 6978
rect 8275 6964 8291 6978
rect 8329 6974 8335 6976
rect 8342 6974 8450 6990
rect 8457 6974 8463 6976
rect 8471 6974 8486 6990
rect 8552 6984 8571 6987
rect 8193 6962 8291 6964
rect 8318 6962 8486 6974
rect 8501 6964 8517 6978
rect 8552 6965 8574 6984
rect 8584 6978 8600 6979
rect 8583 6976 8600 6978
rect 8584 6971 8600 6976
rect 8574 6964 8580 6965
rect 8583 6964 8612 6971
rect 8501 6963 8612 6964
rect 8501 6962 8618 6963
rect 8177 6954 8228 6962
rect 8275 6954 8309 6962
rect 8177 6942 8202 6954
rect 8209 6942 8228 6954
rect 8282 6952 8309 6954
rect 8318 6952 8539 6962
rect 8574 6959 8580 6962
rect 8282 6948 8539 6952
rect 8177 6934 8228 6942
rect 8275 6934 8539 6948
rect 8583 6954 8618 6962
rect 8129 6886 8148 6920
rect 8193 6926 8222 6934
rect 8193 6920 8210 6926
rect 8193 6918 8227 6920
rect 8275 6918 8291 6934
rect 8292 6924 8500 6934
rect 8501 6924 8517 6934
rect 8565 6930 8580 6945
rect 8583 6942 8584 6954
rect 8591 6942 8618 6954
rect 8583 6934 8618 6942
rect 8583 6933 8612 6934
rect 8303 6920 8517 6924
rect 8318 6918 8517 6920
rect 8552 6920 8565 6930
rect 8583 6920 8600 6933
rect 8552 6918 8600 6920
rect 8194 6914 8227 6918
rect 8190 6912 8227 6914
rect 8190 6911 8257 6912
rect 8190 6906 8221 6911
rect 8227 6906 8257 6911
rect 8190 6902 8257 6906
rect 8163 6899 8257 6902
rect 8163 6892 8212 6899
rect 8163 6886 8193 6892
rect 8212 6887 8217 6892
rect 8129 6870 8209 6886
rect 8221 6878 8257 6899
rect 8318 6894 8507 6918
rect 8552 6917 8599 6918
rect 8565 6912 8599 6917
rect 8333 6891 8507 6894
rect 8326 6888 8507 6891
rect 8535 6911 8599 6912
rect 8129 6868 8148 6870
rect 8163 6868 8197 6870
rect 8129 6852 8209 6868
rect 8129 6846 8148 6852
rect 7845 6820 7948 6830
rect 7799 6818 7948 6820
rect 7969 6818 8004 6830
rect 7638 6816 7800 6818
rect 7650 6796 7669 6816
rect 7684 6814 7714 6816
rect 7533 6788 7574 6796
rect 7656 6792 7669 6796
rect 7721 6800 7800 6816
rect 7832 6816 8004 6818
rect 7832 6800 7911 6816
rect 7918 6814 7948 6816
rect 7496 6778 7525 6788
rect 7539 6778 7568 6788
rect 7583 6778 7613 6792
rect 7656 6778 7699 6792
rect 7721 6788 7911 6800
rect 7976 6796 7982 6816
rect 7706 6778 7736 6788
rect 7737 6778 7895 6788
rect 7899 6778 7929 6788
rect 7933 6778 7963 6792
rect 7991 6778 8004 6816
rect 8076 6830 8105 6846
rect 8119 6830 8148 6846
rect 8163 6836 8193 6852
rect 8221 6830 8227 6878
rect 8230 6872 8249 6878
rect 8264 6872 8294 6880
rect 8230 6864 8294 6872
rect 8230 6848 8310 6864
rect 8326 6857 8388 6888
rect 8404 6857 8466 6888
rect 8535 6886 8584 6911
rect 8599 6886 8629 6902
rect 8498 6872 8528 6880
rect 8535 6878 8645 6886
rect 8498 6864 8543 6872
rect 8230 6846 8249 6848
rect 8264 6846 8310 6848
rect 8230 6830 8310 6846
rect 8337 6844 8372 6857
rect 8413 6854 8450 6857
rect 8413 6852 8455 6854
rect 8342 6841 8372 6844
rect 8351 6837 8358 6841
rect 8358 6836 8359 6837
rect 8317 6830 8327 6836
rect 8076 6822 8111 6830
rect 8076 6796 8077 6822
rect 8084 6796 8111 6822
rect 8019 6778 8049 6792
rect 8076 6788 8111 6796
rect 8113 6822 8154 6830
rect 8113 6796 8128 6822
rect 8135 6796 8154 6822
rect 8218 6818 8249 6830
rect 8264 6818 8367 6830
rect 8379 6820 8405 6846
rect 8420 6841 8450 6852
rect 8482 6848 8544 6864
rect 8482 6846 8528 6848
rect 8482 6830 8544 6846
rect 8556 6830 8562 6878
rect 8565 6870 8645 6878
rect 8565 6868 8584 6870
rect 8599 6868 8633 6870
rect 8565 6852 8645 6868
rect 8565 6830 8584 6852
rect 8599 6836 8629 6852
rect 8657 6846 8663 6920
rect 8666 6846 8685 6990
rect 8700 6846 8706 6990
rect 8715 6920 8728 6990
rect 8780 6986 8802 6990
rect 8773 6964 8802 6978
rect 8855 6964 8871 6978
rect 8909 6974 8915 6976
rect 8922 6974 9030 6990
rect 9037 6974 9043 6976
rect 9051 6974 9066 6990
rect 9132 6984 9151 6987
rect 8773 6962 8871 6964
rect 8898 6962 9066 6974
rect 9081 6964 9097 6978
rect 9132 6965 9154 6984
rect 9164 6978 9180 6979
rect 9163 6976 9180 6978
rect 9164 6971 9180 6976
rect 9154 6964 9160 6965
rect 9163 6964 9192 6971
rect 9081 6963 9192 6964
rect 9081 6962 9198 6963
rect 8757 6954 8808 6962
rect 8855 6954 8889 6962
rect 8757 6942 8782 6954
rect 8789 6942 8808 6954
rect 8862 6952 8889 6954
rect 8898 6952 9119 6962
rect 9154 6959 9160 6962
rect 8862 6948 9119 6952
rect 8757 6934 8808 6942
rect 8855 6934 9119 6948
rect 9163 6954 9198 6962
rect 8709 6886 8728 6920
rect 8773 6926 8802 6934
rect 8773 6920 8790 6926
rect 8773 6918 8807 6920
rect 8855 6918 8871 6934
rect 8872 6924 9080 6934
rect 9081 6924 9097 6934
rect 9145 6930 9160 6945
rect 9163 6942 9164 6954
rect 9171 6942 9198 6954
rect 9163 6934 9198 6942
rect 9163 6933 9192 6934
rect 8883 6920 9097 6924
rect 8898 6918 9097 6920
rect 9132 6920 9145 6930
rect 9163 6920 9180 6933
rect 9132 6918 9180 6920
rect 8774 6914 8807 6918
rect 8770 6912 8807 6914
rect 8770 6911 8837 6912
rect 8770 6906 8801 6911
rect 8807 6906 8837 6911
rect 8770 6902 8837 6906
rect 8743 6899 8837 6902
rect 8743 6892 8792 6899
rect 8743 6886 8773 6892
rect 8792 6887 8797 6892
rect 8709 6870 8789 6886
rect 8801 6878 8837 6899
rect 8898 6894 9087 6918
rect 9132 6917 9179 6918
rect 9145 6912 9179 6917
rect 8913 6891 9087 6894
rect 8906 6888 9087 6891
rect 9115 6911 9179 6912
rect 8709 6868 8728 6870
rect 8743 6868 8777 6870
rect 8709 6852 8789 6868
rect 8709 6846 8728 6852
rect 8425 6820 8528 6830
rect 8379 6818 8528 6820
rect 8549 6818 8584 6830
rect 8218 6816 8380 6818
rect 8230 6796 8249 6816
rect 8264 6814 8294 6816
rect 8113 6788 8154 6796
rect 8236 6792 8249 6796
rect 8301 6800 8380 6816
rect 8412 6816 8584 6818
rect 8412 6800 8491 6816
rect 8498 6814 8528 6816
rect 8076 6778 8105 6788
rect 8119 6778 8148 6788
rect 8163 6778 8193 6792
rect 8236 6778 8279 6792
rect 8301 6788 8491 6800
rect 8556 6796 8562 6816
rect 8286 6778 8316 6788
rect 8317 6778 8475 6788
rect 8479 6778 8509 6788
rect 8513 6778 8543 6792
rect 8571 6778 8584 6816
rect 8656 6830 8685 6846
rect 8699 6830 8728 6846
rect 8743 6836 8773 6852
rect 8801 6830 8807 6878
rect 8810 6872 8829 6878
rect 8844 6872 8874 6880
rect 8810 6864 8874 6872
rect 8810 6848 8890 6864
rect 8906 6857 8968 6888
rect 8984 6857 9046 6888
rect 9115 6886 9164 6911
rect 9179 6886 9209 6902
rect 9078 6872 9108 6880
rect 9115 6878 9225 6886
rect 9078 6864 9123 6872
rect 8810 6846 8829 6848
rect 8844 6846 8890 6848
rect 8810 6830 8890 6846
rect 8917 6844 8952 6857
rect 8993 6854 9030 6857
rect 8993 6852 9035 6854
rect 8922 6841 8952 6844
rect 8931 6837 8938 6841
rect 8938 6836 8939 6837
rect 8897 6830 8907 6836
rect 8656 6822 8691 6830
rect 8656 6796 8657 6822
rect 8664 6796 8691 6822
rect 8599 6778 8629 6792
rect 8656 6788 8691 6796
rect 8693 6822 8734 6830
rect 8693 6796 8708 6822
rect 8715 6796 8734 6822
rect 8798 6818 8829 6830
rect 8844 6818 8947 6830
rect 8959 6820 8985 6846
rect 9000 6841 9030 6852
rect 9062 6848 9124 6864
rect 9062 6846 9108 6848
rect 9062 6830 9124 6846
rect 9136 6830 9142 6878
rect 9145 6870 9225 6878
rect 9145 6868 9164 6870
rect 9179 6868 9213 6870
rect 9145 6852 9225 6868
rect 9145 6830 9164 6852
rect 9179 6836 9209 6852
rect 9237 6846 9243 6920
rect 9246 6846 9265 6990
rect 9280 6846 9286 6990
rect 9295 6920 9308 6990
rect 9360 6986 9382 6990
rect 9353 6964 9382 6978
rect 9435 6964 9451 6978
rect 9489 6974 9495 6976
rect 9502 6974 9610 6990
rect 9617 6974 9623 6976
rect 9631 6974 9646 6990
rect 9712 6984 9731 6987
rect 9353 6962 9451 6964
rect 9478 6962 9646 6974
rect 9661 6964 9677 6978
rect 9712 6965 9734 6984
rect 9744 6978 9760 6979
rect 9743 6976 9760 6978
rect 9744 6971 9760 6976
rect 9734 6964 9740 6965
rect 9743 6964 9772 6971
rect 9661 6963 9772 6964
rect 9661 6962 9778 6963
rect 9337 6954 9388 6962
rect 9435 6954 9469 6962
rect 9337 6942 9362 6954
rect 9369 6942 9388 6954
rect 9442 6952 9469 6954
rect 9478 6952 9699 6962
rect 9734 6959 9740 6962
rect 9442 6948 9699 6952
rect 9337 6934 9388 6942
rect 9435 6934 9699 6948
rect 9743 6954 9778 6962
rect 9289 6886 9308 6920
rect 9353 6926 9382 6934
rect 9353 6920 9370 6926
rect 9353 6918 9387 6920
rect 9435 6918 9451 6934
rect 9452 6924 9660 6934
rect 9661 6924 9677 6934
rect 9725 6930 9740 6945
rect 9743 6942 9744 6954
rect 9751 6942 9778 6954
rect 9743 6934 9778 6942
rect 9743 6933 9772 6934
rect 9463 6920 9677 6924
rect 9478 6918 9677 6920
rect 9712 6920 9725 6930
rect 9743 6920 9760 6933
rect 9712 6918 9760 6920
rect 9354 6914 9387 6918
rect 9350 6912 9387 6914
rect 9350 6911 9417 6912
rect 9350 6906 9381 6911
rect 9387 6906 9417 6911
rect 9350 6902 9417 6906
rect 9323 6899 9417 6902
rect 9323 6892 9372 6899
rect 9323 6886 9353 6892
rect 9372 6887 9377 6892
rect 9289 6870 9369 6886
rect 9381 6878 9417 6899
rect 9478 6894 9667 6918
rect 9712 6917 9759 6918
rect 9725 6912 9759 6917
rect 9493 6891 9667 6894
rect 9486 6888 9667 6891
rect 9695 6911 9759 6912
rect 9289 6868 9308 6870
rect 9323 6868 9357 6870
rect 9289 6852 9369 6868
rect 9289 6846 9308 6852
rect 9005 6820 9108 6830
rect 8959 6818 9108 6820
rect 9129 6818 9164 6830
rect 8798 6816 8960 6818
rect 8810 6796 8829 6816
rect 8844 6814 8874 6816
rect 8693 6788 8734 6796
rect 8816 6792 8829 6796
rect 8881 6800 8960 6816
rect 8992 6816 9164 6818
rect 8992 6800 9071 6816
rect 9078 6814 9108 6816
rect 8656 6778 8685 6788
rect 8699 6778 8728 6788
rect 8743 6778 8773 6792
rect 8816 6778 8859 6792
rect 8881 6788 9071 6800
rect 9136 6796 9142 6816
rect 8866 6778 8896 6788
rect 8897 6778 9055 6788
rect 9059 6778 9089 6788
rect 9093 6778 9123 6792
rect 9151 6778 9164 6816
rect 9236 6830 9265 6846
rect 9279 6830 9308 6846
rect 9323 6836 9353 6852
rect 9381 6830 9387 6878
rect 9390 6872 9409 6878
rect 9424 6872 9454 6880
rect 9390 6864 9454 6872
rect 9390 6848 9470 6864
rect 9486 6857 9548 6888
rect 9564 6857 9626 6888
rect 9695 6886 9744 6911
rect 9759 6886 9789 6902
rect 9658 6872 9688 6880
rect 9695 6878 9805 6886
rect 9658 6864 9703 6872
rect 9390 6846 9409 6848
rect 9424 6846 9470 6848
rect 9390 6830 9470 6846
rect 9497 6844 9532 6857
rect 9573 6854 9610 6857
rect 9573 6852 9615 6854
rect 9502 6841 9532 6844
rect 9511 6837 9518 6841
rect 9518 6836 9519 6837
rect 9477 6830 9487 6836
rect 9236 6822 9271 6830
rect 9236 6796 9237 6822
rect 9244 6796 9271 6822
rect 9179 6778 9209 6792
rect 9236 6788 9271 6796
rect 9273 6822 9314 6830
rect 9273 6796 9288 6822
rect 9295 6796 9314 6822
rect 9378 6818 9409 6830
rect 9424 6818 9527 6830
rect 9539 6820 9565 6846
rect 9580 6841 9610 6852
rect 9642 6848 9704 6864
rect 9642 6846 9688 6848
rect 9642 6830 9704 6846
rect 9716 6830 9722 6878
rect 9725 6870 9805 6878
rect 9725 6868 9744 6870
rect 9759 6868 9793 6870
rect 9725 6852 9805 6868
rect 9725 6830 9744 6852
rect 9759 6836 9789 6852
rect 9817 6846 9823 6920
rect 9826 6846 9845 6990
rect 9860 6846 9866 6990
rect 9875 6920 9888 6990
rect 9940 6986 9962 6990
rect 9933 6964 9962 6978
rect 10015 6964 10031 6978
rect 10069 6974 10075 6976
rect 10082 6974 10190 6990
rect 10197 6974 10203 6976
rect 10211 6974 10226 6990
rect 10292 6984 10311 6987
rect 9933 6962 10031 6964
rect 10058 6962 10226 6974
rect 10241 6964 10257 6978
rect 10292 6965 10314 6984
rect 10324 6978 10340 6979
rect 10323 6976 10340 6978
rect 10324 6971 10340 6976
rect 10314 6964 10320 6965
rect 10323 6964 10352 6971
rect 10241 6963 10352 6964
rect 10241 6962 10358 6963
rect 9917 6954 9968 6962
rect 10015 6954 10049 6962
rect 9917 6942 9942 6954
rect 9949 6942 9968 6954
rect 10022 6952 10049 6954
rect 10058 6952 10279 6962
rect 10314 6959 10320 6962
rect 10022 6948 10279 6952
rect 9917 6934 9968 6942
rect 10015 6934 10279 6948
rect 10323 6954 10358 6962
rect 9869 6886 9888 6920
rect 9933 6926 9962 6934
rect 9933 6920 9950 6926
rect 9933 6918 9967 6920
rect 10015 6918 10031 6934
rect 10032 6924 10240 6934
rect 10241 6924 10257 6934
rect 10305 6930 10320 6945
rect 10323 6942 10324 6954
rect 10331 6942 10358 6954
rect 10323 6934 10358 6942
rect 10323 6933 10352 6934
rect 10043 6920 10257 6924
rect 10058 6918 10257 6920
rect 10292 6920 10305 6930
rect 10323 6920 10340 6933
rect 10292 6918 10340 6920
rect 9934 6914 9967 6918
rect 9930 6912 9967 6914
rect 9930 6911 9997 6912
rect 9930 6906 9961 6911
rect 9967 6906 9997 6911
rect 9930 6902 9997 6906
rect 9903 6899 9997 6902
rect 9903 6892 9952 6899
rect 9903 6886 9933 6892
rect 9952 6887 9957 6892
rect 9869 6870 9949 6886
rect 9961 6878 9997 6899
rect 10058 6894 10247 6918
rect 10292 6917 10339 6918
rect 10305 6912 10339 6917
rect 10073 6891 10247 6894
rect 10066 6888 10247 6891
rect 10275 6911 10339 6912
rect 9869 6868 9888 6870
rect 9903 6868 9937 6870
rect 9869 6852 9949 6868
rect 9869 6846 9888 6852
rect 9585 6820 9688 6830
rect 9539 6818 9688 6820
rect 9709 6818 9744 6830
rect 9378 6816 9540 6818
rect 9390 6796 9409 6816
rect 9424 6814 9454 6816
rect 9273 6788 9314 6796
rect 9396 6792 9409 6796
rect 9461 6800 9540 6816
rect 9572 6816 9744 6818
rect 9572 6800 9651 6816
rect 9658 6814 9688 6816
rect 9236 6778 9265 6788
rect 9279 6778 9308 6788
rect 9323 6778 9353 6792
rect 9396 6778 9439 6792
rect 9461 6788 9651 6800
rect 9716 6796 9722 6816
rect 9446 6778 9476 6788
rect 9477 6778 9635 6788
rect 9639 6778 9669 6788
rect 9673 6778 9703 6792
rect 9731 6778 9744 6816
rect 9816 6830 9845 6846
rect 9859 6830 9888 6846
rect 9903 6836 9933 6852
rect 9961 6830 9967 6878
rect 9970 6872 9989 6878
rect 10004 6872 10034 6880
rect 9970 6864 10034 6872
rect 9970 6848 10050 6864
rect 10066 6857 10128 6888
rect 10144 6857 10206 6888
rect 10275 6886 10324 6911
rect 10339 6886 10369 6902
rect 10238 6872 10268 6880
rect 10275 6878 10385 6886
rect 10238 6864 10283 6872
rect 9970 6846 9989 6848
rect 10004 6846 10050 6848
rect 9970 6830 10050 6846
rect 10077 6844 10112 6857
rect 10153 6854 10190 6857
rect 10153 6852 10195 6854
rect 10082 6841 10112 6844
rect 10091 6837 10098 6841
rect 10098 6836 10099 6837
rect 10057 6830 10067 6836
rect 9816 6822 9851 6830
rect 9816 6796 9817 6822
rect 9824 6796 9851 6822
rect 9759 6778 9789 6792
rect 9816 6788 9851 6796
rect 9853 6822 9894 6830
rect 9853 6796 9868 6822
rect 9875 6796 9894 6822
rect 9958 6818 9989 6830
rect 10004 6818 10107 6830
rect 10119 6820 10145 6846
rect 10160 6841 10190 6852
rect 10222 6848 10284 6864
rect 10222 6846 10268 6848
rect 10222 6830 10284 6846
rect 10296 6830 10302 6878
rect 10305 6870 10385 6878
rect 10305 6868 10324 6870
rect 10339 6868 10373 6870
rect 10305 6852 10385 6868
rect 10305 6830 10324 6852
rect 10339 6836 10369 6852
rect 10397 6846 10403 6920
rect 10406 6846 10425 6990
rect 10440 6846 10446 6990
rect 10455 6920 10468 6990
rect 10520 6986 10542 6990
rect 10513 6964 10542 6978
rect 10595 6964 10611 6978
rect 10649 6974 10655 6976
rect 10662 6974 10770 6990
rect 10777 6974 10783 6976
rect 10791 6974 10806 6990
rect 10872 6984 10891 6987
rect 10513 6962 10611 6964
rect 10638 6962 10806 6974
rect 10821 6964 10837 6978
rect 10872 6965 10894 6984
rect 10904 6978 10920 6979
rect 10903 6976 10920 6978
rect 10904 6971 10920 6976
rect 10894 6964 10900 6965
rect 10903 6964 10932 6971
rect 10821 6963 10932 6964
rect 10821 6962 10938 6963
rect 10497 6954 10548 6962
rect 10595 6954 10629 6962
rect 10497 6942 10522 6954
rect 10529 6942 10548 6954
rect 10602 6952 10629 6954
rect 10638 6952 10859 6962
rect 10894 6959 10900 6962
rect 10602 6948 10859 6952
rect 10497 6934 10548 6942
rect 10595 6934 10859 6948
rect 10903 6954 10938 6962
rect 10449 6886 10468 6920
rect 10513 6926 10542 6934
rect 10513 6920 10530 6926
rect 10513 6918 10547 6920
rect 10595 6918 10611 6934
rect 10612 6924 10820 6934
rect 10821 6924 10837 6934
rect 10885 6930 10900 6945
rect 10903 6942 10904 6954
rect 10911 6942 10938 6954
rect 10903 6934 10938 6942
rect 10903 6933 10932 6934
rect 10623 6920 10837 6924
rect 10638 6918 10837 6920
rect 10872 6920 10885 6930
rect 10903 6920 10920 6933
rect 10872 6918 10920 6920
rect 10514 6914 10547 6918
rect 10510 6912 10547 6914
rect 10510 6911 10577 6912
rect 10510 6906 10541 6911
rect 10547 6906 10577 6911
rect 10510 6902 10577 6906
rect 10483 6899 10577 6902
rect 10483 6892 10532 6899
rect 10483 6886 10513 6892
rect 10532 6887 10537 6892
rect 10449 6870 10529 6886
rect 10541 6878 10577 6899
rect 10638 6894 10827 6918
rect 10872 6917 10919 6918
rect 10885 6912 10919 6917
rect 10653 6891 10827 6894
rect 10646 6888 10827 6891
rect 10855 6911 10919 6912
rect 10449 6868 10468 6870
rect 10483 6868 10517 6870
rect 10449 6852 10529 6868
rect 10449 6846 10468 6852
rect 10165 6820 10268 6830
rect 10119 6818 10268 6820
rect 10289 6818 10324 6830
rect 9958 6816 10120 6818
rect 9970 6796 9989 6816
rect 10004 6814 10034 6816
rect 9853 6788 9894 6796
rect 9976 6792 9989 6796
rect 10041 6800 10120 6816
rect 10152 6816 10324 6818
rect 10152 6800 10231 6816
rect 10238 6814 10268 6816
rect 9816 6778 9845 6788
rect 9859 6778 9888 6788
rect 9903 6778 9933 6792
rect 9976 6778 10019 6792
rect 10041 6788 10231 6800
rect 10296 6796 10302 6816
rect 10026 6778 10056 6788
rect 10057 6778 10215 6788
rect 10219 6778 10249 6788
rect 10253 6778 10283 6792
rect 10311 6778 10324 6816
rect 10396 6830 10425 6846
rect 10439 6830 10468 6846
rect 10483 6836 10513 6852
rect 10541 6830 10547 6878
rect 10550 6872 10569 6878
rect 10584 6872 10614 6880
rect 10550 6864 10614 6872
rect 10550 6848 10630 6864
rect 10646 6857 10708 6888
rect 10724 6857 10786 6888
rect 10855 6886 10904 6911
rect 10919 6886 10949 6902
rect 10818 6872 10848 6880
rect 10855 6878 10965 6886
rect 10818 6864 10863 6872
rect 10550 6846 10569 6848
rect 10584 6846 10630 6848
rect 10550 6830 10630 6846
rect 10657 6844 10692 6857
rect 10733 6854 10770 6857
rect 10733 6852 10775 6854
rect 10662 6841 10692 6844
rect 10671 6837 10678 6841
rect 10678 6836 10679 6837
rect 10637 6830 10647 6836
rect 10396 6822 10431 6830
rect 10396 6796 10397 6822
rect 10404 6796 10431 6822
rect 10339 6778 10369 6792
rect 10396 6788 10431 6796
rect 10433 6822 10474 6830
rect 10433 6796 10448 6822
rect 10455 6796 10474 6822
rect 10538 6818 10569 6830
rect 10584 6818 10687 6830
rect 10699 6820 10725 6846
rect 10740 6841 10770 6852
rect 10802 6848 10864 6864
rect 10802 6846 10848 6848
rect 10802 6830 10864 6846
rect 10876 6830 10882 6878
rect 10885 6870 10965 6878
rect 10885 6868 10904 6870
rect 10919 6868 10953 6870
rect 10885 6852 10965 6868
rect 10885 6830 10904 6852
rect 10919 6836 10949 6852
rect 10977 6846 10983 6920
rect 10986 6846 11005 6990
rect 11020 6846 11026 6990
rect 11035 6920 11048 6990
rect 11100 6986 11122 6990
rect 11093 6964 11122 6978
rect 11175 6964 11191 6978
rect 11229 6974 11235 6976
rect 11242 6974 11350 6990
rect 11357 6974 11363 6976
rect 11371 6974 11386 6990
rect 11452 6984 11471 6987
rect 11093 6962 11191 6964
rect 11218 6962 11386 6974
rect 11401 6964 11417 6978
rect 11452 6965 11474 6984
rect 11484 6978 11500 6979
rect 11483 6976 11500 6978
rect 11484 6971 11500 6976
rect 11474 6964 11480 6965
rect 11483 6964 11512 6971
rect 11401 6963 11512 6964
rect 11401 6962 11518 6963
rect 11077 6954 11128 6962
rect 11175 6954 11209 6962
rect 11077 6942 11102 6954
rect 11109 6942 11128 6954
rect 11182 6952 11209 6954
rect 11218 6952 11439 6962
rect 11474 6959 11480 6962
rect 11182 6948 11439 6952
rect 11077 6934 11128 6942
rect 11175 6934 11439 6948
rect 11483 6954 11518 6962
rect 11029 6886 11048 6920
rect 11093 6926 11122 6934
rect 11093 6920 11110 6926
rect 11093 6918 11127 6920
rect 11175 6918 11191 6934
rect 11192 6924 11400 6934
rect 11401 6924 11417 6934
rect 11465 6930 11480 6945
rect 11483 6942 11484 6954
rect 11491 6942 11518 6954
rect 11483 6934 11518 6942
rect 11483 6933 11512 6934
rect 11203 6920 11417 6924
rect 11218 6918 11417 6920
rect 11452 6920 11465 6930
rect 11483 6920 11500 6933
rect 11452 6918 11500 6920
rect 11094 6914 11127 6918
rect 11090 6912 11127 6914
rect 11090 6911 11157 6912
rect 11090 6906 11121 6911
rect 11127 6906 11157 6911
rect 11090 6902 11157 6906
rect 11063 6899 11157 6902
rect 11063 6892 11112 6899
rect 11063 6886 11093 6892
rect 11112 6887 11117 6892
rect 11029 6870 11109 6886
rect 11121 6878 11157 6899
rect 11218 6894 11407 6918
rect 11452 6917 11499 6918
rect 11465 6912 11499 6917
rect 11233 6891 11407 6894
rect 11226 6888 11407 6891
rect 11435 6911 11499 6912
rect 11029 6868 11048 6870
rect 11063 6868 11097 6870
rect 11029 6852 11109 6868
rect 11029 6846 11048 6852
rect 10745 6820 10848 6830
rect 10699 6818 10848 6820
rect 10869 6818 10904 6830
rect 10538 6816 10700 6818
rect 10550 6796 10569 6816
rect 10584 6814 10614 6816
rect 10433 6788 10474 6796
rect 10556 6792 10569 6796
rect 10621 6800 10700 6816
rect 10732 6816 10904 6818
rect 10732 6800 10811 6816
rect 10818 6814 10848 6816
rect 10396 6778 10425 6788
rect 10439 6778 10468 6788
rect 10483 6778 10513 6792
rect 10556 6778 10599 6792
rect 10621 6788 10811 6800
rect 10876 6796 10882 6816
rect 10606 6778 10636 6788
rect 10637 6778 10795 6788
rect 10799 6778 10829 6788
rect 10833 6778 10863 6792
rect 10891 6778 10904 6816
rect 10976 6830 11005 6846
rect 11019 6830 11048 6846
rect 11063 6836 11093 6852
rect 11121 6830 11127 6878
rect 11130 6872 11149 6878
rect 11164 6872 11194 6880
rect 11130 6864 11194 6872
rect 11130 6848 11210 6864
rect 11226 6857 11288 6888
rect 11304 6857 11366 6888
rect 11435 6886 11484 6911
rect 11499 6886 11529 6902
rect 11398 6872 11428 6880
rect 11435 6878 11545 6886
rect 11398 6864 11443 6872
rect 11130 6846 11149 6848
rect 11164 6846 11210 6848
rect 11130 6830 11210 6846
rect 11237 6844 11272 6857
rect 11313 6854 11350 6857
rect 11313 6852 11355 6854
rect 11242 6841 11272 6844
rect 11251 6837 11258 6841
rect 11258 6836 11259 6837
rect 11217 6830 11227 6836
rect 10976 6822 11011 6830
rect 10976 6796 10977 6822
rect 10984 6796 11011 6822
rect 10919 6778 10949 6792
rect 10976 6788 11011 6796
rect 11013 6822 11054 6830
rect 11013 6796 11028 6822
rect 11035 6796 11054 6822
rect 11118 6818 11149 6830
rect 11164 6818 11267 6830
rect 11279 6820 11305 6846
rect 11320 6841 11350 6852
rect 11382 6848 11444 6864
rect 11382 6846 11428 6848
rect 11382 6830 11444 6846
rect 11456 6830 11462 6878
rect 11465 6870 11545 6878
rect 11465 6868 11484 6870
rect 11499 6868 11533 6870
rect 11465 6852 11545 6868
rect 11465 6830 11484 6852
rect 11499 6836 11529 6852
rect 11557 6846 11563 6920
rect 11566 6846 11585 6990
rect 11600 6846 11606 6990
rect 11615 6920 11628 6990
rect 11680 6986 11702 6990
rect 11673 6964 11702 6978
rect 11755 6964 11771 6978
rect 11809 6974 11815 6976
rect 11822 6974 11930 6990
rect 11937 6974 11943 6976
rect 11951 6974 11966 6990
rect 12032 6984 12051 6987
rect 11673 6962 11771 6964
rect 11798 6962 11966 6974
rect 11981 6964 11997 6978
rect 12032 6965 12054 6984
rect 12064 6978 12080 6979
rect 12063 6976 12080 6978
rect 12064 6971 12080 6976
rect 12054 6964 12060 6965
rect 12063 6964 12092 6971
rect 11981 6963 12092 6964
rect 11981 6962 12098 6963
rect 11657 6954 11708 6962
rect 11755 6954 11789 6962
rect 11657 6942 11682 6954
rect 11689 6942 11708 6954
rect 11762 6952 11789 6954
rect 11798 6952 12019 6962
rect 12054 6959 12060 6962
rect 11762 6948 12019 6952
rect 11657 6934 11708 6942
rect 11755 6934 12019 6948
rect 12063 6954 12098 6962
rect 11609 6886 11628 6920
rect 11673 6926 11702 6934
rect 11673 6920 11690 6926
rect 11673 6918 11707 6920
rect 11755 6918 11771 6934
rect 11772 6924 11980 6934
rect 11981 6924 11997 6934
rect 12045 6930 12060 6945
rect 12063 6942 12064 6954
rect 12071 6942 12098 6954
rect 12063 6934 12098 6942
rect 12063 6933 12092 6934
rect 11783 6920 11997 6924
rect 11798 6918 11997 6920
rect 12032 6920 12045 6930
rect 12063 6920 12080 6933
rect 12032 6918 12080 6920
rect 11674 6914 11707 6918
rect 11670 6912 11707 6914
rect 11670 6911 11737 6912
rect 11670 6906 11701 6911
rect 11707 6906 11737 6911
rect 11670 6902 11737 6906
rect 11643 6899 11737 6902
rect 11643 6892 11692 6899
rect 11643 6886 11673 6892
rect 11692 6887 11697 6892
rect 11609 6870 11689 6886
rect 11701 6878 11737 6899
rect 11798 6894 11987 6918
rect 12032 6917 12079 6918
rect 12045 6912 12079 6917
rect 11813 6891 11987 6894
rect 11806 6888 11987 6891
rect 12015 6911 12079 6912
rect 11609 6868 11628 6870
rect 11643 6868 11677 6870
rect 11609 6852 11689 6868
rect 11609 6846 11628 6852
rect 11325 6820 11428 6830
rect 11279 6818 11428 6820
rect 11449 6818 11484 6830
rect 11118 6816 11280 6818
rect 11130 6796 11149 6816
rect 11164 6814 11194 6816
rect 11013 6788 11054 6796
rect 11136 6792 11149 6796
rect 11201 6800 11280 6816
rect 11312 6816 11484 6818
rect 11312 6800 11391 6816
rect 11398 6814 11428 6816
rect 10976 6778 11005 6788
rect 11019 6778 11048 6788
rect 11063 6778 11093 6792
rect 11136 6778 11179 6792
rect 11201 6788 11391 6800
rect 11456 6796 11462 6816
rect 11186 6778 11216 6788
rect 11217 6778 11375 6788
rect 11379 6778 11409 6788
rect 11413 6778 11443 6792
rect 11471 6778 11484 6816
rect 11556 6830 11585 6846
rect 11599 6830 11628 6846
rect 11643 6836 11673 6852
rect 11701 6830 11707 6878
rect 11710 6872 11729 6878
rect 11744 6872 11774 6880
rect 11710 6864 11774 6872
rect 11710 6848 11790 6864
rect 11806 6857 11868 6888
rect 11884 6857 11946 6888
rect 12015 6886 12064 6911
rect 12079 6886 12109 6902
rect 11978 6872 12008 6880
rect 12015 6878 12125 6886
rect 11978 6864 12023 6872
rect 11710 6846 11729 6848
rect 11744 6846 11790 6848
rect 11710 6830 11790 6846
rect 11817 6844 11852 6857
rect 11893 6854 11930 6857
rect 11893 6852 11935 6854
rect 11822 6841 11852 6844
rect 11831 6837 11838 6841
rect 11838 6836 11839 6837
rect 11797 6830 11807 6836
rect 11556 6822 11591 6830
rect 11556 6796 11557 6822
rect 11564 6796 11591 6822
rect 11499 6778 11529 6792
rect 11556 6788 11591 6796
rect 11593 6822 11634 6830
rect 11593 6796 11608 6822
rect 11615 6796 11634 6822
rect 11698 6818 11729 6830
rect 11744 6818 11847 6830
rect 11859 6820 11885 6846
rect 11900 6841 11930 6852
rect 11962 6848 12024 6864
rect 11962 6846 12008 6848
rect 11962 6830 12024 6846
rect 12036 6830 12042 6878
rect 12045 6870 12125 6878
rect 12045 6868 12064 6870
rect 12079 6868 12113 6870
rect 12045 6852 12125 6868
rect 12045 6830 12064 6852
rect 12079 6836 12109 6852
rect 12137 6846 12143 6920
rect 12146 6846 12165 6990
rect 12180 6846 12186 6990
rect 12195 6920 12208 6990
rect 12260 6986 12282 6990
rect 12253 6964 12282 6978
rect 12335 6964 12351 6978
rect 12389 6974 12395 6976
rect 12402 6974 12510 6990
rect 12517 6974 12523 6976
rect 12531 6974 12546 6990
rect 12612 6984 12631 6987
rect 12253 6962 12351 6964
rect 12378 6962 12546 6974
rect 12561 6964 12577 6978
rect 12612 6965 12634 6984
rect 12644 6978 12660 6979
rect 12643 6976 12660 6978
rect 12644 6971 12660 6976
rect 12634 6964 12640 6965
rect 12643 6964 12672 6971
rect 12561 6963 12672 6964
rect 12561 6962 12678 6963
rect 12237 6954 12288 6962
rect 12335 6954 12369 6962
rect 12237 6942 12262 6954
rect 12269 6942 12288 6954
rect 12342 6952 12369 6954
rect 12378 6952 12599 6962
rect 12634 6959 12640 6962
rect 12342 6948 12599 6952
rect 12237 6934 12288 6942
rect 12335 6934 12599 6948
rect 12643 6954 12678 6962
rect 12189 6886 12208 6920
rect 12253 6926 12282 6934
rect 12253 6920 12270 6926
rect 12253 6918 12287 6920
rect 12335 6918 12351 6934
rect 12352 6924 12560 6934
rect 12561 6924 12577 6934
rect 12625 6930 12640 6945
rect 12643 6942 12644 6954
rect 12651 6942 12678 6954
rect 12643 6934 12678 6942
rect 12643 6933 12672 6934
rect 12363 6920 12577 6924
rect 12378 6918 12577 6920
rect 12612 6920 12625 6930
rect 12643 6920 12660 6933
rect 12612 6918 12660 6920
rect 12254 6914 12287 6918
rect 12250 6912 12287 6914
rect 12250 6911 12317 6912
rect 12250 6906 12281 6911
rect 12287 6906 12317 6911
rect 12250 6902 12317 6906
rect 12223 6899 12317 6902
rect 12223 6892 12272 6899
rect 12223 6886 12253 6892
rect 12272 6887 12277 6892
rect 12189 6870 12269 6886
rect 12281 6878 12317 6899
rect 12378 6894 12567 6918
rect 12612 6917 12659 6918
rect 12625 6912 12659 6917
rect 12393 6891 12567 6894
rect 12386 6888 12567 6891
rect 12595 6911 12659 6912
rect 12189 6868 12208 6870
rect 12223 6868 12257 6870
rect 12189 6852 12269 6868
rect 12189 6846 12208 6852
rect 11905 6820 12008 6830
rect 11859 6818 12008 6820
rect 12029 6818 12064 6830
rect 11698 6816 11860 6818
rect 11710 6796 11729 6816
rect 11744 6814 11774 6816
rect 11593 6788 11634 6796
rect 11716 6792 11729 6796
rect 11781 6800 11860 6816
rect 11892 6816 12064 6818
rect 11892 6800 11971 6816
rect 11978 6814 12008 6816
rect 11556 6778 11585 6788
rect 11599 6778 11628 6788
rect 11643 6778 11673 6792
rect 11716 6778 11759 6792
rect 11781 6788 11971 6800
rect 12036 6796 12042 6816
rect 11766 6778 11796 6788
rect 11797 6778 11955 6788
rect 11959 6778 11989 6788
rect 11993 6778 12023 6792
rect 12051 6778 12064 6816
rect 12136 6830 12165 6846
rect 12179 6830 12208 6846
rect 12223 6836 12253 6852
rect 12281 6830 12287 6878
rect 12290 6872 12309 6878
rect 12324 6872 12354 6880
rect 12290 6864 12354 6872
rect 12290 6848 12370 6864
rect 12386 6857 12448 6888
rect 12464 6857 12526 6888
rect 12595 6886 12644 6911
rect 12659 6886 12689 6902
rect 12558 6872 12588 6880
rect 12595 6878 12705 6886
rect 12558 6864 12603 6872
rect 12290 6846 12309 6848
rect 12324 6846 12370 6848
rect 12290 6830 12370 6846
rect 12397 6844 12432 6857
rect 12473 6854 12510 6857
rect 12473 6852 12515 6854
rect 12402 6841 12432 6844
rect 12411 6837 12418 6841
rect 12418 6836 12419 6837
rect 12377 6830 12387 6836
rect 12136 6822 12171 6830
rect 12136 6796 12137 6822
rect 12144 6796 12171 6822
rect 12079 6778 12109 6792
rect 12136 6788 12171 6796
rect 12173 6822 12214 6830
rect 12173 6796 12188 6822
rect 12195 6796 12214 6822
rect 12278 6818 12309 6830
rect 12324 6818 12427 6830
rect 12439 6820 12465 6846
rect 12480 6841 12510 6852
rect 12542 6848 12604 6864
rect 12542 6846 12588 6848
rect 12542 6830 12604 6846
rect 12616 6830 12622 6878
rect 12625 6870 12705 6878
rect 12625 6868 12644 6870
rect 12659 6868 12693 6870
rect 12625 6852 12705 6868
rect 12625 6830 12644 6852
rect 12659 6836 12689 6852
rect 12717 6846 12723 6920
rect 12726 6846 12745 6990
rect 12760 6846 12766 6990
rect 12775 6920 12788 6990
rect 12840 6986 12862 6990
rect 12833 6964 12862 6978
rect 12915 6964 12931 6978
rect 12969 6974 12975 6976
rect 12982 6974 13090 6990
rect 13097 6974 13103 6976
rect 13111 6974 13126 6990
rect 13192 6984 13211 6987
rect 12833 6962 12931 6964
rect 12958 6962 13126 6974
rect 13141 6964 13157 6978
rect 13192 6965 13214 6984
rect 13224 6978 13240 6979
rect 13223 6976 13240 6978
rect 13224 6971 13240 6976
rect 13214 6964 13220 6965
rect 13223 6964 13252 6971
rect 13141 6963 13252 6964
rect 13141 6962 13258 6963
rect 12817 6954 12868 6962
rect 12915 6954 12949 6962
rect 12817 6942 12842 6954
rect 12849 6942 12868 6954
rect 12922 6952 12949 6954
rect 12958 6952 13179 6962
rect 13214 6959 13220 6962
rect 12922 6948 13179 6952
rect 12817 6934 12868 6942
rect 12915 6934 13179 6948
rect 13223 6954 13258 6962
rect 12769 6886 12788 6920
rect 12833 6926 12862 6934
rect 12833 6920 12850 6926
rect 12833 6918 12867 6920
rect 12915 6918 12931 6934
rect 12932 6924 13140 6934
rect 13141 6924 13157 6934
rect 13205 6930 13220 6945
rect 13223 6942 13224 6954
rect 13231 6942 13258 6954
rect 13223 6934 13258 6942
rect 13223 6933 13252 6934
rect 12943 6920 13157 6924
rect 12958 6918 13157 6920
rect 13192 6920 13205 6930
rect 13223 6920 13240 6933
rect 13192 6918 13240 6920
rect 12834 6914 12867 6918
rect 12830 6912 12867 6914
rect 12830 6911 12897 6912
rect 12830 6906 12861 6911
rect 12867 6906 12897 6911
rect 12830 6902 12897 6906
rect 12803 6899 12897 6902
rect 12803 6892 12852 6899
rect 12803 6886 12833 6892
rect 12852 6887 12857 6892
rect 12769 6870 12849 6886
rect 12861 6878 12897 6899
rect 12958 6894 13147 6918
rect 13192 6917 13239 6918
rect 13205 6912 13239 6917
rect 12973 6891 13147 6894
rect 12966 6888 13147 6891
rect 13175 6911 13239 6912
rect 12769 6868 12788 6870
rect 12803 6868 12837 6870
rect 12769 6852 12849 6868
rect 12769 6846 12788 6852
rect 12485 6820 12588 6830
rect 12439 6818 12588 6820
rect 12609 6818 12644 6830
rect 12278 6816 12440 6818
rect 12290 6796 12309 6816
rect 12324 6814 12354 6816
rect 12173 6788 12214 6796
rect 12296 6792 12309 6796
rect 12361 6800 12440 6816
rect 12472 6816 12644 6818
rect 12472 6800 12551 6816
rect 12558 6814 12588 6816
rect 12136 6778 12165 6788
rect 12179 6778 12208 6788
rect 12223 6778 12253 6792
rect 12296 6778 12339 6792
rect 12361 6788 12551 6800
rect 12616 6796 12622 6816
rect 12346 6778 12376 6788
rect 12377 6778 12535 6788
rect 12539 6778 12569 6788
rect 12573 6778 12603 6792
rect 12631 6778 12644 6816
rect 12716 6830 12745 6846
rect 12759 6830 12788 6846
rect 12803 6836 12833 6852
rect 12861 6830 12867 6878
rect 12870 6872 12889 6878
rect 12904 6872 12934 6880
rect 12870 6864 12934 6872
rect 12870 6848 12950 6864
rect 12966 6857 13028 6888
rect 13044 6857 13106 6888
rect 13175 6886 13224 6911
rect 13239 6886 13269 6902
rect 13138 6872 13168 6880
rect 13175 6878 13285 6886
rect 13138 6864 13183 6872
rect 12870 6846 12889 6848
rect 12904 6846 12950 6848
rect 12870 6830 12950 6846
rect 12977 6844 13012 6857
rect 13053 6854 13090 6857
rect 13053 6852 13095 6854
rect 12982 6841 13012 6844
rect 12991 6837 12998 6841
rect 12998 6836 12999 6837
rect 12957 6830 12967 6836
rect 12716 6822 12751 6830
rect 12716 6796 12717 6822
rect 12724 6796 12751 6822
rect 12659 6778 12689 6792
rect 12716 6788 12751 6796
rect 12753 6822 12794 6830
rect 12753 6796 12768 6822
rect 12775 6796 12794 6822
rect 12858 6818 12889 6830
rect 12904 6818 13007 6830
rect 13019 6820 13045 6846
rect 13060 6841 13090 6852
rect 13122 6848 13184 6864
rect 13122 6846 13168 6848
rect 13122 6830 13184 6846
rect 13196 6830 13202 6878
rect 13205 6870 13285 6878
rect 13205 6868 13224 6870
rect 13239 6868 13273 6870
rect 13205 6852 13285 6868
rect 13205 6830 13224 6852
rect 13239 6836 13269 6852
rect 13297 6846 13303 6920
rect 13306 6846 13325 6990
rect 13340 6846 13346 6990
rect 13355 6920 13368 6990
rect 13420 6986 13442 6990
rect 13413 6964 13442 6978
rect 13495 6964 13511 6978
rect 13549 6974 13555 6976
rect 13562 6974 13670 6990
rect 13677 6974 13683 6976
rect 13691 6974 13706 6990
rect 13772 6984 13791 6987
rect 13413 6962 13511 6964
rect 13538 6962 13706 6974
rect 13721 6964 13737 6978
rect 13772 6965 13794 6984
rect 13804 6978 13820 6979
rect 13803 6976 13820 6978
rect 13804 6971 13820 6976
rect 13794 6964 13800 6965
rect 13803 6964 13832 6971
rect 13721 6963 13832 6964
rect 13721 6962 13838 6963
rect 13397 6954 13448 6962
rect 13495 6954 13529 6962
rect 13397 6942 13422 6954
rect 13429 6942 13448 6954
rect 13502 6952 13529 6954
rect 13538 6952 13759 6962
rect 13794 6959 13800 6962
rect 13502 6948 13759 6952
rect 13397 6934 13448 6942
rect 13495 6934 13759 6948
rect 13803 6954 13838 6962
rect 13349 6886 13368 6920
rect 13413 6926 13442 6934
rect 13413 6920 13430 6926
rect 13413 6918 13447 6920
rect 13495 6918 13511 6934
rect 13512 6924 13720 6934
rect 13721 6924 13737 6934
rect 13785 6930 13800 6945
rect 13803 6942 13804 6954
rect 13811 6942 13838 6954
rect 13803 6934 13838 6942
rect 13803 6933 13832 6934
rect 13523 6920 13737 6924
rect 13538 6918 13737 6920
rect 13772 6920 13785 6930
rect 13803 6920 13820 6933
rect 13772 6918 13820 6920
rect 13414 6914 13447 6918
rect 13410 6912 13447 6914
rect 13410 6911 13477 6912
rect 13410 6906 13441 6911
rect 13447 6906 13477 6911
rect 13410 6902 13477 6906
rect 13383 6899 13477 6902
rect 13383 6892 13432 6899
rect 13383 6886 13413 6892
rect 13432 6887 13437 6892
rect 13349 6870 13429 6886
rect 13441 6878 13477 6899
rect 13538 6894 13727 6918
rect 13772 6917 13819 6918
rect 13785 6912 13819 6917
rect 13553 6891 13727 6894
rect 13546 6888 13727 6891
rect 13755 6911 13819 6912
rect 13349 6868 13368 6870
rect 13383 6868 13417 6870
rect 13349 6852 13429 6868
rect 13349 6846 13368 6852
rect 13065 6820 13168 6830
rect 13019 6818 13168 6820
rect 13189 6818 13224 6830
rect 12858 6816 13020 6818
rect 12870 6796 12889 6816
rect 12904 6814 12934 6816
rect 12753 6788 12794 6796
rect 12876 6792 12889 6796
rect 12941 6800 13020 6816
rect 13052 6816 13224 6818
rect 13052 6800 13131 6816
rect 13138 6814 13168 6816
rect 12716 6778 12745 6788
rect 12759 6778 12788 6788
rect 12803 6778 12833 6792
rect 12876 6778 12919 6792
rect 12941 6788 13131 6800
rect 13196 6796 13202 6816
rect 12926 6778 12956 6788
rect 12957 6778 13115 6788
rect 13119 6778 13149 6788
rect 13153 6778 13183 6792
rect 13211 6778 13224 6816
rect 13296 6830 13325 6846
rect 13339 6830 13368 6846
rect 13383 6836 13413 6852
rect 13441 6830 13447 6878
rect 13450 6872 13469 6878
rect 13484 6872 13514 6880
rect 13450 6864 13514 6872
rect 13450 6848 13530 6864
rect 13546 6857 13608 6888
rect 13624 6857 13686 6888
rect 13755 6886 13804 6911
rect 13819 6886 13849 6902
rect 13718 6872 13748 6880
rect 13755 6878 13865 6886
rect 13718 6864 13763 6872
rect 13450 6846 13469 6848
rect 13484 6846 13530 6848
rect 13450 6830 13530 6846
rect 13557 6844 13592 6857
rect 13633 6854 13670 6857
rect 13633 6852 13675 6854
rect 13562 6841 13592 6844
rect 13571 6837 13578 6841
rect 13578 6836 13579 6837
rect 13537 6830 13547 6836
rect 13296 6822 13331 6830
rect 13296 6796 13297 6822
rect 13304 6796 13331 6822
rect 13239 6778 13269 6792
rect 13296 6788 13331 6796
rect 13333 6822 13374 6830
rect 13333 6796 13348 6822
rect 13355 6796 13374 6822
rect 13438 6818 13469 6830
rect 13484 6818 13587 6830
rect 13599 6820 13625 6846
rect 13640 6841 13670 6852
rect 13702 6848 13764 6864
rect 13702 6846 13748 6848
rect 13702 6830 13764 6846
rect 13776 6830 13782 6878
rect 13785 6870 13865 6878
rect 13785 6868 13804 6870
rect 13819 6868 13853 6870
rect 13785 6852 13865 6868
rect 13785 6830 13804 6852
rect 13819 6836 13849 6852
rect 13877 6846 13883 6920
rect 13886 6846 13905 6990
rect 13920 6846 13926 6990
rect 13935 6920 13948 6990
rect 14000 6986 14022 6990
rect 13993 6964 14022 6978
rect 14075 6964 14091 6978
rect 14129 6974 14135 6976
rect 14142 6974 14250 6990
rect 14257 6974 14263 6976
rect 14271 6974 14286 6990
rect 14352 6984 14371 6987
rect 13993 6962 14091 6964
rect 14118 6962 14286 6974
rect 14301 6964 14317 6978
rect 14352 6965 14374 6984
rect 14384 6978 14400 6979
rect 14383 6976 14400 6978
rect 14384 6971 14400 6976
rect 14374 6964 14380 6965
rect 14383 6964 14412 6971
rect 14301 6963 14412 6964
rect 14301 6962 14418 6963
rect 13977 6954 14028 6962
rect 14075 6954 14109 6962
rect 13977 6942 14002 6954
rect 14009 6942 14028 6954
rect 14082 6952 14109 6954
rect 14118 6952 14339 6962
rect 14374 6959 14380 6962
rect 14082 6948 14339 6952
rect 13977 6934 14028 6942
rect 14075 6934 14339 6948
rect 14383 6954 14418 6962
rect 13929 6886 13948 6920
rect 13993 6926 14022 6934
rect 13993 6920 14010 6926
rect 13993 6918 14027 6920
rect 14075 6918 14091 6934
rect 14092 6924 14300 6934
rect 14301 6924 14317 6934
rect 14365 6930 14380 6945
rect 14383 6942 14384 6954
rect 14391 6942 14418 6954
rect 14383 6934 14418 6942
rect 14383 6933 14412 6934
rect 14103 6920 14317 6924
rect 14118 6918 14317 6920
rect 14352 6920 14365 6930
rect 14383 6920 14400 6933
rect 14352 6918 14400 6920
rect 13994 6914 14027 6918
rect 13990 6912 14027 6914
rect 13990 6911 14057 6912
rect 13990 6906 14021 6911
rect 14027 6906 14057 6911
rect 13990 6902 14057 6906
rect 13963 6899 14057 6902
rect 13963 6892 14012 6899
rect 13963 6886 13993 6892
rect 14012 6887 14017 6892
rect 13929 6870 14009 6886
rect 14021 6878 14057 6899
rect 14118 6894 14307 6918
rect 14352 6917 14399 6918
rect 14365 6912 14399 6917
rect 14133 6891 14307 6894
rect 14126 6888 14307 6891
rect 14335 6911 14399 6912
rect 13929 6868 13948 6870
rect 13963 6868 13997 6870
rect 13929 6852 14009 6868
rect 13929 6846 13948 6852
rect 13645 6820 13748 6830
rect 13599 6818 13748 6820
rect 13769 6818 13804 6830
rect 13438 6816 13600 6818
rect 13450 6796 13469 6816
rect 13484 6814 13514 6816
rect 13333 6788 13374 6796
rect 13456 6792 13469 6796
rect 13521 6800 13600 6816
rect 13632 6816 13804 6818
rect 13632 6800 13711 6816
rect 13718 6814 13748 6816
rect 13296 6778 13325 6788
rect 13339 6778 13368 6788
rect 13383 6778 13413 6792
rect 13456 6778 13499 6792
rect 13521 6788 13711 6800
rect 13776 6796 13782 6816
rect 13506 6778 13536 6788
rect 13537 6778 13695 6788
rect 13699 6778 13729 6788
rect 13733 6778 13763 6792
rect 13791 6778 13804 6816
rect 13876 6830 13905 6846
rect 13919 6830 13948 6846
rect 13963 6836 13993 6852
rect 14021 6830 14027 6878
rect 14030 6872 14049 6878
rect 14064 6872 14094 6880
rect 14030 6864 14094 6872
rect 14030 6848 14110 6864
rect 14126 6857 14188 6888
rect 14204 6857 14266 6888
rect 14335 6886 14384 6911
rect 14399 6886 14429 6902
rect 14298 6872 14328 6880
rect 14335 6878 14445 6886
rect 14298 6864 14343 6872
rect 14030 6846 14049 6848
rect 14064 6846 14110 6848
rect 14030 6830 14110 6846
rect 14137 6844 14172 6857
rect 14213 6854 14250 6857
rect 14213 6852 14255 6854
rect 14142 6841 14172 6844
rect 14151 6837 14158 6841
rect 14158 6836 14159 6837
rect 14117 6830 14127 6836
rect 13876 6822 13911 6830
rect 13876 6796 13877 6822
rect 13884 6796 13911 6822
rect 13819 6778 13849 6792
rect 13876 6788 13911 6796
rect 13913 6822 13954 6830
rect 13913 6796 13928 6822
rect 13935 6796 13954 6822
rect 14018 6818 14049 6830
rect 14064 6818 14167 6830
rect 14179 6820 14205 6846
rect 14220 6841 14250 6852
rect 14282 6848 14344 6864
rect 14282 6846 14328 6848
rect 14282 6830 14344 6846
rect 14356 6830 14362 6878
rect 14365 6870 14445 6878
rect 14365 6868 14384 6870
rect 14399 6868 14433 6870
rect 14365 6852 14445 6868
rect 14365 6830 14384 6852
rect 14399 6836 14429 6852
rect 14457 6846 14463 6920
rect 14466 6846 14485 6990
rect 14500 6846 14506 6990
rect 14515 6920 14528 6990
rect 14580 6986 14602 6990
rect 14573 6964 14602 6978
rect 14655 6964 14671 6978
rect 14709 6974 14715 6976
rect 14722 6974 14830 6990
rect 14837 6974 14843 6976
rect 14851 6974 14866 6990
rect 14932 6984 14951 6987
rect 14573 6962 14671 6964
rect 14698 6962 14866 6974
rect 14881 6964 14897 6978
rect 14932 6965 14954 6984
rect 14964 6978 14980 6979
rect 14963 6976 14980 6978
rect 14964 6971 14980 6976
rect 14954 6964 14960 6965
rect 14963 6964 14992 6971
rect 14881 6963 14992 6964
rect 14881 6962 14998 6963
rect 14557 6954 14608 6962
rect 14655 6954 14689 6962
rect 14557 6942 14582 6954
rect 14589 6942 14608 6954
rect 14662 6952 14689 6954
rect 14698 6952 14919 6962
rect 14954 6959 14960 6962
rect 14662 6948 14919 6952
rect 14557 6934 14608 6942
rect 14655 6934 14919 6948
rect 14963 6954 14998 6962
rect 14509 6886 14528 6920
rect 14573 6926 14602 6934
rect 14573 6920 14590 6926
rect 14573 6918 14607 6920
rect 14655 6918 14671 6934
rect 14672 6924 14880 6934
rect 14881 6924 14897 6934
rect 14945 6930 14960 6945
rect 14963 6942 14964 6954
rect 14971 6942 14998 6954
rect 14963 6934 14998 6942
rect 14963 6933 14992 6934
rect 14683 6920 14897 6924
rect 14698 6918 14897 6920
rect 14932 6920 14945 6930
rect 14963 6920 14980 6933
rect 14932 6918 14980 6920
rect 14574 6914 14607 6918
rect 14570 6912 14607 6914
rect 14570 6911 14637 6912
rect 14570 6906 14601 6911
rect 14607 6906 14637 6911
rect 14570 6902 14637 6906
rect 14543 6899 14637 6902
rect 14543 6892 14592 6899
rect 14543 6886 14573 6892
rect 14592 6887 14597 6892
rect 14509 6870 14589 6886
rect 14601 6878 14637 6899
rect 14698 6894 14887 6918
rect 14932 6917 14979 6918
rect 14945 6912 14979 6917
rect 14713 6891 14887 6894
rect 14706 6888 14887 6891
rect 14915 6911 14979 6912
rect 14509 6868 14528 6870
rect 14543 6868 14577 6870
rect 14509 6852 14589 6868
rect 14509 6846 14528 6852
rect 14225 6820 14328 6830
rect 14179 6818 14328 6820
rect 14349 6818 14384 6830
rect 14018 6816 14180 6818
rect 14030 6796 14049 6816
rect 14064 6814 14094 6816
rect 13913 6788 13954 6796
rect 14036 6792 14049 6796
rect 14101 6800 14180 6816
rect 14212 6816 14384 6818
rect 14212 6800 14291 6816
rect 14298 6814 14328 6816
rect 13876 6778 13905 6788
rect 13919 6778 13948 6788
rect 13963 6778 13993 6792
rect 14036 6778 14079 6792
rect 14101 6788 14291 6800
rect 14356 6796 14362 6816
rect 14086 6778 14116 6788
rect 14117 6778 14275 6788
rect 14279 6778 14309 6788
rect 14313 6778 14343 6792
rect 14371 6778 14384 6816
rect 14456 6830 14485 6846
rect 14499 6830 14528 6846
rect 14543 6836 14573 6852
rect 14601 6830 14607 6878
rect 14610 6872 14629 6878
rect 14644 6872 14674 6880
rect 14610 6864 14674 6872
rect 14610 6848 14690 6864
rect 14706 6857 14768 6888
rect 14784 6857 14846 6888
rect 14915 6886 14964 6911
rect 14979 6886 15009 6902
rect 14878 6872 14908 6880
rect 14915 6878 15025 6886
rect 14878 6864 14923 6872
rect 14610 6846 14629 6848
rect 14644 6846 14690 6848
rect 14610 6830 14690 6846
rect 14717 6844 14752 6857
rect 14793 6854 14830 6857
rect 14793 6852 14835 6854
rect 14722 6841 14752 6844
rect 14731 6837 14738 6841
rect 14738 6836 14739 6837
rect 14697 6830 14707 6836
rect 14456 6822 14491 6830
rect 14456 6796 14457 6822
rect 14464 6796 14491 6822
rect 14399 6778 14429 6792
rect 14456 6788 14491 6796
rect 14493 6822 14534 6830
rect 14493 6796 14508 6822
rect 14515 6796 14534 6822
rect 14598 6818 14629 6830
rect 14644 6818 14747 6830
rect 14759 6820 14785 6846
rect 14800 6841 14830 6852
rect 14862 6848 14924 6864
rect 14862 6846 14908 6848
rect 14862 6830 14924 6846
rect 14936 6830 14942 6878
rect 14945 6870 15025 6878
rect 14945 6868 14964 6870
rect 14979 6868 15013 6870
rect 14945 6852 15025 6868
rect 14945 6830 14964 6852
rect 14979 6836 15009 6852
rect 15037 6846 15043 6920
rect 15046 6846 15065 6990
rect 15080 6846 15086 6990
rect 15095 6920 15108 6990
rect 15160 6986 15182 6990
rect 15153 6964 15182 6978
rect 15235 6964 15251 6978
rect 15289 6974 15295 6976
rect 15302 6974 15410 6990
rect 15417 6974 15423 6976
rect 15431 6974 15446 6990
rect 15512 6984 15531 6987
rect 15153 6962 15251 6964
rect 15278 6962 15446 6974
rect 15461 6964 15477 6978
rect 15512 6965 15534 6984
rect 15544 6978 15560 6979
rect 15543 6976 15560 6978
rect 15544 6971 15560 6976
rect 15534 6964 15540 6965
rect 15543 6964 15572 6971
rect 15461 6963 15572 6964
rect 15461 6962 15578 6963
rect 15137 6954 15188 6962
rect 15235 6954 15269 6962
rect 15137 6942 15162 6954
rect 15169 6942 15188 6954
rect 15242 6952 15269 6954
rect 15278 6952 15499 6962
rect 15534 6959 15540 6962
rect 15242 6948 15499 6952
rect 15137 6934 15188 6942
rect 15235 6934 15499 6948
rect 15543 6954 15578 6962
rect 15089 6886 15108 6920
rect 15153 6926 15182 6934
rect 15153 6920 15170 6926
rect 15153 6918 15187 6920
rect 15235 6918 15251 6934
rect 15252 6924 15460 6934
rect 15461 6924 15477 6934
rect 15525 6930 15540 6945
rect 15543 6942 15544 6954
rect 15551 6942 15578 6954
rect 15543 6934 15578 6942
rect 15543 6933 15572 6934
rect 15263 6920 15477 6924
rect 15278 6918 15477 6920
rect 15512 6920 15525 6930
rect 15543 6920 15560 6933
rect 15512 6918 15560 6920
rect 15154 6914 15187 6918
rect 15150 6912 15187 6914
rect 15150 6911 15217 6912
rect 15150 6906 15181 6911
rect 15187 6906 15217 6911
rect 15150 6902 15217 6906
rect 15123 6899 15217 6902
rect 15123 6892 15172 6899
rect 15123 6886 15153 6892
rect 15172 6887 15177 6892
rect 15089 6870 15169 6886
rect 15181 6878 15217 6899
rect 15278 6894 15467 6918
rect 15512 6917 15559 6918
rect 15525 6912 15559 6917
rect 15293 6891 15467 6894
rect 15286 6888 15467 6891
rect 15495 6911 15559 6912
rect 15089 6868 15108 6870
rect 15123 6868 15157 6870
rect 15089 6852 15169 6868
rect 15089 6846 15108 6852
rect 14805 6820 14908 6830
rect 14759 6818 14908 6820
rect 14929 6818 14964 6830
rect 14598 6816 14760 6818
rect 14610 6796 14629 6816
rect 14644 6814 14674 6816
rect 14493 6788 14534 6796
rect 14616 6792 14629 6796
rect 14681 6800 14760 6816
rect 14792 6816 14964 6818
rect 14792 6800 14871 6816
rect 14878 6814 14908 6816
rect 14456 6778 14485 6788
rect 14499 6778 14528 6788
rect 14543 6778 14573 6792
rect 14616 6778 14659 6792
rect 14681 6788 14871 6800
rect 14936 6796 14942 6816
rect 14666 6778 14696 6788
rect 14697 6778 14855 6788
rect 14859 6778 14889 6788
rect 14893 6778 14923 6792
rect 14951 6778 14964 6816
rect 15036 6830 15065 6846
rect 15079 6830 15108 6846
rect 15123 6836 15153 6852
rect 15181 6830 15187 6878
rect 15190 6872 15209 6878
rect 15224 6872 15254 6880
rect 15190 6864 15254 6872
rect 15190 6848 15270 6864
rect 15286 6857 15348 6888
rect 15364 6857 15426 6888
rect 15495 6886 15544 6911
rect 15559 6886 15589 6902
rect 15458 6872 15488 6880
rect 15495 6878 15605 6886
rect 15458 6864 15503 6872
rect 15190 6846 15209 6848
rect 15224 6846 15270 6848
rect 15190 6830 15270 6846
rect 15297 6844 15332 6857
rect 15373 6854 15410 6857
rect 15373 6852 15415 6854
rect 15302 6841 15332 6844
rect 15311 6837 15318 6841
rect 15318 6836 15319 6837
rect 15277 6830 15287 6836
rect 15036 6822 15071 6830
rect 15036 6796 15037 6822
rect 15044 6796 15071 6822
rect 14979 6778 15009 6792
rect 15036 6788 15071 6796
rect 15073 6822 15114 6830
rect 15073 6796 15088 6822
rect 15095 6796 15114 6822
rect 15178 6818 15209 6830
rect 15224 6818 15327 6830
rect 15339 6820 15365 6846
rect 15380 6841 15410 6852
rect 15442 6848 15504 6864
rect 15442 6846 15488 6848
rect 15442 6830 15504 6846
rect 15516 6830 15522 6878
rect 15525 6870 15605 6878
rect 15525 6868 15544 6870
rect 15559 6868 15593 6870
rect 15525 6852 15605 6868
rect 15525 6830 15544 6852
rect 15559 6836 15589 6852
rect 15617 6846 15623 6920
rect 15626 6846 15645 6990
rect 15660 6846 15666 6990
rect 15675 6920 15688 6990
rect 15740 6986 15762 6990
rect 15733 6964 15762 6978
rect 15815 6964 15831 6978
rect 15869 6974 15875 6976
rect 15882 6974 15990 6990
rect 15997 6974 16003 6976
rect 16011 6974 16026 6990
rect 16092 6984 16111 6987
rect 15733 6962 15831 6964
rect 15858 6962 16026 6974
rect 16041 6964 16057 6978
rect 16092 6965 16114 6984
rect 16124 6978 16140 6979
rect 16123 6976 16140 6978
rect 16124 6971 16140 6976
rect 16114 6964 16120 6965
rect 16123 6964 16152 6971
rect 16041 6963 16152 6964
rect 16041 6962 16158 6963
rect 15717 6954 15768 6962
rect 15815 6954 15849 6962
rect 15717 6942 15742 6954
rect 15749 6942 15768 6954
rect 15822 6952 15849 6954
rect 15858 6952 16079 6962
rect 16114 6959 16120 6962
rect 15822 6948 16079 6952
rect 15717 6934 15768 6942
rect 15815 6934 16079 6948
rect 16123 6954 16158 6962
rect 15669 6886 15688 6920
rect 15733 6926 15762 6934
rect 15733 6920 15750 6926
rect 15733 6918 15767 6920
rect 15815 6918 15831 6934
rect 15832 6924 16040 6934
rect 16041 6924 16057 6934
rect 16105 6930 16120 6945
rect 16123 6942 16124 6954
rect 16131 6942 16158 6954
rect 16123 6934 16158 6942
rect 16123 6933 16152 6934
rect 15843 6920 16057 6924
rect 15858 6918 16057 6920
rect 16092 6920 16105 6930
rect 16123 6920 16140 6933
rect 16092 6918 16140 6920
rect 15734 6914 15767 6918
rect 15730 6912 15767 6914
rect 15730 6911 15797 6912
rect 15730 6906 15761 6911
rect 15767 6906 15797 6911
rect 15730 6902 15797 6906
rect 15703 6899 15797 6902
rect 15703 6892 15752 6899
rect 15703 6886 15733 6892
rect 15752 6887 15757 6892
rect 15669 6870 15749 6886
rect 15761 6878 15797 6899
rect 15858 6894 16047 6918
rect 16092 6917 16139 6918
rect 16105 6912 16139 6917
rect 15873 6891 16047 6894
rect 15866 6888 16047 6891
rect 16075 6911 16139 6912
rect 15669 6868 15688 6870
rect 15703 6868 15737 6870
rect 15669 6852 15749 6868
rect 15669 6846 15688 6852
rect 15385 6820 15488 6830
rect 15339 6818 15488 6820
rect 15509 6818 15544 6830
rect 15178 6816 15340 6818
rect 15190 6796 15209 6816
rect 15224 6814 15254 6816
rect 15073 6788 15114 6796
rect 15196 6792 15209 6796
rect 15261 6800 15340 6816
rect 15372 6816 15544 6818
rect 15372 6800 15451 6816
rect 15458 6814 15488 6816
rect 15036 6778 15065 6788
rect 15079 6778 15108 6788
rect 15123 6778 15153 6792
rect 15196 6778 15239 6792
rect 15261 6788 15451 6800
rect 15516 6796 15522 6816
rect 15246 6778 15276 6788
rect 15277 6778 15435 6788
rect 15439 6778 15469 6788
rect 15473 6778 15503 6792
rect 15531 6778 15544 6816
rect 15616 6830 15645 6846
rect 15659 6830 15688 6846
rect 15703 6836 15733 6852
rect 15761 6830 15767 6878
rect 15770 6872 15789 6878
rect 15804 6872 15834 6880
rect 15770 6864 15834 6872
rect 15770 6848 15850 6864
rect 15866 6857 15928 6888
rect 15944 6857 16006 6888
rect 16075 6886 16124 6911
rect 16139 6886 16169 6902
rect 16038 6872 16068 6880
rect 16075 6878 16185 6886
rect 16038 6864 16083 6872
rect 15770 6846 15789 6848
rect 15804 6846 15850 6848
rect 15770 6830 15850 6846
rect 15877 6844 15912 6857
rect 15953 6854 15990 6857
rect 15953 6852 15995 6854
rect 15882 6841 15912 6844
rect 15891 6837 15898 6841
rect 15898 6836 15899 6837
rect 15857 6830 15867 6836
rect 15616 6822 15651 6830
rect 15616 6796 15617 6822
rect 15624 6796 15651 6822
rect 15559 6778 15589 6792
rect 15616 6788 15651 6796
rect 15653 6822 15694 6830
rect 15653 6796 15668 6822
rect 15675 6796 15694 6822
rect 15758 6818 15789 6830
rect 15804 6818 15907 6830
rect 15919 6820 15945 6846
rect 15960 6841 15990 6852
rect 16022 6848 16084 6864
rect 16022 6846 16068 6848
rect 16022 6830 16084 6846
rect 16096 6830 16102 6878
rect 16105 6870 16185 6878
rect 16105 6868 16124 6870
rect 16139 6868 16173 6870
rect 16105 6852 16185 6868
rect 16105 6830 16124 6852
rect 16139 6836 16169 6852
rect 16197 6846 16203 6920
rect 16206 6846 16225 6990
rect 16240 6846 16246 6990
rect 16255 6920 16268 6990
rect 16320 6986 16342 6990
rect 16313 6964 16342 6978
rect 16395 6964 16411 6978
rect 16449 6974 16455 6976
rect 16462 6974 16570 6990
rect 16577 6974 16583 6976
rect 16591 6974 16606 6990
rect 16672 6984 16691 6987
rect 16313 6962 16411 6964
rect 16438 6962 16606 6974
rect 16621 6964 16637 6978
rect 16672 6965 16694 6984
rect 16704 6978 16720 6979
rect 16703 6976 16720 6978
rect 16704 6971 16720 6976
rect 16694 6964 16700 6965
rect 16703 6964 16732 6971
rect 16621 6963 16732 6964
rect 16621 6962 16738 6963
rect 16297 6954 16348 6962
rect 16395 6954 16429 6962
rect 16297 6942 16322 6954
rect 16329 6942 16348 6954
rect 16402 6952 16429 6954
rect 16438 6952 16659 6962
rect 16694 6959 16700 6962
rect 16402 6948 16659 6952
rect 16297 6934 16348 6942
rect 16395 6934 16659 6948
rect 16703 6954 16738 6962
rect 16249 6886 16268 6920
rect 16313 6926 16342 6934
rect 16313 6920 16330 6926
rect 16313 6918 16347 6920
rect 16395 6918 16411 6934
rect 16412 6924 16620 6934
rect 16621 6924 16637 6934
rect 16685 6930 16700 6945
rect 16703 6942 16704 6954
rect 16711 6942 16738 6954
rect 16703 6934 16738 6942
rect 16703 6933 16732 6934
rect 16423 6920 16637 6924
rect 16438 6918 16637 6920
rect 16672 6920 16685 6930
rect 16703 6920 16720 6933
rect 16672 6918 16720 6920
rect 16314 6914 16347 6918
rect 16310 6912 16347 6914
rect 16310 6911 16377 6912
rect 16310 6906 16341 6911
rect 16347 6906 16377 6911
rect 16310 6902 16377 6906
rect 16283 6899 16377 6902
rect 16283 6892 16332 6899
rect 16283 6886 16313 6892
rect 16332 6887 16337 6892
rect 16249 6870 16329 6886
rect 16341 6878 16377 6899
rect 16438 6894 16627 6918
rect 16672 6917 16719 6918
rect 16685 6912 16719 6917
rect 16453 6891 16627 6894
rect 16446 6888 16627 6891
rect 16655 6911 16719 6912
rect 16249 6868 16268 6870
rect 16283 6868 16317 6870
rect 16249 6852 16329 6868
rect 16249 6846 16268 6852
rect 15965 6820 16068 6830
rect 15919 6818 16068 6820
rect 16089 6818 16124 6830
rect 15758 6816 15920 6818
rect 15770 6796 15789 6816
rect 15804 6814 15834 6816
rect 15653 6788 15694 6796
rect 15776 6792 15789 6796
rect 15841 6800 15920 6816
rect 15952 6816 16124 6818
rect 15952 6800 16031 6816
rect 16038 6814 16068 6816
rect 15616 6778 15645 6788
rect 15659 6778 15688 6788
rect 15703 6778 15733 6792
rect 15776 6778 15819 6792
rect 15841 6788 16031 6800
rect 16096 6796 16102 6816
rect 15826 6778 15856 6788
rect 15857 6778 16015 6788
rect 16019 6778 16049 6788
rect 16053 6778 16083 6792
rect 16111 6778 16124 6816
rect 16196 6830 16225 6846
rect 16239 6830 16268 6846
rect 16283 6836 16313 6852
rect 16341 6830 16347 6878
rect 16350 6872 16369 6878
rect 16384 6872 16414 6880
rect 16350 6864 16414 6872
rect 16350 6848 16430 6864
rect 16446 6857 16508 6888
rect 16524 6857 16586 6888
rect 16655 6886 16704 6911
rect 16719 6886 16749 6902
rect 16618 6872 16648 6880
rect 16655 6878 16765 6886
rect 16618 6864 16663 6872
rect 16350 6846 16369 6848
rect 16384 6846 16430 6848
rect 16350 6830 16430 6846
rect 16457 6844 16492 6857
rect 16533 6854 16570 6857
rect 16533 6852 16575 6854
rect 16462 6841 16492 6844
rect 16471 6837 16478 6841
rect 16478 6836 16479 6837
rect 16437 6830 16447 6836
rect 16196 6822 16231 6830
rect 16196 6796 16197 6822
rect 16204 6796 16231 6822
rect 16139 6778 16169 6792
rect 16196 6788 16231 6796
rect 16233 6822 16274 6830
rect 16233 6796 16248 6822
rect 16255 6796 16274 6822
rect 16338 6818 16369 6830
rect 16384 6818 16487 6830
rect 16499 6820 16525 6846
rect 16540 6841 16570 6852
rect 16602 6848 16664 6864
rect 16602 6846 16648 6848
rect 16602 6830 16664 6846
rect 16676 6830 16682 6878
rect 16685 6870 16765 6878
rect 16685 6868 16704 6870
rect 16719 6868 16753 6870
rect 16685 6852 16765 6868
rect 16685 6830 16704 6852
rect 16719 6836 16749 6852
rect 16777 6846 16783 6920
rect 16786 6846 16805 6990
rect 16820 6846 16826 6990
rect 16835 6920 16848 6990
rect 16900 6986 16922 6990
rect 16893 6964 16922 6978
rect 16975 6964 16991 6978
rect 17029 6974 17035 6976
rect 17042 6974 17150 6990
rect 17157 6974 17163 6976
rect 17171 6974 17186 6990
rect 17252 6984 17271 6987
rect 16893 6962 16991 6964
rect 17018 6962 17186 6974
rect 17201 6964 17217 6978
rect 17252 6965 17274 6984
rect 17284 6978 17300 6979
rect 17283 6976 17300 6978
rect 17284 6971 17300 6976
rect 17274 6964 17280 6965
rect 17283 6964 17312 6971
rect 17201 6963 17312 6964
rect 17201 6962 17318 6963
rect 16877 6954 16928 6962
rect 16975 6954 17009 6962
rect 16877 6942 16902 6954
rect 16909 6942 16928 6954
rect 16982 6952 17009 6954
rect 17018 6952 17239 6962
rect 17274 6959 17280 6962
rect 16982 6948 17239 6952
rect 16877 6934 16928 6942
rect 16975 6934 17239 6948
rect 17283 6954 17318 6962
rect 16829 6886 16848 6920
rect 16893 6926 16922 6934
rect 16893 6920 16910 6926
rect 16893 6918 16927 6920
rect 16975 6918 16991 6934
rect 16992 6924 17200 6934
rect 17201 6924 17217 6934
rect 17265 6930 17280 6945
rect 17283 6942 17284 6954
rect 17291 6942 17318 6954
rect 17283 6934 17318 6942
rect 17283 6933 17312 6934
rect 17003 6920 17217 6924
rect 17018 6918 17217 6920
rect 17252 6920 17265 6930
rect 17283 6920 17300 6933
rect 17252 6918 17300 6920
rect 16894 6914 16927 6918
rect 16890 6912 16927 6914
rect 16890 6911 16957 6912
rect 16890 6906 16921 6911
rect 16927 6906 16957 6911
rect 16890 6902 16957 6906
rect 16863 6899 16957 6902
rect 16863 6892 16912 6899
rect 16863 6886 16893 6892
rect 16912 6887 16917 6892
rect 16829 6870 16909 6886
rect 16921 6878 16957 6899
rect 17018 6894 17207 6918
rect 17252 6917 17299 6918
rect 17265 6912 17299 6917
rect 17033 6891 17207 6894
rect 17026 6888 17207 6891
rect 17235 6911 17299 6912
rect 16829 6868 16848 6870
rect 16863 6868 16897 6870
rect 16829 6852 16909 6868
rect 16829 6846 16848 6852
rect 16545 6820 16648 6830
rect 16499 6818 16648 6820
rect 16669 6818 16704 6830
rect 16338 6816 16500 6818
rect 16350 6796 16369 6816
rect 16384 6814 16414 6816
rect 16233 6788 16274 6796
rect 16356 6792 16369 6796
rect 16421 6800 16500 6816
rect 16532 6816 16704 6818
rect 16532 6800 16611 6816
rect 16618 6814 16648 6816
rect 16196 6778 16225 6788
rect 16239 6778 16268 6788
rect 16283 6778 16313 6792
rect 16356 6778 16399 6792
rect 16421 6788 16611 6800
rect 16676 6796 16682 6816
rect 16406 6778 16436 6788
rect 16437 6778 16595 6788
rect 16599 6778 16629 6788
rect 16633 6778 16663 6792
rect 16691 6778 16704 6816
rect 16776 6830 16805 6846
rect 16819 6830 16848 6846
rect 16863 6836 16893 6852
rect 16921 6830 16927 6878
rect 16930 6872 16949 6878
rect 16964 6872 16994 6880
rect 16930 6864 16994 6872
rect 16930 6848 17010 6864
rect 17026 6857 17088 6888
rect 17104 6857 17166 6888
rect 17235 6886 17284 6911
rect 17299 6886 17329 6902
rect 17198 6872 17228 6880
rect 17235 6878 17345 6886
rect 17198 6864 17243 6872
rect 16930 6846 16949 6848
rect 16964 6846 17010 6848
rect 16930 6830 17010 6846
rect 17037 6844 17072 6857
rect 17113 6854 17150 6857
rect 17113 6852 17155 6854
rect 17042 6841 17072 6844
rect 17051 6837 17058 6841
rect 17058 6836 17059 6837
rect 17017 6830 17027 6836
rect 16776 6822 16811 6830
rect 16776 6796 16777 6822
rect 16784 6796 16811 6822
rect 16719 6778 16749 6792
rect 16776 6788 16811 6796
rect 16813 6822 16854 6830
rect 16813 6796 16828 6822
rect 16835 6796 16854 6822
rect 16918 6818 16949 6830
rect 16964 6818 17067 6830
rect 17079 6820 17105 6846
rect 17120 6841 17150 6852
rect 17182 6848 17244 6864
rect 17182 6846 17228 6848
rect 17182 6830 17244 6846
rect 17256 6830 17262 6878
rect 17265 6870 17345 6878
rect 17265 6868 17284 6870
rect 17299 6868 17333 6870
rect 17265 6852 17345 6868
rect 17265 6830 17284 6852
rect 17299 6836 17329 6852
rect 17357 6846 17363 6920
rect 17366 6846 17385 6990
rect 17400 6846 17406 6990
rect 17415 6920 17428 6990
rect 17480 6986 17502 6990
rect 17473 6964 17502 6978
rect 17555 6964 17571 6978
rect 17609 6974 17615 6976
rect 17622 6974 17730 6990
rect 17737 6974 17743 6976
rect 17751 6974 17766 6990
rect 17832 6984 17851 6987
rect 17473 6962 17571 6964
rect 17598 6962 17766 6974
rect 17781 6964 17797 6978
rect 17832 6965 17854 6984
rect 17864 6978 17880 6979
rect 17863 6976 17880 6978
rect 17864 6971 17880 6976
rect 17854 6964 17860 6965
rect 17863 6964 17892 6971
rect 17781 6963 17892 6964
rect 17781 6962 17898 6963
rect 17457 6954 17508 6962
rect 17555 6954 17589 6962
rect 17457 6942 17482 6954
rect 17489 6942 17508 6954
rect 17562 6952 17589 6954
rect 17598 6952 17819 6962
rect 17854 6959 17860 6962
rect 17562 6948 17819 6952
rect 17457 6934 17508 6942
rect 17555 6934 17819 6948
rect 17863 6954 17898 6962
rect 17409 6886 17428 6920
rect 17473 6926 17502 6934
rect 17473 6920 17490 6926
rect 17473 6918 17507 6920
rect 17555 6918 17571 6934
rect 17572 6924 17780 6934
rect 17781 6924 17797 6934
rect 17845 6930 17860 6945
rect 17863 6942 17864 6954
rect 17871 6942 17898 6954
rect 17863 6934 17898 6942
rect 17863 6933 17892 6934
rect 17583 6920 17797 6924
rect 17598 6918 17797 6920
rect 17832 6920 17845 6930
rect 17863 6920 17880 6933
rect 17832 6918 17880 6920
rect 17474 6914 17507 6918
rect 17470 6912 17507 6914
rect 17470 6911 17537 6912
rect 17470 6906 17501 6911
rect 17507 6906 17537 6911
rect 17470 6902 17537 6906
rect 17443 6899 17537 6902
rect 17443 6892 17492 6899
rect 17443 6886 17473 6892
rect 17492 6887 17497 6892
rect 17409 6870 17489 6886
rect 17501 6878 17537 6899
rect 17598 6894 17787 6918
rect 17832 6917 17879 6918
rect 17845 6912 17879 6917
rect 17613 6891 17787 6894
rect 17606 6888 17787 6891
rect 17815 6911 17879 6912
rect 17409 6868 17428 6870
rect 17443 6868 17477 6870
rect 17409 6852 17489 6868
rect 17409 6846 17428 6852
rect 17125 6820 17228 6830
rect 17079 6818 17228 6820
rect 17249 6818 17284 6830
rect 16918 6816 17080 6818
rect 16930 6796 16949 6816
rect 16964 6814 16994 6816
rect 16813 6788 16854 6796
rect 16936 6792 16949 6796
rect 17001 6800 17080 6816
rect 17112 6816 17284 6818
rect 17112 6800 17191 6816
rect 17198 6814 17228 6816
rect 16776 6778 16805 6788
rect 16819 6778 16848 6788
rect 16863 6778 16893 6792
rect 16936 6778 16979 6792
rect 17001 6788 17191 6800
rect 17256 6796 17262 6816
rect 16986 6778 17016 6788
rect 17017 6778 17175 6788
rect 17179 6778 17209 6788
rect 17213 6778 17243 6792
rect 17271 6778 17284 6816
rect 17356 6830 17385 6846
rect 17399 6830 17428 6846
rect 17443 6836 17473 6852
rect 17501 6830 17507 6878
rect 17510 6872 17529 6878
rect 17544 6872 17574 6880
rect 17510 6864 17574 6872
rect 17510 6848 17590 6864
rect 17606 6857 17668 6888
rect 17684 6857 17746 6888
rect 17815 6886 17864 6911
rect 17879 6886 17909 6902
rect 17778 6872 17808 6880
rect 17815 6878 17925 6886
rect 17778 6864 17823 6872
rect 17510 6846 17529 6848
rect 17544 6846 17590 6848
rect 17510 6830 17590 6846
rect 17617 6844 17652 6857
rect 17693 6854 17730 6857
rect 17693 6852 17735 6854
rect 17622 6841 17652 6844
rect 17631 6837 17638 6841
rect 17638 6836 17639 6837
rect 17597 6830 17607 6836
rect 17356 6822 17391 6830
rect 17356 6796 17357 6822
rect 17364 6796 17391 6822
rect 17299 6778 17329 6792
rect 17356 6788 17391 6796
rect 17393 6822 17434 6830
rect 17393 6796 17408 6822
rect 17415 6796 17434 6822
rect 17498 6818 17529 6830
rect 17544 6818 17647 6830
rect 17659 6820 17685 6846
rect 17700 6841 17730 6852
rect 17762 6848 17824 6864
rect 17762 6846 17808 6848
rect 17762 6830 17824 6846
rect 17836 6830 17842 6878
rect 17845 6870 17925 6878
rect 17845 6868 17864 6870
rect 17879 6868 17913 6870
rect 17845 6852 17925 6868
rect 17845 6830 17864 6852
rect 17879 6836 17909 6852
rect 17937 6846 17943 6920
rect 17946 6846 17965 6990
rect 17980 6846 17986 6990
rect 17995 6920 18008 6990
rect 18060 6986 18082 6990
rect 18053 6964 18082 6978
rect 18135 6964 18151 6978
rect 18189 6974 18195 6976
rect 18202 6974 18310 6990
rect 18317 6974 18323 6976
rect 18331 6974 18346 6990
rect 18412 6984 18431 6987
rect 18053 6962 18151 6964
rect 18178 6962 18346 6974
rect 18361 6964 18377 6978
rect 18412 6965 18434 6984
rect 18444 6978 18460 6979
rect 18443 6976 18460 6978
rect 18444 6971 18460 6976
rect 18434 6964 18440 6965
rect 18443 6964 18472 6971
rect 18361 6963 18472 6964
rect 18361 6962 18478 6963
rect 18037 6954 18088 6962
rect 18135 6954 18169 6962
rect 18037 6942 18062 6954
rect 18069 6942 18088 6954
rect 18142 6952 18169 6954
rect 18178 6952 18399 6962
rect 18434 6959 18440 6962
rect 18142 6948 18399 6952
rect 18037 6934 18088 6942
rect 18135 6934 18399 6948
rect 18443 6954 18478 6962
rect 17989 6886 18008 6920
rect 18053 6926 18082 6934
rect 18053 6920 18070 6926
rect 18053 6918 18087 6920
rect 18135 6918 18151 6934
rect 18152 6924 18360 6934
rect 18361 6924 18377 6934
rect 18425 6930 18440 6945
rect 18443 6942 18444 6954
rect 18451 6942 18478 6954
rect 18443 6934 18478 6942
rect 18443 6933 18472 6934
rect 18163 6920 18377 6924
rect 18178 6918 18377 6920
rect 18412 6920 18425 6930
rect 18443 6920 18460 6933
rect 18412 6918 18460 6920
rect 18054 6914 18087 6918
rect 18050 6912 18087 6914
rect 18050 6911 18117 6912
rect 18050 6906 18081 6911
rect 18087 6906 18117 6911
rect 18050 6902 18117 6906
rect 18023 6899 18117 6902
rect 18023 6892 18072 6899
rect 18023 6886 18053 6892
rect 18072 6887 18077 6892
rect 17989 6870 18069 6886
rect 18081 6878 18117 6899
rect 18178 6894 18367 6918
rect 18412 6917 18459 6918
rect 18425 6912 18459 6917
rect 18193 6891 18367 6894
rect 18186 6888 18367 6891
rect 18395 6911 18459 6912
rect 17989 6868 18008 6870
rect 18023 6868 18057 6870
rect 17989 6852 18069 6868
rect 17989 6846 18008 6852
rect 17705 6820 17808 6830
rect 17659 6818 17808 6820
rect 17829 6818 17864 6830
rect 17498 6816 17660 6818
rect 17510 6796 17529 6816
rect 17544 6814 17574 6816
rect 17393 6788 17434 6796
rect 17516 6792 17529 6796
rect 17581 6800 17660 6816
rect 17692 6816 17864 6818
rect 17692 6800 17771 6816
rect 17778 6814 17808 6816
rect 17356 6778 17385 6788
rect 17399 6778 17428 6788
rect 17443 6778 17473 6792
rect 17516 6778 17559 6792
rect 17581 6788 17771 6800
rect 17836 6796 17842 6816
rect 17566 6778 17596 6788
rect 17597 6778 17755 6788
rect 17759 6778 17789 6788
rect 17793 6778 17823 6792
rect 17851 6778 17864 6816
rect 17936 6830 17965 6846
rect 17979 6830 18008 6846
rect 18023 6836 18053 6852
rect 18081 6830 18087 6878
rect 18090 6872 18109 6878
rect 18124 6872 18154 6880
rect 18090 6864 18154 6872
rect 18090 6848 18170 6864
rect 18186 6857 18248 6888
rect 18264 6857 18326 6888
rect 18395 6886 18444 6911
rect 18459 6886 18489 6902
rect 18358 6872 18388 6880
rect 18395 6878 18505 6886
rect 18358 6864 18403 6872
rect 18090 6846 18109 6848
rect 18124 6846 18170 6848
rect 18090 6830 18170 6846
rect 18197 6844 18232 6857
rect 18273 6854 18310 6857
rect 18273 6852 18315 6854
rect 18202 6841 18232 6844
rect 18211 6837 18218 6841
rect 18218 6836 18219 6837
rect 18177 6830 18187 6836
rect 17936 6822 17971 6830
rect 17936 6796 17937 6822
rect 17944 6796 17971 6822
rect 17879 6778 17909 6792
rect 17936 6788 17971 6796
rect 17973 6822 18014 6830
rect 17973 6796 17988 6822
rect 17995 6796 18014 6822
rect 18078 6818 18109 6830
rect 18124 6818 18227 6830
rect 18239 6820 18265 6846
rect 18280 6841 18310 6852
rect 18342 6848 18404 6864
rect 18342 6846 18388 6848
rect 18342 6830 18404 6846
rect 18416 6830 18422 6878
rect 18425 6870 18505 6878
rect 18425 6868 18444 6870
rect 18459 6868 18493 6870
rect 18425 6852 18505 6868
rect 18425 6830 18444 6852
rect 18459 6836 18489 6852
rect 18517 6846 18523 6920
rect 18532 6846 18545 6990
rect 18285 6820 18388 6830
rect 18239 6818 18388 6820
rect 18409 6818 18444 6830
rect 18078 6816 18240 6818
rect 18090 6796 18109 6816
rect 18124 6814 18154 6816
rect 17973 6788 18014 6796
rect 18096 6792 18109 6796
rect 18161 6800 18240 6816
rect 18272 6816 18444 6818
rect 18272 6800 18351 6816
rect 18358 6814 18388 6816
rect 17936 6778 17965 6788
rect 17979 6778 18008 6788
rect 18023 6778 18053 6792
rect 18096 6778 18139 6792
rect 18161 6788 18351 6800
rect 18416 6796 18422 6816
rect 18146 6778 18176 6788
rect 18177 6778 18335 6788
rect 18339 6778 18369 6788
rect 18373 6778 18403 6792
rect 18431 6778 18444 6816
rect 18516 6830 18545 6846
rect 18516 6822 18551 6830
rect 18516 6796 18517 6822
rect 18524 6796 18551 6822
rect 18459 6778 18489 6792
rect 18516 6788 18551 6796
rect 18516 6778 18545 6788
rect -1 6772 18545 6778
rect 0 6764 18545 6772
rect 15 6734 28 6764
rect 43 6750 73 6764
rect 116 6750 159 6764
rect 166 6750 386 6764
rect 393 6750 423 6764
rect 83 6736 98 6748
rect 117 6736 130 6750
rect 198 6746 351 6750
rect 80 6734 102 6736
rect 180 6734 372 6746
rect 451 6734 464 6764
rect 479 6750 509 6764
rect 546 6734 565 6764
rect 580 6734 586 6764
rect 595 6734 608 6764
rect 623 6750 653 6764
rect 696 6750 739 6764
rect 746 6750 966 6764
rect 973 6750 1003 6764
rect 663 6736 678 6748
rect 697 6736 710 6750
rect 778 6746 931 6750
rect 660 6734 682 6736
rect 760 6734 952 6746
rect 1031 6734 1044 6764
rect 1059 6750 1089 6764
rect 1126 6734 1145 6764
rect 1160 6734 1166 6764
rect 1175 6734 1188 6764
rect 1203 6750 1233 6764
rect 1276 6750 1319 6764
rect 1326 6750 1546 6764
rect 1553 6750 1583 6764
rect 1243 6736 1258 6748
rect 1277 6736 1290 6750
rect 1358 6746 1511 6750
rect 1240 6734 1262 6736
rect 1340 6734 1532 6746
rect 1611 6734 1624 6764
rect 1639 6750 1669 6764
rect 1706 6734 1725 6764
rect 1740 6734 1746 6764
rect 1755 6734 1768 6764
rect 1783 6750 1813 6764
rect 1856 6750 1899 6764
rect 1906 6750 2126 6764
rect 2133 6750 2163 6764
rect 1823 6736 1838 6748
rect 1857 6736 1870 6750
rect 1938 6746 2091 6750
rect 1820 6734 1842 6736
rect 1920 6734 2112 6746
rect 2191 6734 2204 6764
rect 2219 6750 2249 6764
rect 2286 6734 2305 6764
rect 2320 6734 2326 6764
rect 2335 6734 2348 6764
rect 2363 6750 2393 6764
rect 2436 6750 2479 6764
rect 2486 6750 2706 6764
rect 2713 6750 2743 6764
rect 2403 6736 2418 6748
rect 2437 6736 2450 6750
rect 2518 6746 2671 6750
rect 2400 6734 2422 6736
rect 2500 6734 2692 6746
rect 2771 6734 2784 6764
rect 2799 6750 2829 6764
rect 2866 6734 2885 6764
rect 2900 6734 2906 6764
rect 2915 6734 2928 6764
rect 2943 6750 2973 6764
rect 3016 6750 3059 6764
rect 3066 6750 3286 6764
rect 3293 6750 3323 6764
rect 2983 6736 2998 6748
rect 3017 6736 3030 6750
rect 3098 6746 3251 6750
rect 2980 6734 3002 6736
rect 3080 6734 3272 6746
rect 3351 6734 3364 6764
rect 3379 6750 3409 6764
rect 3446 6734 3465 6764
rect 3480 6734 3486 6764
rect 3495 6734 3508 6764
rect 3523 6750 3553 6764
rect 3596 6750 3639 6764
rect 3646 6750 3866 6764
rect 3873 6750 3903 6764
rect 3563 6736 3578 6748
rect 3597 6736 3610 6750
rect 3678 6746 3831 6750
rect 3560 6734 3582 6736
rect 3660 6734 3852 6746
rect 3931 6734 3944 6764
rect 3959 6750 3989 6764
rect 4026 6734 4045 6764
rect 4060 6734 4066 6764
rect 4075 6734 4088 6764
rect 4103 6750 4133 6764
rect 4176 6750 4219 6764
rect 4226 6750 4446 6764
rect 4453 6750 4483 6764
rect 4143 6736 4158 6748
rect 4177 6736 4190 6750
rect 4258 6746 4411 6750
rect 4140 6734 4162 6736
rect 4240 6734 4432 6746
rect 4511 6734 4524 6764
rect 4539 6750 4569 6764
rect 4606 6734 4625 6764
rect 4640 6734 4646 6764
rect 4655 6734 4668 6764
rect 4683 6750 4713 6764
rect 4756 6750 4799 6764
rect 4806 6750 5026 6764
rect 5033 6750 5063 6764
rect 4723 6736 4738 6748
rect 4757 6736 4770 6750
rect 4838 6746 4991 6750
rect 4720 6734 4742 6736
rect 4820 6734 5012 6746
rect 5091 6734 5104 6764
rect 5119 6750 5149 6764
rect 5186 6734 5205 6764
rect 5220 6734 5226 6764
rect 5235 6734 5248 6764
rect 5263 6750 5293 6764
rect 5336 6750 5379 6764
rect 5386 6750 5606 6764
rect 5613 6750 5643 6764
rect 5303 6736 5318 6748
rect 5337 6736 5350 6750
rect 5418 6746 5571 6750
rect 5300 6734 5322 6736
rect 5400 6734 5592 6746
rect 5671 6734 5684 6764
rect 5699 6750 5729 6764
rect 5766 6734 5785 6764
rect 5800 6734 5806 6764
rect 5815 6734 5828 6764
rect 5843 6750 5873 6764
rect 5916 6750 5959 6764
rect 5966 6750 6186 6764
rect 6193 6750 6223 6764
rect 5883 6736 5898 6748
rect 5917 6736 5930 6750
rect 5998 6746 6151 6750
rect 5880 6734 5902 6736
rect 5980 6734 6172 6746
rect 6251 6734 6264 6764
rect 6279 6750 6309 6764
rect 6346 6734 6365 6764
rect 6380 6734 6386 6764
rect 6395 6734 6408 6764
rect 6423 6750 6453 6764
rect 6496 6750 6539 6764
rect 6546 6750 6766 6764
rect 6773 6750 6803 6764
rect 6463 6736 6478 6748
rect 6497 6736 6510 6750
rect 6578 6746 6731 6750
rect 6460 6734 6482 6736
rect 6560 6734 6752 6746
rect 6831 6734 6844 6764
rect 6859 6750 6889 6764
rect 6926 6734 6945 6764
rect 6960 6734 6966 6764
rect 6975 6734 6988 6764
rect 7003 6750 7033 6764
rect 7076 6750 7119 6764
rect 7126 6750 7346 6764
rect 7353 6750 7383 6764
rect 7043 6736 7058 6748
rect 7077 6736 7090 6750
rect 7158 6746 7311 6750
rect 7040 6734 7062 6736
rect 7140 6734 7332 6746
rect 7411 6734 7424 6764
rect 7439 6750 7469 6764
rect 7506 6734 7525 6764
rect 7540 6734 7546 6764
rect 7555 6734 7568 6764
rect 7583 6750 7613 6764
rect 7656 6750 7699 6764
rect 7706 6750 7926 6764
rect 7933 6750 7963 6764
rect 7623 6736 7638 6748
rect 7657 6736 7670 6750
rect 7738 6746 7891 6750
rect 7620 6734 7642 6736
rect 7720 6734 7912 6746
rect 7991 6734 8004 6764
rect 8019 6750 8049 6764
rect 8086 6734 8105 6764
rect 8120 6734 8126 6764
rect 8135 6734 8148 6764
rect 8163 6750 8193 6764
rect 8236 6750 8279 6764
rect 8286 6750 8506 6764
rect 8513 6750 8543 6764
rect 8203 6736 8218 6748
rect 8237 6736 8250 6750
rect 8318 6746 8471 6750
rect 8200 6734 8222 6736
rect 8300 6734 8492 6746
rect 8571 6734 8584 6764
rect 8599 6750 8629 6764
rect 8666 6734 8685 6764
rect 8700 6734 8706 6764
rect 8715 6734 8728 6764
rect 8743 6750 8773 6764
rect 8816 6750 8859 6764
rect 8866 6750 9086 6764
rect 9093 6750 9123 6764
rect 8783 6736 8798 6748
rect 8817 6736 8830 6750
rect 8898 6746 9051 6750
rect 8780 6734 8802 6736
rect 8880 6734 9072 6746
rect 9151 6734 9164 6764
rect 9179 6750 9209 6764
rect 9246 6734 9265 6764
rect 9280 6734 9286 6764
rect 9295 6734 9308 6764
rect 9323 6750 9353 6764
rect 9396 6750 9439 6764
rect 9446 6750 9666 6764
rect 9673 6750 9703 6764
rect 9363 6736 9378 6748
rect 9397 6736 9410 6750
rect 9478 6746 9631 6750
rect 9360 6734 9382 6736
rect 9460 6734 9652 6746
rect 9731 6734 9744 6764
rect 9759 6750 9789 6764
rect 9826 6734 9845 6764
rect 9860 6734 9866 6764
rect 9875 6734 9888 6764
rect 9903 6750 9933 6764
rect 9976 6750 10019 6764
rect 10026 6750 10246 6764
rect 10253 6750 10283 6764
rect 9943 6736 9958 6748
rect 9977 6736 9990 6750
rect 10058 6746 10211 6750
rect 9940 6734 9962 6736
rect 10040 6734 10232 6746
rect 10311 6734 10324 6764
rect 10339 6750 10369 6764
rect 10406 6734 10425 6764
rect 10440 6734 10446 6764
rect 10455 6734 10468 6764
rect 10483 6750 10513 6764
rect 10556 6750 10599 6764
rect 10606 6750 10826 6764
rect 10833 6750 10863 6764
rect 10523 6736 10538 6748
rect 10557 6736 10570 6750
rect 10638 6746 10791 6750
rect 10520 6734 10542 6736
rect 10620 6734 10812 6746
rect 10891 6734 10904 6764
rect 10919 6750 10949 6764
rect 10986 6734 11005 6764
rect 11020 6734 11026 6764
rect 11035 6734 11048 6764
rect 11063 6750 11093 6764
rect 11136 6750 11179 6764
rect 11186 6750 11406 6764
rect 11413 6750 11443 6764
rect 11103 6736 11118 6748
rect 11137 6736 11150 6750
rect 11218 6746 11371 6750
rect 11100 6734 11122 6736
rect 11200 6734 11392 6746
rect 11471 6734 11484 6764
rect 11499 6750 11529 6764
rect 11566 6734 11585 6764
rect 11600 6734 11606 6764
rect 11615 6734 11628 6764
rect 11643 6750 11673 6764
rect 11716 6750 11759 6764
rect 11766 6750 11986 6764
rect 11993 6750 12023 6764
rect 11683 6736 11698 6748
rect 11717 6736 11730 6750
rect 11798 6746 11951 6750
rect 11680 6734 11702 6736
rect 11780 6734 11972 6746
rect 12051 6734 12064 6764
rect 12079 6750 12109 6764
rect 12146 6734 12165 6764
rect 12180 6734 12186 6764
rect 12195 6734 12208 6764
rect 12223 6750 12253 6764
rect 12296 6750 12339 6764
rect 12346 6750 12566 6764
rect 12573 6750 12603 6764
rect 12263 6736 12278 6748
rect 12297 6736 12310 6750
rect 12378 6746 12531 6750
rect 12260 6734 12282 6736
rect 12360 6734 12552 6746
rect 12631 6734 12644 6764
rect 12659 6750 12689 6764
rect 12726 6734 12745 6764
rect 12760 6734 12766 6764
rect 12775 6734 12788 6764
rect 12803 6750 12833 6764
rect 12876 6750 12919 6764
rect 12926 6750 13146 6764
rect 13153 6750 13183 6764
rect 12843 6736 12858 6748
rect 12877 6736 12890 6750
rect 12958 6746 13111 6750
rect 12840 6734 12862 6736
rect 12940 6734 13132 6746
rect 13211 6734 13224 6764
rect 13239 6750 13269 6764
rect 13306 6734 13325 6764
rect 13340 6734 13346 6764
rect 13355 6734 13368 6764
rect 13383 6750 13413 6764
rect 13456 6750 13499 6764
rect 13506 6750 13726 6764
rect 13733 6750 13763 6764
rect 13423 6736 13438 6748
rect 13457 6736 13470 6750
rect 13538 6746 13691 6750
rect 13420 6734 13442 6736
rect 13520 6734 13712 6746
rect 13791 6734 13804 6764
rect 13819 6750 13849 6764
rect 13886 6734 13905 6764
rect 13920 6734 13926 6764
rect 13935 6734 13948 6764
rect 13963 6750 13993 6764
rect 14036 6750 14079 6764
rect 14086 6750 14306 6764
rect 14313 6750 14343 6764
rect 14003 6736 14018 6748
rect 14037 6736 14050 6750
rect 14118 6746 14271 6750
rect 14000 6734 14022 6736
rect 14100 6734 14292 6746
rect 14371 6734 14384 6764
rect 14399 6750 14429 6764
rect 14466 6734 14485 6764
rect 14500 6734 14506 6764
rect 14515 6734 14528 6764
rect 14543 6750 14573 6764
rect 14616 6750 14659 6764
rect 14666 6750 14886 6764
rect 14893 6750 14923 6764
rect 14583 6736 14598 6748
rect 14617 6736 14630 6750
rect 14698 6746 14851 6750
rect 14580 6734 14602 6736
rect 14680 6734 14872 6746
rect 14951 6734 14964 6764
rect 14979 6750 15009 6764
rect 15046 6734 15065 6764
rect 15080 6734 15086 6764
rect 15095 6734 15108 6764
rect 15123 6750 15153 6764
rect 15196 6750 15239 6764
rect 15246 6750 15466 6764
rect 15473 6750 15503 6764
rect 15163 6736 15178 6748
rect 15197 6736 15210 6750
rect 15278 6746 15431 6750
rect 15160 6734 15182 6736
rect 15260 6734 15452 6746
rect 15531 6734 15544 6764
rect 15559 6750 15589 6764
rect 15626 6734 15645 6764
rect 15660 6734 15666 6764
rect 15675 6734 15688 6764
rect 15703 6750 15733 6764
rect 15776 6750 15819 6764
rect 15826 6750 16046 6764
rect 16053 6750 16083 6764
rect 15743 6736 15758 6748
rect 15777 6736 15790 6750
rect 15858 6746 16011 6750
rect 15740 6734 15762 6736
rect 15840 6734 16032 6746
rect 16111 6734 16124 6764
rect 16139 6750 16169 6764
rect 16206 6734 16225 6764
rect 16240 6734 16246 6764
rect 16255 6734 16268 6764
rect 16283 6750 16313 6764
rect 16356 6750 16399 6764
rect 16406 6750 16626 6764
rect 16633 6750 16663 6764
rect 16323 6736 16338 6748
rect 16357 6736 16370 6750
rect 16438 6746 16591 6750
rect 16320 6734 16342 6736
rect 16420 6734 16612 6746
rect 16691 6734 16704 6764
rect 16719 6750 16749 6764
rect 16786 6734 16805 6764
rect 16820 6734 16826 6764
rect 16835 6734 16848 6764
rect 16863 6750 16893 6764
rect 16936 6750 16979 6764
rect 16986 6750 17206 6764
rect 17213 6750 17243 6764
rect 16903 6736 16918 6748
rect 16937 6736 16950 6750
rect 17018 6746 17171 6750
rect 16900 6734 16922 6736
rect 17000 6734 17192 6746
rect 17271 6734 17284 6764
rect 17299 6750 17329 6764
rect 17366 6734 17385 6764
rect 17400 6734 17406 6764
rect 17415 6734 17428 6764
rect 17443 6750 17473 6764
rect 17516 6750 17559 6764
rect 17566 6750 17786 6764
rect 17793 6750 17823 6764
rect 17483 6736 17498 6748
rect 17517 6736 17530 6750
rect 17598 6746 17751 6750
rect 17480 6734 17502 6736
rect 17580 6734 17772 6746
rect 17851 6734 17864 6764
rect 17879 6750 17909 6764
rect 17946 6734 17965 6764
rect 17980 6734 17986 6764
rect 17995 6734 18008 6764
rect 18023 6750 18053 6764
rect 18096 6750 18139 6764
rect 18146 6750 18366 6764
rect 18373 6750 18403 6764
rect 18063 6736 18078 6748
rect 18097 6736 18110 6750
rect 18178 6746 18331 6750
rect 18060 6734 18082 6736
rect 18160 6734 18352 6746
rect 18431 6734 18444 6764
rect 18459 6750 18489 6764
rect 18532 6734 18545 6764
rect 0 6720 18545 6734
rect 15 6650 28 6720
rect 80 6716 102 6720
rect 73 6694 102 6708
rect 155 6694 171 6708
rect 209 6704 215 6706
rect 222 6704 330 6720
rect 337 6704 343 6706
rect 351 6704 366 6720
rect 432 6714 451 6717
rect 73 6692 171 6694
rect 198 6692 366 6704
rect 381 6694 397 6708
rect 432 6695 454 6714
rect 464 6708 480 6709
rect 463 6706 480 6708
rect 464 6701 480 6706
rect 454 6694 460 6695
rect 463 6694 492 6701
rect 381 6693 492 6694
rect 381 6692 498 6693
rect 57 6684 108 6692
rect 155 6684 189 6692
rect 57 6672 82 6684
rect 89 6672 108 6684
rect 162 6682 189 6684
rect 198 6682 419 6692
rect 454 6689 460 6692
rect 162 6678 419 6682
rect 57 6664 108 6672
rect 155 6664 419 6678
rect 463 6684 498 6692
rect 9 6616 28 6650
rect 73 6656 102 6664
rect 73 6650 90 6656
rect 73 6648 107 6650
rect 155 6648 171 6664
rect 172 6654 380 6664
rect 381 6654 397 6664
rect 445 6660 460 6675
rect 463 6672 464 6684
rect 471 6672 498 6684
rect 463 6664 498 6672
rect 463 6663 492 6664
rect 183 6650 397 6654
rect 198 6648 397 6650
rect 432 6650 445 6660
rect 463 6650 480 6663
rect 432 6648 480 6650
rect 74 6644 107 6648
rect 70 6642 107 6644
rect 70 6641 137 6642
rect 70 6636 101 6641
rect 107 6636 137 6641
rect 70 6632 137 6636
rect 43 6629 137 6632
rect 43 6622 92 6629
rect 43 6616 73 6622
rect 92 6617 97 6622
rect 9 6600 89 6616
rect 101 6608 137 6629
rect 198 6624 387 6648
rect 432 6647 479 6648
rect 445 6642 479 6647
rect 213 6621 387 6624
rect 206 6618 387 6621
rect 415 6641 479 6642
rect 9 6598 28 6600
rect 43 6598 77 6600
rect 9 6582 89 6598
rect 9 6576 28 6582
rect -1 6560 28 6576
rect 43 6566 73 6582
rect 101 6560 107 6608
rect 110 6602 129 6608
rect 144 6602 174 6610
rect 110 6594 174 6602
rect 110 6578 190 6594
rect 206 6587 268 6618
rect 284 6587 346 6618
rect 415 6616 464 6641
rect 479 6616 509 6632
rect 378 6602 408 6610
rect 415 6608 525 6616
rect 378 6594 423 6602
rect 110 6576 129 6578
rect 144 6576 190 6578
rect 110 6560 190 6576
rect 217 6574 252 6587
rect 293 6584 330 6587
rect 293 6582 335 6584
rect 222 6571 252 6574
rect 231 6567 238 6571
rect 238 6566 239 6567
rect 197 6560 207 6566
rect -7 6552 34 6560
rect -7 6526 8 6552
rect 15 6526 34 6552
rect 98 6548 129 6560
rect 144 6548 247 6560
rect 259 6550 285 6576
rect 300 6571 330 6582
rect 362 6578 424 6594
rect 362 6576 408 6578
rect 362 6560 424 6576
rect 436 6560 442 6608
rect 445 6600 525 6608
rect 445 6598 464 6600
rect 479 6598 513 6600
rect 445 6582 525 6598
rect 445 6560 464 6582
rect 479 6566 509 6582
rect 537 6576 543 6650
rect 546 6576 565 6720
rect 580 6576 586 6720
rect 595 6650 608 6720
rect 660 6716 682 6720
rect 653 6694 682 6708
rect 735 6694 751 6708
rect 789 6704 795 6706
rect 802 6704 910 6720
rect 917 6704 923 6706
rect 931 6704 946 6720
rect 1012 6714 1031 6717
rect 653 6692 751 6694
rect 778 6692 946 6704
rect 961 6694 977 6708
rect 1012 6695 1034 6714
rect 1044 6708 1060 6709
rect 1043 6706 1060 6708
rect 1044 6701 1060 6706
rect 1034 6694 1040 6695
rect 1043 6694 1072 6701
rect 961 6693 1072 6694
rect 961 6692 1078 6693
rect 637 6684 688 6692
rect 735 6684 769 6692
rect 637 6672 662 6684
rect 669 6672 688 6684
rect 742 6682 769 6684
rect 778 6682 999 6692
rect 1034 6689 1040 6692
rect 742 6678 999 6682
rect 637 6664 688 6672
rect 735 6664 999 6678
rect 1043 6684 1078 6692
rect 589 6616 608 6650
rect 653 6656 682 6664
rect 653 6650 670 6656
rect 653 6648 687 6650
rect 735 6648 751 6664
rect 752 6654 960 6664
rect 961 6654 977 6664
rect 1025 6660 1040 6675
rect 1043 6672 1044 6684
rect 1051 6672 1078 6684
rect 1043 6664 1078 6672
rect 1043 6663 1072 6664
rect 763 6650 977 6654
rect 778 6648 977 6650
rect 1012 6650 1025 6660
rect 1043 6650 1060 6663
rect 1012 6648 1060 6650
rect 654 6644 687 6648
rect 650 6642 687 6644
rect 650 6641 717 6642
rect 650 6636 681 6641
rect 687 6636 717 6641
rect 650 6632 717 6636
rect 623 6629 717 6632
rect 623 6622 672 6629
rect 623 6616 653 6622
rect 672 6617 677 6622
rect 589 6600 669 6616
rect 681 6608 717 6629
rect 778 6624 967 6648
rect 1012 6647 1059 6648
rect 1025 6642 1059 6647
rect 793 6621 967 6624
rect 786 6618 967 6621
rect 995 6641 1059 6642
rect 589 6598 608 6600
rect 623 6598 657 6600
rect 589 6582 669 6598
rect 589 6576 608 6582
rect 305 6550 408 6560
rect 259 6548 408 6550
rect 429 6548 464 6560
rect 98 6546 260 6548
rect 110 6526 129 6546
rect 144 6544 174 6546
rect -7 6518 34 6526
rect 116 6522 129 6526
rect 181 6530 260 6546
rect 292 6546 464 6548
rect 292 6530 371 6546
rect 378 6544 408 6546
rect -1 6508 28 6518
rect 43 6508 73 6522
rect 116 6508 159 6522
rect 181 6518 371 6530
rect 436 6526 442 6546
rect 166 6508 196 6518
rect 197 6508 355 6518
rect 359 6508 389 6518
rect 393 6508 423 6522
rect 451 6508 464 6546
rect 536 6560 565 6576
rect 579 6560 608 6576
rect 623 6566 653 6582
rect 681 6560 687 6608
rect 690 6602 709 6608
rect 724 6602 754 6610
rect 690 6594 754 6602
rect 690 6578 770 6594
rect 786 6587 848 6618
rect 864 6587 926 6618
rect 995 6616 1044 6641
rect 1059 6616 1089 6632
rect 958 6602 988 6610
rect 995 6608 1105 6616
rect 958 6594 1003 6602
rect 690 6576 709 6578
rect 724 6576 770 6578
rect 690 6560 770 6576
rect 797 6574 832 6587
rect 873 6584 910 6587
rect 873 6582 915 6584
rect 802 6571 832 6574
rect 811 6567 818 6571
rect 818 6566 819 6567
rect 777 6560 787 6566
rect 536 6552 571 6560
rect 536 6526 537 6552
rect 544 6526 571 6552
rect 479 6508 509 6522
rect 536 6518 571 6526
rect 573 6552 614 6560
rect 573 6526 588 6552
rect 595 6526 614 6552
rect 678 6548 709 6560
rect 724 6548 827 6560
rect 839 6550 865 6576
rect 880 6571 910 6582
rect 942 6578 1004 6594
rect 942 6576 988 6578
rect 942 6560 1004 6576
rect 1016 6560 1022 6608
rect 1025 6600 1105 6608
rect 1025 6598 1044 6600
rect 1059 6598 1093 6600
rect 1025 6582 1105 6598
rect 1025 6560 1044 6582
rect 1059 6566 1089 6582
rect 1117 6576 1123 6650
rect 1126 6576 1145 6720
rect 1160 6576 1166 6720
rect 1175 6650 1188 6720
rect 1240 6716 1262 6720
rect 1233 6694 1262 6708
rect 1315 6694 1331 6708
rect 1369 6704 1375 6706
rect 1382 6704 1490 6720
rect 1497 6704 1503 6706
rect 1511 6704 1526 6720
rect 1592 6714 1611 6717
rect 1233 6692 1331 6694
rect 1358 6692 1526 6704
rect 1541 6694 1557 6708
rect 1592 6695 1614 6714
rect 1624 6708 1640 6709
rect 1623 6706 1640 6708
rect 1624 6701 1640 6706
rect 1614 6694 1620 6695
rect 1623 6694 1652 6701
rect 1541 6693 1652 6694
rect 1541 6692 1658 6693
rect 1217 6684 1268 6692
rect 1315 6684 1349 6692
rect 1217 6672 1242 6684
rect 1249 6672 1268 6684
rect 1322 6682 1349 6684
rect 1358 6682 1579 6692
rect 1614 6689 1620 6692
rect 1322 6678 1579 6682
rect 1217 6664 1268 6672
rect 1315 6664 1579 6678
rect 1623 6684 1658 6692
rect 1169 6616 1188 6650
rect 1233 6656 1262 6664
rect 1233 6650 1250 6656
rect 1233 6648 1267 6650
rect 1315 6648 1331 6664
rect 1332 6654 1540 6664
rect 1541 6654 1557 6664
rect 1605 6660 1620 6675
rect 1623 6672 1624 6684
rect 1631 6672 1658 6684
rect 1623 6664 1658 6672
rect 1623 6663 1652 6664
rect 1343 6650 1557 6654
rect 1358 6648 1557 6650
rect 1592 6650 1605 6660
rect 1623 6650 1640 6663
rect 1592 6648 1640 6650
rect 1234 6644 1267 6648
rect 1230 6642 1267 6644
rect 1230 6641 1297 6642
rect 1230 6636 1261 6641
rect 1267 6636 1297 6641
rect 1230 6632 1297 6636
rect 1203 6629 1297 6632
rect 1203 6622 1252 6629
rect 1203 6616 1233 6622
rect 1252 6617 1257 6622
rect 1169 6600 1249 6616
rect 1261 6608 1297 6629
rect 1358 6624 1547 6648
rect 1592 6647 1639 6648
rect 1605 6642 1639 6647
rect 1373 6621 1547 6624
rect 1366 6618 1547 6621
rect 1575 6641 1639 6642
rect 1169 6598 1188 6600
rect 1203 6598 1237 6600
rect 1169 6582 1249 6598
rect 1169 6576 1188 6582
rect 885 6550 988 6560
rect 839 6548 988 6550
rect 1009 6548 1044 6560
rect 678 6546 840 6548
rect 690 6526 709 6546
rect 724 6544 754 6546
rect 573 6518 614 6526
rect 696 6522 709 6526
rect 761 6530 840 6546
rect 872 6546 1044 6548
rect 872 6530 951 6546
rect 958 6544 988 6546
rect 536 6508 565 6518
rect 579 6508 608 6518
rect 623 6508 653 6522
rect 696 6508 739 6522
rect 761 6518 951 6530
rect 1016 6526 1022 6546
rect 746 6508 776 6518
rect 777 6508 935 6518
rect 939 6508 969 6518
rect 973 6508 1003 6522
rect 1031 6508 1044 6546
rect 1116 6560 1145 6576
rect 1159 6560 1188 6576
rect 1203 6566 1233 6582
rect 1261 6560 1267 6608
rect 1270 6602 1289 6608
rect 1304 6602 1334 6610
rect 1270 6594 1334 6602
rect 1270 6578 1350 6594
rect 1366 6587 1428 6618
rect 1444 6587 1506 6618
rect 1575 6616 1624 6641
rect 1639 6616 1669 6632
rect 1538 6602 1568 6610
rect 1575 6608 1685 6616
rect 1538 6594 1583 6602
rect 1270 6576 1289 6578
rect 1304 6576 1350 6578
rect 1270 6560 1350 6576
rect 1377 6574 1412 6587
rect 1453 6584 1490 6587
rect 1453 6582 1495 6584
rect 1382 6571 1412 6574
rect 1391 6567 1398 6571
rect 1398 6566 1399 6567
rect 1357 6560 1367 6566
rect 1116 6552 1151 6560
rect 1116 6526 1117 6552
rect 1124 6526 1151 6552
rect 1059 6508 1089 6522
rect 1116 6518 1151 6526
rect 1153 6552 1194 6560
rect 1153 6526 1168 6552
rect 1175 6526 1194 6552
rect 1258 6548 1289 6560
rect 1304 6548 1407 6560
rect 1419 6550 1445 6576
rect 1460 6571 1490 6582
rect 1522 6578 1584 6594
rect 1522 6576 1568 6578
rect 1522 6560 1584 6576
rect 1596 6560 1602 6608
rect 1605 6600 1685 6608
rect 1605 6598 1624 6600
rect 1639 6598 1673 6600
rect 1605 6582 1685 6598
rect 1605 6560 1624 6582
rect 1639 6566 1669 6582
rect 1697 6576 1703 6650
rect 1706 6576 1725 6720
rect 1740 6576 1746 6720
rect 1755 6650 1768 6720
rect 1820 6716 1842 6720
rect 1813 6694 1842 6708
rect 1895 6694 1911 6708
rect 1949 6704 1955 6706
rect 1962 6704 2070 6720
rect 2077 6704 2083 6706
rect 2091 6704 2106 6720
rect 2172 6714 2191 6717
rect 1813 6692 1911 6694
rect 1938 6692 2106 6704
rect 2121 6694 2137 6708
rect 2172 6695 2194 6714
rect 2204 6708 2220 6709
rect 2203 6706 2220 6708
rect 2204 6701 2220 6706
rect 2194 6694 2200 6695
rect 2203 6694 2232 6701
rect 2121 6693 2232 6694
rect 2121 6692 2238 6693
rect 1797 6684 1848 6692
rect 1895 6684 1929 6692
rect 1797 6672 1822 6684
rect 1829 6672 1848 6684
rect 1902 6682 1929 6684
rect 1938 6682 2159 6692
rect 2194 6689 2200 6692
rect 1902 6678 2159 6682
rect 1797 6664 1848 6672
rect 1895 6664 2159 6678
rect 2203 6684 2238 6692
rect 1749 6616 1768 6650
rect 1813 6656 1842 6664
rect 1813 6650 1830 6656
rect 1813 6648 1847 6650
rect 1895 6648 1911 6664
rect 1912 6654 2120 6664
rect 2121 6654 2137 6664
rect 2185 6660 2200 6675
rect 2203 6672 2204 6684
rect 2211 6672 2238 6684
rect 2203 6664 2238 6672
rect 2203 6663 2232 6664
rect 1923 6650 2137 6654
rect 1938 6648 2137 6650
rect 2172 6650 2185 6660
rect 2203 6650 2220 6663
rect 2172 6648 2220 6650
rect 1814 6644 1847 6648
rect 1810 6642 1847 6644
rect 1810 6641 1877 6642
rect 1810 6636 1841 6641
rect 1847 6636 1877 6641
rect 1810 6632 1877 6636
rect 1783 6629 1877 6632
rect 1783 6622 1832 6629
rect 1783 6616 1813 6622
rect 1832 6617 1837 6622
rect 1749 6600 1829 6616
rect 1841 6608 1877 6629
rect 1938 6624 2127 6648
rect 2172 6647 2219 6648
rect 2185 6642 2219 6647
rect 1953 6621 2127 6624
rect 1946 6618 2127 6621
rect 2155 6641 2219 6642
rect 1749 6598 1768 6600
rect 1783 6598 1817 6600
rect 1749 6582 1829 6598
rect 1749 6576 1768 6582
rect 1465 6550 1568 6560
rect 1419 6548 1568 6550
rect 1589 6548 1624 6560
rect 1258 6546 1420 6548
rect 1270 6526 1289 6546
rect 1304 6544 1334 6546
rect 1153 6518 1194 6526
rect 1276 6522 1289 6526
rect 1341 6530 1420 6546
rect 1452 6546 1624 6548
rect 1452 6530 1531 6546
rect 1538 6544 1568 6546
rect 1116 6508 1145 6518
rect 1159 6508 1188 6518
rect 1203 6508 1233 6522
rect 1276 6508 1319 6522
rect 1341 6518 1531 6530
rect 1596 6526 1602 6546
rect 1326 6508 1356 6518
rect 1357 6508 1515 6518
rect 1519 6508 1549 6518
rect 1553 6508 1583 6522
rect 1611 6508 1624 6546
rect 1696 6560 1725 6576
rect 1739 6560 1768 6576
rect 1783 6566 1813 6582
rect 1841 6560 1847 6608
rect 1850 6602 1869 6608
rect 1884 6602 1914 6610
rect 1850 6594 1914 6602
rect 1850 6578 1930 6594
rect 1946 6587 2008 6618
rect 2024 6587 2086 6618
rect 2155 6616 2204 6641
rect 2219 6616 2249 6632
rect 2118 6602 2148 6610
rect 2155 6608 2265 6616
rect 2118 6594 2163 6602
rect 1850 6576 1869 6578
rect 1884 6576 1930 6578
rect 1850 6560 1930 6576
rect 1957 6574 1992 6587
rect 2033 6584 2070 6587
rect 2033 6582 2075 6584
rect 1962 6571 1992 6574
rect 1971 6567 1978 6571
rect 1978 6566 1979 6567
rect 1937 6560 1947 6566
rect 1696 6552 1731 6560
rect 1696 6526 1697 6552
rect 1704 6526 1731 6552
rect 1639 6508 1669 6522
rect 1696 6518 1731 6526
rect 1733 6552 1774 6560
rect 1733 6526 1748 6552
rect 1755 6526 1774 6552
rect 1838 6548 1869 6560
rect 1884 6548 1987 6560
rect 1999 6550 2025 6576
rect 2040 6571 2070 6582
rect 2102 6578 2164 6594
rect 2102 6576 2148 6578
rect 2102 6560 2164 6576
rect 2176 6560 2182 6608
rect 2185 6600 2265 6608
rect 2185 6598 2204 6600
rect 2219 6598 2253 6600
rect 2185 6582 2265 6598
rect 2185 6560 2204 6582
rect 2219 6566 2249 6582
rect 2277 6576 2283 6650
rect 2286 6576 2305 6720
rect 2320 6576 2326 6720
rect 2335 6650 2348 6720
rect 2400 6716 2422 6720
rect 2393 6694 2422 6708
rect 2475 6694 2491 6708
rect 2529 6704 2535 6706
rect 2542 6704 2650 6720
rect 2657 6704 2663 6706
rect 2671 6704 2686 6720
rect 2752 6714 2771 6717
rect 2393 6692 2491 6694
rect 2518 6692 2686 6704
rect 2701 6694 2717 6708
rect 2752 6695 2774 6714
rect 2784 6708 2800 6709
rect 2783 6706 2800 6708
rect 2784 6701 2800 6706
rect 2774 6694 2780 6695
rect 2783 6694 2812 6701
rect 2701 6693 2812 6694
rect 2701 6692 2818 6693
rect 2377 6684 2428 6692
rect 2475 6684 2509 6692
rect 2377 6672 2402 6684
rect 2409 6672 2428 6684
rect 2482 6682 2509 6684
rect 2518 6682 2739 6692
rect 2774 6689 2780 6692
rect 2482 6678 2739 6682
rect 2377 6664 2428 6672
rect 2475 6664 2739 6678
rect 2783 6684 2818 6692
rect 2329 6616 2348 6650
rect 2393 6656 2422 6664
rect 2393 6650 2410 6656
rect 2393 6648 2427 6650
rect 2475 6648 2491 6664
rect 2492 6654 2700 6664
rect 2701 6654 2717 6664
rect 2765 6660 2780 6675
rect 2783 6672 2784 6684
rect 2791 6672 2818 6684
rect 2783 6664 2818 6672
rect 2783 6663 2812 6664
rect 2503 6650 2717 6654
rect 2518 6648 2717 6650
rect 2752 6650 2765 6660
rect 2783 6650 2800 6663
rect 2752 6648 2800 6650
rect 2394 6644 2427 6648
rect 2390 6642 2427 6644
rect 2390 6641 2457 6642
rect 2390 6636 2421 6641
rect 2427 6636 2457 6641
rect 2390 6632 2457 6636
rect 2363 6629 2457 6632
rect 2363 6622 2412 6629
rect 2363 6616 2393 6622
rect 2412 6617 2417 6622
rect 2329 6600 2409 6616
rect 2421 6608 2457 6629
rect 2518 6624 2707 6648
rect 2752 6647 2799 6648
rect 2765 6642 2799 6647
rect 2533 6621 2707 6624
rect 2526 6618 2707 6621
rect 2735 6641 2799 6642
rect 2329 6598 2348 6600
rect 2363 6598 2397 6600
rect 2329 6582 2409 6598
rect 2329 6576 2348 6582
rect 2045 6550 2148 6560
rect 1999 6548 2148 6550
rect 2169 6548 2204 6560
rect 1838 6546 2000 6548
rect 1850 6526 1869 6546
rect 1884 6544 1914 6546
rect 1733 6518 1774 6526
rect 1856 6522 1869 6526
rect 1921 6530 2000 6546
rect 2032 6546 2204 6548
rect 2032 6530 2111 6546
rect 2118 6544 2148 6546
rect 1696 6508 1725 6518
rect 1739 6508 1768 6518
rect 1783 6508 1813 6522
rect 1856 6508 1899 6522
rect 1921 6518 2111 6530
rect 2176 6526 2182 6546
rect 1906 6508 1936 6518
rect 1937 6508 2095 6518
rect 2099 6508 2129 6518
rect 2133 6508 2163 6522
rect 2191 6508 2204 6546
rect 2276 6560 2305 6576
rect 2319 6560 2348 6576
rect 2363 6566 2393 6582
rect 2421 6560 2427 6608
rect 2430 6602 2449 6608
rect 2464 6602 2494 6610
rect 2430 6594 2494 6602
rect 2430 6578 2510 6594
rect 2526 6587 2588 6618
rect 2604 6587 2666 6618
rect 2735 6616 2784 6641
rect 2799 6616 2829 6632
rect 2698 6602 2728 6610
rect 2735 6608 2845 6616
rect 2698 6594 2743 6602
rect 2430 6576 2449 6578
rect 2464 6576 2510 6578
rect 2430 6560 2510 6576
rect 2537 6574 2572 6587
rect 2613 6584 2650 6587
rect 2613 6582 2655 6584
rect 2542 6571 2572 6574
rect 2551 6567 2558 6571
rect 2558 6566 2559 6567
rect 2517 6560 2527 6566
rect 2276 6552 2311 6560
rect 2276 6526 2277 6552
rect 2284 6526 2311 6552
rect 2219 6508 2249 6522
rect 2276 6518 2311 6526
rect 2313 6552 2354 6560
rect 2313 6526 2328 6552
rect 2335 6526 2354 6552
rect 2418 6548 2449 6560
rect 2464 6548 2567 6560
rect 2579 6550 2605 6576
rect 2620 6571 2650 6582
rect 2682 6578 2744 6594
rect 2682 6576 2728 6578
rect 2682 6560 2744 6576
rect 2756 6560 2762 6608
rect 2765 6600 2845 6608
rect 2765 6598 2784 6600
rect 2799 6598 2833 6600
rect 2765 6582 2845 6598
rect 2765 6560 2784 6582
rect 2799 6566 2829 6582
rect 2857 6576 2863 6650
rect 2866 6576 2885 6720
rect 2900 6576 2906 6720
rect 2915 6650 2928 6720
rect 2980 6716 3002 6720
rect 2973 6694 3002 6708
rect 3055 6694 3071 6708
rect 3109 6704 3115 6706
rect 3122 6704 3230 6720
rect 3237 6704 3243 6706
rect 3251 6704 3266 6720
rect 3332 6714 3351 6717
rect 2973 6692 3071 6694
rect 3098 6692 3266 6704
rect 3281 6694 3297 6708
rect 3332 6695 3354 6714
rect 3364 6708 3380 6709
rect 3363 6706 3380 6708
rect 3364 6701 3380 6706
rect 3354 6694 3360 6695
rect 3363 6694 3392 6701
rect 3281 6693 3392 6694
rect 3281 6692 3398 6693
rect 2957 6684 3008 6692
rect 3055 6684 3089 6692
rect 2957 6672 2982 6684
rect 2989 6672 3008 6684
rect 3062 6682 3089 6684
rect 3098 6682 3319 6692
rect 3354 6689 3360 6692
rect 3062 6678 3319 6682
rect 2957 6664 3008 6672
rect 3055 6664 3319 6678
rect 3363 6684 3398 6692
rect 2909 6616 2928 6650
rect 2973 6656 3002 6664
rect 2973 6650 2990 6656
rect 2973 6648 3007 6650
rect 3055 6648 3071 6664
rect 3072 6654 3280 6664
rect 3281 6654 3297 6664
rect 3345 6660 3360 6675
rect 3363 6672 3364 6684
rect 3371 6672 3398 6684
rect 3363 6664 3398 6672
rect 3363 6663 3392 6664
rect 3083 6650 3297 6654
rect 3098 6648 3297 6650
rect 3332 6650 3345 6660
rect 3363 6650 3380 6663
rect 3332 6648 3380 6650
rect 2974 6644 3007 6648
rect 2970 6642 3007 6644
rect 2970 6641 3037 6642
rect 2970 6636 3001 6641
rect 3007 6636 3037 6641
rect 2970 6632 3037 6636
rect 2943 6629 3037 6632
rect 2943 6622 2992 6629
rect 2943 6616 2973 6622
rect 2992 6617 2997 6622
rect 2909 6600 2989 6616
rect 3001 6608 3037 6629
rect 3098 6624 3287 6648
rect 3332 6647 3379 6648
rect 3345 6642 3379 6647
rect 3113 6621 3287 6624
rect 3106 6618 3287 6621
rect 3315 6641 3379 6642
rect 2909 6598 2928 6600
rect 2943 6598 2977 6600
rect 2909 6582 2989 6598
rect 2909 6576 2928 6582
rect 2625 6550 2728 6560
rect 2579 6548 2728 6550
rect 2749 6548 2784 6560
rect 2418 6546 2580 6548
rect 2430 6526 2449 6546
rect 2464 6544 2494 6546
rect 2313 6518 2354 6526
rect 2436 6522 2449 6526
rect 2501 6530 2580 6546
rect 2612 6546 2784 6548
rect 2612 6530 2691 6546
rect 2698 6544 2728 6546
rect 2276 6508 2305 6518
rect 2319 6508 2348 6518
rect 2363 6508 2393 6522
rect 2436 6508 2479 6522
rect 2501 6518 2691 6530
rect 2756 6526 2762 6546
rect 2486 6508 2516 6518
rect 2517 6508 2675 6518
rect 2679 6508 2709 6518
rect 2713 6508 2743 6522
rect 2771 6508 2784 6546
rect 2856 6560 2885 6576
rect 2899 6560 2928 6576
rect 2943 6566 2973 6582
rect 3001 6560 3007 6608
rect 3010 6602 3029 6608
rect 3044 6602 3074 6610
rect 3010 6594 3074 6602
rect 3010 6578 3090 6594
rect 3106 6587 3168 6618
rect 3184 6587 3246 6618
rect 3315 6616 3364 6641
rect 3379 6616 3409 6632
rect 3278 6602 3308 6610
rect 3315 6608 3425 6616
rect 3278 6594 3323 6602
rect 3010 6576 3029 6578
rect 3044 6576 3090 6578
rect 3010 6560 3090 6576
rect 3117 6574 3152 6587
rect 3193 6584 3230 6587
rect 3193 6582 3235 6584
rect 3122 6571 3152 6574
rect 3131 6567 3138 6571
rect 3138 6566 3139 6567
rect 3097 6560 3107 6566
rect 2856 6552 2891 6560
rect 2856 6526 2857 6552
rect 2864 6526 2891 6552
rect 2799 6508 2829 6522
rect 2856 6518 2891 6526
rect 2893 6552 2934 6560
rect 2893 6526 2908 6552
rect 2915 6526 2934 6552
rect 2998 6548 3029 6560
rect 3044 6548 3147 6560
rect 3159 6550 3185 6576
rect 3200 6571 3230 6582
rect 3262 6578 3324 6594
rect 3262 6576 3308 6578
rect 3262 6560 3324 6576
rect 3336 6560 3342 6608
rect 3345 6600 3425 6608
rect 3345 6598 3364 6600
rect 3379 6598 3413 6600
rect 3345 6582 3425 6598
rect 3345 6560 3364 6582
rect 3379 6566 3409 6582
rect 3437 6576 3443 6650
rect 3446 6576 3465 6720
rect 3480 6576 3486 6720
rect 3495 6650 3508 6720
rect 3560 6716 3582 6720
rect 3553 6694 3582 6708
rect 3635 6694 3651 6708
rect 3689 6704 3695 6706
rect 3702 6704 3810 6720
rect 3817 6704 3823 6706
rect 3831 6704 3846 6720
rect 3912 6714 3931 6717
rect 3553 6692 3651 6694
rect 3678 6692 3846 6704
rect 3861 6694 3877 6708
rect 3912 6695 3934 6714
rect 3944 6708 3960 6709
rect 3943 6706 3960 6708
rect 3944 6701 3960 6706
rect 3934 6694 3940 6695
rect 3943 6694 3972 6701
rect 3861 6693 3972 6694
rect 3861 6692 3978 6693
rect 3537 6684 3588 6692
rect 3635 6684 3669 6692
rect 3537 6672 3562 6684
rect 3569 6672 3588 6684
rect 3642 6682 3669 6684
rect 3678 6682 3899 6692
rect 3934 6689 3940 6692
rect 3642 6678 3899 6682
rect 3537 6664 3588 6672
rect 3635 6664 3899 6678
rect 3943 6684 3978 6692
rect 3489 6616 3508 6650
rect 3553 6656 3582 6664
rect 3553 6650 3570 6656
rect 3553 6648 3587 6650
rect 3635 6648 3651 6664
rect 3652 6654 3860 6664
rect 3861 6654 3877 6664
rect 3925 6660 3940 6675
rect 3943 6672 3944 6684
rect 3951 6672 3978 6684
rect 3943 6664 3978 6672
rect 3943 6663 3972 6664
rect 3663 6650 3877 6654
rect 3678 6648 3877 6650
rect 3912 6650 3925 6660
rect 3943 6650 3960 6663
rect 3912 6648 3960 6650
rect 3554 6644 3587 6648
rect 3550 6642 3587 6644
rect 3550 6641 3617 6642
rect 3550 6636 3581 6641
rect 3587 6636 3617 6641
rect 3550 6632 3617 6636
rect 3523 6629 3617 6632
rect 3523 6622 3572 6629
rect 3523 6616 3553 6622
rect 3572 6617 3577 6622
rect 3489 6600 3569 6616
rect 3581 6608 3617 6629
rect 3678 6624 3867 6648
rect 3912 6647 3959 6648
rect 3925 6642 3959 6647
rect 3693 6621 3867 6624
rect 3686 6618 3867 6621
rect 3895 6641 3959 6642
rect 3489 6598 3508 6600
rect 3523 6598 3557 6600
rect 3489 6582 3569 6598
rect 3489 6576 3508 6582
rect 3205 6550 3308 6560
rect 3159 6548 3308 6550
rect 3329 6548 3364 6560
rect 2998 6546 3160 6548
rect 3010 6526 3029 6546
rect 3044 6544 3074 6546
rect 2893 6518 2934 6526
rect 3016 6522 3029 6526
rect 3081 6530 3160 6546
rect 3192 6546 3364 6548
rect 3192 6530 3271 6546
rect 3278 6544 3308 6546
rect 2856 6508 2885 6518
rect 2899 6508 2928 6518
rect 2943 6508 2973 6522
rect 3016 6508 3059 6522
rect 3081 6518 3271 6530
rect 3336 6526 3342 6546
rect 3066 6508 3096 6518
rect 3097 6508 3255 6518
rect 3259 6508 3289 6518
rect 3293 6508 3323 6522
rect 3351 6508 3364 6546
rect 3436 6560 3465 6576
rect 3479 6560 3508 6576
rect 3523 6566 3553 6582
rect 3581 6560 3587 6608
rect 3590 6602 3609 6608
rect 3624 6602 3654 6610
rect 3590 6594 3654 6602
rect 3590 6578 3670 6594
rect 3686 6587 3748 6618
rect 3764 6587 3826 6618
rect 3895 6616 3944 6641
rect 3959 6616 3989 6632
rect 3858 6602 3888 6610
rect 3895 6608 4005 6616
rect 3858 6594 3903 6602
rect 3590 6576 3609 6578
rect 3624 6576 3670 6578
rect 3590 6560 3670 6576
rect 3697 6574 3732 6587
rect 3773 6584 3810 6587
rect 3773 6582 3815 6584
rect 3702 6571 3732 6574
rect 3711 6567 3718 6571
rect 3718 6566 3719 6567
rect 3677 6560 3687 6566
rect 3436 6552 3471 6560
rect 3436 6526 3437 6552
rect 3444 6526 3471 6552
rect 3379 6508 3409 6522
rect 3436 6518 3471 6526
rect 3473 6552 3514 6560
rect 3473 6526 3488 6552
rect 3495 6526 3514 6552
rect 3578 6548 3609 6560
rect 3624 6548 3727 6560
rect 3739 6550 3765 6576
rect 3780 6571 3810 6582
rect 3842 6578 3904 6594
rect 3842 6576 3888 6578
rect 3842 6560 3904 6576
rect 3916 6560 3922 6608
rect 3925 6600 4005 6608
rect 3925 6598 3944 6600
rect 3959 6598 3993 6600
rect 3925 6582 4005 6598
rect 3925 6560 3944 6582
rect 3959 6566 3989 6582
rect 4017 6576 4023 6650
rect 4026 6576 4045 6720
rect 4060 6576 4066 6720
rect 4075 6650 4088 6720
rect 4140 6716 4162 6720
rect 4133 6694 4162 6708
rect 4215 6694 4231 6708
rect 4269 6704 4275 6706
rect 4282 6704 4390 6720
rect 4397 6704 4403 6706
rect 4411 6704 4426 6720
rect 4492 6714 4511 6717
rect 4133 6692 4231 6694
rect 4258 6692 4426 6704
rect 4441 6694 4457 6708
rect 4492 6695 4514 6714
rect 4524 6708 4540 6709
rect 4523 6706 4540 6708
rect 4524 6701 4540 6706
rect 4514 6694 4520 6695
rect 4523 6694 4552 6701
rect 4441 6693 4552 6694
rect 4441 6692 4558 6693
rect 4117 6684 4168 6692
rect 4215 6684 4249 6692
rect 4117 6672 4142 6684
rect 4149 6672 4168 6684
rect 4222 6682 4249 6684
rect 4258 6682 4479 6692
rect 4514 6689 4520 6692
rect 4222 6678 4479 6682
rect 4117 6664 4168 6672
rect 4215 6664 4479 6678
rect 4523 6684 4558 6692
rect 4069 6616 4088 6650
rect 4133 6656 4162 6664
rect 4133 6650 4150 6656
rect 4133 6648 4167 6650
rect 4215 6648 4231 6664
rect 4232 6654 4440 6664
rect 4441 6654 4457 6664
rect 4505 6660 4520 6675
rect 4523 6672 4524 6684
rect 4531 6672 4558 6684
rect 4523 6664 4558 6672
rect 4523 6663 4552 6664
rect 4243 6650 4457 6654
rect 4258 6648 4457 6650
rect 4492 6650 4505 6660
rect 4523 6650 4540 6663
rect 4492 6648 4540 6650
rect 4134 6644 4167 6648
rect 4130 6642 4167 6644
rect 4130 6641 4197 6642
rect 4130 6636 4161 6641
rect 4167 6636 4197 6641
rect 4130 6632 4197 6636
rect 4103 6629 4197 6632
rect 4103 6622 4152 6629
rect 4103 6616 4133 6622
rect 4152 6617 4157 6622
rect 4069 6600 4149 6616
rect 4161 6608 4197 6629
rect 4258 6624 4447 6648
rect 4492 6647 4539 6648
rect 4505 6642 4539 6647
rect 4273 6621 4447 6624
rect 4266 6618 4447 6621
rect 4475 6641 4539 6642
rect 4069 6598 4088 6600
rect 4103 6598 4137 6600
rect 4069 6582 4149 6598
rect 4069 6576 4088 6582
rect 3785 6550 3888 6560
rect 3739 6548 3888 6550
rect 3909 6548 3944 6560
rect 3578 6546 3740 6548
rect 3590 6526 3609 6546
rect 3624 6544 3654 6546
rect 3473 6518 3514 6526
rect 3596 6522 3609 6526
rect 3661 6530 3740 6546
rect 3772 6546 3944 6548
rect 3772 6530 3851 6546
rect 3858 6544 3888 6546
rect 3436 6508 3465 6518
rect 3479 6508 3508 6518
rect 3523 6508 3553 6522
rect 3596 6508 3639 6522
rect 3661 6518 3851 6530
rect 3916 6526 3922 6546
rect 3646 6508 3676 6518
rect 3677 6508 3835 6518
rect 3839 6508 3869 6518
rect 3873 6508 3903 6522
rect 3931 6508 3944 6546
rect 4016 6560 4045 6576
rect 4059 6560 4088 6576
rect 4103 6566 4133 6582
rect 4161 6560 4167 6608
rect 4170 6602 4189 6608
rect 4204 6602 4234 6610
rect 4170 6594 4234 6602
rect 4170 6578 4250 6594
rect 4266 6587 4328 6618
rect 4344 6587 4406 6618
rect 4475 6616 4524 6641
rect 4539 6616 4569 6632
rect 4438 6602 4468 6610
rect 4475 6608 4585 6616
rect 4438 6594 4483 6602
rect 4170 6576 4189 6578
rect 4204 6576 4250 6578
rect 4170 6560 4250 6576
rect 4277 6574 4312 6587
rect 4353 6584 4390 6587
rect 4353 6582 4395 6584
rect 4282 6571 4312 6574
rect 4291 6567 4298 6571
rect 4298 6566 4299 6567
rect 4257 6560 4267 6566
rect 4016 6552 4051 6560
rect 4016 6526 4017 6552
rect 4024 6526 4051 6552
rect 3959 6508 3989 6522
rect 4016 6518 4051 6526
rect 4053 6552 4094 6560
rect 4053 6526 4068 6552
rect 4075 6526 4094 6552
rect 4158 6548 4189 6560
rect 4204 6548 4307 6560
rect 4319 6550 4345 6576
rect 4360 6571 4390 6582
rect 4422 6578 4484 6594
rect 4422 6576 4468 6578
rect 4422 6560 4484 6576
rect 4496 6560 4502 6608
rect 4505 6600 4585 6608
rect 4505 6598 4524 6600
rect 4539 6598 4573 6600
rect 4505 6582 4585 6598
rect 4505 6560 4524 6582
rect 4539 6566 4569 6582
rect 4597 6576 4603 6650
rect 4606 6576 4625 6720
rect 4640 6576 4646 6720
rect 4655 6650 4668 6720
rect 4720 6716 4742 6720
rect 4713 6694 4742 6708
rect 4795 6694 4811 6708
rect 4849 6704 4855 6706
rect 4862 6704 4970 6720
rect 4977 6704 4983 6706
rect 4991 6704 5006 6720
rect 5072 6714 5091 6717
rect 4713 6692 4811 6694
rect 4838 6692 5006 6704
rect 5021 6694 5037 6708
rect 5072 6695 5094 6714
rect 5104 6708 5120 6709
rect 5103 6706 5120 6708
rect 5104 6701 5120 6706
rect 5094 6694 5100 6695
rect 5103 6694 5132 6701
rect 5021 6693 5132 6694
rect 5021 6692 5138 6693
rect 4697 6684 4748 6692
rect 4795 6684 4829 6692
rect 4697 6672 4722 6684
rect 4729 6672 4748 6684
rect 4802 6682 4829 6684
rect 4838 6682 5059 6692
rect 5094 6689 5100 6692
rect 4802 6678 5059 6682
rect 4697 6664 4748 6672
rect 4795 6664 5059 6678
rect 5103 6684 5138 6692
rect 4649 6616 4668 6650
rect 4713 6656 4742 6664
rect 4713 6650 4730 6656
rect 4713 6648 4747 6650
rect 4795 6648 4811 6664
rect 4812 6654 5020 6664
rect 5021 6654 5037 6664
rect 5085 6660 5100 6675
rect 5103 6672 5104 6684
rect 5111 6672 5138 6684
rect 5103 6664 5138 6672
rect 5103 6663 5132 6664
rect 4823 6650 5037 6654
rect 4838 6648 5037 6650
rect 5072 6650 5085 6660
rect 5103 6650 5120 6663
rect 5072 6648 5120 6650
rect 4714 6644 4747 6648
rect 4710 6642 4747 6644
rect 4710 6641 4777 6642
rect 4710 6636 4741 6641
rect 4747 6636 4777 6641
rect 4710 6632 4777 6636
rect 4683 6629 4777 6632
rect 4683 6622 4732 6629
rect 4683 6616 4713 6622
rect 4732 6617 4737 6622
rect 4649 6600 4729 6616
rect 4741 6608 4777 6629
rect 4838 6624 5027 6648
rect 5072 6647 5119 6648
rect 5085 6642 5119 6647
rect 4853 6621 5027 6624
rect 4846 6618 5027 6621
rect 5055 6641 5119 6642
rect 4649 6598 4668 6600
rect 4683 6598 4717 6600
rect 4649 6582 4729 6598
rect 4649 6576 4668 6582
rect 4365 6550 4468 6560
rect 4319 6548 4468 6550
rect 4489 6548 4524 6560
rect 4158 6546 4320 6548
rect 4170 6526 4189 6546
rect 4204 6544 4234 6546
rect 4053 6518 4094 6526
rect 4176 6522 4189 6526
rect 4241 6530 4320 6546
rect 4352 6546 4524 6548
rect 4352 6530 4431 6546
rect 4438 6544 4468 6546
rect 4016 6508 4045 6518
rect 4059 6508 4088 6518
rect 4103 6508 4133 6522
rect 4176 6508 4219 6522
rect 4241 6518 4431 6530
rect 4496 6526 4502 6546
rect 4226 6508 4256 6518
rect 4257 6508 4415 6518
rect 4419 6508 4449 6518
rect 4453 6508 4483 6522
rect 4511 6508 4524 6546
rect 4596 6560 4625 6576
rect 4639 6560 4668 6576
rect 4683 6566 4713 6582
rect 4741 6560 4747 6608
rect 4750 6602 4769 6608
rect 4784 6602 4814 6610
rect 4750 6594 4814 6602
rect 4750 6578 4830 6594
rect 4846 6587 4908 6618
rect 4924 6587 4986 6618
rect 5055 6616 5104 6641
rect 5119 6616 5149 6632
rect 5018 6602 5048 6610
rect 5055 6608 5165 6616
rect 5018 6594 5063 6602
rect 4750 6576 4769 6578
rect 4784 6576 4830 6578
rect 4750 6560 4830 6576
rect 4857 6574 4892 6587
rect 4933 6584 4970 6587
rect 4933 6582 4975 6584
rect 4862 6571 4892 6574
rect 4871 6567 4878 6571
rect 4878 6566 4879 6567
rect 4837 6560 4847 6566
rect 4596 6552 4631 6560
rect 4596 6526 4597 6552
rect 4604 6526 4631 6552
rect 4539 6508 4569 6522
rect 4596 6518 4631 6526
rect 4633 6552 4674 6560
rect 4633 6526 4648 6552
rect 4655 6526 4674 6552
rect 4738 6548 4769 6560
rect 4784 6548 4887 6560
rect 4899 6550 4925 6576
rect 4940 6571 4970 6582
rect 5002 6578 5064 6594
rect 5002 6576 5048 6578
rect 5002 6560 5064 6576
rect 5076 6560 5082 6608
rect 5085 6600 5165 6608
rect 5085 6598 5104 6600
rect 5119 6598 5153 6600
rect 5085 6582 5165 6598
rect 5085 6560 5104 6582
rect 5119 6566 5149 6582
rect 5177 6576 5183 6650
rect 5186 6576 5205 6720
rect 5220 6576 5226 6720
rect 5235 6650 5248 6720
rect 5300 6716 5322 6720
rect 5293 6694 5322 6708
rect 5375 6694 5391 6708
rect 5429 6704 5435 6706
rect 5442 6704 5550 6720
rect 5557 6704 5563 6706
rect 5571 6704 5586 6720
rect 5652 6714 5671 6717
rect 5293 6692 5391 6694
rect 5418 6692 5586 6704
rect 5601 6694 5617 6708
rect 5652 6695 5674 6714
rect 5684 6708 5700 6709
rect 5683 6706 5700 6708
rect 5684 6701 5700 6706
rect 5674 6694 5680 6695
rect 5683 6694 5712 6701
rect 5601 6693 5712 6694
rect 5601 6692 5718 6693
rect 5277 6684 5328 6692
rect 5375 6684 5409 6692
rect 5277 6672 5302 6684
rect 5309 6672 5328 6684
rect 5382 6682 5409 6684
rect 5418 6682 5639 6692
rect 5674 6689 5680 6692
rect 5382 6678 5639 6682
rect 5277 6664 5328 6672
rect 5375 6664 5639 6678
rect 5683 6684 5718 6692
rect 5229 6616 5248 6650
rect 5293 6656 5322 6664
rect 5293 6650 5310 6656
rect 5293 6648 5327 6650
rect 5375 6648 5391 6664
rect 5392 6654 5600 6664
rect 5601 6654 5617 6664
rect 5665 6660 5680 6675
rect 5683 6672 5684 6684
rect 5691 6672 5718 6684
rect 5683 6664 5718 6672
rect 5683 6663 5712 6664
rect 5403 6650 5617 6654
rect 5418 6648 5617 6650
rect 5652 6650 5665 6660
rect 5683 6650 5700 6663
rect 5652 6648 5700 6650
rect 5294 6644 5327 6648
rect 5290 6642 5327 6644
rect 5290 6641 5357 6642
rect 5290 6636 5321 6641
rect 5327 6636 5357 6641
rect 5290 6632 5357 6636
rect 5263 6629 5357 6632
rect 5263 6622 5312 6629
rect 5263 6616 5293 6622
rect 5312 6617 5317 6622
rect 5229 6600 5309 6616
rect 5321 6608 5357 6629
rect 5418 6624 5607 6648
rect 5652 6647 5699 6648
rect 5665 6642 5699 6647
rect 5433 6621 5607 6624
rect 5426 6618 5607 6621
rect 5635 6641 5699 6642
rect 5229 6598 5248 6600
rect 5263 6598 5297 6600
rect 5229 6582 5309 6598
rect 5229 6576 5248 6582
rect 4945 6550 5048 6560
rect 4899 6548 5048 6550
rect 5069 6548 5104 6560
rect 4738 6546 4900 6548
rect 4750 6526 4769 6546
rect 4784 6544 4814 6546
rect 4633 6518 4674 6526
rect 4756 6522 4769 6526
rect 4821 6530 4900 6546
rect 4932 6546 5104 6548
rect 4932 6530 5011 6546
rect 5018 6544 5048 6546
rect 4596 6508 4625 6518
rect 4639 6508 4668 6518
rect 4683 6508 4713 6522
rect 4756 6508 4799 6522
rect 4821 6518 5011 6530
rect 5076 6526 5082 6546
rect 4806 6508 4836 6518
rect 4837 6508 4995 6518
rect 4999 6508 5029 6518
rect 5033 6508 5063 6522
rect 5091 6508 5104 6546
rect 5176 6560 5205 6576
rect 5219 6560 5248 6576
rect 5263 6566 5293 6582
rect 5321 6560 5327 6608
rect 5330 6602 5349 6608
rect 5364 6602 5394 6610
rect 5330 6594 5394 6602
rect 5330 6578 5410 6594
rect 5426 6587 5488 6618
rect 5504 6587 5566 6618
rect 5635 6616 5684 6641
rect 5699 6616 5729 6632
rect 5598 6602 5628 6610
rect 5635 6608 5745 6616
rect 5598 6594 5643 6602
rect 5330 6576 5349 6578
rect 5364 6576 5410 6578
rect 5330 6560 5410 6576
rect 5437 6574 5472 6587
rect 5513 6584 5550 6587
rect 5513 6582 5555 6584
rect 5442 6571 5472 6574
rect 5451 6567 5458 6571
rect 5458 6566 5459 6567
rect 5417 6560 5427 6566
rect 5176 6552 5211 6560
rect 5176 6526 5177 6552
rect 5184 6526 5211 6552
rect 5119 6508 5149 6522
rect 5176 6518 5211 6526
rect 5213 6552 5254 6560
rect 5213 6526 5228 6552
rect 5235 6526 5254 6552
rect 5318 6548 5349 6560
rect 5364 6548 5467 6560
rect 5479 6550 5505 6576
rect 5520 6571 5550 6582
rect 5582 6578 5644 6594
rect 5582 6576 5628 6578
rect 5582 6560 5644 6576
rect 5656 6560 5662 6608
rect 5665 6600 5745 6608
rect 5665 6598 5684 6600
rect 5699 6598 5733 6600
rect 5665 6582 5745 6598
rect 5665 6560 5684 6582
rect 5699 6566 5729 6582
rect 5757 6576 5763 6650
rect 5766 6576 5785 6720
rect 5800 6576 5806 6720
rect 5815 6650 5828 6720
rect 5880 6716 5902 6720
rect 5873 6694 5902 6708
rect 5955 6694 5971 6708
rect 6009 6704 6015 6706
rect 6022 6704 6130 6720
rect 6137 6704 6143 6706
rect 6151 6704 6166 6720
rect 6232 6714 6251 6717
rect 5873 6692 5971 6694
rect 5998 6692 6166 6704
rect 6181 6694 6197 6708
rect 6232 6695 6254 6714
rect 6264 6708 6280 6709
rect 6263 6706 6280 6708
rect 6264 6701 6280 6706
rect 6254 6694 6260 6695
rect 6263 6694 6292 6701
rect 6181 6693 6292 6694
rect 6181 6692 6298 6693
rect 5857 6684 5908 6692
rect 5955 6684 5989 6692
rect 5857 6672 5882 6684
rect 5889 6672 5908 6684
rect 5962 6682 5989 6684
rect 5998 6682 6219 6692
rect 6254 6689 6260 6692
rect 5962 6678 6219 6682
rect 5857 6664 5908 6672
rect 5955 6664 6219 6678
rect 6263 6684 6298 6692
rect 5809 6616 5828 6650
rect 5873 6656 5902 6664
rect 5873 6650 5890 6656
rect 5873 6648 5907 6650
rect 5955 6648 5971 6664
rect 5972 6654 6180 6664
rect 6181 6654 6197 6664
rect 6245 6660 6260 6675
rect 6263 6672 6264 6684
rect 6271 6672 6298 6684
rect 6263 6664 6298 6672
rect 6263 6663 6292 6664
rect 5983 6650 6197 6654
rect 5998 6648 6197 6650
rect 6232 6650 6245 6660
rect 6263 6650 6280 6663
rect 6232 6648 6280 6650
rect 5874 6644 5907 6648
rect 5870 6642 5907 6644
rect 5870 6641 5937 6642
rect 5870 6636 5901 6641
rect 5907 6636 5937 6641
rect 5870 6632 5937 6636
rect 5843 6629 5937 6632
rect 5843 6622 5892 6629
rect 5843 6616 5873 6622
rect 5892 6617 5897 6622
rect 5809 6600 5889 6616
rect 5901 6608 5937 6629
rect 5998 6624 6187 6648
rect 6232 6647 6279 6648
rect 6245 6642 6279 6647
rect 6013 6621 6187 6624
rect 6006 6618 6187 6621
rect 6215 6641 6279 6642
rect 5809 6598 5828 6600
rect 5843 6598 5877 6600
rect 5809 6582 5889 6598
rect 5809 6576 5828 6582
rect 5525 6550 5628 6560
rect 5479 6548 5628 6550
rect 5649 6548 5684 6560
rect 5318 6546 5480 6548
rect 5330 6526 5349 6546
rect 5364 6544 5394 6546
rect 5213 6518 5254 6526
rect 5336 6522 5349 6526
rect 5401 6530 5480 6546
rect 5512 6546 5684 6548
rect 5512 6530 5591 6546
rect 5598 6544 5628 6546
rect 5176 6508 5205 6518
rect 5219 6508 5248 6518
rect 5263 6508 5293 6522
rect 5336 6508 5379 6522
rect 5401 6518 5591 6530
rect 5656 6526 5662 6546
rect 5386 6508 5416 6518
rect 5417 6508 5575 6518
rect 5579 6508 5609 6518
rect 5613 6508 5643 6522
rect 5671 6508 5684 6546
rect 5756 6560 5785 6576
rect 5799 6560 5828 6576
rect 5843 6566 5873 6582
rect 5901 6560 5907 6608
rect 5910 6602 5929 6608
rect 5944 6602 5974 6610
rect 5910 6594 5974 6602
rect 5910 6578 5990 6594
rect 6006 6587 6068 6618
rect 6084 6587 6146 6618
rect 6215 6616 6264 6641
rect 6279 6616 6309 6632
rect 6178 6602 6208 6610
rect 6215 6608 6325 6616
rect 6178 6594 6223 6602
rect 5910 6576 5929 6578
rect 5944 6576 5990 6578
rect 5910 6560 5990 6576
rect 6017 6574 6052 6587
rect 6093 6584 6130 6587
rect 6093 6582 6135 6584
rect 6022 6571 6052 6574
rect 6031 6567 6038 6571
rect 6038 6566 6039 6567
rect 5997 6560 6007 6566
rect 5756 6552 5791 6560
rect 5756 6526 5757 6552
rect 5764 6526 5791 6552
rect 5699 6508 5729 6522
rect 5756 6518 5791 6526
rect 5793 6552 5834 6560
rect 5793 6526 5808 6552
rect 5815 6526 5834 6552
rect 5898 6548 5929 6560
rect 5944 6548 6047 6560
rect 6059 6550 6085 6576
rect 6100 6571 6130 6582
rect 6162 6578 6224 6594
rect 6162 6576 6208 6578
rect 6162 6560 6224 6576
rect 6236 6560 6242 6608
rect 6245 6600 6325 6608
rect 6245 6598 6264 6600
rect 6279 6598 6313 6600
rect 6245 6582 6325 6598
rect 6245 6560 6264 6582
rect 6279 6566 6309 6582
rect 6337 6576 6343 6650
rect 6346 6576 6365 6720
rect 6380 6576 6386 6720
rect 6395 6650 6408 6720
rect 6460 6716 6482 6720
rect 6453 6694 6482 6708
rect 6535 6694 6551 6708
rect 6589 6704 6595 6706
rect 6602 6704 6710 6720
rect 6717 6704 6723 6706
rect 6731 6704 6746 6720
rect 6812 6714 6831 6717
rect 6453 6692 6551 6694
rect 6578 6692 6746 6704
rect 6761 6694 6777 6708
rect 6812 6695 6834 6714
rect 6844 6708 6860 6709
rect 6843 6706 6860 6708
rect 6844 6701 6860 6706
rect 6834 6694 6840 6695
rect 6843 6694 6872 6701
rect 6761 6693 6872 6694
rect 6761 6692 6878 6693
rect 6437 6684 6488 6692
rect 6535 6684 6569 6692
rect 6437 6672 6462 6684
rect 6469 6672 6488 6684
rect 6542 6682 6569 6684
rect 6578 6682 6799 6692
rect 6834 6689 6840 6692
rect 6542 6678 6799 6682
rect 6437 6664 6488 6672
rect 6535 6664 6799 6678
rect 6843 6684 6878 6692
rect 6389 6616 6408 6650
rect 6453 6656 6482 6664
rect 6453 6650 6470 6656
rect 6453 6648 6487 6650
rect 6535 6648 6551 6664
rect 6552 6654 6760 6664
rect 6761 6654 6777 6664
rect 6825 6660 6840 6675
rect 6843 6672 6844 6684
rect 6851 6672 6878 6684
rect 6843 6664 6878 6672
rect 6843 6663 6872 6664
rect 6563 6650 6777 6654
rect 6578 6648 6777 6650
rect 6812 6650 6825 6660
rect 6843 6650 6860 6663
rect 6812 6648 6860 6650
rect 6454 6644 6487 6648
rect 6450 6642 6487 6644
rect 6450 6641 6517 6642
rect 6450 6636 6481 6641
rect 6487 6636 6517 6641
rect 6450 6632 6517 6636
rect 6423 6629 6517 6632
rect 6423 6622 6472 6629
rect 6423 6616 6453 6622
rect 6472 6617 6477 6622
rect 6389 6600 6469 6616
rect 6481 6608 6517 6629
rect 6578 6624 6767 6648
rect 6812 6647 6859 6648
rect 6825 6642 6859 6647
rect 6593 6621 6767 6624
rect 6586 6618 6767 6621
rect 6795 6641 6859 6642
rect 6389 6598 6408 6600
rect 6423 6598 6457 6600
rect 6389 6582 6469 6598
rect 6389 6576 6408 6582
rect 6105 6550 6208 6560
rect 6059 6548 6208 6550
rect 6229 6548 6264 6560
rect 5898 6546 6060 6548
rect 5910 6526 5929 6546
rect 5944 6544 5974 6546
rect 5793 6518 5834 6526
rect 5916 6522 5929 6526
rect 5981 6530 6060 6546
rect 6092 6546 6264 6548
rect 6092 6530 6171 6546
rect 6178 6544 6208 6546
rect 5756 6508 5785 6518
rect 5799 6508 5828 6518
rect 5843 6508 5873 6522
rect 5916 6508 5959 6522
rect 5981 6518 6171 6530
rect 6236 6526 6242 6546
rect 5966 6508 5996 6518
rect 5997 6508 6155 6518
rect 6159 6508 6189 6518
rect 6193 6508 6223 6522
rect 6251 6508 6264 6546
rect 6336 6560 6365 6576
rect 6379 6560 6408 6576
rect 6423 6566 6453 6582
rect 6481 6560 6487 6608
rect 6490 6602 6509 6608
rect 6524 6602 6554 6610
rect 6490 6594 6554 6602
rect 6490 6578 6570 6594
rect 6586 6587 6648 6618
rect 6664 6587 6726 6618
rect 6795 6616 6844 6641
rect 6859 6616 6889 6632
rect 6758 6602 6788 6610
rect 6795 6608 6905 6616
rect 6758 6594 6803 6602
rect 6490 6576 6509 6578
rect 6524 6576 6570 6578
rect 6490 6560 6570 6576
rect 6597 6574 6632 6587
rect 6673 6584 6710 6587
rect 6673 6582 6715 6584
rect 6602 6571 6632 6574
rect 6611 6567 6618 6571
rect 6618 6566 6619 6567
rect 6577 6560 6587 6566
rect 6336 6552 6371 6560
rect 6336 6526 6337 6552
rect 6344 6526 6371 6552
rect 6279 6508 6309 6522
rect 6336 6518 6371 6526
rect 6373 6552 6414 6560
rect 6373 6526 6388 6552
rect 6395 6526 6414 6552
rect 6478 6548 6509 6560
rect 6524 6548 6627 6560
rect 6639 6550 6665 6576
rect 6680 6571 6710 6582
rect 6742 6578 6804 6594
rect 6742 6576 6788 6578
rect 6742 6560 6804 6576
rect 6816 6560 6822 6608
rect 6825 6600 6905 6608
rect 6825 6598 6844 6600
rect 6859 6598 6893 6600
rect 6825 6582 6905 6598
rect 6825 6560 6844 6582
rect 6859 6566 6889 6582
rect 6917 6576 6923 6650
rect 6926 6576 6945 6720
rect 6960 6576 6966 6720
rect 6975 6650 6988 6720
rect 7040 6716 7062 6720
rect 7033 6694 7062 6708
rect 7115 6694 7131 6708
rect 7169 6704 7175 6706
rect 7182 6704 7290 6720
rect 7297 6704 7303 6706
rect 7311 6704 7326 6720
rect 7392 6714 7411 6717
rect 7033 6692 7131 6694
rect 7158 6692 7326 6704
rect 7341 6694 7357 6708
rect 7392 6695 7414 6714
rect 7424 6708 7440 6709
rect 7423 6706 7440 6708
rect 7424 6701 7440 6706
rect 7414 6694 7420 6695
rect 7423 6694 7452 6701
rect 7341 6693 7452 6694
rect 7341 6692 7458 6693
rect 7017 6684 7068 6692
rect 7115 6684 7149 6692
rect 7017 6672 7042 6684
rect 7049 6672 7068 6684
rect 7122 6682 7149 6684
rect 7158 6682 7379 6692
rect 7414 6689 7420 6692
rect 7122 6678 7379 6682
rect 7017 6664 7068 6672
rect 7115 6664 7379 6678
rect 7423 6684 7458 6692
rect 6969 6616 6988 6650
rect 7033 6656 7062 6664
rect 7033 6650 7050 6656
rect 7033 6648 7067 6650
rect 7115 6648 7131 6664
rect 7132 6654 7340 6664
rect 7341 6654 7357 6664
rect 7405 6660 7420 6675
rect 7423 6672 7424 6684
rect 7431 6672 7458 6684
rect 7423 6664 7458 6672
rect 7423 6663 7452 6664
rect 7143 6650 7357 6654
rect 7158 6648 7357 6650
rect 7392 6650 7405 6660
rect 7423 6650 7440 6663
rect 7392 6648 7440 6650
rect 7034 6644 7067 6648
rect 7030 6642 7067 6644
rect 7030 6641 7097 6642
rect 7030 6636 7061 6641
rect 7067 6636 7097 6641
rect 7030 6632 7097 6636
rect 7003 6629 7097 6632
rect 7003 6622 7052 6629
rect 7003 6616 7033 6622
rect 7052 6617 7057 6622
rect 6969 6600 7049 6616
rect 7061 6608 7097 6629
rect 7158 6624 7347 6648
rect 7392 6647 7439 6648
rect 7405 6642 7439 6647
rect 7173 6621 7347 6624
rect 7166 6618 7347 6621
rect 7375 6641 7439 6642
rect 6969 6598 6988 6600
rect 7003 6598 7037 6600
rect 6969 6582 7049 6598
rect 6969 6576 6988 6582
rect 6685 6550 6788 6560
rect 6639 6548 6788 6550
rect 6809 6548 6844 6560
rect 6478 6546 6640 6548
rect 6490 6526 6509 6546
rect 6524 6544 6554 6546
rect 6373 6518 6414 6526
rect 6496 6522 6509 6526
rect 6561 6530 6640 6546
rect 6672 6546 6844 6548
rect 6672 6530 6751 6546
rect 6758 6544 6788 6546
rect 6336 6508 6365 6518
rect 6379 6508 6408 6518
rect 6423 6508 6453 6522
rect 6496 6508 6539 6522
rect 6561 6518 6751 6530
rect 6816 6526 6822 6546
rect 6546 6508 6576 6518
rect 6577 6508 6735 6518
rect 6739 6508 6769 6518
rect 6773 6508 6803 6522
rect 6831 6508 6844 6546
rect 6916 6560 6945 6576
rect 6959 6560 6988 6576
rect 7003 6566 7033 6582
rect 7061 6560 7067 6608
rect 7070 6602 7089 6608
rect 7104 6602 7134 6610
rect 7070 6594 7134 6602
rect 7070 6578 7150 6594
rect 7166 6587 7228 6618
rect 7244 6587 7306 6618
rect 7375 6616 7424 6641
rect 7439 6616 7469 6632
rect 7338 6602 7368 6610
rect 7375 6608 7485 6616
rect 7338 6594 7383 6602
rect 7070 6576 7089 6578
rect 7104 6576 7150 6578
rect 7070 6560 7150 6576
rect 7177 6574 7212 6587
rect 7253 6584 7290 6587
rect 7253 6582 7295 6584
rect 7182 6571 7212 6574
rect 7191 6567 7198 6571
rect 7198 6566 7199 6567
rect 7157 6560 7167 6566
rect 6916 6552 6951 6560
rect 6916 6526 6917 6552
rect 6924 6526 6951 6552
rect 6859 6508 6889 6522
rect 6916 6518 6951 6526
rect 6953 6552 6994 6560
rect 6953 6526 6968 6552
rect 6975 6526 6994 6552
rect 7058 6548 7089 6560
rect 7104 6548 7207 6560
rect 7219 6550 7245 6576
rect 7260 6571 7290 6582
rect 7322 6578 7384 6594
rect 7322 6576 7368 6578
rect 7322 6560 7384 6576
rect 7396 6560 7402 6608
rect 7405 6600 7485 6608
rect 7405 6598 7424 6600
rect 7439 6598 7473 6600
rect 7405 6582 7485 6598
rect 7405 6560 7424 6582
rect 7439 6566 7469 6582
rect 7497 6576 7503 6650
rect 7506 6576 7525 6720
rect 7540 6576 7546 6720
rect 7555 6650 7568 6720
rect 7620 6716 7642 6720
rect 7613 6694 7642 6708
rect 7695 6694 7711 6708
rect 7749 6704 7755 6706
rect 7762 6704 7870 6720
rect 7877 6704 7883 6706
rect 7891 6704 7906 6720
rect 7972 6714 7991 6717
rect 7613 6692 7711 6694
rect 7738 6692 7906 6704
rect 7921 6694 7937 6708
rect 7972 6695 7994 6714
rect 8004 6708 8020 6709
rect 8003 6706 8020 6708
rect 8004 6701 8020 6706
rect 7994 6694 8000 6695
rect 8003 6694 8032 6701
rect 7921 6693 8032 6694
rect 7921 6692 8038 6693
rect 7597 6684 7648 6692
rect 7695 6684 7729 6692
rect 7597 6672 7622 6684
rect 7629 6672 7648 6684
rect 7702 6682 7729 6684
rect 7738 6682 7959 6692
rect 7994 6689 8000 6692
rect 7702 6678 7959 6682
rect 7597 6664 7648 6672
rect 7695 6664 7959 6678
rect 8003 6684 8038 6692
rect 7549 6616 7568 6650
rect 7613 6656 7642 6664
rect 7613 6650 7630 6656
rect 7613 6648 7647 6650
rect 7695 6648 7711 6664
rect 7712 6654 7920 6664
rect 7921 6654 7937 6664
rect 7985 6660 8000 6675
rect 8003 6672 8004 6684
rect 8011 6672 8038 6684
rect 8003 6664 8038 6672
rect 8003 6663 8032 6664
rect 7723 6650 7937 6654
rect 7738 6648 7937 6650
rect 7972 6650 7985 6660
rect 8003 6650 8020 6663
rect 7972 6648 8020 6650
rect 7614 6644 7647 6648
rect 7610 6642 7647 6644
rect 7610 6641 7677 6642
rect 7610 6636 7641 6641
rect 7647 6636 7677 6641
rect 7610 6632 7677 6636
rect 7583 6629 7677 6632
rect 7583 6622 7632 6629
rect 7583 6616 7613 6622
rect 7632 6617 7637 6622
rect 7549 6600 7629 6616
rect 7641 6608 7677 6629
rect 7738 6624 7927 6648
rect 7972 6647 8019 6648
rect 7985 6642 8019 6647
rect 7753 6621 7927 6624
rect 7746 6618 7927 6621
rect 7955 6641 8019 6642
rect 7549 6598 7568 6600
rect 7583 6598 7617 6600
rect 7549 6582 7629 6598
rect 7549 6576 7568 6582
rect 7265 6550 7368 6560
rect 7219 6548 7368 6550
rect 7389 6548 7424 6560
rect 7058 6546 7220 6548
rect 7070 6526 7089 6546
rect 7104 6544 7134 6546
rect 6953 6518 6994 6526
rect 7076 6522 7089 6526
rect 7141 6530 7220 6546
rect 7252 6546 7424 6548
rect 7252 6530 7331 6546
rect 7338 6544 7368 6546
rect 6916 6508 6945 6518
rect 6959 6508 6988 6518
rect 7003 6508 7033 6522
rect 7076 6508 7119 6522
rect 7141 6518 7331 6530
rect 7396 6526 7402 6546
rect 7126 6508 7156 6518
rect 7157 6508 7315 6518
rect 7319 6508 7349 6518
rect 7353 6508 7383 6522
rect 7411 6508 7424 6546
rect 7496 6560 7525 6576
rect 7539 6560 7568 6576
rect 7583 6566 7613 6582
rect 7641 6560 7647 6608
rect 7650 6602 7669 6608
rect 7684 6602 7714 6610
rect 7650 6594 7714 6602
rect 7650 6578 7730 6594
rect 7746 6587 7808 6618
rect 7824 6587 7886 6618
rect 7955 6616 8004 6641
rect 8019 6616 8049 6632
rect 7918 6602 7948 6610
rect 7955 6608 8065 6616
rect 7918 6594 7963 6602
rect 7650 6576 7669 6578
rect 7684 6576 7730 6578
rect 7650 6560 7730 6576
rect 7757 6574 7792 6587
rect 7833 6584 7870 6587
rect 7833 6582 7875 6584
rect 7762 6571 7792 6574
rect 7771 6567 7778 6571
rect 7778 6566 7779 6567
rect 7737 6560 7747 6566
rect 7496 6552 7531 6560
rect 7496 6526 7497 6552
rect 7504 6526 7531 6552
rect 7439 6508 7469 6522
rect 7496 6518 7531 6526
rect 7533 6552 7574 6560
rect 7533 6526 7548 6552
rect 7555 6526 7574 6552
rect 7638 6548 7669 6560
rect 7684 6548 7787 6560
rect 7799 6550 7825 6576
rect 7840 6571 7870 6582
rect 7902 6578 7964 6594
rect 7902 6576 7948 6578
rect 7902 6560 7964 6576
rect 7976 6560 7982 6608
rect 7985 6600 8065 6608
rect 7985 6598 8004 6600
rect 8019 6598 8053 6600
rect 7985 6582 8065 6598
rect 7985 6560 8004 6582
rect 8019 6566 8049 6582
rect 8077 6576 8083 6650
rect 8086 6576 8105 6720
rect 8120 6576 8126 6720
rect 8135 6650 8148 6720
rect 8200 6716 8222 6720
rect 8193 6694 8222 6708
rect 8275 6694 8291 6708
rect 8329 6704 8335 6706
rect 8342 6704 8450 6720
rect 8457 6704 8463 6706
rect 8471 6704 8486 6720
rect 8552 6714 8571 6717
rect 8193 6692 8291 6694
rect 8318 6692 8486 6704
rect 8501 6694 8517 6708
rect 8552 6695 8574 6714
rect 8584 6708 8600 6709
rect 8583 6706 8600 6708
rect 8584 6701 8600 6706
rect 8574 6694 8580 6695
rect 8583 6694 8612 6701
rect 8501 6693 8612 6694
rect 8501 6692 8618 6693
rect 8177 6684 8228 6692
rect 8275 6684 8309 6692
rect 8177 6672 8202 6684
rect 8209 6672 8228 6684
rect 8282 6682 8309 6684
rect 8318 6682 8539 6692
rect 8574 6689 8580 6692
rect 8282 6678 8539 6682
rect 8177 6664 8228 6672
rect 8275 6664 8539 6678
rect 8583 6684 8618 6692
rect 8129 6616 8148 6650
rect 8193 6656 8222 6664
rect 8193 6650 8210 6656
rect 8193 6648 8227 6650
rect 8275 6648 8291 6664
rect 8292 6654 8500 6664
rect 8501 6654 8517 6664
rect 8565 6660 8580 6675
rect 8583 6672 8584 6684
rect 8591 6672 8618 6684
rect 8583 6664 8618 6672
rect 8583 6663 8612 6664
rect 8303 6650 8517 6654
rect 8318 6648 8517 6650
rect 8552 6650 8565 6660
rect 8583 6650 8600 6663
rect 8552 6648 8600 6650
rect 8194 6644 8227 6648
rect 8190 6642 8227 6644
rect 8190 6641 8257 6642
rect 8190 6636 8221 6641
rect 8227 6636 8257 6641
rect 8190 6632 8257 6636
rect 8163 6629 8257 6632
rect 8163 6622 8212 6629
rect 8163 6616 8193 6622
rect 8212 6617 8217 6622
rect 8129 6600 8209 6616
rect 8221 6608 8257 6629
rect 8318 6624 8507 6648
rect 8552 6647 8599 6648
rect 8565 6642 8599 6647
rect 8333 6621 8507 6624
rect 8326 6618 8507 6621
rect 8535 6641 8599 6642
rect 8129 6598 8148 6600
rect 8163 6598 8197 6600
rect 8129 6582 8209 6598
rect 8129 6576 8148 6582
rect 7845 6550 7948 6560
rect 7799 6548 7948 6550
rect 7969 6548 8004 6560
rect 7638 6546 7800 6548
rect 7650 6526 7669 6546
rect 7684 6544 7714 6546
rect 7533 6518 7574 6526
rect 7656 6522 7669 6526
rect 7721 6530 7800 6546
rect 7832 6546 8004 6548
rect 7832 6530 7911 6546
rect 7918 6544 7948 6546
rect 7496 6508 7525 6518
rect 7539 6508 7568 6518
rect 7583 6508 7613 6522
rect 7656 6508 7699 6522
rect 7721 6518 7911 6530
rect 7976 6526 7982 6546
rect 7706 6508 7736 6518
rect 7737 6508 7895 6518
rect 7899 6508 7929 6518
rect 7933 6508 7963 6522
rect 7991 6508 8004 6546
rect 8076 6560 8105 6576
rect 8119 6560 8148 6576
rect 8163 6566 8193 6582
rect 8221 6560 8227 6608
rect 8230 6602 8249 6608
rect 8264 6602 8294 6610
rect 8230 6594 8294 6602
rect 8230 6578 8310 6594
rect 8326 6587 8388 6618
rect 8404 6587 8466 6618
rect 8535 6616 8584 6641
rect 8599 6616 8629 6632
rect 8498 6602 8528 6610
rect 8535 6608 8645 6616
rect 8498 6594 8543 6602
rect 8230 6576 8249 6578
rect 8264 6576 8310 6578
rect 8230 6560 8310 6576
rect 8337 6574 8372 6587
rect 8413 6584 8450 6587
rect 8413 6582 8455 6584
rect 8342 6571 8372 6574
rect 8351 6567 8358 6571
rect 8358 6566 8359 6567
rect 8317 6560 8327 6566
rect 8076 6552 8111 6560
rect 8076 6526 8077 6552
rect 8084 6526 8111 6552
rect 8019 6508 8049 6522
rect 8076 6518 8111 6526
rect 8113 6552 8154 6560
rect 8113 6526 8128 6552
rect 8135 6526 8154 6552
rect 8218 6548 8249 6560
rect 8264 6548 8367 6560
rect 8379 6550 8405 6576
rect 8420 6571 8450 6582
rect 8482 6578 8544 6594
rect 8482 6576 8528 6578
rect 8482 6560 8544 6576
rect 8556 6560 8562 6608
rect 8565 6600 8645 6608
rect 8565 6598 8584 6600
rect 8599 6598 8633 6600
rect 8565 6582 8645 6598
rect 8565 6560 8584 6582
rect 8599 6566 8629 6582
rect 8657 6576 8663 6650
rect 8666 6576 8685 6720
rect 8700 6576 8706 6720
rect 8715 6650 8728 6720
rect 8780 6716 8802 6720
rect 8773 6694 8802 6708
rect 8855 6694 8871 6708
rect 8909 6704 8915 6706
rect 8922 6704 9030 6720
rect 9037 6704 9043 6706
rect 9051 6704 9066 6720
rect 9132 6714 9151 6717
rect 8773 6692 8871 6694
rect 8898 6692 9066 6704
rect 9081 6694 9097 6708
rect 9132 6695 9154 6714
rect 9164 6708 9180 6709
rect 9163 6706 9180 6708
rect 9164 6701 9180 6706
rect 9154 6694 9160 6695
rect 9163 6694 9192 6701
rect 9081 6693 9192 6694
rect 9081 6692 9198 6693
rect 8757 6684 8808 6692
rect 8855 6684 8889 6692
rect 8757 6672 8782 6684
rect 8789 6672 8808 6684
rect 8862 6682 8889 6684
rect 8898 6682 9119 6692
rect 9154 6689 9160 6692
rect 8862 6678 9119 6682
rect 8757 6664 8808 6672
rect 8855 6664 9119 6678
rect 9163 6684 9198 6692
rect 8709 6616 8728 6650
rect 8773 6656 8802 6664
rect 8773 6650 8790 6656
rect 8773 6648 8807 6650
rect 8855 6648 8871 6664
rect 8872 6654 9080 6664
rect 9081 6654 9097 6664
rect 9145 6660 9160 6675
rect 9163 6672 9164 6684
rect 9171 6672 9198 6684
rect 9163 6664 9198 6672
rect 9163 6663 9192 6664
rect 8883 6650 9097 6654
rect 8898 6648 9097 6650
rect 9132 6650 9145 6660
rect 9163 6650 9180 6663
rect 9132 6648 9180 6650
rect 8774 6644 8807 6648
rect 8770 6642 8807 6644
rect 8770 6641 8837 6642
rect 8770 6636 8801 6641
rect 8807 6636 8837 6641
rect 8770 6632 8837 6636
rect 8743 6629 8837 6632
rect 8743 6622 8792 6629
rect 8743 6616 8773 6622
rect 8792 6617 8797 6622
rect 8709 6600 8789 6616
rect 8801 6608 8837 6629
rect 8898 6624 9087 6648
rect 9132 6647 9179 6648
rect 9145 6642 9179 6647
rect 8913 6621 9087 6624
rect 8906 6618 9087 6621
rect 9115 6641 9179 6642
rect 8709 6598 8728 6600
rect 8743 6598 8777 6600
rect 8709 6582 8789 6598
rect 8709 6576 8728 6582
rect 8425 6550 8528 6560
rect 8379 6548 8528 6550
rect 8549 6548 8584 6560
rect 8218 6546 8380 6548
rect 8230 6526 8249 6546
rect 8264 6544 8294 6546
rect 8113 6518 8154 6526
rect 8236 6522 8249 6526
rect 8301 6530 8380 6546
rect 8412 6546 8584 6548
rect 8412 6530 8491 6546
rect 8498 6544 8528 6546
rect 8076 6508 8105 6518
rect 8119 6508 8148 6518
rect 8163 6508 8193 6522
rect 8236 6508 8279 6522
rect 8301 6518 8491 6530
rect 8556 6526 8562 6546
rect 8286 6508 8316 6518
rect 8317 6508 8475 6518
rect 8479 6508 8509 6518
rect 8513 6508 8543 6522
rect 8571 6508 8584 6546
rect 8656 6560 8685 6576
rect 8699 6560 8728 6576
rect 8743 6566 8773 6582
rect 8801 6560 8807 6608
rect 8810 6602 8829 6608
rect 8844 6602 8874 6610
rect 8810 6594 8874 6602
rect 8810 6578 8890 6594
rect 8906 6587 8968 6618
rect 8984 6587 9046 6618
rect 9115 6616 9164 6641
rect 9179 6616 9209 6632
rect 9078 6602 9108 6610
rect 9115 6608 9225 6616
rect 9078 6594 9123 6602
rect 8810 6576 8829 6578
rect 8844 6576 8890 6578
rect 8810 6560 8890 6576
rect 8917 6574 8952 6587
rect 8993 6584 9030 6587
rect 8993 6582 9035 6584
rect 8922 6571 8952 6574
rect 8931 6567 8938 6571
rect 8938 6566 8939 6567
rect 8897 6560 8907 6566
rect 8656 6552 8691 6560
rect 8656 6526 8657 6552
rect 8664 6526 8691 6552
rect 8599 6508 8629 6522
rect 8656 6518 8691 6526
rect 8693 6552 8734 6560
rect 8693 6526 8708 6552
rect 8715 6526 8734 6552
rect 8798 6548 8829 6560
rect 8844 6548 8947 6560
rect 8959 6550 8985 6576
rect 9000 6571 9030 6582
rect 9062 6578 9124 6594
rect 9062 6576 9108 6578
rect 9062 6560 9124 6576
rect 9136 6560 9142 6608
rect 9145 6600 9225 6608
rect 9145 6598 9164 6600
rect 9179 6598 9213 6600
rect 9145 6582 9225 6598
rect 9145 6560 9164 6582
rect 9179 6566 9209 6582
rect 9237 6576 9243 6650
rect 9246 6576 9265 6720
rect 9280 6576 9286 6720
rect 9295 6650 9308 6720
rect 9360 6716 9382 6720
rect 9353 6694 9382 6708
rect 9435 6694 9451 6708
rect 9489 6704 9495 6706
rect 9502 6704 9610 6720
rect 9617 6704 9623 6706
rect 9631 6704 9646 6720
rect 9712 6714 9731 6717
rect 9353 6692 9451 6694
rect 9478 6692 9646 6704
rect 9661 6694 9677 6708
rect 9712 6695 9734 6714
rect 9744 6708 9760 6709
rect 9743 6706 9760 6708
rect 9744 6701 9760 6706
rect 9734 6694 9740 6695
rect 9743 6694 9772 6701
rect 9661 6693 9772 6694
rect 9661 6692 9778 6693
rect 9337 6684 9388 6692
rect 9435 6684 9469 6692
rect 9337 6672 9362 6684
rect 9369 6672 9388 6684
rect 9442 6682 9469 6684
rect 9478 6682 9699 6692
rect 9734 6689 9740 6692
rect 9442 6678 9699 6682
rect 9337 6664 9388 6672
rect 9435 6664 9699 6678
rect 9743 6684 9778 6692
rect 9289 6616 9308 6650
rect 9353 6656 9382 6664
rect 9353 6650 9370 6656
rect 9353 6648 9387 6650
rect 9435 6648 9451 6664
rect 9452 6654 9660 6664
rect 9661 6654 9677 6664
rect 9725 6660 9740 6675
rect 9743 6672 9744 6684
rect 9751 6672 9778 6684
rect 9743 6664 9778 6672
rect 9743 6663 9772 6664
rect 9463 6650 9677 6654
rect 9478 6648 9677 6650
rect 9712 6650 9725 6660
rect 9743 6650 9760 6663
rect 9712 6648 9760 6650
rect 9354 6644 9387 6648
rect 9350 6642 9387 6644
rect 9350 6641 9417 6642
rect 9350 6636 9381 6641
rect 9387 6636 9417 6641
rect 9350 6632 9417 6636
rect 9323 6629 9417 6632
rect 9323 6622 9372 6629
rect 9323 6616 9353 6622
rect 9372 6617 9377 6622
rect 9289 6600 9369 6616
rect 9381 6608 9417 6629
rect 9478 6624 9667 6648
rect 9712 6647 9759 6648
rect 9725 6642 9759 6647
rect 9493 6621 9667 6624
rect 9486 6618 9667 6621
rect 9695 6641 9759 6642
rect 9289 6598 9308 6600
rect 9323 6598 9357 6600
rect 9289 6582 9369 6598
rect 9289 6576 9308 6582
rect 9005 6550 9108 6560
rect 8959 6548 9108 6550
rect 9129 6548 9164 6560
rect 8798 6546 8960 6548
rect 8810 6526 8829 6546
rect 8844 6544 8874 6546
rect 8693 6518 8734 6526
rect 8816 6522 8829 6526
rect 8881 6530 8960 6546
rect 8992 6546 9164 6548
rect 8992 6530 9071 6546
rect 9078 6544 9108 6546
rect 8656 6508 8685 6518
rect 8699 6508 8728 6518
rect 8743 6508 8773 6522
rect 8816 6508 8859 6522
rect 8881 6518 9071 6530
rect 9136 6526 9142 6546
rect 8866 6508 8896 6518
rect 8897 6508 9055 6518
rect 9059 6508 9089 6518
rect 9093 6508 9123 6522
rect 9151 6508 9164 6546
rect 9236 6560 9265 6576
rect 9279 6560 9308 6576
rect 9323 6566 9353 6582
rect 9381 6560 9387 6608
rect 9390 6602 9409 6608
rect 9424 6602 9454 6610
rect 9390 6594 9454 6602
rect 9390 6578 9470 6594
rect 9486 6587 9548 6618
rect 9564 6587 9626 6618
rect 9695 6616 9744 6641
rect 9759 6616 9789 6632
rect 9658 6602 9688 6610
rect 9695 6608 9805 6616
rect 9658 6594 9703 6602
rect 9390 6576 9409 6578
rect 9424 6576 9470 6578
rect 9390 6560 9470 6576
rect 9497 6574 9532 6587
rect 9573 6584 9610 6587
rect 9573 6582 9615 6584
rect 9502 6571 9532 6574
rect 9511 6567 9518 6571
rect 9518 6566 9519 6567
rect 9477 6560 9487 6566
rect 9236 6552 9271 6560
rect 9236 6526 9237 6552
rect 9244 6526 9271 6552
rect 9179 6508 9209 6522
rect 9236 6518 9271 6526
rect 9273 6552 9314 6560
rect 9273 6526 9288 6552
rect 9295 6526 9314 6552
rect 9378 6548 9409 6560
rect 9424 6548 9527 6560
rect 9539 6550 9565 6576
rect 9580 6571 9610 6582
rect 9642 6578 9704 6594
rect 9642 6576 9688 6578
rect 9642 6560 9704 6576
rect 9716 6560 9722 6608
rect 9725 6600 9805 6608
rect 9725 6598 9744 6600
rect 9759 6598 9793 6600
rect 9725 6582 9805 6598
rect 9725 6560 9744 6582
rect 9759 6566 9789 6582
rect 9817 6576 9823 6650
rect 9826 6576 9845 6720
rect 9860 6576 9866 6720
rect 9875 6650 9888 6720
rect 9940 6716 9962 6720
rect 9933 6694 9962 6708
rect 10015 6694 10031 6708
rect 10069 6704 10075 6706
rect 10082 6704 10190 6720
rect 10197 6704 10203 6706
rect 10211 6704 10226 6720
rect 10292 6714 10311 6717
rect 9933 6692 10031 6694
rect 10058 6692 10226 6704
rect 10241 6694 10257 6708
rect 10292 6695 10314 6714
rect 10324 6708 10340 6709
rect 10323 6706 10340 6708
rect 10324 6701 10340 6706
rect 10314 6694 10320 6695
rect 10323 6694 10352 6701
rect 10241 6693 10352 6694
rect 10241 6692 10358 6693
rect 9917 6684 9968 6692
rect 10015 6684 10049 6692
rect 9917 6672 9942 6684
rect 9949 6672 9968 6684
rect 10022 6682 10049 6684
rect 10058 6682 10279 6692
rect 10314 6689 10320 6692
rect 10022 6678 10279 6682
rect 9917 6664 9968 6672
rect 10015 6664 10279 6678
rect 10323 6684 10358 6692
rect 9869 6616 9888 6650
rect 9933 6656 9962 6664
rect 9933 6650 9950 6656
rect 9933 6648 9967 6650
rect 10015 6648 10031 6664
rect 10032 6654 10240 6664
rect 10241 6654 10257 6664
rect 10305 6660 10320 6675
rect 10323 6672 10324 6684
rect 10331 6672 10358 6684
rect 10323 6664 10358 6672
rect 10323 6663 10352 6664
rect 10043 6650 10257 6654
rect 10058 6648 10257 6650
rect 10292 6650 10305 6660
rect 10323 6650 10340 6663
rect 10292 6648 10340 6650
rect 9934 6644 9967 6648
rect 9930 6642 9967 6644
rect 9930 6641 9997 6642
rect 9930 6636 9961 6641
rect 9967 6636 9997 6641
rect 9930 6632 9997 6636
rect 9903 6629 9997 6632
rect 9903 6622 9952 6629
rect 9903 6616 9933 6622
rect 9952 6617 9957 6622
rect 9869 6600 9949 6616
rect 9961 6608 9997 6629
rect 10058 6624 10247 6648
rect 10292 6647 10339 6648
rect 10305 6642 10339 6647
rect 10073 6621 10247 6624
rect 10066 6618 10247 6621
rect 10275 6641 10339 6642
rect 9869 6598 9888 6600
rect 9903 6598 9937 6600
rect 9869 6582 9949 6598
rect 9869 6576 9888 6582
rect 9585 6550 9688 6560
rect 9539 6548 9688 6550
rect 9709 6548 9744 6560
rect 9378 6546 9540 6548
rect 9390 6526 9409 6546
rect 9424 6544 9454 6546
rect 9273 6518 9314 6526
rect 9396 6522 9409 6526
rect 9461 6530 9540 6546
rect 9572 6546 9744 6548
rect 9572 6530 9651 6546
rect 9658 6544 9688 6546
rect 9236 6508 9265 6518
rect 9279 6508 9308 6518
rect 9323 6508 9353 6522
rect 9396 6508 9439 6522
rect 9461 6518 9651 6530
rect 9716 6526 9722 6546
rect 9446 6508 9476 6518
rect 9477 6508 9635 6518
rect 9639 6508 9669 6518
rect 9673 6508 9703 6522
rect 9731 6508 9744 6546
rect 9816 6560 9845 6576
rect 9859 6560 9888 6576
rect 9903 6566 9933 6582
rect 9961 6560 9967 6608
rect 9970 6602 9989 6608
rect 10004 6602 10034 6610
rect 9970 6594 10034 6602
rect 9970 6578 10050 6594
rect 10066 6587 10128 6618
rect 10144 6587 10206 6618
rect 10275 6616 10324 6641
rect 10339 6616 10369 6632
rect 10238 6602 10268 6610
rect 10275 6608 10385 6616
rect 10238 6594 10283 6602
rect 9970 6576 9989 6578
rect 10004 6576 10050 6578
rect 9970 6560 10050 6576
rect 10077 6574 10112 6587
rect 10153 6584 10190 6587
rect 10153 6582 10195 6584
rect 10082 6571 10112 6574
rect 10091 6567 10098 6571
rect 10098 6566 10099 6567
rect 10057 6560 10067 6566
rect 9816 6552 9851 6560
rect 9816 6526 9817 6552
rect 9824 6526 9851 6552
rect 9759 6508 9789 6522
rect 9816 6518 9851 6526
rect 9853 6552 9894 6560
rect 9853 6526 9868 6552
rect 9875 6526 9894 6552
rect 9958 6548 9989 6560
rect 10004 6548 10107 6560
rect 10119 6550 10145 6576
rect 10160 6571 10190 6582
rect 10222 6578 10284 6594
rect 10222 6576 10268 6578
rect 10222 6560 10284 6576
rect 10296 6560 10302 6608
rect 10305 6600 10385 6608
rect 10305 6598 10324 6600
rect 10339 6598 10373 6600
rect 10305 6582 10385 6598
rect 10305 6560 10324 6582
rect 10339 6566 10369 6582
rect 10397 6576 10403 6650
rect 10406 6576 10425 6720
rect 10440 6576 10446 6720
rect 10455 6650 10468 6720
rect 10520 6716 10542 6720
rect 10513 6694 10542 6708
rect 10595 6694 10611 6708
rect 10649 6704 10655 6706
rect 10662 6704 10770 6720
rect 10777 6704 10783 6706
rect 10791 6704 10806 6720
rect 10872 6714 10891 6717
rect 10513 6692 10611 6694
rect 10638 6692 10806 6704
rect 10821 6694 10837 6708
rect 10872 6695 10894 6714
rect 10904 6708 10920 6709
rect 10903 6706 10920 6708
rect 10904 6701 10920 6706
rect 10894 6694 10900 6695
rect 10903 6694 10932 6701
rect 10821 6693 10932 6694
rect 10821 6692 10938 6693
rect 10497 6684 10548 6692
rect 10595 6684 10629 6692
rect 10497 6672 10522 6684
rect 10529 6672 10548 6684
rect 10602 6682 10629 6684
rect 10638 6682 10859 6692
rect 10894 6689 10900 6692
rect 10602 6678 10859 6682
rect 10497 6664 10548 6672
rect 10595 6664 10859 6678
rect 10903 6684 10938 6692
rect 10449 6616 10468 6650
rect 10513 6656 10542 6664
rect 10513 6650 10530 6656
rect 10513 6648 10547 6650
rect 10595 6648 10611 6664
rect 10612 6654 10820 6664
rect 10821 6654 10837 6664
rect 10885 6660 10900 6675
rect 10903 6672 10904 6684
rect 10911 6672 10938 6684
rect 10903 6664 10938 6672
rect 10903 6663 10932 6664
rect 10623 6650 10837 6654
rect 10638 6648 10837 6650
rect 10872 6650 10885 6660
rect 10903 6650 10920 6663
rect 10872 6648 10920 6650
rect 10514 6644 10547 6648
rect 10510 6642 10547 6644
rect 10510 6641 10577 6642
rect 10510 6636 10541 6641
rect 10547 6636 10577 6641
rect 10510 6632 10577 6636
rect 10483 6629 10577 6632
rect 10483 6622 10532 6629
rect 10483 6616 10513 6622
rect 10532 6617 10537 6622
rect 10449 6600 10529 6616
rect 10541 6608 10577 6629
rect 10638 6624 10827 6648
rect 10872 6647 10919 6648
rect 10885 6642 10919 6647
rect 10653 6621 10827 6624
rect 10646 6618 10827 6621
rect 10855 6641 10919 6642
rect 10449 6598 10468 6600
rect 10483 6598 10517 6600
rect 10449 6582 10529 6598
rect 10449 6576 10468 6582
rect 10165 6550 10268 6560
rect 10119 6548 10268 6550
rect 10289 6548 10324 6560
rect 9958 6546 10120 6548
rect 9970 6526 9989 6546
rect 10004 6544 10034 6546
rect 9853 6518 9894 6526
rect 9976 6522 9989 6526
rect 10041 6530 10120 6546
rect 10152 6546 10324 6548
rect 10152 6530 10231 6546
rect 10238 6544 10268 6546
rect 9816 6508 9845 6518
rect 9859 6508 9888 6518
rect 9903 6508 9933 6522
rect 9976 6508 10019 6522
rect 10041 6518 10231 6530
rect 10296 6526 10302 6546
rect 10026 6508 10056 6518
rect 10057 6508 10215 6518
rect 10219 6508 10249 6518
rect 10253 6508 10283 6522
rect 10311 6508 10324 6546
rect 10396 6560 10425 6576
rect 10439 6560 10468 6576
rect 10483 6566 10513 6582
rect 10541 6560 10547 6608
rect 10550 6602 10569 6608
rect 10584 6602 10614 6610
rect 10550 6594 10614 6602
rect 10550 6578 10630 6594
rect 10646 6587 10708 6618
rect 10724 6587 10786 6618
rect 10855 6616 10904 6641
rect 10919 6616 10949 6632
rect 10818 6602 10848 6610
rect 10855 6608 10965 6616
rect 10818 6594 10863 6602
rect 10550 6576 10569 6578
rect 10584 6576 10630 6578
rect 10550 6560 10630 6576
rect 10657 6574 10692 6587
rect 10733 6584 10770 6587
rect 10733 6582 10775 6584
rect 10662 6571 10692 6574
rect 10671 6567 10678 6571
rect 10678 6566 10679 6567
rect 10637 6560 10647 6566
rect 10396 6552 10431 6560
rect 10396 6526 10397 6552
rect 10404 6526 10431 6552
rect 10339 6508 10369 6522
rect 10396 6518 10431 6526
rect 10433 6552 10474 6560
rect 10433 6526 10448 6552
rect 10455 6526 10474 6552
rect 10538 6548 10569 6560
rect 10584 6548 10687 6560
rect 10699 6550 10725 6576
rect 10740 6571 10770 6582
rect 10802 6578 10864 6594
rect 10802 6576 10848 6578
rect 10802 6560 10864 6576
rect 10876 6560 10882 6608
rect 10885 6600 10965 6608
rect 10885 6598 10904 6600
rect 10919 6598 10953 6600
rect 10885 6582 10965 6598
rect 10885 6560 10904 6582
rect 10919 6566 10949 6582
rect 10977 6576 10983 6650
rect 10986 6576 11005 6720
rect 11020 6576 11026 6720
rect 11035 6650 11048 6720
rect 11100 6716 11122 6720
rect 11093 6694 11122 6708
rect 11175 6694 11191 6708
rect 11229 6704 11235 6706
rect 11242 6704 11350 6720
rect 11357 6704 11363 6706
rect 11371 6704 11386 6720
rect 11452 6714 11471 6717
rect 11093 6692 11191 6694
rect 11218 6692 11386 6704
rect 11401 6694 11417 6708
rect 11452 6695 11474 6714
rect 11484 6708 11500 6709
rect 11483 6706 11500 6708
rect 11484 6701 11500 6706
rect 11474 6694 11480 6695
rect 11483 6694 11512 6701
rect 11401 6693 11512 6694
rect 11401 6692 11518 6693
rect 11077 6684 11128 6692
rect 11175 6684 11209 6692
rect 11077 6672 11102 6684
rect 11109 6672 11128 6684
rect 11182 6682 11209 6684
rect 11218 6682 11439 6692
rect 11474 6689 11480 6692
rect 11182 6678 11439 6682
rect 11077 6664 11128 6672
rect 11175 6664 11439 6678
rect 11483 6684 11518 6692
rect 11029 6616 11048 6650
rect 11093 6656 11122 6664
rect 11093 6650 11110 6656
rect 11093 6648 11127 6650
rect 11175 6648 11191 6664
rect 11192 6654 11400 6664
rect 11401 6654 11417 6664
rect 11465 6660 11480 6675
rect 11483 6672 11484 6684
rect 11491 6672 11518 6684
rect 11483 6664 11518 6672
rect 11483 6663 11512 6664
rect 11203 6650 11417 6654
rect 11218 6648 11417 6650
rect 11452 6650 11465 6660
rect 11483 6650 11500 6663
rect 11452 6648 11500 6650
rect 11094 6644 11127 6648
rect 11090 6642 11127 6644
rect 11090 6641 11157 6642
rect 11090 6636 11121 6641
rect 11127 6636 11157 6641
rect 11090 6632 11157 6636
rect 11063 6629 11157 6632
rect 11063 6622 11112 6629
rect 11063 6616 11093 6622
rect 11112 6617 11117 6622
rect 11029 6600 11109 6616
rect 11121 6608 11157 6629
rect 11218 6624 11407 6648
rect 11452 6647 11499 6648
rect 11465 6642 11499 6647
rect 11233 6621 11407 6624
rect 11226 6618 11407 6621
rect 11435 6641 11499 6642
rect 11029 6598 11048 6600
rect 11063 6598 11097 6600
rect 11029 6582 11109 6598
rect 11029 6576 11048 6582
rect 10745 6550 10848 6560
rect 10699 6548 10848 6550
rect 10869 6548 10904 6560
rect 10538 6546 10700 6548
rect 10550 6526 10569 6546
rect 10584 6544 10614 6546
rect 10433 6518 10474 6526
rect 10556 6522 10569 6526
rect 10621 6530 10700 6546
rect 10732 6546 10904 6548
rect 10732 6530 10811 6546
rect 10818 6544 10848 6546
rect 10396 6508 10425 6518
rect 10439 6508 10468 6518
rect 10483 6508 10513 6522
rect 10556 6508 10599 6522
rect 10621 6518 10811 6530
rect 10876 6526 10882 6546
rect 10606 6508 10636 6518
rect 10637 6508 10795 6518
rect 10799 6508 10829 6518
rect 10833 6508 10863 6522
rect 10891 6508 10904 6546
rect 10976 6560 11005 6576
rect 11019 6560 11048 6576
rect 11063 6566 11093 6582
rect 11121 6560 11127 6608
rect 11130 6602 11149 6608
rect 11164 6602 11194 6610
rect 11130 6594 11194 6602
rect 11130 6578 11210 6594
rect 11226 6587 11288 6618
rect 11304 6587 11366 6618
rect 11435 6616 11484 6641
rect 11499 6616 11529 6632
rect 11398 6602 11428 6610
rect 11435 6608 11545 6616
rect 11398 6594 11443 6602
rect 11130 6576 11149 6578
rect 11164 6576 11210 6578
rect 11130 6560 11210 6576
rect 11237 6574 11272 6587
rect 11313 6584 11350 6587
rect 11313 6582 11355 6584
rect 11242 6571 11272 6574
rect 11251 6567 11258 6571
rect 11258 6566 11259 6567
rect 11217 6560 11227 6566
rect 10976 6552 11011 6560
rect 10976 6526 10977 6552
rect 10984 6526 11011 6552
rect 10919 6508 10949 6522
rect 10976 6518 11011 6526
rect 11013 6552 11054 6560
rect 11013 6526 11028 6552
rect 11035 6526 11054 6552
rect 11118 6548 11149 6560
rect 11164 6548 11267 6560
rect 11279 6550 11305 6576
rect 11320 6571 11350 6582
rect 11382 6578 11444 6594
rect 11382 6576 11428 6578
rect 11382 6560 11444 6576
rect 11456 6560 11462 6608
rect 11465 6600 11545 6608
rect 11465 6598 11484 6600
rect 11499 6598 11533 6600
rect 11465 6582 11545 6598
rect 11465 6560 11484 6582
rect 11499 6566 11529 6582
rect 11557 6576 11563 6650
rect 11566 6576 11585 6720
rect 11600 6576 11606 6720
rect 11615 6650 11628 6720
rect 11680 6716 11702 6720
rect 11673 6694 11702 6708
rect 11755 6694 11771 6708
rect 11809 6704 11815 6706
rect 11822 6704 11930 6720
rect 11937 6704 11943 6706
rect 11951 6704 11966 6720
rect 12032 6714 12051 6717
rect 11673 6692 11771 6694
rect 11798 6692 11966 6704
rect 11981 6694 11997 6708
rect 12032 6695 12054 6714
rect 12064 6708 12080 6709
rect 12063 6706 12080 6708
rect 12064 6701 12080 6706
rect 12054 6694 12060 6695
rect 12063 6694 12092 6701
rect 11981 6693 12092 6694
rect 11981 6692 12098 6693
rect 11657 6684 11708 6692
rect 11755 6684 11789 6692
rect 11657 6672 11682 6684
rect 11689 6672 11708 6684
rect 11762 6682 11789 6684
rect 11798 6682 12019 6692
rect 12054 6689 12060 6692
rect 11762 6678 12019 6682
rect 11657 6664 11708 6672
rect 11755 6664 12019 6678
rect 12063 6684 12098 6692
rect 11609 6616 11628 6650
rect 11673 6656 11702 6664
rect 11673 6650 11690 6656
rect 11673 6648 11707 6650
rect 11755 6648 11771 6664
rect 11772 6654 11980 6664
rect 11981 6654 11997 6664
rect 12045 6660 12060 6675
rect 12063 6672 12064 6684
rect 12071 6672 12098 6684
rect 12063 6664 12098 6672
rect 12063 6663 12092 6664
rect 11783 6650 11997 6654
rect 11798 6648 11997 6650
rect 12032 6650 12045 6660
rect 12063 6650 12080 6663
rect 12032 6648 12080 6650
rect 11674 6644 11707 6648
rect 11670 6642 11707 6644
rect 11670 6641 11737 6642
rect 11670 6636 11701 6641
rect 11707 6636 11737 6641
rect 11670 6632 11737 6636
rect 11643 6629 11737 6632
rect 11643 6622 11692 6629
rect 11643 6616 11673 6622
rect 11692 6617 11697 6622
rect 11609 6600 11689 6616
rect 11701 6608 11737 6629
rect 11798 6624 11987 6648
rect 12032 6647 12079 6648
rect 12045 6642 12079 6647
rect 11813 6621 11987 6624
rect 11806 6618 11987 6621
rect 12015 6641 12079 6642
rect 11609 6598 11628 6600
rect 11643 6598 11677 6600
rect 11609 6582 11689 6598
rect 11609 6576 11628 6582
rect 11325 6550 11428 6560
rect 11279 6548 11428 6550
rect 11449 6548 11484 6560
rect 11118 6546 11280 6548
rect 11130 6526 11149 6546
rect 11164 6544 11194 6546
rect 11013 6518 11054 6526
rect 11136 6522 11149 6526
rect 11201 6530 11280 6546
rect 11312 6546 11484 6548
rect 11312 6530 11391 6546
rect 11398 6544 11428 6546
rect 10976 6508 11005 6518
rect 11019 6508 11048 6518
rect 11063 6508 11093 6522
rect 11136 6508 11179 6522
rect 11201 6518 11391 6530
rect 11456 6526 11462 6546
rect 11186 6508 11216 6518
rect 11217 6508 11375 6518
rect 11379 6508 11409 6518
rect 11413 6508 11443 6522
rect 11471 6508 11484 6546
rect 11556 6560 11585 6576
rect 11599 6560 11628 6576
rect 11643 6566 11673 6582
rect 11701 6560 11707 6608
rect 11710 6602 11729 6608
rect 11744 6602 11774 6610
rect 11710 6594 11774 6602
rect 11710 6578 11790 6594
rect 11806 6587 11868 6618
rect 11884 6587 11946 6618
rect 12015 6616 12064 6641
rect 12079 6616 12109 6632
rect 11978 6602 12008 6610
rect 12015 6608 12125 6616
rect 11978 6594 12023 6602
rect 11710 6576 11729 6578
rect 11744 6576 11790 6578
rect 11710 6560 11790 6576
rect 11817 6574 11852 6587
rect 11893 6584 11930 6587
rect 11893 6582 11935 6584
rect 11822 6571 11852 6574
rect 11831 6567 11838 6571
rect 11838 6566 11839 6567
rect 11797 6560 11807 6566
rect 11556 6552 11591 6560
rect 11556 6526 11557 6552
rect 11564 6526 11591 6552
rect 11499 6508 11529 6522
rect 11556 6518 11591 6526
rect 11593 6552 11634 6560
rect 11593 6526 11608 6552
rect 11615 6526 11634 6552
rect 11698 6548 11729 6560
rect 11744 6548 11847 6560
rect 11859 6550 11885 6576
rect 11900 6571 11930 6582
rect 11962 6578 12024 6594
rect 11962 6576 12008 6578
rect 11962 6560 12024 6576
rect 12036 6560 12042 6608
rect 12045 6600 12125 6608
rect 12045 6598 12064 6600
rect 12079 6598 12113 6600
rect 12045 6582 12125 6598
rect 12045 6560 12064 6582
rect 12079 6566 12109 6582
rect 12137 6576 12143 6650
rect 12146 6576 12165 6720
rect 12180 6576 12186 6720
rect 12195 6650 12208 6720
rect 12260 6716 12282 6720
rect 12253 6694 12282 6708
rect 12335 6694 12351 6708
rect 12389 6704 12395 6706
rect 12402 6704 12510 6720
rect 12517 6704 12523 6706
rect 12531 6704 12546 6720
rect 12612 6714 12631 6717
rect 12253 6692 12351 6694
rect 12378 6692 12546 6704
rect 12561 6694 12577 6708
rect 12612 6695 12634 6714
rect 12644 6708 12660 6709
rect 12643 6706 12660 6708
rect 12644 6701 12660 6706
rect 12634 6694 12640 6695
rect 12643 6694 12672 6701
rect 12561 6693 12672 6694
rect 12561 6692 12678 6693
rect 12237 6684 12288 6692
rect 12335 6684 12369 6692
rect 12237 6672 12262 6684
rect 12269 6672 12288 6684
rect 12342 6682 12369 6684
rect 12378 6682 12599 6692
rect 12634 6689 12640 6692
rect 12342 6678 12599 6682
rect 12237 6664 12288 6672
rect 12335 6664 12599 6678
rect 12643 6684 12678 6692
rect 12189 6616 12208 6650
rect 12253 6656 12282 6664
rect 12253 6650 12270 6656
rect 12253 6648 12287 6650
rect 12335 6648 12351 6664
rect 12352 6654 12560 6664
rect 12561 6654 12577 6664
rect 12625 6660 12640 6675
rect 12643 6672 12644 6684
rect 12651 6672 12678 6684
rect 12643 6664 12678 6672
rect 12643 6663 12672 6664
rect 12363 6650 12577 6654
rect 12378 6648 12577 6650
rect 12612 6650 12625 6660
rect 12643 6650 12660 6663
rect 12612 6648 12660 6650
rect 12254 6644 12287 6648
rect 12250 6642 12287 6644
rect 12250 6641 12317 6642
rect 12250 6636 12281 6641
rect 12287 6636 12317 6641
rect 12250 6632 12317 6636
rect 12223 6629 12317 6632
rect 12223 6622 12272 6629
rect 12223 6616 12253 6622
rect 12272 6617 12277 6622
rect 12189 6600 12269 6616
rect 12281 6608 12317 6629
rect 12378 6624 12567 6648
rect 12612 6647 12659 6648
rect 12625 6642 12659 6647
rect 12393 6621 12567 6624
rect 12386 6618 12567 6621
rect 12595 6641 12659 6642
rect 12189 6598 12208 6600
rect 12223 6598 12257 6600
rect 12189 6582 12269 6598
rect 12189 6576 12208 6582
rect 11905 6550 12008 6560
rect 11859 6548 12008 6550
rect 12029 6548 12064 6560
rect 11698 6546 11860 6548
rect 11710 6526 11729 6546
rect 11744 6544 11774 6546
rect 11593 6518 11634 6526
rect 11716 6522 11729 6526
rect 11781 6530 11860 6546
rect 11892 6546 12064 6548
rect 11892 6530 11971 6546
rect 11978 6544 12008 6546
rect 11556 6508 11585 6518
rect 11599 6508 11628 6518
rect 11643 6508 11673 6522
rect 11716 6508 11759 6522
rect 11781 6518 11971 6530
rect 12036 6526 12042 6546
rect 11766 6508 11796 6518
rect 11797 6508 11955 6518
rect 11959 6508 11989 6518
rect 11993 6508 12023 6522
rect 12051 6508 12064 6546
rect 12136 6560 12165 6576
rect 12179 6560 12208 6576
rect 12223 6566 12253 6582
rect 12281 6560 12287 6608
rect 12290 6602 12309 6608
rect 12324 6602 12354 6610
rect 12290 6594 12354 6602
rect 12290 6578 12370 6594
rect 12386 6587 12448 6618
rect 12464 6587 12526 6618
rect 12595 6616 12644 6641
rect 12659 6616 12689 6632
rect 12558 6602 12588 6610
rect 12595 6608 12705 6616
rect 12558 6594 12603 6602
rect 12290 6576 12309 6578
rect 12324 6576 12370 6578
rect 12290 6560 12370 6576
rect 12397 6574 12432 6587
rect 12473 6584 12510 6587
rect 12473 6582 12515 6584
rect 12402 6571 12432 6574
rect 12411 6567 12418 6571
rect 12418 6566 12419 6567
rect 12377 6560 12387 6566
rect 12136 6552 12171 6560
rect 12136 6526 12137 6552
rect 12144 6526 12171 6552
rect 12079 6508 12109 6522
rect 12136 6518 12171 6526
rect 12173 6552 12214 6560
rect 12173 6526 12188 6552
rect 12195 6526 12214 6552
rect 12278 6548 12309 6560
rect 12324 6548 12427 6560
rect 12439 6550 12465 6576
rect 12480 6571 12510 6582
rect 12542 6578 12604 6594
rect 12542 6576 12588 6578
rect 12542 6560 12604 6576
rect 12616 6560 12622 6608
rect 12625 6600 12705 6608
rect 12625 6598 12644 6600
rect 12659 6598 12693 6600
rect 12625 6582 12705 6598
rect 12625 6560 12644 6582
rect 12659 6566 12689 6582
rect 12717 6576 12723 6650
rect 12726 6576 12745 6720
rect 12760 6576 12766 6720
rect 12775 6650 12788 6720
rect 12840 6716 12862 6720
rect 12833 6694 12862 6708
rect 12915 6694 12931 6708
rect 12969 6704 12975 6706
rect 12982 6704 13090 6720
rect 13097 6704 13103 6706
rect 13111 6704 13126 6720
rect 13192 6714 13211 6717
rect 12833 6692 12931 6694
rect 12958 6692 13126 6704
rect 13141 6694 13157 6708
rect 13192 6695 13214 6714
rect 13224 6708 13240 6709
rect 13223 6706 13240 6708
rect 13224 6701 13240 6706
rect 13214 6694 13220 6695
rect 13223 6694 13252 6701
rect 13141 6693 13252 6694
rect 13141 6692 13258 6693
rect 12817 6684 12868 6692
rect 12915 6684 12949 6692
rect 12817 6672 12842 6684
rect 12849 6672 12868 6684
rect 12922 6682 12949 6684
rect 12958 6682 13179 6692
rect 13214 6689 13220 6692
rect 12922 6678 13179 6682
rect 12817 6664 12868 6672
rect 12915 6664 13179 6678
rect 13223 6684 13258 6692
rect 12769 6616 12788 6650
rect 12833 6656 12862 6664
rect 12833 6650 12850 6656
rect 12833 6648 12867 6650
rect 12915 6648 12931 6664
rect 12932 6654 13140 6664
rect 13141 6654 13157 6664
rect 13205 6660 13220 6675
rect 13223 6672 13224 6684
rect 13231 6672 13258 6684
rect 13223 6664 13258 6672
rect 13223 6663 13252 6664
rect 12943 6650 13157 6654
rect 12958 6648 13157 6650
rect 13192 6650 13205 6660
rect 13223 6650 13240 6663
rect 13192 6648 13240 6650
rect 12834 6644 12867 6648
rect 12830 6642 12867 6644
rect 12830 6641 12897 6642
rect 12830 6636 12861 6641
rect 12867 6636 12897 6641
rect 12830 6632 12897 6636
rect 12803 6629 12897 6632
rect 12803 6622 12852 6629
rect 12803 6616 12833 6622
rect 12852 6617 12857 6622
rect 12769 6600 12849 6616
rect 12861 6608 12897 6629
rect 12958 6624 13147 6648
rect 13192 6647 13239 6648
rect 13205 6642 13239 6647
rect 12973 6621 13147 6624
rect 12966 6618 13147 6621
rect 13175 6641 13239 6642
rect 12769 6598 12788 6600
rect 12803 6598 12837 6600
rect 12769 6582 12849 6598
rect 12769 6576 12788 6582
rect 12485 6550 12588 6560
rect 12439 6548 12588 6550
rect 12609 6548 12644 6560
rect 12278 6546 12440 6548
rect 12290 6526 12309 6546
rect 12324 6544 12354 6546
rect 12173 6518 12214 6526
rect 12296 6522 12309 6526
rect 12361 6530 12440 6546
rect 12472 6546 12644 6548
rect 12472 6530 12551 6546
rect 12558 6544 12588 6546
rect 12136 6508 12165 6518
rect 12179 6508 12208 6518
rect 12223 6508 12253 6522
rect 12296 6508 12339 6522
rect 12361 6518 12551 6530
rect 12616 6526 12622 6546
rect 12346 6508 12376 6518
rect 12377 6508 12535 6518
rect 12539 6508 12569 6518
rect 12573 6508 12603 6522
rect 12631 6508 12644 6546
rect 12716 6560 12745 6576
rect 12759 6560 12788 6576
rect 12803 6566 12833 6582
rect 12861 6560 12867 6608
rect 12870 6602 12889 6608
rect 12904 6602 12934 6610
rect 12870 6594 12934 6602
rect 12870 6578 12950 6594
rect 12966 6587 13028 6618
rect 13044 6587 13106 6618
rect 13175 6616 13224 6641
rect 13239 6616 13269 6632
rect 13138 6602 13168 6610
rect 13175 6608 13285 6616
rect 13138 6594 13183 6602
rect 12870 6576 12889 6578
rect 12904 6576 12950 6578
rect 12870 6560 12950 6576
rect 12977 6574 13012 6587
rect 13053 6584 13090 6587
rect 13053 6582 13095 6584
rect 12982 6571 13012 6574
rect 12991 6567 12998 6571
rect 12998 6566 12999 6567
rect 12957 6560 12967 6566
rect 12716 6552 12751 6560
rect 12716 6526 12717 6552
rect 12724 6526 12751 6552
rect 12659 6508 12689 6522
rect 12716 6518 12751 6526
rect 12753 6552 12794 6560
rect 12753 6526 12768 6552
rect 12775 6526 12794 6552
rect 12858 6548 12889 6560
rect 12904 6548 13007 6560
rect 13019 6550 13045 6576
rect 13060 6571 13090 6582
rect 13122 6578 13184 6594
rect 13122 6576 13168 6578
rect 13122 6560 13184 6576
rect 13196 6560 13202 6608
rect 13205 6600 13285 6608
rect 13205 6598 13224 6600
rect 13239 6598 13273 6600
rect 13205 6582 13285 6598
rect 13205 6560 13224 6582
rect 13239 6566 13269 6582
rect 13297 6576 13303 6650
rect 13306 6576 13325 6720
rect 13340 6576 13346 6720
rect 13355 6650 13368 6720
rect 13420 6716 13442 6720
rect 13413 6694 13442 6708
rect 13495 6694 13511 6708
rect 13549 6704 13555 6706
rect 13562 6704 13670 6720
rect 13677 6704 13683 6706
rect 13691 6704 13706 6720
rect 13772 6714 13791 6717
rect 13413 6692 13511 6694
rect 13538 6692 13706 6704
rect 13721 6694 13737 6708
rect 13772 6695 13794 6714
rect 13804 6708 13820 6709
rect 13803 6706 13820 6708
rect 13804 6701 13820 6706
rect 13794 6694 13800 6695
rect 13803 6694 13832 6701
rect 13721 6693 13832 6694
rect 13721 6692 13838 6693
rect 13397 6684 13448 6692
rect 13495 6684 13529 6692
rect 13397 6672 13422 6684
rect 13429 6672 13448 6684
rect 13502 6682 13529 6684
rect 13538 6682 13759 6692
rect 13794 6689 13800 6692
rect 13502 6678 13759 6682
rect 13397 6664 13448 6672
rect 13495 6664 13759 6678
rect 13803 6684 13838 6692
rect 13349 6616 13368 6650
rect 13413 6656 13442 6664
rect 13413 6650 13430 6656
rect 13413 6648 13447 6650
rect 13495 6648 13511 6664
rect 13512 6654 13720 6664
rect 13721 6654 13737 6664
rect 13785 6660 13800 6675
rect 13803 6672 13804 6684
rect 13811 6672 13838 6684
rect 13803 6664 13838 6672
rect 13803 6663 13832 6664
rect 13523 6650 13737 6654
rect 13538 6648 13737 6650
rect 13772 6650 13785 6660
rect 13803 6650 13820 6663
rect 13772 6648 13820 6650
rect 13414 6644 13447 6648
rect 13410 6642 13447 6644
rect 13410 6641 13477 6642
rect 13410 6636 13441 6641
rect 13447 6636 13477 6641
rect 13410 6632 13477 6636
rect 13383 6629 13477 6632
rect 13383 6622 13432 6629
rect 13383 6616 13413 6622
rect 13432 6617 13437 6622
rect 13349 6600 13429 6616
rect 13441 6608 13477 6629
rect 13538 6624 13727 6648
rect 13772 6647 13819 6648
rect 13785 6642 13819 6647
rect 13553 6621 13727 6624
rect 13546 6618 13727 6621
rect 13755 6641 13819 6642
rect 13349 6598 13368 6600
rect 13383 6598 13417 6600
rect 13349 6582 13429 6598
rect 13349 6576 13368 6582
rect 13065 6550 13168 6560
rect 13019 6548 13168 6550
rect 13189 6548 13224 6560
rect 12858 6546 13020 6548
rect 12870 6526 12889 6546
rect 12904 6544 12934 6546
rect 12753 6518 12794 6526
rect 12876 6522 12889 6526
rect 12941 6530 13020 6546
rect 13052 6546 13224 6548
rect 13052 6530 13131 6546
rect 13138 6544 13168 6546
rect 12716 6508 12745 6518
rect 12759 6508 12788 6518
rect 12803 6508 12833 6522
rect 12876 6508 12919 6522
rect 12941 6518 13131 6530
rect 13196 6526 13202 6546
rect 12926 6508 12956 6518
rect 12957 6508 13115 6518
rect 13119 6508 13149 6518
rect 13153 6508 13183 6522
rect 13211 6508 13224 6546
rect 13296 6560 13325 6576
rect 13339 6560 13368 6576
rect 13383 6566 13413 6582
rect 13441 6560 13447 6608
rect 13450 6602 13469 6608
rect 13484 6602 13514 6610
rect 13450 6594 13514 6602
rect 13450 6578 13530 6594
rect 13546 6587 13608 6618
rect 13624 6587 13686 6618
rect 13755 6616 13804 6641
rect 13819 6616 13849 6632
rect 13718 6602 13748 6610
rect 13755 6608 13865 6616
rect 13718 6594 13763 6602
rect 13450 6576 13469 6578
rect 13484 6576 13530 6578
rect 13450 6560 13530 6576
rect 13557 6574 13592 6587
rect 13633 6584 13670 6587
rect 13633 6582 13675 6584
rect 13562 6571 13592 6574
rect 13571 6567 13578 6571
rect 13578 6566 13579 6567
rect 13537 6560 13547 6566
rect 13296 6552 13331 6560
rect 13296 6526 13297 6552
rect 13304 6526 13331 6552
rect 13239 6508 13269 6522
rect 13296 6518 13331 6526
rect 13333 6552 13374 6560
rect 13333 6526 13348 6552
rect 13355 6526 13374 6552
rect 13438 6548 13469 6560
rect 13484 6548 13587 6560
rect 13599 6550 13625 6576
rect 13640 6571 13670 6582
rect 13702 6578 13764 6594
rect 13702 6576 13748 6578
rect 13702 6560 13764 6576
rect 13776 6560 13782 6608
rect 13785 6600 13865 6608
rect 13785 6598 13804 6600
rect 13819 6598 13853 6600
rect 13785 6582 13865 6598
rect 13785 6560 13804 6582
rect 13819 6566 13849 6582
rect 13877 6576 13883 6650
rect 13886 6576 13905 6720
rect 13920 6576 13926 6720
rect 13935 6650 13948 6720
rect 14000 6716 14022 6720
rect 13993 6694 14022 6708
rect 14075 6694 14091 6708
rect 14129 6704 14135 6706
rect 14142 6704 14250 6720
rect 14257 6704 14263 6706
rect 14271 6704 14286 6720
rect 14352 6714 14371 6717
rect 13993 6692 14091 6694
rect 14118 6692 14286 6704
rect 14301 6694 14317 6708
rect 14352 6695 14374 6714
rect 14384 6708 14400 6709
rect 14383 6706 14400 6708
rect 14384 6701 14400 6706
rect 14374 6694 14380 6695
rect 14383 6694 14412 6701
rect 14301 6693 14412 6694
rect 14301 6692 14418 6693
rect 13977 6684 14028 6692
rect 14075 6684 14109 6692
rect 13977 6672 14002 6684
rect 14009 6672 14028 6684
rect 14082 6682 14109 6684
rect 14118 6682 14339 6692
rect 14374 6689 14380 6692
rect 14082 6678 14339 6682
rect 13977 6664 14028 6672
rect 14075 6664 14339 6678
rect 14383 6684 14418 6692
rect 13929 6616 13948 6650
rect 13993 6656 14022 6664
rect 13993 6650 14010 6656
rect 13993 6648 14027 6650
rect 14075 6648 14091 6664
rect 14092 6654 14300 6664
rect 14301 6654 14317 6664
rect 14365 6660 14380 6675
rect 14383 6672 14384 6684
rect 14391 6672 14418 6684
rect 14383 6664 14418 6672
rect 14383 6663 14412 6664
rect 14103 6650 14317 6654
rect 14118 6648 14317 6650
rect 14352 6650 14365 6660
rect 14383 6650 14400 6663
rect 14352 6648 14400 6650
rect 13994 6644 14027 6648
rect 13990 6642 14027 6644
rect 13990 6641 14057 6642
rect 13990 6636 14021 6641
rect 14027 6636 14057 6641
rect 13990 6632 14057 6636
rect 13963 6629 14057 6632
rect 13963 6622 14012 6629
rect 13963 6616 13993 6622
rect 14012 6617 14017 6622
rect 13929 6600 14009 6616
rect 14021 6608 14057 6629
rect 14118 6624 14307 6648
rect 14352 6647 14399 6648
rect 14365 6642 14399 6647
rect 14133 6621 14307 6624
rect 14126 6618 14307 6621
rect 14335 6641 14399 6642
rect 13929 6598 13948 6600
rect 13963 6598 13997 6600
rect 13929 6582 14009 6598
rect 13929 6576 13948 6582
rect 13645 6550 13748 6560
rect 13599 6548 13748 6550
rect 13769 6548 13804 6560
rect 13438 6546 13600 6548
rect 13450 6526 13469 6546
rect 13484 6544 13514 6546
rect 13333 6518 13374 6526
rect 13456 6522 13469 6526
rect 13521 6530 13600 6546
rect 13632 6546 13804 6548
rect 13632 6530 13711 6546
rect 13718 6544 13748 6546
rect 13296 6508 13325 6518
rect 13339 6508 13368 6518
rect 13383 6508 13413 6522
rect 13456 6508 13499 6522
rect 13521 6518 13711 6530
rect 13776 6526 13782 6546
rect 13506 6508 13536 6518
rect 13537 6508 13695 6518
rect 13699 6508 13729 6518
rect 13733 6508 13763 6522
rect 13791 6508 13804 6546
rect 13876 6560 13905 6576
rect 13919 6560 13948 6576
rect 13963 6566 13993 6582
rect 14021 6560 14027 6608
rect 14030 6602 14049 6608
rect 14064 6602 14094 6610
rect 14030 6594 14094 6602
rect 14030 6578 14110 6594
rect 14126 6587 14188 6618
rect 14204 6587 14266 6618
rect 14335 6616 14384 6641
rect 14399 6616 14429 6632
rect 14298 6602 14328 6610
rect 14335 6608 14445 6616
rect 14298 6594 14343 6602
rect 14030 6576 14049 6578
rect 14064 6576 14110 6578
rect 14030 6560 14110 6576
rect 14137 6574 14172 6587
rect 14213 6584 14250 6587
rect 14213 6582 14255 6584
rect 14142 6571 14172 6574
rect 14151 6567 14158 6571
rect 14158 6566 14159 6567
rect 14117 6560 14127 6566
rect 13876 6552 13911 6560
rect 13876 6526 13877 6552
rect 13884 6526 13911 6552
rect 13819 6508 13849 6522
rect 13876 6518 13911 6526
rect 13913 6552 13954 6560
rect 13913 6526 13928 6552
rect 13935 6526 13954 6552
rect 14018 6548 14049 6560
rect 14064 6548 14167 6560
rect 14179 6550 14205 6576
rect 14220 6571 14250 6582
rect 14282 6578 14344 6594
rect 14282 6576 14328 6578
rect 14282 6560 14344 6576
rect 14356 6560 14362 6608
rect 14365 6600 14445 6608
rect 14365 6598 14384 6600
rect 14399 6598 14433 6600
rect 14365 6582 14445 6598
rect 14365 6560 14384 6582
rect 14399 6566 14429 6582
rect 14457 6576 14463 6650
rect 14466 6576 14485 6720
rect 14500 6576 14506 6720
rect 14515 6650 14528 6720
rect 14580 6716 14602 6720
rect 14573 6694 14602 6708
rect 14655 6694 14671 6708
rect 14709 6704 14715 6706
rect 14722 6704 14830 6720
rect 14837 6704 14843 6706
rect 14851 6704 14866 6720
rect 14932 6714 14951 6717
rect 14573 6692 14671 6694
rect 14698 6692 14866 6704
rect 14881 6694 14897 6708
rect 14932 6695 14954 6714
rect 14964 6708 14980 6709
rect 14963 6706 14980 6708
rect 14964 6701 14980 6706
rect 14954 6694 14960 6695
rect 14963 6694 14992 6701
rect 14881 6693 14992 6694
rect 14881 6692 14998 6693
rect 14557 6684 14608 6692
rect 14655 6684 14689 6692
rect 14557 6672 14582 6684
rect 14589 6672 14608 6684
rect 14662 6682 14689 6684
rect 14698 6682 14919 6692
rect 14954 6689 14960 6692
rect 14662 6678 14919 6682
rect 14557 6664 14608 6672
rect 14655 6664 14919 6678
rect 14963 6684 14998 6692
rect 14509 6616 14528 6650
rect 14573 6656 14602 6664
rect 14573 6650 14590 6656
rect 14573 6648 14607 6650
rect 14655 6648 14671 6664
rect 14672 6654 14880 6664
rect 14881 6654 14897 6664
rect 14945 6660 14960 6675
rect 14963 6672 14964 6684
rect 14971 6672 14998 6684
rect 14963 6664 14998 6672
rect 14963 6663 14992 6664
rect 14683 6650 14897 6654
rect 14698 6648 14897 6650
rect 14932 6650 14945 6660
rect 14963 6650 14980 6663
rect 14932 6648 14980 6650
rect 14574 6644 14607 6648
rect 14570 6642 14607 6644
rect 14570 6641 14637 6642
rect 14570 6636 14601 6641
rect 14607 6636 14637 6641
rect 14570 6632 14637 6636
rect 14543 6629 14637 6632
rect 14543 6622 14592 6629
rect 14543 6616 14573 6622
rect 14592 6617 14597 6622
rect 14509 6600 14589 6616
rect 14601 6608 14637 6629
rect 14698 6624 14887 6648
rect 14932 6647 14979 6648
rect 14945 6642 14979 6647
rect 14713 6621 14887 6624
rect 14706 6618 14887 6621
rect 14915 6641 14979 6642
rect 14509 6598 14528 6600
rect 14543 6598 14577 6600
rect 14509 6582 14589 6598
rect 14509 6576 14528 6582
rect 14225 6550 14328 6560
rect 14179 6548 14328 6550
rect 14349 6548 14384 6560
rect 14018 6546 14180 6548
rect 14030 6526 14049 6546
rect 14064 6544 14094 6546
rect 13913 6518 13954 6526
rect 14036 6522 14049 6526
rect 14101 6530 14180 6546
rect 14212 6546 14384 6548
rect 14212 6530 14291 6546
rect 14298 6544 14328 6546
rect 13876 6508 13905 6518
rect 13919 6508 13948 6518
rect 13963 6508 13993 6522
rect 14036 6508 14079 6522
rect 14101 6518 14291 6530
rect 14356 6526 14362 6546
rect 14086 6508 14116 6518
rect 14117 6508 14275 6518
rect 14279 6508 14309 6518
rect 14313 6508 14343 6522
rect 14371 6508 14384 6546
rect 14456 6560 14485 6576
rect 14499 6560 14528 6576
rect 14543 6566 14573 6582
rect 14601 6560 14607 6608
rect 14610 6602 14629 6608
rect 14644 6602 14674 6610
rect 14610 6594 14674 6602
rect 14610 6578 14690 6594
rect 14706 6587 14768 6618
rect 14784 6587 14846 6618
rect 14915 6616 14964 6641
rect 14979 6616 15009 6632
rect 14878 6602 14908 6610
rect 14915 6608 15025 6616
rect 14878 6594 14923 6602
rect 14610 6576 14629 6578
rect 14644 6576 14690 6578
rect 14610 6560 14690 6576
rect 14717 6574 14752 6587
rect 14793 6584 14830 6587
rect 14793 6582 14835 6584
rect 14722 6571 14752 6574
rect 14731 6567 14738 6571
rect 14738 6566 14739 6567
rect 14697 6560 14707 6566
rect 14456 6552 14491 6560
rect 14456 6526 14457 6552
rect 14464 6526 14491 6552
rect 14399 6508 14429 6522
rect 14456 6518 14491 6526
rect 14493 6552 14534 6560
rect 14493 6526 14508 6552
rect 14515 6526 14534 6552
rect 14598 6548 14629 6560
rect 14644 6548 14747 6560
rect 14759 6550 14785 6576
rect 14800 6571 14830 6582
rect 14862 6578 14924 6594
rect 14862 6576 14908 6578
rect 14862 6560 14924 6576
rect 14936 6560 14942 6608
rect 14945 6600 15025 6608
rect 14945 6598 14964 6600
rect 14979 6598 15013 6600
rect 14945 6582 15025 6598
rect 14945 6560 14964 6582
rect 14979 6566 15009 6582
rect 15037 6576 15043 6650
rect 15046 6576 15065 6720
rect 15080 6576 15086 6720
rect 15095 6650 15108 6720
rect 15160 6716 15182 6720
rect 15153 6694 15182 6708
rect 15235 6694 15251 6708
rect 15289 6704 15295 6706
rect 15302 6704 15410 6720
rect 15417 6704 15423 6706
rect 15431 6704 15446 6720
rect 15512 6714 15531 6717
rect 15153 6692 15251 6694
rect 15278 6692 15446 6704
rect 15461 6694 15477 6708
rect 15512 6695 15534 6714
rect 15544 6708 15560 6709
rect 15543 6706 15560 6708
rect 15544 6701 15560 6706
rect 15534 6694 15540 6695
rect 15543 6694 15572 6701
rect 15461 6693 15572 6694
rect 15461 6692 15578 6693
rect 15137 6684 15188 6692
rect 15235 6684 15269 6692
rect 15137 6672 15162 6684
rect 15169 6672 15188 6684
rect 15242 6682 15269 6684
rect 15278 6682 15499 6692
rect 15534 6689 15540 6692
rect 15242 6678 15499 6682
rect 15137 6664 15188 6672
rect 15235 6664 15499 6678
rect 15543 6684 15578 6692
rect 15089 6616 15108 6650
rect 15153 6656 15182 6664
rect 15153 6650 15170 6656
rect 15153 6648 15187 6650
rect 15235 6648 15251 6664
rect 15252 6654 15460 6664
rect 15461 6654 15477 6664
rect 15525 6660 15540 6675
rect 15543 6672 15544 6684
rect 15551 6672 15578 6684
rect 15543 6664 15578 6672
rect 15543 6663 15572 6664
rect 15263 6650 15477 6654
rect 15278 6648 15477 6650
rect 15512 6650 15525 6660
rect 15543 6650 15560 6663
rect 15512 6648 15560 6650
rect 15154 6644 15187 6648
rect 15150 6642 15187 6644
rect 15150 6641 15217 6642
rect 15150 6636 15181 6641
rect 15187 6636 15217 6641
rect 15150 6632 15217 6636
rect 15123 6629 15217 6632
rect 15123 6622 15172 6629
rect 15123 6616 15153 6622
rect 15172 6617 15177 6622
rect 15089 6600 15169 6616
rect 15181 6608 15217 6629
rect 15278 6624 15467 6648
rect 15512 6647 15559 6648
rect 15525 6642 15559 6647
rect 15293 6621 15467 6624
rect 15286 6618 15467 6621
rect 15495 6641 15559 6642
rect 15089 6598 15108 6600
rect 15123 6598 15157 6600
rect 15089 6582 15169 6598
rect 15089 6576 15108 6582
rect 14805 6550 14908 6560
rect 14759 6548 14908 6550
rect 14929 6548 14964 6560
rect 14598 6546 14760 6548
rect 14610 6526 14629 6546
rect 14644 6544 14674 6546
rect 14493 6518 14534 6526
rect 14616 6522 14629 6526
rect 14681 6530 14760 6546
rect 14792 6546 14964 6548
rect 14792 6530 14871 6546
rect 14878 6544 14908 6546
rect 14456 6508 14485 6518
rect 14499 6508 14528 6518
rect 14543 6508 14573 6522
rect 14616 6508 14659 6522
rect 14681 6518 14871 6530
rect 14936 6526 14942 6546
rect 14666 6508 14696 6518
rect 14697 6508 14855 6518
rect 14859 6508 14889 6518
rect 14893 6508 14923 6522
rect 14951 6508 14964 6546
rect 15036 6560 15065 6576
rect 15079 6560 15108 6576
rect 15123 6566 15153 6582
rect 15181 6560 15187 6608
rect 15190 6602 15209 6608
rect 15224 6602 15254 6610
rect 15190 6594 15254 6602
rect 15190 6578 15270 6594
rect 15286 6587 15348 6618
rect 15364 6587 15426 6618
rect 15495 6616 15544 6641
rect 15559 6616 15589 6632
rect 15458 6602 15488 6610
rect 15495 6608 15605 6616
rect 15458 6594 15503 6602
rect 15190 6576 15209 6578
rect 15224 6576 15270 6578
rect 15190 6560 15270 6576
rect 15297 6574 15332 6587
rect 15373 6584 15410 6587
rect 15373 6582 15415 6584
rect 15302 6571 15332 6574
rect 15311 6567 15318 6571
rect 15318 6566 15319 6567
rect 15277 6560 15287 6566
rect 15036 6552 15071 6560
rect 15036 6526 15037 6552
rect 15044 6526 15071 6552
rect 14979 6508 15009 6522
rect 15036 6518 15071 6526
rect 15073 6552 15114 6560
rect 15073 6526 15088 6552
rect 15095 6526 15114 6552
rect 15178 6548 15209 6560
rect 15224 6548 15327 6560
rect 15339 6550 15365 6576
rect 15380 6571 15410 6582
rect 15442 6578 15504 6594
rect 15442 6576 15488 6578
rect 15442 6560 15504 6576
rect 15516 6560 15522 6608
rect 15525 6600 15605 6608
rect 15525 6598 15544 6600
rect 15559 6598 15593 6600
rect 15525 6582 15605 6598
rect 15525 6560 15544 6582
rect 15559 6566 15589 6582
rect 15617 6576 15623 6650
rect 15626 6576 15645 6720
rect 15660 6576 15666 6720
rect 15675 6650 15688 6720
rect 15740 6716 15762 6720
rect 15733 6694 15762 6708
rect 15815 6694 15831 6708
rect 15869 6704 15875 6706
rect 15882 6704 15990 6720
rect 15997 6704 16003 6706
rect 16011 6704 16026 6720
rect 16092 6714 16111 6717
rect 15733 6692 15831 6694
rect 15858 6692 16026 6704
rect 16041 6694 16057 6708
rect 16092 6695 16114 6714
rect 16124 6708 16140 6709
rect 16123 6706 16140 6708
rect 16124 6701 16140 6706
rect 16114 6694 16120 6695
rect 16123 6694 16152 6701
rect 16041 6693 16152 6694
rect 16041 6692 16158 6693
rect 15717 6684 15768 6692
rect 15815 6684 15849 6692
rect 15717 6672 15742 6684
rect 15749 6672 15768 6684
rect 15822 6682 15849 6684
rect 15858 6682 16079 6692
rect 16114 6689 16120 6692
rect 15822 6678 16079 6682
rect 15717 6664 15768 6672
rect 15815 6664 16079 6678
rect 16123 6684 16158 6692
rect 15669 6616 15688 6650
rect 15733 6656 15762 6664
rect 15733 6650 15750 6656
rect 15733 6648 15767 6650
rect 15815 6648 15831 6664
rect 15832 6654 16040 6664
rect 16041 6654 16057 6664
rect 16105 6660 16120 6675
rect 16123 6672 16124 6684
rect 16131 6672 16158 6684
rect 16123 6664 16158 6672
rect 16123 6663 16152 6664
rect 15843 6650 16057 6654
rect 15858 6648 16057 6650
rect 16092 6650 16105 6660
rect 16123 6650 16140 6663
rect 16092 6648 16140 6650
rect 15734 6644 15767 6648
rect 15730 6642 15767 6644
rect 15730 6641 15797 6642
rect 15730 6636 15761 6641
rect 15767 6636 15797 6641
rect 15730 6632 15797 6636
rect 15703 6629 15797 6632
rect 15703 6622 15752 6629
rect 15703 6616 15733 6622
rect 15752 6617 15757 6622
rect 15669 6600 15749 6616
rect 15761 6608 15797 6629
rect 15858 6624 16047 6648
rect 16092 6647 16139 6648
rect 16105 6642 16139 6647
rect 15873 6621 16047 6624
rect 15866 6618 16047 6621
rect 16075 6641 16139 6642
rect 15669 6598 15688 6600
rect 15703 6598 15737 6600
rect 15669 6582 15749 6598
rect 15669 6576 15688 6582
rect 15385 6550 15488 6560
rect 15339 6548 15488 6550
rect 15509 6548 15544 6560
rect 15178 6546 15340 6548
rect 15190 6526 15209 6546
rect 15224 6544 15254 6546
rect 15073 6518 15114 6526
rect 15196 6522 15209 6526
rect 15261 6530 15340 6546
rect 15372 6546 15544 6548
rect 15372 6530 15451 6546
rect 15458 6544 15488 6546
rect 15036 6508 15065 6518
rect 15079 6508 15108 6518
rect 15123 6508 15153 6522
rect 15196 6508 15239 6522
rect 15261 6518 15451 6530
rect 15516 6526 15522 6546
rect 15246 6508 15276 6518
rect 15277 6508 15435 6518
rect 15439 6508 15469 6518
rect 15473 6508 15503 6522
rect 15531 6508 15544 6546
rect 15616 6560 15645 6576
rect 15659 6560 15688 6576
rect 15703 6566 15733 6582
rect 15761 6560 15767 6608
rect 15770 6602 15789 6608
rect 15804 6602 15834 6610
rect 15770 6594 15834 6602
rect 15770 6578 15850 6594
rect 15866 6587 15928 6618
rect 15944 6587 16006 6618
rect 16075 6616 16124 6641
rect 16139 6616 16169 6632
rect 16038 6602 16068 6610
rect 16075 6608 16185 6616
rect 16038 6594 16083 6602
rect 15770 6576 15789 6578
rect 15804 6576 15850 6578
rect 15770 6560 15850 6576
rect 15877 6574 15912 6587
rect 15953 6584 15990 6587
rect 15953 6582 15995 6584
rect 15882 6571 15912 6574
rect 15891 6567 15898 6571
rect 15898 6566 15899 6567
rect 15857 6560 15867 6566
rect 15616 6552 15651 6560
rect 15616 6526 15617 6552
rect 15624 6526 15651 6552
rect 15559 6508 15589 6522
rect 15616 6518 15651 6526
rect 15653 6552 15694 6560
rect 15653 6526 15668 6552
rect 15675 6526 15694 6552
rect 15758 6548 15789 6560
rect 15804 6548 15907 6560
rect 15919 6550 15945 6576
rect 15960 6571 15990 6582
rect 16022 6578 16084 6594
rect 16022 6576 16068 6578
rect 16022 6560 16084 6576
rect 16096 6560 16102 6608
rect 16105 6600 16185 6608
rect 16105 6598 16124 6600
rect 16139 6598 16173 6600
rect 16105 6582 16185 6598
rect 16105 6560 16124 6582
rect 16139 6566 16169 6582
rect 16197 6576 16203 6650
rect 16206 6576 16225 6720
rect 16240 6576 16246 6720
rect 16255 6650 16268 6720
rect 16320 6716 16342 6720
rect 16313 6694 16342 6708
rect 16395 6694 16411 6708
rect 16449 6704 16455 6706
rect 16462 6704 16570 6720
rect 16577 6704 16583 6706
rect 16591 6704 16606 6720
rect 16672 6714 16691 6717
rect 16313 6692 16411 6694
rect 16438 6692 16606 6704
rect 16621 6694 16637 6708
rect 16672 6695 16694 6714
rect 16704 6708 16720 6709
rect 16703 6706 16720 6708
rect 16704 6701 16720 6706
rect 16694 6694 16700 6695
rect 16703 6694 16732 6701
rect 16621 6693 16732 6694
rect 16621 6692 16738 6693
rect 16297 6684 16348 6692
rect 16395 6684 16429 6692
rect 16297 6672 16322 6684
rect 16329 6672 16348 6684
rect 16402 6682 16429 6684
rect 16438 6682 16659 6692
rect 16694 6689 16700 6692
rect 16402 6678 16659 6682
rect 16297 6664 16348 6672
rect 16395 6664 16659 6678
rect 16703 6684 16738 6692
rect 16249 6616 16268 6650
rect 16313 6656 16342 6664
rect 16313 6650 16330 6656
rect 16313 6648 16347 6650
rect 16395 6648 16411 6664
rect 16412 6654 16620 6664
rect 16621 6654 16637 6664
rect 16685 6660 16700 6675
rect 16703 6672 16704 6684
rect 16711 6672 16738 6684
rect 16703 6664 16738 6672
rect 16703 6663 16732 6664
rect 16423 6650 16637 6654
rect 16438 6648 16637 6650
rect 16672 6650 16685 6660
rect 16703 6650 16720 6663
rect 16672 6648 16720 6650
rect 16314 6644 16347 6648
rect 16310 6642 16347 6644
rect 16310 6641 16377 6642
rect 16310 6636 16341 6641
rect 16347 6636 16377 6641
rect 16310 6632 16377 6636
rect 16283 6629 16377 6632
rect 16283 6622 16332 6629
rect 16283 6616 16313 6622
rect 16332 6617 16337 6622
rect 16249 6600 16329 6616
rect 16341 6608 16377 6629
rect 16438 6624 16627 6648
rect 16672 6647 16719 6648
rect 16685 6642 16719 6647
rect 16453 6621 16627 6624
rect 16446 6618 16627 6621
rect 16655 6641 16719 6642
rect 16249 6598 16268 6600
rect 16283 6598 16317 6600
rect 16249 6582 16329 6598
rect 16249 6576 16268 6582
rect 15965 6550 16068 6560
rect 15919 6548 16068 6550
rect 16089 6548 16124 6560
rect 15758 6546 15920 6548
rect 15770 6526 15789 6546
rect 15804 6544 15834 6546
rect 15653 6518 15694 6526
rect 15776 6522 15789 6526
rect 15841 6530 15920 6546
rect 15952 6546 16124 6548
rect 15952 6530 16031 6546
rect 16038 6544 16068 6546
rect 15616 6508 15645 6518
rect 15659 6508 15688 6518
rect 15703 6508 15733 6522
rect 15776 6508 15819 6522
rect 15841 6518 16031 6530
rect 16096 6526 16102 6546
rect 15826 6508 15856 6518
rect 15857 6508 16015 6518
rect 16019 6508 16049 6518
rect 16053 6508 16083 6522
rect 16111 6508 16124 6546
rect 16196 6560 16225 6576
rect 16239 6560 16268 6576
rect 16283 6566 16313 6582
rect 16341 6560 16347 6608
rect 16350 6602 16369 6608
rect 16384 6602 16414 6610
rect 16350 6594 16414 6602
rect 16350 6578 16430 6594
rect 16446 6587 16508 6618
rect 16524 6587 16586 6618
rect 16655 6616 16704 6641
rect 16719 6616 16749 6632
rect 16618 6602 16648 6610
rect 16655 6608 16765 6616
rect 16618 6594 16663 6602
rect 16350 6576 16369 6578
rect 16384 6576 16430 6578
rect 16350 6560 16430 6576
rect 16457 6574 16492 6587
rect 16533 6584 16570 6587
rect 16533 6582 16575 6584
rect 16462 6571 16492 6574
rect 16471 6567 16478 6571
rect 16478 6566 16479 6567
rect 16437 6560 16447 6566
rect 16196 6552 16231 6560
rect 16196 6526 16197 6552
rect 16204 6526 16231 6552
rect 16139 6508 16169 6522
rect 16196 6518 16231 6526
rect 16233 6552 16274 6560
rect 16233 6526 16248 6552
rect 16255 6526 16274 6552
rect 16338 6548 16369 6560
rect 16384 6548 16487 6560
rect 16499 6550 16525 6576
rect 16540 6571 16570 6582
rect 16602 6578 16664 6594
rect 16602 6576 16648 6578
rect 16602 6560 16664 6576
rect 16676 6560 16682 6608
rect 16685 6600 16765 6608
rect 16685 6598 16704 6600
rect 16719 6598 16753 6600
rect 16685 6582 16765 6598
rect 16685 6560 16704 6582
rect 16719 6566 16749 6582
rect 16777 6576 16783 6650
rect 16786 6576 16805 6720
rect 16820 6576 16826 6720
rect 16835 6650 16848 6720
rect 16900 6716 16922 6720
rect 16893 6694 16922 6708
rect 16975 6694 16991 6708
rect 17029 6704 17035 6706
rect 17042 6704 17150 6720
rect 17157 6704 17163 6706
rect 17171 6704 17186 6720
rect 17252 6714 17271 6717
rect 16893 6692 16991 6694
rect 17018 6692 17186 6704
rect 17201 6694 17217 6708
rect 17252 6695 17274 6714
rect 17284 6708 17300 6709
rect 17283 6706 17300 6708
rect 17284 6701 17300 6706
rect 17274 6694 17280 6695
rect 17283 6694 17312 6701
rect 17201 6693 17312 6694
rect 17201 6692 17318 6693
rect 16877 6684 16928 6692
rect 16975 6684 17009 6692
rect 16877 6672 16902 6684
rect 16909 6672 16928 6684
rect 16982 6682 17009 6684
rect 17018 6682 17239 6692
rect 17274 6689 17280 6692
rect 16982 6678 17239 6682
rect 16877 6664 16928 6672
rect 16975 6664 17239 6678
rect 17283 6684 17318 6692
rect 16829 6616 16848 6650
rect 16893 6656 16922 6664
rect 16893 6650 16910 6656
rect 16893 6648 16927 6650
rect 16975 6648 16991 6664
rect 16992 6654 17200 6664
rect 17201 6654 17217 6664
rect 17265 6660 17280 6675
rect 17283 6672 17284 6684
rect 17291 6672 17318 6684
rect 17283 6664 17318 6672
rect 17283 6663 17312 6664
rect 17003 6650 17217 6654
rect 17018 6648 17217 6650
rect 17252 6650 17265 6660
rect 17283 6650 17300 6663
rect 17252 6648 17300 6650
rect 16894 6644 16927 6648
rect 16890 6642 16927 6644
rect 16890 6641 16957 6642
rect 16890 6636 16921 6641
rect 16927 6636 16957 6641
rect 16890 6632 16957 6636
rect 16863 6629 16957 6632
rect 16863 6622 16912 6629
rect 16863 6616 16893 6622
rect 16912 6617 16917 6622
rect 16829 6600 16909 6616
rect 16921 6608 16957 6629
rect 17018 6624 17207 6648
rect 17252 6647 17299 6648
rect 17265 6642 17299 6647
rect 17033 6621 17207 6624
rect 17026 6618 17207 6621
rect 17235 6641 17299 6642
rect 16829 6598 16848 6600
rect 16863 6598 16897 6600
rect 16829 6582 16909 6598
rect 16829 6576 16848 6582
rect 16545 6550 16648 6560
rect 16499 6548 16648 6550
rect 16669 6548 16704 6560
rect 16338 6546 16500 6548
rect 16350 6526 16369 6546
rect 16384 6544 16414 6546
rect 16233 6518 16274 6526
rect 16356 6522 16369 6526
rect 16421 6530 16500 6546
rect 16532 6546 16704 6548
rect 16532 6530 16611 6546
rect 16618 6544 16648 6546
rect 16196 6508 16225 6518
rect 16239 6508 16268 6518
rect 16283 6508 16313 6522
rect 16356 6508 16399 6522
rect 16421 6518 16611 6530
rect 16676 6526 16682 6546
rect 16406 6508 16436 6518
rect 16437 6508 16595 6518
rect 16599 6508 16629 6518
rect 16633 6508 16663 6522
rect 16691 6508 16704 6546
rect 16776 6560 16805 6576
rect 16819 6560 16848 6576
rect 16863 6566 16893 6582
rect 16921 6560 16927 6608
rect 16930 6602 16949 6608
rect 16964 6602 16994 6610
rect 16930 6594 16994 6602
rect 16930 6578 17010 6594
rect 17026 6587 17088 6618
rect 17104 6587 17166 6618
rect 17235 6616 17284 6641
rect 17299 6616 17329 6632
rect 17198 6602 17228 6610
rect 17235 6608 17345 6616
rect 17198 6594 17243 6602
rect 16930 6576 16949 6578
rect 16964 6576 17010 6578
rect 16930 6560 17010 6576
rect 17037 6574 17072 6587
rect 17113 6584 17150 6587
rect 17113 6582 17155 6584
rect 17042 6571 17072 6574
rect 17051 6567 17058 6571
rect 17058 6566 17059 6567
rect 17017 6560 17027 6566
rect 16776 6552 16811 6560
rect 16776 6526 16777 6552
rect 16784 6526 16811 6552
rect 16719 6508 16749 6522
rect 16776 6518 16811 6526
rect 16813 6552 16854 6560
rect 16813 6526 16828 6552
rect 16835 6526 16854 6552
rect 16918 6548 16949 6560
rect 16964 6548 17067 6560
rect 17079 6550 17105 6576
rect 17120 6571 17150 6582
rect 17182 6578 17244 6594
rect 17182 6576 17228 6578
rect 17182 6560 17244 6576
rect 17256 6560 17262 6608
rect 17265 6600 17345 6608
rect 17265 6598 17284 6600
rect 17299 6598 17333 6600
rect 17265 6582 17345 6598
rect 17265 6560 17284 6582
rect 17299 6566 17329 6582
rect 17357 6576 17363 6650
rect 17366 6576 17385 6720
rect 17400 6576 17406 6720
rect 17415 6650 17428 6720
rect 17480 6716 17502 6720
rect 17473 6694 17502 6708
rect 17555 6694 17571 6708
rect 17609 6704 17615 6706
rect 17622 6704 17730 6720
rect 17737 6704 17743 6706
rect 17751 6704 17766 6720
rect 17832 6714 17851 6717
rect 17473 6692 17571 6694
rect 17598 6692 17766 6704
rect 17781 6694 17797 6708
rect 17832 6695 17854 6714
rect 17864 6708 17880 6709
rect 17863 6706 17880 6708
rect 17864 6701 17880 6706
rect 17854 6694 17860 6695
rect 17863 6694 17892 6701
rect 17781 6693 17892 6694
rect 17781 6692 17898 6693
rect 17457 6684 17508 6692
rect 17555 6684 17589 6692
rect 17457 6672 17482 6684
rect 17489 6672 17508 6684
rect 17562 6682 17589 6684
rect 17598 6682 17819 6692
rect 17854 6689 17860 6692
rect 17562 6678 17819 6682
rect 17457 6664 17508 6672
rect 17555 6664 17819 6678
rect 17863 6684 17898 6692
rect 17409 6616 17428 6650
rect 17473 6656 17502 6664
rect 17473 6650 17490 6656
rect 17473 6648 17507 6650
rect 17555 6648 17571 6664
rect 17572 6654 17780 6664
rect 17781 6654 17797 6664
rect 17845 6660 17860 6675
rect 17863 6672 17864 6684
rect 17871 6672 17898 6684
rect 17863 6664 17898 6672
rect 17863 6663 17892 6664
rect 17583 6650 17797 6654
rect 17598 6648 17797 6650
rect 17832 6650 17845 6660
rect 17863 6650 17880 6663
rect 17832 6648 17880 6650
rect 17474 6644 17507 6648
rect 17470 6642 17507 6644
rect 17470 6641 17537 6642
rect 17470 6636 17501 6641
rect 17507 6636 17537 6641
rect 17470 6632 17537 6636
rect 17443 6629 17537 6632
rect 17443 6622 17492 6629
rect 17443 6616 17473 6622
rect 17492 6617 17497 6622
rect 17409 6600 17489 6616
rect 17501 6608 17537 6629
rect 17598 6624 17787 6648
rect 17832 6647 17879 6648
rect 17845 6642 17879 6647
rect 17613 6621 17787 6624
rect 17606 6618 17787 6621
rect 17815 6641 17879 6642
rect 17409 6598 17428 6600
rect 17443 6598 17477 6600
rect 17409 6582 17489 6598
rect 17409 6576 17428 6582
rect 17125 6550 17228 6560
rect 17079 6548 17228 6550
rect 17249 6548 17284 6560
rect 16918 6546 17080 6548
rect 16930 6526 16949 6546
rect 16964 6544 16994 6546
rect 16813 6518 16854 6526
rect 16936 6522 16949 6526
rect 17001 6530 17080 6546
rect 17112 6546 17284 6548
rect 17112 6530 17191 6546
rect 17198 6544 17228 6546
rect 16776 6508 16805 6518
rect 16819 6508 16848 6518
rect 16863 6508 16893 6522
rect 16936 6508 16979 6522
rect 17001 6518 17191 6530
rect 17256 6526 17262 6546
rect 16986 6508 17016 6518
rect 17017 6508 17175 6518
rect 17179 6508 17209 6518
rect 17213 6508 17243 6522
rect 17271 6508 17284 6546
rect 17356 6560 17385 6576
rect 17399 6560 17428 6576
rect 17443 6566 17473 6582
rect 17501 6560 17507 6608
rect 17510 6602 17529 6608
rect 17544 6602 17574 6610
rect 17510 6594 17574 6602
rect 17510 6578 17590 6594
rect 17606 6587 17668 6618
rect 17684 6587 17746 6618
rect 17815 6616 17864 6641
rect 17879 6616 17909 6632
rect 17778 6602 17808 6610
rect 17815 6608 17925 6616
rect 17778 6594 17823 6602
rect 17510 6576 17529 6578
rect 17544 6576 17590 6578
rect 17510 6560 17590 6576
rect 17617 6574 17652 6587
rect 17693 6584 17730 6587
rect 17693 6582 17735 6584
rect 17622 6571 17652 6574
rect 17631 6567 17638 6571
rect 17638 6566 17639 6567
rect 17597 6560 17607 6566
rect 17356 6552 17391 6560
rect 17356 6526 17357 6552
rect 17364 6526 17391 6552
rect 17299 6508 17329 6522
rect 17356 6518 17391 6526
rect 17393 6552 17434 6560
rect 17393 6526 17408 6552
rect 17415 6526 17434 6552
rect 17498 6548 17529 6560
rect 17544 6548 17647 6560
rect 17659 6550 17685 6576
rect 17700 6571 17730 6582
rect 17762 6578 17824 6594
rect 17762 6576 17808 6578
rect 17762 6560 17824 6576
rect 17836 6560 17842 6608
rect 17845 6600 17925 6608
rect 17845 6598 17864 6600
rect 17879 6598 17913 6600
rect 17845 6582 17925 6598
rect 17845 6560 17864 6582
rect 17879 6566 17909 6582
rect 17937 6576 17943 6650
rect 17946 6576 17965 6720
rect 17980 6576 17986 6720
rect 17995 6650 18008 6720
rect 18060 6716 18082 6720
rect 18053 6694 18082 6708
rect 18135 6694 18151 6708
rect 18189 6704 18195 6706
rect 18202 6704 18310 6720
rect 18317 6704 18323 6706
rect 18331 6704 18346 6720
rect 18412 6714 18431 6717
rect 18053 6692 18151 6694
rect 18178 6692 18346 6704
rect 18361 6694 18377 6708
rect 18412 6695 18434 6714
rect 18444 6708 18460 6709
rect 18443 6706 18460 6708
rect 18444 6701 18460 6706
rect 18434 6694 18440 6695
rect 18443 6694 18472 6701
rect 18361 6693 18472 6694
rect 18361 6692 18478 6693
rect 18037 6684 18088 6692
rect 18135 6684 18169 6692
rect 18037 6672 18062 6684
rect 18069 6672 18088 6684
rect 18142 6682 18169 6684
rect 18178 6682 18399 6692
rect 18434 6689 18440 6692
rect 18142 6678 18399 6682
rect 18037 6664 18088 6672
rect 18135 6664 18399 6678
rect 18443 6684 18478 6692
rect 17989 6616 18008 6650
rect 18053 6656 18082 6664
rect 18053 6650 18070 6656
rect 18053 6648 18087 6650
rect 18135 6648 18151 6664
rect 18152 6654 18360 6664
rect 18361 6654 18377 6664
rect 18425 6660 18440 6675
rect 18443 6672 18444 6684
rect 18451 6672 18478 6684
rect 18443 6664 18478 6672
rect 18443 6663 18472 6664
rect 18163 6650 18377 6654
rect 18178 6648 18377 6650
rect 18412 6650 18425 6660
rect 18443 6650 18460 6663
rect 18412 6648 18460 6650
rect 18054 6644 18087 6648
rect 18050 6642 18087 6644
rect 18050 6641 18117 6642
rect 18050 6636 18081 6641
rect 18087 6636 18117 6641
rect 18050 6632 18117 6636
rect 18023 6629 18117 6632
rect 18023 6622 18072 6629
rect 18023 6616 18053 6622
rect 18072 6617 18077 6622
rect 17989 6600 18069 6616
rect 18081 6608 18117 6629
rect 18178 6624 18367 6648
rect 18412 6647 18459 6648
rect 18425 6642 18459 6647
rect 18193 6621 18367 6624
rect 18186 6618 18367 6621
rect 18395 6641 18459 6642
rect 17989 6598 18008 6600
rect 18023 6598 18057 6600
rect 17989 6582 18069 6598
rect 17989 6576 18008 6582
rect 17705 6550 17808 6560
rect 17659 6548 17808 6550
rect 17829 6548 17864 6560
rect 17498 6546 17660 6548
rect 17510 6526 17529 6546
rect 17544 6544 17574 6546
rect 17393 6518 17434 6526
rect 17516 6522 17529 6526
rect 17581 6530 17660 6546
rect 17692 6546 17864 6548
rect 17692 6530 17771 6546
rect 17778 6544 17808 6546
rect 17356 6508 17385 6518
rect 17399 6508 17428 6518
rect 17443 6508 17473 6522
rect 17516 6508 17559 6522
rect 17581 6518 17771 6530
rect 17836 6526 17842 6546
rect 17566 6508 17596 6518
rect 17597 6508 17755 6518
rect 17759 6508 17789 6518
rect 17793 6508 17823 6522
rect 17851 6508 17864 6546
rect 17936 6560 17965 6576
rect 17979 6560 18008 6576
rect 18023 6566 18053 6582
rect 18081 6560 18087 6608
rect 18090 6602 18109 6608
rect 18124 6602 18154 6610
rect 18090 6594 18154 6602
rect 18090 6578 18170 6594
rect 18186 6587 18248 6618
rect 18264 6587 18326 6618
rect 18395 6616 18444 6641
rect 18459 6616 18489 6632
rect 18358 6602 18388 6610
rect 18395 6608 18505 6616
rect 18358 6594 18403 6602
rect 18090 6576 18109 6578
rect 18124 6576 18170 6578
rect 18090 6560 18170 6576
rect 18197 6574 18232 6587
rect 18273 6584 18310 6587
rect 18273 6582 18315 6584
rect 18202 6571 18232 6574
rect 18211 6567 18218 6571
rect 18218 6566 18219 6567
rect 18177 6560 18187 6566
rect 17936 6552 17971 6560
rect 17936 6526 17937 6552
rect 17944 6526 17971 6552
rect 17879 6508 17909 6522
rect 17936 6518 17971 6526
rect 17973 6552 18014 6560
rect 17973 6526 17988 6552
rect 17995 6526 18014 6552
rect 18078 6548 18109 6560
rect 18124 6548 18227 6560
rect 18239 6550 18265 6576
rect 18280 6571 18310 6582
rect 18342 6578 18404 6594
rect 18342 6576 18388 6578
rect 18342 6560 18404 6576
rect 18416 6560 18422 6608
rect 18425 6600 18505 6608
rect 18425 6598 18444 6600
rect 18459 6598 18493 6600
rect 18425 6582 18505 6598
rect 18425 6560 18444 6582
rect 18459 6566 18489 6582
rect 18517 6576 18523 6650
rect 18532 6576 18545 6720
rect 18285 6550 18388 6560
rect 18239 6548 18388 6550
rect 18409 6548 18444 6560
rect 18078 6546 18240 6548
rect 18090 6526 18109 6546
rect 18124 6544 18154 6546
rect 17973 6518 18014 6526
rect 18096 6522 18109 6526
rect 18161 6530 18240 6546
rect 18272 6546 18444 6548
rect 18272 6530 18351 6546
rect 18358 6544 18388 6546
rect 17936 6508 17965 6518
rect 17979 6508 18008 6518
rect 18023 6508 18053 6522
rect 18096 6508 18139 6522
rect 18161 6518 18351 6530
rect 18416 6526 18422 6546
rect 18146 6508 18176 6518
rect 18177 6508 18335 6518
rect 18339 6508 18369 6518
rect 18373 6508 18403 6522
rect 18431 6508 18444 6546
rect 18516 6560 18545 6576
rect 18516 6552 18551 6560
rect 18516 6526 18517 6552
rect 18524 6526 18551 6552
rect 18459 6508 18489 6522
rect 18516 6518 18551 6526
rect 18516 6508 18545 6518
rect -1 6502 18545 6508
rect 0 6494 18545 6502
rect 15 6464 28 6494
rect 43 6480 73 6494
rect 116 6480 159 6494
rect 166 6480 386 6494
rect 393 6480 423 6494
rect 83 6466 98 6478
rect 117 6466 130 6480
rect 198 6476 351 6480
rect 80 6464 102 6466
rect 180 6464 372 6476
rect 451 6464 464 6494
rect 479 6480 509 6494
rect 546 6464 565 6494
rect 580 6464 586 6494
rect 595 6464 608 6494
rect 623 6480 653 6494
rect 696 6480 739 6494
rect 746 6480 966 6494
rect 973 6480 1003 6494
rect 663 6466 678 6478
rect 697 6466 710 6480
rect 778 6476 931 6480
rect 660 6464 682 6466
rect 760 6464 952 6476
rect 1031 6464 1044 6494
rect 1059 6480 1089 6494
rect 1126 6464 1145 6494
rect 1160 6464 1166 6494
rect 1175 6464 1188 6494
rect 1203 6480 1233 6494
rect 1276 6480 1319 6494
rect 1326 6480 1546 6494
rect 1553 6480 1583 6494
rect 1243 6466 1258 6478
rect 1277 6466 1290 6480
rect 1358 6476 1511 6480
rect 1240 6464 1262 6466
rect 1340 6464 1532 6476
rect 1611 6464 1624 6494
rect 1639 6480 1669 6494
rect 1706 6464 1725 6494
rect 1740 6464 1746 6494
rect 1755 6464 1768 6494
rect 1783 6480 1813 6494
rect 1856 6480 1899 6494
rect 1906 6480 2126 6494
rect 2133 6480 2163 6494
rect 1823 6466 1838 6478
rect 1857 6466 1870 6480
rect 1938 6476 2091 6480
rect 1820 6464 1842 6466
rect 1920 6464 2112 6476
rect 2191 6464 2204 6494
rect 2219 6480 2249 6494
rect 2286 6464 2305 6494
rect 2320 6464 2326 6494
rect 2335 6464 2348 6494
rect 2363 6480 2393 6494
rect 2436 6480 2479 6494
rect 2486 6480 2706 6494
rect 2713 6480 2743 6494
rect 2403 6466 2418 6478
rect 2437 6466 2450 6480
rect 2518 6476 2671 6480
rect 2400 6464 2422 6466
rect 2500 6464 2692 6476
rect 2771 6464 2784 6494
rect 2799 6480 2829 6494
rect 2866 6464 2885 6494
rect 2900 6464 2906 6494
rect 2915 6464 2928 6494
rect 2943 6480 2973 6494
rect 3016 6480 3059 6494
rect 3066 6480 3286 6494
rect 3293 6480 3323 6494
rect 2983 6466 2998 6478
rect 3017 6466 3030 6480
rect 3098 6476 3251 6480
rect 2980 6464 3002 6466
rect 3080 6464 3272 6476
rect 3351 6464 3364 6494
rect 3379 6480 3409 6494
rect 3446 6464 3465 6494
rect 3480 6464 3486 6494
rect 3495 6464 3508 6494
rect 3523 6480 3553 6494
rect 3596 6480 3639 6494
rect 3646 6480 3866 6494
rect 3873 6480 3903 6494
rect 3563 6466 3578 6478
rect 3597 6466 3610 6480
rect 3678 6476 3831 6480
rect 3560 6464 3582 6466
rect 3660 6464 3852 6476
rect 3931 6464 3944 6494
rect 3959 6480 3989 6494
rect 4026 6464 4045 6494
rect 4060 6464 4066 6494
rect 4075 6464 4088 6494
rect 4103 6480 4133 6494
rect 4176 6480 4219 6494
rect 4226 6480 4446 6494
rect 4453 6480 4483 6494
rect 4143 6466 4158 6478
rect 4177 6466 4190 6480
rect 4258 6476 4411 6480
rect 4140 6464 4162 6466
rect 4240 6464 4432 6476
rect 4511 6464 4524 6494
rect 4539 6480 4569 6494
rect 4606 6464 4625 6494
rect 4640 6464 4646 6494
rect 4655 6464 4668 6494
rect 4683 6480 4713 6494
rect 4756 6480 4799 6494
rect 4806 6480 5026 6494
rect 5033 6480 5063 6494
rect 4723 6466 4738 6478
rect 4757 6466 4770 6480
rect 4838 6476 4991 6480
rect 4720 6464 4742 6466
rect 4820 6464 5012 6476
rect 5091 6464 5104 6494
rect 5119 6480 5149 6494
rect 5186 6464 5205 6494
rect 5220 6464 5226 6494
rect 5235 6464 5248 6494
rect 5263 6480 5293 6494
rect 5336 6480 5379 6494
rect 5386 6480 5606 6494
rect 5613 6480 5643 6494
rect 5303 6466 5318 6478
rect 5337 6466 5350 6480
rect 5418 6476 5571 6480
rect 5300 6464 5322 6466
rect 5400 6464 5592 6476
rect 5671 6464 5684 6494
rect 5699 6480 5729 6494
rect 5766 6464 5785 6494
rect 5800 6464 5806 6494
rect 5815 6464 5828 6494
rect 5843 6480 5873 6494
rect 5916 6480 5959 6494
rect 5966 6480 6186 6494
rect 6193 6480 6223 6494
rect 5883 6466 5898 6478
rect 5917 6466 5930 6480
rect 5998 6476 6151 6480
rect 5880 6464 5902 6466
rect 5980 6464 6172 6476
rect 6251 6464 6264 6494
rect 6279 6480 6309 6494
rect 6346 6464 6365 6494
rect 6380 6464 6386 6494
rect 6395 6464 6408 6494
rect 6423 6480 6453 6494
rect 6496 6480 6539 6494
rect 6546 6480 6766 6494
rect 6773 6480 6803 6494
rect 6463 6466 6478 6478
rect 6497 6466 6510 6480
rect 6578 6476 6731 6480
rect 6460 6464 6482 6466
rect 6560 6464 6752 6476
rect 6831 6464 6844 6494
rect 6859 6480 6889 6494
rect 6926 6464 6945 6494
rect 6960 6464 6966 6494
rect 6975 6464 6988 6494
rect 7003 6480 7033 6494
rect 7076 6480 7119 6494
rect 7126 6480 7346 6494
rect 7353 6480 7383 6494
rect 7043 6466 7058 6478
rect 7077 6466 7090 6480
rect 7158 6476 7311 6480
rect 7040 6464 7062 6466
rect 7140 6464 7332 6476
rect 7411 6464 7424 6494
rect 7439 6480 7469 6494
rect 7506 6464 7525 6494
rect 7540 6464 7546 6494
rect 7555 6464 7568 6494
rect 7583 6480 7613 6494
rect 7656 6480 7699 6494
rect 7706 6480 7926 6494
rect 7933 6480 7963 6494
rect 7623 6466 7638 6478
rect 7657 6466 7670 6480
rect 7738 6476 7891 6480
rect 7620 6464 7642 6466
rect 7720 6464 7912 6476
rect 7991 6464 8004 6494
rect 8019 6480 8049 6494
rect 8086 6464 8105 6494
rect 8120 6464 8126 6494
rect 8135 6464 8148 6494
rect 8163 6480 8193 6494
rect 8236 6480 8279 6494
rect 8286 6480 8506 6494
rect 8513 6480 8543 6494
rect 8203 6466 8218 6478
rect 8237 6466 8250 6480
rect 8318 6476 8471 6480
rect 8200 6464 8222 6466
rect 8300 6464 8492 6476
rect 8571 6464 8584 6494
rect 8599 6480 8629 6494
rect 8666 6464 8685 6494
rect 8700 6464 8706 6494
rect 8715 6464 8728 6494
rect 8743 6480 8773 6494
rect 8816 6480 8859 6494
rect 8866 6480 9086 6494
rect 9093 6480 9123 6494
rect 8783 6466 8798 6478
rect 8817 6466 8830 6480
rect 8898 6476 9051 6480
rect 8780 6464 8802 6466
rect 8880 6464 9072 6476
rect 9151 6464 9164 6494
rect 9179 6480 9209 6494
rect 9246 6464 9265 6494
rect 9280 6464 9286 6494
rect 9295 6464 9308 6494
rect 9323 6480 9353 6494
rect 9396 6480 9439 6494
rect 9446 6480 9666 6494
rect 9673 6480 9703 6494
rect 9363 6466 9378 6478
rect 9397 6466 9410 6480
rect 9478 6476 9631 6480
rect 9360 6464 9382 6466
rect 9460 6464 9652 6476
rect 9731 6464 9744 6494
rect 9759 6480 9789 6494
rect 9826 6464 9845 6494
rect 9860 6464 9866 6494
rect 9875 6464 9888 6494
rect 9903 6480 9933 6494
rect 9976 6480 10019 6494
rect 10026 6480 10246 6494
rect 10253 6480 10283 6494
rect 9943 6466 9958 6478
rect 9977 6466 9990 6480
rect 10058 6476 10211 6480
rect 9940 6464 9962 6466
rect 10040 6464 10232 6476
rect 10311 6464 10324 6494
rect 10339 6480 10369 6494
rect 10406 6464 10425 6494
rect 10440 6464 10446 6494
rect 10455 6464 10468 6494
rect 10483 6480 10513 6494
rect 10556 6480 10599 6494
rect 10606 6480 10826 6494
rect 10833 6480 10863 6494
rect 10523 6466 10538 6478
rect 10557 6466 10570 6480
rect 10638 6476 10791 6480
rect 10520 6464 10542 6466
rect 10620 6464 10812 6476
rect 10891 6464 10904 6494
rect 10919 6480 10949 6494
rect 10986 6464 11005 6494
rect 11020 6464 11026 6494
rect 11035 6464 11048 6494
rect 11063 6480 11093 6494
rect 11136 6480 11179 6494
rect 11186 6480 11406 6494
rect 11413 6480 11443 6494
rect 11103 6466 11118 6478
rect 11137 6466 11150 6480
rect 11218 6476 11371 6480
rect 11100 6464 11122 6466
rect 11200 6464 11392 6476
rect 11471 6464 11484 6494
rect 11499 6480 11529 6494
rect 11566 6464 11585 6494
rect 11600 6464 11606 6494
rect 11615 6464 11628 6494
rect 11643 6480 11673 6494
rect 11716 6480 11759 6494
rect 11766 6480 11986 6494
rect 11993 6480 12023 6494
rect 11683 6466 11698 6478
rect 11717 6466 11730 6480
rect 11798 6476 11951 6480
rect 11680 6464 11702 6466
rect 11780 6464 11972 6476
rect 12051 6464 12064 6494
rect 12079 6480 12109 6494
rect 12146 6464 12165 6494
rect 12180 6464 12186 6494
rect 12195 6464 12208 6494
rect 12223 6480 12253 6494
rect 12296 6480 12339 6494
rect 12346 6480 12566 6494
rect 12573 6480 12603 6494
rect 12263 6466 12278 6478
rect 12297 6466 12310 6480
rect 12378 6476 12531 6480
rect 12260 6464 12282 6466
rect 12360 6464 12552 6476
rect 12631 6464 12644 6494
rect 12659 6480 12689 6494
rect 12726 6464 12745 6494
rect 12760 6464 12766 6494
rect 12775 6464 12788 6494
rect 12803 6480 12833 6494
rect 12876 6480 12919 6494
rect 12926 6480 13146 6494
rect 13153 6480 13183 6494
rect 12843 6466 12858 6478
rect 12877 6466 12890 6480
rect 12958 6476 13111 6480
rect 12840 6464 12862 6466
rect 12940 6464 13132 6476
rect 13211 6464 13224 6494
rect 13239 6480 13269 6494
rect 13306 6464 13325 6494
rect 13340 6464 13346 6494
rect 13355 6464 13368 6494
rect 13383 6480 13413 6494
rect 13456 6480 13499 6494
rect 13506 6480 13726 6494
rect 13733 6480 13763 6494
rect 13423 6466 13438 6478
rect 13457 6466 13470 6480
rect 13538 6476 13691 6480
rect 13420 6464 13442 6466
rect 13520 6464 13712 6476
rect 13791 6464 13804 6494
rect 13819 6480 13849 6494
rect 13886 6464 13905 6494
rect 13920 6464 13926 6494
rect 13935 6464 13948 6494
rect 13963 6480 13993 6494
rect 14036 6480 14079 6494
rect 14086 6480 14306 6494
rect 14313 6480 14343 6494
rect 14003 6466 14018 6478
rect 14037 6466 14050 6480
rect 14118 6476 14271 6480
rect 14000 6464 14022 6466
rect 14100 6464 14292 6476
rect 14371 6464 14384 6494
rect 14399 6480 14429 6494
rect 14466 6464 14485 6494
rect 14500 6464 14506 6494
rect 14515 6464 14528 6494
rect 14543 6480 14573 6494
rect 14616 6480 14659 6494
rect 14666 6480 14886 6494
rect 14893 6480 14923 6494
rect 14583 6466 14598 6478
rect 14617 6466 14630 6480
rect 14698 6476 14851 6480
rect 14580 6464 14602 6466
rect 14680 6464 14872 6476
rect 14951 6464 14964 6494
rect 14979 6480 15009 6494
rect 15046 6464 15065 6494
rect 15080 6464 15086 6494
rect 15095 6464 15108 6494
rect 15123 6480 15153 6494
rect 15196 6480 15239 6494
rect 15246 6480 15466 6494
rect 15473 6480 15503 6494
rect 15163 6466 15178 6478
rect 15197 6466 15210 6480
rect 15278 6476 15431 6480
rect 15160 6464 15182 6466
rect 15260 6464 15452 6476
rect 15531 6464 15544 6494
rect 15559 6480 15589 6494
rect 15626 6464 15645 6494
rect 15660 6464 15666 6494
rect 15675 6464 15688 6494
rect 15703 6480 15733 6494
rect 15776 6480 15819 6494
rect 15826 6480 16046 6494
rect 16053 6480 16083 6494
rect 15743 6466 15758 6478
rect 15777 6466 15790 6480
rect 15858 6476 16011 6480
rect 15740 6464 15762 6466
rect 15840 6464 16032 6476
rect 16111 6464 16124 6494
rect 16139 6480 16169 6494
rect 16206 6464 16225 6494
rect 16240 6464 16246 6494
rect 16255 6464 16268 6494
rect 16283 6480 16313 6494
rect 16356 6480 16399 6494
rect 16406 6480 16626 6494
rect 16633 6480 16663 6494
rect 16323 6466 16338 6478
rect 16357 6466 16370 6480
rect 16438 6476 16591 6480
rect 16320 6464 16342 6466
rect 16420 6464 16612 6476
rect 16691 6464 16704 6494
rect 16719 6480 16749 6494
rect 16786 6464 16805 6494
rect 16820 6464 16826 6494
rect 16835 6464 16848 6494
rect 16863 6480 16893 6494
rect 16936 6480 16979 6494
rect 16986 6480 17206 6494
rect 17213 6480 17243 6494
rect 16903 6466 16918 6478
rect 16937 6466 16950 6480
rect 17018 6476 17171 6480
rect 16900 6464 16922 6466
rect 17000 6464 17192 6476
rect 17271 6464 17284 6494
rect 17299 6480 17329 6494
rect 17366 6464 17385 6494
rect 17400 6464 17406 6494
rect 17415 6464 17428 6494
rect 17443 6480 17473 6494
rect 17516 6480 17559 6494
rect 17566 6480 17786 6494
rect 17793 6480 17823 6494
rect 17483 6466 17498 6478
rect 17517 6466 17530 6480
rect 17598 6476 17751 6480
rect 17480 6464 17502 6466
rect 17580 6464 17772 6476
rect 17851 6464 17864 6494
rect 17879 6480 17909 6494
rect 17946 6464 17965 6494
rect 17980 6464 17986 6494
rect 17995 6464 18008 6494
rect 18023 6480 18053 6494
rect 18096 6480 18139 6494
rect 18146 6480 18366 6494
rect 18373 6480 18403 6494
rect 18063 6466 18078 6478
rect 18097 6466 18110 6480
rect 18178 6476 18331 6480
rect 18060 6464 18082 6466
rect 18160 6464 18352 6476
rect 18431 6464 18444 6494
rect 18459 6480 18489 6494
rect 18532 6464 18545 6494
rect 0 6450 18545 6464
rect 15 6380 28 6450
rect 80 6446 102 6450
rect 73 6424 102 6438
rect 155 6424 171 6438
rect 209 6434 215 6436
rect 222 6434 330 6450
rect 337 6434 343 6436
rect 351 6434 366 6450
rect 432 6444 451 6447
rect 73 6422 171 6424
rect 198 6422 366 6434
rect 381 6424 397 6438
rect 432 6425 454 6444
rect 464 6438 480 6439
rect 463 6436 480 6438
rect 464 6431 480 6436
rect 454 6424 460 6425
rect 463 6424 492 6431
rect 381 6423 492 6424
rect 381 6422 498 6423
rect 57 6414 108 6422
rect 155 6414 189 6422
rect 57 6402 82 6414
rect 89 6402 108 6414
rect 162 6412 189 6414
rect 198 6412 419 6422
rect 454 6419 460 6422
rect 162 6408 419 6412
rect 57 6394 108 6402
rect 155 6394 419 6408
rect 463 6414 498 6422
rect 9 6346 28 6380
rect 73 6386 102 6394
rect 73 6380 90 6386
rect 73 6378 107 6380
rect 155 6378 171 6394
rect 172 6384 380 6394
rect 381 6384 397 6394
rect 445 6390 460 6405
rect 463 6402 464 6414
rect 471 6402 498 6414
rect 463 6394 498 6402
rect 463 6393 492 6394
rect 183 6380 397 6384
rect 198 6378 397 6380
rect 432 6380 445 6390
rect 463 6380 480 6393
rect 432 6378 480 6380
rect 74 6374 107 6378
rect 70 6372 107 6374
rect 70 6371 137 6372
rect 70 6366 101 6371
rect 107 6366 137 6371
rect 70 6362 137 6366
rect 43 6359 137 6362
rect 43 6352 92 6359
rect 43 6346 73 6352
rect 92 6347 97 6352
rect 9 6330 89 6346
rect 101 6338 137 6359
rect 198 6354 387 6378
rect 432 6377 479 6378
rect 445 6372 479 6377
rect 213 6351 387 6354
rect 206 6348 387 6351
rect 415 6371 479 6372
rect 9 6328 28 6330
rect 43 6328 77 6330
rect 9 6312 89 6328
rect 9 6306 28 6312
rect -1 6290 28 6306
rect 43 6296 73 6312
rect 101 6290 107 6338
rect 110 6332 129 6338
rect 144 6332 174 6340
rect 110 6324 174 6332
rect 110 6308 190 6324
rect 206 6317 268 6348
rect 284 6317 346 6348
rect 415 6346 464 6371
rect 479 6346 509 6362
rect 378 6332 408 6340
rect 415 6338 525 6346
rect 378 6324 423 6332
rect 110 6306 129 6308
rect 144 6306 190 6308
rect 110 6290 190 6306
rect 217 6304 252 6317
rect 293 6314 330 6317
rect 293 6312 335 6314
rect 222 6301 252 6304
rect 231 6297 238 6301
rect 238 6296 239 6297
rect 197 6290 207 6296
rect -7 6282 34 6290
rect -7 6256 8 6282
rect 15 6256 34 6282
rect 98 6278 129 6290
rect 144 6278 247 6290
rect 259 6280 285 6306
rect 300 6301 330 6312
rect 362 6308 424 6324
rect 362 6306 408 6308
rect 362 6290 424 6306
rect 436 6290 442 6338
rect 445 6330 525 6338
rect 445 6328 464 6330
rect 479 6328 513 6330
rect 445 6312 525 6328
rect 445 6290 464 6312
rect 479 6296 509 6312
rect 537 6306 543 6380
rect 546 6306 565 6450
rect 580 6306 586 6450
rect 595 6380 608 6450
rect 660 6446 682 6450
rect 653 6424 682 6438
rect 735 6424 751 6438
rect 789 6434 795 6436
rect 802 6434 910 6450
rect 917 6434 923 6436
rect 931 6434 946 6450
rect 1012 6444 1031 6447
rect 653 6422 751 6424
rect 778 6422 946 6434
rect 961 6424 977 6438
rect 1012 6425 1034 6444
rect 1044 6438 1060 6439
rect 1043 6436 1060 6438
rect 1044 6431 1060 6436
rect 1034 6424 1040 6425
rect 1043 6424 1072 6431
rect 961 6423 1072 6424
rect 961 6422 1078 6423
rect 637 6414 688 6422
rect 735 6414 769 6422
rect 637 6402 662 6414
rect 669 6402 688 6414
rect 742 6412 769 6414
rect 778 6412 999 6422
rect 1034 6419 1040 6422
rect 742 6408 999 6412
rect 637 6394 688 6402
rect 735 6394 999 6408
rect 1043 6414 1078 6422
rect 589 6346 608 6380
rect 653 6386 682 6394
rect 653 6380 670 6386
rect 653 6378 687 6380
rect 735 6378 751 6394
rect 752 6384 960 6394
rect 961 6384 977 6394
rect 1025 6390 1040 6405
rect 1043 6402 1044 6414
rect 1051 6402 1078 6414
rect 1043 6394 1078 6402
rect 1043 6393 1072 6394
rect 763 6380 977 6384
rect 778 6378 977 6380
rect 1012 6380 1025 6390
rect 1043 6380 1060 6393
rect 1012 6378 1060 6380
rect 654 6374 687 6378
rect 650 6372 687 6374
rect 650 6371 717 6372
rect 650 6366 681 6371
rect 687 6366 717 6371
rect 650 6362 717 6366
rect 623 6359 717 6362
rect 623 6352 672 6359
rect 623 6346 653 6352
rect 672 6347 677 6352
rect 589 6330 669 6346
rect 681 6338 717 6359
rect 778 6354 967 6378
rect 1012 6377 1059 6378
rect 1025 6372 1059 6377
rect 793 6351 967 6354
rect 786 6348 967 6351
rect 995 6371 1059 6372
rect 589 6328 608 6330
rect 623 6328 657 6330
rect 589 6312 669 6328
rect 589 6306 608 6312
rect 305 6280 408 6290
rect 259 6278 408 6280
rect 429 6278 464 6290
rect 98 6276 260 6278
rect 110 6256 129 6276
rect 144 6274 174 6276
rect -7 6248 34 6256
rect 116 6252 129 6256
rect 181 6260 260 6276
rect 292 6276 464 6278
rect 292 6260 371 6276
rect 378 6274 408 6276
rect -1 6238 28 6248
rect 43 6238 73 6252
rect 116 6238 159 6252
rect 181 6248 371 6260
rect 436 6256 442 6276
rect 166 6238 196 6248
rect 197 6238 355 6248
rect 359 6238 389 6248
rect 393 6238 423 6252
rect 451 6238 464 6276
rect 536 6290 565 6306
rect 579 6290 608 6306
rect 623 6296 653 6312
rect 681 6290 687 6338
rect 690 6332 709 6338
rect 724 6332 754 6340
rect 690 6324 754 6332
rect 690 6308 770 6324
rect 786 6317 848 6348
rect 864 6317 926 6348
rect 995 6346 1044 6371
rect 1059 6346 1089 6362
rect 958 6332 988 6340
rect 995 6338 1105 6346
rect 958 6324 1003 6332
rect 690 6306 709 6308
rect 724 6306 770 6308
rect 690 6290 770 6306
rect 797 6304 832 6317
rect 873 6314 910 6317
rect 873 6312 915 6314
rect 802 6301 832 6304
rect 811 6297 818 6301
rect 818 6296 819 6297
rect 777 6290 787 6296
rect 536 6282 571 6290
rect 536 6256 537 6282
rect 544 6256 571 6282
rect 479 6238 509 6252
rect 536 6248 571 6256
rect 573 6282 614 6290
rect 573 6256 588 6282
rect 595 6256 614 6282
rect 678 6278 709 6290
rect 724 6278 827 6290
rect 839 6280 865 6306
rect 880 6301 910 6312
rect 942 6308 1004 6324
rect 942 6306 988 6308
rect 942 6290 1004 6306
rect 1016 6290 1022 6338
rect 1025 6330 1105 6338
rect 1025 6328 1044 6330
rect 1059 6328 1093 6330
rect 1025 6312 1105 6328
rect 1025 6290 1044 6312
rect 1059 6296 1089 6312
rect 1117 6306 1123 6380
rect 1126 6306 1145 6450
rect 1160 6306 1166 6450
rect 1175 6380 1188 6450
rect 1240 6446 1262 6450
rect 1233 6424 1262 6438
rect 1315 6424 1331 6438
rect 1369 6434 1375 6436
rect 1382 6434 1490 6450
rect 1497 6434 1503 6436
rect 1511 6434 1526 6450
rect 1592 6444 1611 6447
rect 1233 6422 1331 6424
rect 1358 6422 1526 6434
rect 1541 6424 1557 6438
rect 1592 6425 1614 6444
rect 1624 6438 1640 6439
rect 1623 6436 1640 6438
rect 1624 6431 1640 6436
rect 1614 6424 1620 6425
rect 1623 6424 1652 6431
rect 1541 6423 1652 6424
rect 1541 6422 1658 6423
rect 1217 6414 1268 6422
rect 1315 6414 1349 6422
rect 1217 6402 1242 6414
rect 1249 6402 1268 6414
rect 1322 6412 1349 6414
rect 1358 6412 1579 6422
rect 1614 6419 1620 6422
rect 1322 6408 1579 6412
rect 1217 6394 1268 6402
rect 1315 6394 1579 6408
rect 1623 6414 1658 6422
rect 1169 6346 1188 6380
rect 1233 6386 1262 6394
rect 1233 6380 1250 6386
rect 1233 6378 1267 6380
rect 1315 6378 1331 6394
rect 1332 6384 1540 6394
rect 1541 6384 1557 6394
rect 1605 6390 1620 6405
rect 1623 6402 1624 6414
rect 1631 6402 1658 6414
rect 1623 6394 1658 6402
rect 1623 6393 1652 6394
rect 1343 6380 1557 6384
rect 1358 6378 1557 6380
rect 1592 6380 1605 6390
rect 1623 6380 1640 6393
rect 1592 6378 1640 6380
rect 1234 6374 1267 6378
rect 1230 6372 1267 6374
rect 1230 6371 1297 6372
rect 1230 6366 1261 6371
rect 1267 6366 1297 6371
rect 1230 6362 1297 6366
rect 1203 6359 1297 6362
rect 1203 6352 1252 6359
rect 1203 6346 1233 6352
rect 1252 6347 1257 6352
rect 1169 6330 1249 6346
rect 1261 6338 1297 6359
rect 1358 6354 1547 6378
rect 1592 6377 1639 6378
rect 1605 6372 1639 6377
rect 1373 6351 1547 6354
rect 1366 6348 1547 6351
rect 1575 6371 1639 6372
rect 1169 6328 1188 6330
rect 1203 6328 1237 6330
rect 1169 6312 1249 6328
rect 1169 6306 1188 6312
rect 885 6280 988 6290
rect 839 6278 988 6280
rect 1009 6278 1044 6290
rect 678 6276 840 6278
rect 690 6256 709 6276
rect 724 6274 754 6276
rect 573 6248 614 6256
rect 696 6252 709 6256
rect 761 6260 840 6276
rect 872 6276 1044 6278
rect 872 6260 951 6276
rect 958 6274 988 6276
rect 536 6238 565 6248
rect 579 6238 608 6248
rect 623 6238 653 6252
rect 696 6238 739 6252
rect 761 6248 951 6260
rect 1016 6256 1022 6276
rect 746 6238 776 6248
rect 777 6238 935 6248
rect 939 6238 969 6248
rect 973 6238 1003 6252
rect 1031 6238 1044 6276
rect 1116 6290 1145 6306
rect 1159 6290 1188 6306
rect 1203 6296 1233 6312
rect 1261 6290 1267 6338
rect 1270 6332 1289 6338
rect 1304 6332 1334 6340
rect 1270 6324 1334 6332
rect 1270 6308 1350 6324
rect 1366 6317 1428 6348
rect 1444 6317 1506 6348
rect 1575 6346 1624 6371
rect 1639 6346 1669 6362
rect 1538 6332 1568 6340
rect 1575 6338 1685 6346
rect 1538 6324 1583 6332
rect 1270 6306 1289 6308
rect 1304 6306 1350 6308
rect 1270 6290 1350 6306
rect 1377 6304 1412 6317
rect 1453 6314 1490 6317
rect 1453 6312 1495 6314
rect 1382 6301 1412 6304
rect 1391 6297 1398 6301
rect 1398 6296 1399 6297
rect 1357 6290 1367 6296
rect 1116 6282 1151 6290
rect 1116 6256 1117 6282
rect 1124 6256 1151 6282
rect 1059 6238 1089 6252
rect 1116 6248 1151 6256
rect 1153 6282 1194 6290
rect 1153 6256 1168 6282
rect 1175 6256 1194 6282
rect 1258 6278 1289 6290
rect 1304 6278 1407 6290
rect 1419 6280 1445 6306
rect 1460 6301 1490 6312
rect 1522 6308 1584 6324
rect 1522 6306 1568 6308
rect 1522 6290 1584 6306
rect 1596 6290 1602 6338
rect 1605 6330 1685 6338
rect 1605 6328 1624 6330
rect 1639 6328 1673 6330
rect 1605 6312 1685 6328
rect 1605 6290 1624 6312
rect 1639 6296 1669 6312
rect 1697 6306 1703 6380
rect 1706 6306 1725 6450
rect 1740 6306 1746 6450
rect 1755 6380 1768 6450
rect 1820 6446 1842 6450
rect 1813 6424 1842 6438
rect 1895 6424 1911 6438
rect 1949 6434 1955 6436
rect 1962 6434 2070 6450
rect 2077 6434 2083 6436
rect 2091 6434 2106 6450
rect 2172 6444 2191 6447
rect 1813 6422 1911 6424
rect 1938 6422 2106 6434
rect 2121 6424 2137 6438
rect 2172 6425 2194 6444
rect 2204 6438 2220 6439
rect 2203 6436 2220 6438
rect 2204 6431 2220 6436
rect 2194 6424 2200 6425
rect 2203 6424 2232 6431
rect 2121 6423 2232 6424
rect 2121 6422 2238 6423
rect 1797 6414 1848 6422
rect 1895 6414 1929 6422
rect 1797 6402 1822 6414
rect 1829 6402 1848 6414
rect 1902 6412 1929 6414
rect 1938 6412 2159 6422
rect 2194 6419 2200 6422
rect 1902 6408 2159 6412
rect 1797 6394 1848 6402
rect 1895 6394 2159 6408
rect 2203 6414 2238 6422
rect 1749 6346 1768 6380
rect 1813 6386 1842 6394
rect 1813 6380 1830 6386
rect 1813 6378 1847 6380
rect 1895 6378 1911 6394
rect 1912 6384 2120 6394
rect 2121 6384 2137 6394
rect 2185 6390 2200 6405
rect 2203 6402 2204 6414
rect 2211 6402 2238 6414
rect 2203 6394 2238 6402
rect 2203 6393 2232 6394
rect 1923 6380 2137 6384
rect 1938 6378 2137 6380
rect 2172 6380 2185 6390
rect 2203 6380 2220 6393
rect 2172 6378 2220 6380
rect 1814 6374 1847 6378
rect 1810 6372 1847 6374
rect 1810 6371 1877 6372
rect 1810 6366 1841 6371
rect 1847 6366 1877 6371
rect 1810 6362 1877 6366
rect 1783 6359 1877 6362
rect 1783 6352 1832 6359
rect 1783 6346 1813 6352
rect 1832 6347 1837 6352
rect 1749 6330 1829 6346
rect 1841 6338 1877 6359
rect 1938 6354 2127 6378
rect 2172 6377 2219 6378
rect 2185 6372 2219 6377
rect 1953 6351 2127 6354
rect 1946 6348 2127 6351
rect 2155 6371 2219 6372
rect 1749 6328 1768 6330
rect 1783 6328 1817 6330
rect 1749 6312 1829 6328
rect 1749 6306 1768 6312
rect 1465 6280 1568 6290
rect 1419 6278 1568 6280
rect 1589 6278 1624 6290
rect 1258 6276 1420 6278
rect 1270 6256 1289 6276
rect 1304 6274 1334 6276
rect 1153 6248 1194 6256
rect 1276 6252 1289 6256
rect 1341 6260 1420 6276
rect 1452 6276 1624 6278
rect 1452 6260 1531 6276
rect 1538 6274 1568 6276
rect 1116 6238 1145 6248
rect 1159 6238 1188 6248
rect 1203 6238 1233 6252
rect 1276 6238 1319 6252
rect 1341 6248 1531 6260
rect 1596 6256 1602 6276
rect 1326 6238 1356 6248
rect 1357 6238 1515 6248
rect 1519 6238 1549 6248
rect 1553 6238 1583 6252
rect 1611 6238 1624 6276
rect 1696 6290 1725 6306
rect 1739 6290 1768 6306
rect 1783 6296 1813 6312
rect 1841 6290 1847 6338
rect 1850 6332 1869 6338
rect 1884 6332 1914 6340
rect 1850 6324 1914 6332
rect 1850 6308 1930 6324
rect 1946 6317 2008 6348
rect 2024 6317 2086 6348
rect 2155 6346 2204 6371
rect 2219 6346 2249 6362
rect 2118 6332 2148 6340
rect 2155 6338 2265 6346
rect 2118 6324 2163 6332
rect 1850 6306 1869 6308
rect 1884 6306 1930 6308
rect 1850 6290 1930 6306
rect 1957 6304 1992 6317
rect 2033 6314 2070 6317
rect 2033 6312 2075 6314
rect 1962 6301 1992 6304
rect 1971 6297 1978 6301
rect 1978 6296 1979 6297
rect 1937 6290 1947 6296
rect 1696 6282 1731 6290
rect 1696 6256 1697 6282
rect 1704 6256 1731 6282
rect 1639 6238 1669 6252
rect 1696 6248 1731 6256
rect 1733 6282 1774 6290
rect 1733 6256 1748 6282
rect 1755 6256 1774 6282
rect 1838 6278 1869 6290
rect 1884 6278 1987 6290
rect 1999 6280 2025 6306
rect 2040 6301 2070 6312
rect 2102 6308 2164 6324
rect 2102 6306 2148 6308
rect 2102 6290 2164 6306
rect 2176 6290 2182 6338
rect 2185 6330 2265 6338
rect 2185 6328 2204 6330
rect 2219 6328 2253 6330
rect 2185 6312 2265 6328
rect 2185 6290 2204 6312
rect 2219 6296 2249 6312
rect 2277 6306 2283 6380
rect 2286 6306 2305 6450
rect 2320 6306 2326 6450
rect 2335 6380 2348 6450
rect 2400 6446 2422 6450
rect 2393 6424 2422 6438
rect 2475 6424 2491 6438
rect 2529 6434 2535 6436
rect 2542 6434 2650 6450
rect 2657 6434 2663 6436
rect 2671 6434 2686 6450
rect 2752 6444 2771 6447
rect 2393 6422 2491 6424
rect 2518 6422 2686 6434
rect 2701 6424 2717 6438
rect 2752 6425 2774 6444
rect 2784 6438 2800 6439
rect 2783 6436 2800 6438
rect 2784 6431 2800 6436
rect 2774 6424 2780 6425
rect 2783 6424 2812 6431
rect 2701 6423 2812 6424
rect 2701 6422 2818 6423
rect 2377 6414 2428 6422
rect 2475 6414 2509 6422
rect 2377 6402 2402 6414
rect 2409 6402 2428 6414
rect 2482 6412 2509 6414
rect 2518 6412 2739 6422
rect 2774 6419 2780 6422
rect 2482 6408 2739 6412
rect 2377 6394 2428 6402
rect 2475 6394 2739 6408
rect 2783 6414 2818 6422
rect 2329 6346 2348 6380
rect 2393 6386 2422 6394
rect 2393 6380 2410 6386
rect 2393 6378 2427 6380
rect 2475 6378 2491 6394
rect 2492 6384 2700 6394
rect 2701 6384 2717 6394
rect 2765 6390 2780 6405
rect 2783 6402 2784 6414
rect 2791 6402 2818 6414
rect 2783 6394 2818 6402
rect 2783 6393 2812 6394
rect 2503 6380 2717 6384
rect 2518 6378 2717 6380
rect 2752 6380 2765 6390
rect 2783 6380 2800 6393
rect 2752 6378 2800 6380
rect 2394 6374 2427 6378
rect 2390 6372 2427 6374
rect 2390 6371 2457 6372
rect 2390 6366 2421 6371
rect 2427 6366 2457 6371
rect 2390 6362 2457 6366
rect 2363 6359 2457 6362
rect 2363 6352 2412 6359
rect 2363 6346 2393 6352
rect 2412 6347 2417 6352
rect 2329 6330 2409 6346
rect 2421 6338 2457 6359
rect 2518 6354 2707 6378
rect 2752 6377 2799 6378
rect 2765 6372 2799 6377
rect 2533 6351 2707 6354
rect 2526 6348 2707 6351
rect 2735 6371 2799 6372
rect 2329 6328 2348 6330
rect 2363 6328 2397 6330
rect 2329 6312 2409 6328
rect 2329 6306 2348 6312
rect 2045 6280 2148 6290
rect 1999 6278 2148 6280
rect 2169 6278 2204 6290
rect 1838 6276 2000 6278
rect 1850 6256 1869 6276
rect 1884 6274 1914 6276
rect 1733 6248 1774 6256
rect 1856 6252 1869 6256
rect 1921 6260 2000 6276
rect 2032 6276 2204 6278
rect 2032 6260 2111 6276
rect 2118 6274 2148 6276
rect 1696 6238 1725 6248
rect 1739 6238 1768 6248
rect 1783 6238 1813 6252
rect 1856 6238 1899 6252
rect 1921 6248 2111 6260
rect 2176 6256 2182 6276
rect 1906 6238 1936 6248
rect 1937 6238 2095 6248
rect 2099 6238 2129 6248
rect 2133 6238 2163 6252
rect 2191 6238 2204 6276
rect 2276 6290 2305 6306
rect 2319 6290 2348 6306
rect 2363 6296 2393 6312
rect 2421 6290 2427 6338
rect 2430 6332 2449 6338
rect 2464 6332 2494 6340
rect 2430 6324 2494 6332
rect 2430 6308 2510 6324
rect 2526 6317 2588 6348
rect 2604 6317 2666 6348
rect 2735 6346 2784 6371
rect 2799 6346 2829 6362
rect 2698 6332 2728 6340
rect 2735 6338 2845 6346
rect 2698 6324 2743 6332
rect 2430 6306 2449 6308
rect 2464 6306 2510 6308
rect 2430 6290 2510 6306
rect 2537 6304 2572 6317
rect 2613 6314 2650 6317
rect 2613 6312 2655 6314
rect 2542 6301 2572 6304
rect 2551 6297 2558 6301
rect 2558 6296 2559 6297
rect 2517 6290 2527 6296
rect 2276 6282 2311 6290
rect 2276 6256 2277 6282
rect 2284 6256 2311 6282
rect 2219 6238 2249 6252
rect 2276 6248 2311 6256
rect 2313 6282 2354 6290
rect 2313 6256 2328 6282
rect 2335 6256 2354 6282
rect 2418 6278 2449 6290
rect 2464 6278 2567 6290
rect 2579 6280 2605 6306
rect 2620 6301 2650 6312
rect 2682 6308 2744 6324
rect 2682 6306 2728 6308
rect 2682 6290 2744 6306
rect 2756 6290 2762 6338
rect 2765 6330 2845 6338
rect 2765 6328 2784 6330
rect 2799 6328 2833 6330
rect 2765 6312 2845 6328
rect 2765 6290 2784 6312
rect 2799 6296 2829 6312
rect 2857 6306 2863 6380
rect 2866 6306 2885 6450
rect 2900 6306 2906 6450
rect 2915 6380 2928 6450
rect 2980 6446 3002 6450
rect 2973 6424 3002 6438
rect 3055 6424 3071 6438
rect 3109 6434 3115 6436
rect 3122 6434 3230 6450
rect 3237 6434 3243 6436
rect 3251 6434 3266 6450
rect 3332 6444 3351 6447
rect 2973 6422 3071 6424
rect 3098 6422 3266 6434
rect 3281 6424 3297 6438
rect 3332 6425 3354 6444
rect 3364 6438 3380 6439
rect 3363 6436 3380 6438
rect 3364 6431 3380 6436
rect 3354 6424 3360 6425
rect 3363 6424 3392 6431
rect 3281 6423 3392 6424
rect 3281 6422 3398 6423
rect 2957 6414 3008 6422
rect 3055 6414 3089 6422
rect 2957 6402 2982 6414
rect 2989 6402 3008 6414
rect 3062 6412 3089 6414
rect 3098 6412 3319 6422
rect 3354 6419 3360 6422
rect 3062 6408 3319 6412
rect 2957 6394 3008 6402
rect 3055 6394 3319 6408
rect 3363 6414 3398 6422
rect 2909 6346 2928 6380
rect 2973 6386 3002 6394
rect 2973 6380 2990 6386
rect 2973 6378 3007 6380
rect 3055 6378 3071 6394
rect 3072 6384 3280 6394
rect 3281 6384 3297 6394
rect 3345 6390 3360 6405
rect 3363 6402 3364 6414
rect 3371 6402 3398 6414
rect 3363 6394 3398 6402
rect 3363 6393 3392 6394
rect 3083 6380 3297 6384
rect 3098 6378 3297 6380
rect 3332 6380 3345 6390
rect 3363 6380 3380 6393
rect 3332 6378 3380 6380
rect 2974 6374 3007 6378
rect 2970 6372 3007 6374
rect 2970 6371 3037 6372
rect 2970 6366 3001 6371
rect 3007 6366 3037 6371
rect 2970 6362 3037 6366
rect 2943 6359 3037 6362
rect 2943 6352 2992 6359
rect 2943 6346 2973 6352
rect 2992 6347 2997 6352
rect 2909 6330 2989 6346
rect 3001 6338 3037 6359
rect 3098 6354 3287 6378
rect 3332 6377 3379 6378
rect 3345 6372 3379 6377
rect 3113 6351 3287 6354
rect 3106 6348 3287 6351
rect 3315 6371 3379 6372
rect 2909 6328 2928 6330
rect 2943 6328 2977 6330
rect 2909 6312 2989 6328
rect 2909 6306 2928 6312
rect 2625 6280 2728 6290
rect 2579 6278 2728 6280
rect 2749 6278 2784 6290
rect 2418 6276 2580 6278
rect 2430 6256 2449 6276
rect 2464 6274 2494 6276
rect 2313 6248 2354 6256
rect 2436 6252 2449 6256
rect 2501 6260 2580 6276
rect 2612 6276 2784 6278
rect 2612 6260 2691 6276
rect 2698 6274 2728 6276
rect 2276 6238 2305 6248
rect 2319 6238 2348 6248
rect 2363 6238 2393 6252
rect 2436 6238 2479 6252
rect 2501 6248 2691 6260
rect 2756 6256 2762 6276
rect 2486 6238 2516 6248
rect 2517 6238 2675 6248
rect 2679 6238 2709 6248
rect 2713 6238 2743 6252
rect 2771 6238 2784 6276
rect 2856 6290 2885 6306
rect 2899 6290 2928 6306
rect 2943 6296 2973 6312
rect 3001 6290 3007 6338
rect 3010 6332 3029 6338
rect 3044 6332 3074 6340
rect 3010 6324 3074 6332
rect 3010 6308 3090 6324
rect 3106 6317 3168 6348
rect 3184 6317 3246 6348
rect 3315 6346 3364 6371
rect 3379 6346 3409 6362
rect 3278 6332 3308 6340
rect 3315 6338 3425 6346
rect 3278 6324 3323 6332
rect 3010 6306 3029 6308
rect 3044 6306 3090 6308
rect 3010 6290 3090 6306
rect 3117 6304 3152 6317
rect 3193 6314 3230 6317
rect 3193 6312 3235 6314
rect 3122 6301 3152 6304
rect 3131 6297 3138 6301
rect 3138 6296 3139 6297
rect 3097 6290 3107 6296
rect 2856 6282 2891 6290
rect 2856 6256 2857 6282
rect 2864 6256 2891 6282
rect 2799 6238 2829 6252
rect 2856 6248 2891 6256
rect 2893 6282 2934 6290
rect 2893 6256 2908 6282
rect 2915 6256 2934 6282
rect 2998 6278 3029 6290
rect 3044 6278 3147 6290
rect 3159 6280 3185 6306
rect 3200 6301 3230 6312
rect 3262 6308 3324 6324
rect 3262 6306 3308 6308
rect 3262 6290 3324 6306
rect 3336 6290 3342 6338
rect 3345 6330 3425 6338
rect 3345 6328 3364 6330
rect 3379 6328 3413 6330
rect 3345 6312 3425 6328
rect 3345 6290 3364 6312
rect 3379 6296 3409 6312
rect 3437 6306 3443 6380
rect 3446 6306 3465 6450
rect 3480 6306 3486 6450
rect 3495 6380 3508 6450
rect 3560 6446 3582 6450
rect 3553 6424 3582 6438
rect 3635 6424 3651 6438
rect 3689 6434 3695 6436
rect 3702 6434 3810 6450
rect 3817 6434 3823 6436
rect 3831 6434 3846 6450
rect 3912 6444 3931 6447
rect 3553 6422 3651 6424
rect 3678 6422 3846 6434
rect 3861 6424 3877 6438
rect 3912 6425 3934 6444
rect 3944 6438 3960 6439
rect 3943 6436 3960 6438
rect 3944 6431 3960 6436
rect 3934 6424 3940 6425
rect 3943 6424 3972 6431
rect 3861 6423 3972 6424
rect 3861 6422 3978 6423
rect 3537 6414 3588 6422
rect 3635 6414 3669 6422
rect 3537 6402 3562 6414
rect 3569 6402 3588 6414
rect 3642 6412 3669 6414
rect 3678 6412 3899 6422
rect 3934 6419 3940 6422
rect 3642 6408 3899 6412
rect 3537 6394 3588 6402
rect 3635 6394 3899 6408
rect 3943 6414 3978 6422
rect 3489 6346 3508 6380
rect 3553 6386 3582 6394
rect 3553 6380 3570 6386
rect 3553 6378 3587 6380
rect 3635 6378 3651 6394
rect 3652 6384 3860 6394
rect 3861 6384 3877 6394
rect 3925 6390 3940 6405
rect 3943 6402 3944 6414
rect 3951 6402 3978 6414
rect 3943 6394 3978 6402
rect 3943 6393 3972 6394
rect 3663 6380 3877 6384
rect 3678 6378 3877 6380
rect 3912 6380 3925 6390
rect 3943 6380 3960 6393
rect 3912 6378 3960 6380
rect 3554 6374 3587 6378
rect 3550 6372 3587 6374
rect 3550 6371 3617 6372
rect 3550 6366 3581 6371
rect 3587 6366 3617 6371
rect 3550 6362 3617 6366
rect 3523 6359 3617 6362
rect 3523 6352 3572 6359
rect 3523 6346 3553 6352
rect 3572 6347 3577 6352
rect 3489 6330 3569 6346
rect 3581 6338 3617 6359
rect 3678 6354 3867 6378
rect 3912 6377 3959 6378
rect 3925 6372 3959 6377
rect 3693 6351 3867 6354
rect 3686 6348 3867 6351
rect 3895 6371 3959 6372
rect 3489 6328 3508 6330
rect 3523 6328 3557 6330
rect 3489 6312 3569 6328
rect 3489 6306 3508 6312
rect 3205 6280 3308 6290
rect 3159 6278 3308 6280
rect 3329 6278 3364 6290
rect 2998 6276 3160 6278
rect 3010 6256 3029 6276
rect 3044 6274 3074 6276
rect 2893 6248 2934 6256
rect 3016 6252 3029 6256
rect 3081 6260 3160 6276
rect 3192 6276 3364 6278
rect 3192 6260 3271 6276
rect 3278 6274 3308 6276
rect 2856 6238 2885 6248
rect 2899 6238 2928 6248
rect 2943 6238 2973 6252
rect 3016 6238 3059 6252
rect 3081 6248 3271 6260
rect 3336 6256 3342 6276
rect 3066 6238 3096 6248
rect 3097 6238 3255 6248
rect 3259 6238 3289 6248
rect 3293 6238 3323 6252
rect 3351 6238 3364 6276
rect 3436 6290 3465 6306
rect 3479 6290 3508 6306
rect 3523 6296 3553 6312
rect 3581 6290 3587 6338
rect 3590 6332 3609 6338
rect 3624 6332 3654 6340
rect 3590 6324 3654 6332
rect 3590 6308 3670 6324
rect 3686 6317 3748 6348
rect 3764 6317 3826 6348
rect 3895 6346 3944 6371
rect 3959 6346 3989 6362
rect 3858 6332 3888 6340
rect 3895 6338 4005 6346
rect 3858 6324 3903 6332
rect 3590 6306 3609 6308
rect 3624 6306 3670 6308
rect 3590 6290 3670 6306
rect 3697 6304 3732 6317
rect 3773 6314 3810 6317
rect 3773 6312 3815 6314
rect 3702 6301 3732 6304
rect 3711 6297 3718 6301
rect 3718 6296 3719 6297
rect 3677 6290 3687 6296
rect 3436 6282 3471 6290
rect 3436 6256 3437 6282
rect 3444 6256 3471 6282
rect 3379 6238 3409 6252
rect 3436 6248 3471 6256
rect 3473 6282 3514 6290
rect 3473 6256 3488 6282
rect 3495 6256 3514 6282
rect 3578 6278 3609 6290
rect 3624 6278 3727 6290
rect 3739 6280 3765 6306
rect 3780 6301 3810 6312
rect 3842 6308 3904 6324
rect 3842 6306 3888 6308
rect 3842 6290 3904 6306
rect 3916 6290 3922 6338
rect 3925 6330 4005 6338
rect 3925 6328 3944 6330
rect 3959 6328 3993 6330
rect 3925 6312 4005 6328
rect 3925 6290 3944 6312
rect 3959 6296 3989 6312
rect 4017 6306 4023 6380
rect 4026 6306 4045 6450
rect 4060 6306 4066 6450
rect 4075 6380 4088 6450
rect 4140 6446 4162 6450
rect 4133 6424 4162 6438
rect 4215 6424 4231 6438
rect 4269 6434 4275 6436
rect 4282 6434 4390 6450
rect 4397 6434 4403 6436
rect 4411 6434 4426 6450
rect 4492 6444 4511 6447
rect 4133 6422 4231 6424
rect 4258 6422 4426 6434
rect 4441 6424 4457 6438
rect 4492 6425 4514 6444
rect 4524 6438 4540 6439
rect 4523 6436 4540 6438
rect 4524 6431 4540 6436
rect 4514 6424 4520 6425
rect 4523 6424 4552 6431
rect 4441 6423 4552 6424
rect 4441 6422 4558 6423
rect 4117 6414 4168 6422
rect 4215 6414 4249 6422
rect 4117 6402 4142 6414
rect 4149 6402 4168 6414
rect 4222 6412 4249 6414
rect 4258 6412 4479 6422
rect 4514 6419 4520 6422
rect 4222 6408 4479 6412
rect 4117 6394 4168 6402
rect 4215 6394 4479 6408
rect 4523 6414 4558 6422
rect 4069 6346 4088 6380
rect 4133 6386 4162 6394
rect 4133 6380 4150 6386
rect 4133 6378 4167 6380
rect 4215 6378 4231 6394
rect 4232 6384 4440 6394
rect 4441 6384 4457 6394
rect 4505 6390 4520 6405
rect 4523 6402 4524 6414
rect 4531 6402 4558 6414
rect 4523 6394 4558 6402
rect 4523 6393 4552 6394
rect 4243 6380 4457 6384
rect 4258 6378 4457 6380
rect 4492 6380 4505 6390
rect 4523 6380 4540 6393
rect 4492 6378 4540 6380
rect 4134 6374 4167 6378
rect 4130 6372 4167 6374
rect 4130 6371 4197 6372
rect 4130 6366 4161 6371
rect 4167 6366 4197 6371
rect 4130 6362 4197 6366
rect 4103 6359 4197 6362
rect 4103 6352 4152 6359
rect 4103 6346 4133 6352
rect 4152 6347 4157 6352
rect 4069 6330 4149 6346
rect 4161 6338 4197 6359
rect 4258 6354 4447 6378
rect 4492 6377 4539 6378
rect 4505 6372 4539 6377
rect 4273 6351 4447 6354
rect 4266 6348 4447 6351
rect 4475 6371 4539 6372
rect 4069 6328 4088 6330
rect 4103 6328 4137 6330
rect 4069 6312 4149 6328
rect 4069 6306 4088 6312
rect 3785 6280 3888 6290
rect 3739 6278 3888 6280
rect 3909 6278 3944 6290
rect 3578 6276 3740 6278
rect 3590 6256 3609 6276
rect 3624 6274 3654 6276
rect 3473 6248 3514 6256
rect 3596 6252 3609 6256
rect 3661 6260 3740 6276
rect 3772 6276 3944 6278
rect 3772 6260 3851 6276
rect 3858 6274 3888 6276
rect 3436 6238 3465 6248
rect 3479 6238 3508 6248
rect 3523 6238 3553 6252
rect 3596 6238 3639 6252
rect 3661 6248 3851 6260
rect 3916 6256 3922 6276
rect 3646 6238 3676 6248
rect 3677 6238 3835 6248
rect 3839 6238 3869 6248
rect 3873 6238 3903 6252
rect 3931 6238 3944 6276
rect 4016 6290 4045 6306
rect 4059 6290 4088 6306
rect 4103 6296 4133 6312
rect 4161 6290 4167 6338
rect 4170 6332 4189 6338
rect 4204 6332 4234 6340
rect 4170 6324 4234 6332
rect 4170 6308 4250 6324
rect 4266 6317 4328 6348
rect 4344 6317 4406 6348
rect 4475 6346 4524 6371
rect 4539 6346 4569 6362
rect 4438 6332 4468 6340
rect 4475 6338 4585 6346
rect 4438 6324 4483 6332
rect 4170 6306 4189 6308
rect 4204 6306 4250 6308
rect 4170 6290 4250 6306
rect 4277 6304 4312 6317
rect 4353 6314 4390 6317
rect 4353 6312 4395 6314
rect 4282 6301 4312 6304
rect 4291 6297 4298 6301
rect 4298 6296 4299 6297
rect 4257 6290 4267 6296
rect 4016 6282 4051 6290
rect 4016 6256 4017 6282
rect 4024 6256 4051 6282
rect 3959 6238 3989 6252
rect 4016 6248 4051 6256
rect 4053 6282 4094 6290
rect 4053 6256 4068 6282
rect 4075 6256 4094 6282
rect 4158 6278 4189 6290
rect 4204 6278 4307 6290
rect 4319 6280 4345 6306
rect 4360 6301 4390 6312
rect 4422 6308 4484 6324
rect 4422 6306 4468 6308
rect 4422 6290 4484 6306
rect 4496 6290 4502 6338
rect 4505 6330 4585 6338
rect 4505 6328 4524 6330
rect 4539 6328 4573 6330
rect 4505 6312 4585 6328
rect 4505 6290 4524 6312
rect 4539 6296 4569 6312
rect 4597 6306 4603 6380
rect 4606 6306 4625 6450
rect 4640 6306 4646 6450
rect 4655 6380 4668 6450
rect 4720 6446 4742 6450
rect 4713 6424 4742 6438
rect 4795 6424 4811 6438
rect 4849 6434 4855 6436
rect 4862 6434 4970 6450
rect 4977 6434 4983 6436
rect 4991 6434 5006 6450
rect 5072 6444 5091 6447
rect 4713 6422 4811 6424
rect 4838 6422 5006 6434
rect 5021 6424 5037 6438
rect 5072 6425 5094 6444
rect 5104 6438 5120 6439
rect 5103 6436 5120 6438
rect 5104 6431 5120 6436
rect 5094 6424 5100 6425
rect 5103 6424 5132 6431
rect 5021 6423 5132 6424
rect 5021 6422 5138 6423
rect 4697 6414 4748 6422
rect 4795 6414 4829 6422
rect 4697 6402 4722 6414
rect 4729 6402 4748 6414
rect 4802 6412 4829 6414
rect 4838 6412 5059 6422
rect 5094 6419 5100 6422
rect 4802 6408 5059 6412
rect 4697 6394 4748 6402
rect 4795 6394 5059 6408
rect 5103 6414 5138 6422
rect 4649 6346 4668 6380
rect 4713 6386 4742 6394
rect 4713 6380 4730 6386
rect 4713 6378 4747 6380
rect 4795 6378 4811 6394
rect 4812 6384 5020 6394
rect 5021 6384 5037 6394
rect 5085 6390 5100 6405
rect 5103 6402 5104 6414
rect 5111 6402 5138 6414
rect 5103 6394 5138 6402
rect 5103 6393 5132 6394
rect 4823 6380 5037 6384
rect 4838 6378 5037 6380
rect 5072 6380 5085 6390
rect 5103 6380 5120 6393
rect 5072 6378 5120 6380
rect 4714 6374 4747 6378
rect 4710 6372 4747 6374
rect 4710 6371 4777 6372
rect 4710 6366 4741 6371
rect 4747 6366 4777 6371
rect 4710 6362 4777 6366
rect 4683 6359 4777 6362
rect 4683 6352 4732 6359
rect 4683 6346 4713 6352
rect 4732 6347 4737 6352
rect 4649 6330 4729 6346
rect 4741 6338 4777 6359
rect 4838 6354 5027 6378
rect 5072 6377 5119 6378
rect 5085 6372 5119 6377
rect 4853 6351 5027 6354
rect 4846 6348 5027 6351
rect 5055 6371 5119 6372
rect 4649 6328 4668 6330
rect 4683 6328 4717 6330
rect 4649 6312 4729 6328
rect 4649 6306 4668 6312
rect 4365 6280 4468 6290
rect 4319 6278 4468 6280
rect 4489 6278 4524 6290
rect 4158 6276 4320 6278
rect 4170 6256 4189 6276
rect 4204 6274 4234 6276
rect 4053 6248 4094 6256
rect 4176 6252 4189 6256
rect 4241 6260 4320 6276
rect 4352 6276 4524 6278
rect 4352 6260 4431 6276
rect 4438 6274 4468 6276
rect 4016 6238 4045 6248
rect 4059 6238 4088 6248
rect 4103 6238 4133 6252
rect 4176 6238 4219 6252
rect 4241 6248 4431 6260
rect 4496 6256 4502 6276
rect 4226 6238 4256 6248
rect 4257 6238 4415 6248
rect 4419 6238 4449 6248
rect 4453 6238 4483 6252
rect 4511 6238 4524 6276
rect 4596 6290 4625 6306
rect 4639 6290 4668 6306
rect 4683 6296 4713 6312
rect 4741 6290 4747 6338
rect 4750 6332 4769 6338
rect 4784 6332 4814 6340
rect 4750 6324 4814 6332
rect 4750 6308 4830 6324
rect 4846 6317 4908 6348
rect 4924 6317 4986 6348
rect 5055 6346 5104 6371
rect 5119 6346 5149 6362
rect 5018 6332 5048 6340
rect 5055 6338 5165 6346
rect 5018 6324 5063 6332
rect 4750 6306 4769 6308
rect 4784 6306 4830 6308
rect 4750 6290 4830 6306
rect 4857 6304 4892 6317
rect 4933 6314 4970 6317
rect 4933 6312 4975 6314
rect 4862 6301 4892 6304
rect 4871 6297 4878 6301
rect 4878 6296 4879 6297
rect 4837 6290 4847 6296
rect 4596 6282 4631 6290
rect 4596 6256 4597 6282
rect 4604 6256 4631 6282
rect 4539 6238 4569 6252
rect 4596 6248 4631 6256
rect 4633 6282 4674 6290
rect 4633 6256 4648 6282
rect 4655 6256 4674 6282
rect 4738 6278 4769 6290
rect 4784 6278 4887 6290
rect 4899 6280 4925 6306
rect 4940 6301 4970 6312
rect 5002 6308 5064 6324
rect 5002 6306 5048 6308
rect 5002 6290 5064 6306
rect 5076 6290 5082 6338
rect 5085 6330 5165 6338
rect 5085 6328 5104 6330
rect 5119 6328 5153 6330
rect 5085 6312 5165 6328
rect 5085 6290 5104 6312
rect 5119 6296 5149 6312
rect 5177 6306 5183 6380
rect 5186 6306 5205 6450
rect 5220 6306 5226 6450
rect 5235 6380 5248 6450
rect 5300 6446 5322 6450
rect 5293 6424 5322 6438
rect 5375 6424 5391 6438
rect 5429 6434 5435 6436
rect 5442 6434 5550 6450
rect 5557 6434 5563 6436
rect 5571 6434 5586 6450
rect 5652 6444 5671 6447
rect 5293 6422 5391 6424
rect 5418 6422 5586 6434
rect 5601 6424 5617 6438
rect 5652 6425 5674 6444
rect 5684 6438 5700 6439
rect 5683 6436 5700 6438
rect 5684 6431 5700 6436
rect 5674 6424 5680 6425
rect 5683 6424 5712 6431
rect 5601 6423 5712 6424
rect 5601 6422 5718 6423
rect 5277 6414 5328 6422
rect 5375 6414 5409 6422
rect 5277 6402 5302 6414
rect 5309 6402 5328 6414
rect 5382 6412 5409 6414
rect 5418 6412 5639 6422
rect 5674 6419 5680 6422
rect 5382 6408 5639 6412
rect 5277 6394 5328 6402
rect 5375 6394 5639 6408
rect 5683 6414 5718 6422
rect 5229 6346 5248 6380
rect 5293 6386 5322 6394
rect 5293 6380 5310 6386
rect 5293 6378 5327 6380
rect 5375 6378 5391 6394
rect 5392 6384 5600 6394
rect 5601 6384 5617 6394
rect 5665 6390 5680 6405
rect 5683 6402 5684 6414
rect 5691 6402 5718 6414
rect 5683 6394 5718 6402
rect 5683 6393 5712 6394
rect 5403 6380 5617 6384
rect 5418 6378 5617 6380
rect 5652 6380 5665 6390
rect 5683 6380 5700 6393
rect 5652 6378 5700 6380
rect 5294 6374 5327 6378
rect 5290 6372 5327 6374
rect 5290 6371 5357 6372
rect 5290 6366 5321 6371
rect 5327 6366 5357 6371
rect 5290 6362 5357 6366
rect 5263 6359 5357 6362
rect 5263 6352 5312 6359
rect 5263 6346 5293 6352
rect 5312 6347 5317 6352
rect 5229 6330 5309 6346
rect 5321 6338 5357 6359
rect 5418 6354 5607 6378
rect 5652 6377 5699 6378
rect 5665 6372 5699 6377
rect 5433 6351 5607 6354
rect 5426 6348 5607 6351
rect 5635 6371 5699 6372
rect 5229 6328 5248 6330
rect 5263 6328 5297 6330
rect 5229 6312 5309 6328
rect 5229 6306 5248 6312
rect 4945 6280 5048 6290
rect 4899 6278 5048 6280
rect 5069 6278 5104 6290
rect 4738 6276 4900 6278
rect 4750 6256 4769 6276
rect 4784 6274 4814 6276
rect 4633 6248 4674 6256
rect 4756 6252 4769 6256
rect 4821 6260 4900 6276
rect 4932 6276 5104 6278
rect 4932 6260 5011 6276
rect 5018 6274 5048 6276
rect 4596 6238 4625 6248
rect 4639 6238 4668 6248
rect 4683 6238 4713 6252
rect 4756 6238 4799 6252
rect 4821 6248 5011 6260
rect 5076 6256 5082 6276
rect 4806 6238 4836 6248
rect 4837 6238 4995 6248
rect 4999 6238 5029 6248
rect 5033 6238 5063 6252
rect 5091 6238 5104 6276
rect 5176 6290 5205 6306
rect 5219 6290 5248 6306
rect 5263 6296 5293 6312
rect 5321 6290 5327 6338
rect 5330 6332 5349 6338
rect 5364 6332 5394 6340
rect 5330 6324 5394 6332
rect 5330 6308 5410 6324
rect 5426 6317 5488 6348
rect 5504 6317 5566 6348
rect 5635 6346 5684 6371
rect 5699 6346 5729 6362
rect 5598 6332 5628 6340
rect 5635 6338 5745 6346
rect 5598 6324 5643 6332
rect 5330 6306 5349 6308
rect 5364 6306 5410 6308
rect 5330 6290 5410 6306
rect 5437 6304 5472 6317
rect 5513 6314 5550 6317
rect 5513 6312 5555 6314
rect 5442 6301 5472 6304
rect 5451 6297 5458 6301
rect 5458 6296 5459 6297
rect 5417 6290 5427 6296
rect 5176 6282 5211 6290
rect 5176 6256 5177 6282
rect 5184 6256 5211 6282
rect 5119 6238 5149 6252
rect 5176 6248 5211 6256
rect 5213 6282 5254 6290
rect 5213 6256 5228 6282
rect 5235 6256 5254 6282
rect 5318 6278 5349 6290
rect 5364 6278 5467 6290
rect 5479 6280 5505 6306
rect 5520 6301 5550 6312
rect 5582 6308 5644 6324
rect 5582 6306 5628 6308
rect 5582 6290 5644 6306
rect 5656 6290 5662 6338
rect 5665 6330 5745 6338
rect 5665 6328 5684 6330
rect 5699 6328 5733 6330
rect 5665 6312 5745 6328
rect 5665 6290 5684 6312
rect 5699 6296 5729 6312
rect 5757 6306 5763 6380
rect 5766 6306 5785 6450
rect 5800 6306 5806 6450
rect 5815 6380 5828 6450
rect 5880 6446 5902 6450
rect 5873 6424 5902 6438
rect 5955 6424 5971 6438
rect 6009 6434 6015 6436
rect 6022 6434 6130 6450
rect 6137 6434 6143 6436
rect 6151 6434 6166 6450
rect 6232 6444 6251 6447
rect 5873 6422 5971 6424
rect 5998 6422 6166 6434
rect 6181 6424 6197 6438
rect 6232 6425 6254 6444
rect 6264 6438 6280 6439
rect 6263 6436 6280 6438
rect 6264 6431 6280 6436
rect 6254 6424 6260 6425
rect 6263 6424 6292 6431
rect 6181 6423 6292 6424
rect 6181 6422 6298 6423
rect 5857 6414 5908 6422
rect 5955 6414 5989 6422
rect 5857 6402 5882 6414
rect 5889 6402 5908 6414
rect 5962 6412 5989 6414
rect 5998 6412 6219 6422
rect 6254 6419 6260 6422
rect 5962 6408 6219 6412
rect 5857 6394 5908 6402
rect 5955 6394 6219 6408
rect 6263 6414 6298 6422
rect 5809 6346 5828 6380
rect 5873 6386 5902 6394
rect 5873 6380 5890 6386
rect 5873 6378 5907 6380
rect 5955 6378 5971 6394
rect 5972 6384 6180 6394
rect 6181 6384 6197 6394
rect 6245 6390 6260 6405
rect 6263 6402 6264 6414
rect 6271 6402 6298 6414
rect 6263 6394 6298 6402
rect 6263 6393 6292 6394
rect 5983 6380 6197 6384
rect 5998 6378 6197 6380
rect 6232 6380 6245 6390
rect 6263 6380 6280 6393
rect 6232 6378 6280 6380
rect 5874 6374 5907 6378
rect 5870 6372 5907 6374
rect 5870 6371 5937 6372
rect 5870 6366 5901 6371
rect 5907 6366 5937 6371
rect 5870 6362 5937 6366
rect 5843 6359 5937 6362
rect 5843 6352 5892 6359
rect 5843 6346 5873 6352
rect 5892 6347 5897 6352
rect 5809 6330 5889 6346
rect 5901 6338 5937 6359
rect 5998 6354 6187 6378
rect 6232 6377 6279 6378
rect 6245 6372 6279 6377
rect 6013 6351 6187 6354
rect 6006 6348 6187 6351
rect 6215 6371 6279 6372
rect 5809 6328 5828 6330
rect 5843 6328 5877 6330
rect 5809 6312 5889 6328
rect 5809 6306 5828 6312
rect 5525 6280 5628 6290
rect 5479 6278 5628 6280
rect 5649 6278 5684 6290
rect 5318 6276 5480 6278
rect 5330 6256 5349 6276
rect 5364 6274 5394 6276
rect 5213 6248 5254 6256
rect 5336 6252 5349 6256
rect 5401 6260 5480 6276
rect 5512 6276 5684 6278
rect 5512 6260 5591 6276
rect 5598 6274 5628 6276
rect 5176 6238 5205 6248
rect 5219 6238 5248 6248
rect 5263 6238 5293 6252
rect 5336 6238 5379 6252
rect 5401 6248 5591 6260
rect 5656 6256 5662 6276
rect 5386 6238 5416 6248
rect 5417 6238 5575 6248
rect 5579 6238 5609 6248
rect 5613 6238 5643 6252
rect 5671 6238 5684 6276
rect 5756 6290 5785 6306
rect 5799 6290 5828 6306
rect 5843 6296 5873 6312
rect 5901 6290 5907 6338
rect 5910 6332 5929 6338
rect 5944 6332 5974 6340
rect 5910 6324 5974 6332
rect 5910 6308 5990 6324
rect 6006 6317 6068 6348
rect 6084 6317 6146 6348
rect 6215 6346 6264 6371
rect 6279 6346 6309 6362
rect 6178 6332 6208 6340
rect 6215 6338 6325 6346
rect 6178 6324 6223 6332
rect 5910 6306 5929 6308
rect 5944 6306 5990 6308
rect 5910 6290 5990 6306
rect 6017 6304 6052 6317
rect 6093 6314 6130 6317
rect 6093 6312 6135 6314
rect 6022 6301 6052 6304
rect 6031 6297 6038 6301
rect 6038 6296 6039 6297
rect 5997 6290 6007 6296
rect 5756 6282 5791 6290
rect 5756 6256 5757 6282
rect 5764 6256 5791 6282
rect 5699 6238 5729 6252
rect 5756 6248 5791 6256
rect 5793 6282 5834 6290
rect 5793 6256 5808 6282
rect 5815 6256 5834 6282
rect 5898 6278 5929 6290
rect 5944 6278 6047 6290
rect 6059 6280 6085 6306
rect 6100 6301 6130 6312
rect 6162 6308 6224 6324
rect 6162 6306 6208 6308
rect 6162 6290 6224 6306
rect 6236 6290 6242 6338
rect 6245 6330 6325 6338
rect 6245 6328 6264 6330
rect 6279 6328 6313 6330
rect 6245 6312 6325 6328
rect 6245 6290 6264 6312
rect 6279 6296 6309 6312
rect 6337 6306 6343 6380
rect 6346 6306 6365 6450
rect 6380 6306 6386 6450
rect 6395 6380 6408 6450
rect 6460 6446 6482 6450
rect 6453 6424 6482 6438
rect 6535 6424 6551 6438
rect 6589 6434 6595 6436
rect 6602 6434 6710 6450
rect 6717 6434 6723 6436
rect 6731 6434 6746 6450
rect 6812 6444 6831 6447
rect 6453 6422 6551 6424
rect 6578 6422 6746 6434
rect 6761 6424 6777 6438
rect 6812 6425 6834 6444
rect 6844 6438 6860 6439
rect 6843 6436 6860 6438
rect 6844 6431 6860 6436
rect 6834 6424 6840 6425
rect 6843 6424 6872 6431
rect 6761 6423 6872 6424
rect 6761 6422 6878 6423
rect 6437 6414 6488 6422
rect 6535 6414 6569 6422
rect 6437 6402 6462 6414
rect 6469 6402 6488 6414
rect 6542 6412 6569 6414
rect 6578 6412 6799 6422
rect 6834 6419 6840 6422
rect 6542 6408 6799 6412
rect 6437 6394 6488 6402
rect 6535 6394 6799 6408
rect 6843 6414 6878 6422
rect 6389 6346 6408 6380
rect 6453 6386 6482 6394
rect 6453 6380 6470 6386
rect 6453 6378 6487 6380
rect 6535 6378 6551 6394
rect 6552 6384 6760 6394
rect 6761 6384 6777 6394
rect 6825 6390 6840 6405
rect 6843 6402 6844 6414
rect 6851 6402 6878 6414
rect 6843 6394 6878 6402
rect 6843 6393 6872 6394
rect 6563 6380 6777 6384
rect 6578 6378 6777 6380
rect 6812 6380 6825 6390
rect 6843 6380 6860 6393
rect 6812 6378 6860 6380
rect 6454 6374 6487 6378
rect 6450 6372 6487 6374
rect 6450 6371 6517 6372
rect 6450 6366 6481 6371
rect 6487 6366 6517 6371
rect 6450 6362 6517 6366
rect 6423 6359 6517 6362
rect 6423 6352 6472 6359
rect 6423 6346 6453 6352
rect 6472 6347 6477 6352
rect 6389 6330 6469 6346
rect 6481 6338 6517 6359
rect 6578 6354 6767 6378
rect 6812 6377 6859 6378
rect 6825 6372 6859 6377
rect 6593 6351 6767 6354
rect 6586 6348 6767 6351
rect 6795 6371 6859 6372
rect 6389 6328 6408 6330
rect 6423 6328 6457 6330
rect 6389 6312 6469 6328
rect 6389 6306 6408 6312
rect 6105 6280 6208 6290
rect 6059 6278 6208 6280
rect 6229 6278 6264 6290
rect 5898 6276 6060 6278
rect 5910 6256 5929 6276
rect 5944 6274 5974 6276
rect 5793 6248 5834 6256
rect 5916 6252 5929 6256
rect 5981 6260 6060 6276
rect 6092 6276 6264 6278
rect 6092 6260 6171 6276
rect 6178 6274 6208 6276
rect 5756 6238 5785 6248
rect 5799 6238 5828 6248
rect 5843 6238 5873 6252
rect 5916 6238 5959 6252
rect 5981 6248 6171 6260
rect 6236 6256 6242 6276
rect 5966 6238 5996 6248
rect 5997 6238 6155 6248
rect 6159 6238 6189 6248
rect 6193 6238 6223 6252
rect 6251 6238 6264 6276
rect 6336 6290 6365 6306
rect 6379 6290 6408 6306
rect 6423 6296 6453 6312
rect 6481 6290 6487 6338
rect 6490 6332 6509 6338
rect 6524 6332 6554 6340
rect 6490 6324 6554 6332
rect 6490 6308 6570 6324
rect 6586 6317 6648 6348
rect 6664 6317 6726 6348
rect 6795 6346 6844 6371
rect 6859 6346 6889 6362
rect 6758 6332 6788 6340
rect 6795 6338 6905 6346
rect 6758 6324 6803 6332
rect 6490 6306 6509 6308
rect 6524 6306 6570 6308
rect 6490 6290 6570 6306
rect 6597 6304 6632 6317
rect 6673 6314 6710 6317
rect 6673 6312 6715 6314
rect 6602 6301 6632 6304
rect 6611 6297 6618 6301
rect 6618 6296 6619 6297
rect 6577 6290 6587 6296
rect 6336 6282 6371 6290
rect 6336 6256 6337 6282
rect 6344 6256 6371 6282
rect 6279 6238 6309 6252
rect 6336 6248 6371 6256
rect 6373 6282 6414 6290
rect 6373 6256 6388 6282
rect 6395 6256 6414 6282
rect 6478 6278 6509 6290
rect 6524 6278 6627 6290
rect 6639 6280 6665 6306
rect 6680 6301 6710 6312
rect 6742 6308 6804 6324
rect 6742 6306 6788 6308
rect 6742 6290 6804 6306
rect 6816 6290 6822 6338
rect 6825 6330 6905 6338
rect 6825 6328 6844 6330
rect 6859 6328 6893 6330
rect 6825 6312 6905 6328
rect 6825 6290 6844 6312
rect 6859 6296 6889 6312
rect 6917 6306 6923 6380
rect 6926 6306 6945 6450
rect 6960 6306 6966 6450
rect 6975 6380 6988 6450
rect 7040 6446 7062 6450
rect 7033 6424 7062 6438
rect 7115 6424 7131 6438
rect 7169 6434 7175 6436
rect 7182 6434 7290 6450
rect 7297 6434 7303 6436
rect 7311 6434 7326 6450
rect 7392 6444 7411 6447
rect 7033 6422 7131 6424
rect 7158 6422 7326 6434
rect 7341 6424 7357 6438
rect 7392 6425 7414 6444
rect 7424 6438 7440 6439
rect 7423 6436 7440 6438
rect 7424 6431 7440 6436
rect 7414 6424 7420 6425
rect 7423 6424 7452 6431
rect 7341 6423 7452 6424
rect 7341 6422 7458 6423
rect 7017 6414 7068 6422
rect 7115 6414 7149 6422
rect 7017 6402 7042 6414
rect 7049 6402 7068 6414
rect 7122 6412 7149 6414
rect 7158 6412 7379 6422
rect 7414 6419 7420 6422
rect 7122 6408 7379 6412
rect 7017 6394 7068 6402
rect 7115 6394 7379 6408
rect 7423 6414 7458 6422
rect 6969 6346 6988 6380
rect 7033 6386 7062 6394
rect 7033 6380 7050 6386
rect 7033 6378 7067 6380
rect 7115 6378 7131 6394
rect 7132 6384 7340 6394
rect 7341 6384 7357 6394
rect 7405 6390 7420 6405
rect 7423 6402 7424 6414
rect 7431 6402 7458 6414
rect 7423 6394 7458 6402
rect 7423 6393 7452 6394
rect 7143 6380 7357 6384
rect 7158 6378 7357 6380
rect 7392 6380 7405 6390
rect 7423 6380 7440 6393
rect 7392 6378 7440 6380
rect 7034 6374 7067 6378
rect 7030 6372 7067 6374
rect 7030 6371 7097 6372
rect 7030 6366 7061 6371
rect 7067 6366 7097 6371
rect 7030 6362 7097 6366
rect 7003 6359 7097 6362
rect 7003 6352 7052 6359
rect 7003 6346 7033 6352
rect 7052 6347 7057 6352
rect 6969 6330 7049 6346
rect 7061 6338 7097 6359
rect 7158 6354 7347 6378
rect 7392 6377 7439 6378
rect 7405 6372 7439 6377
rect 7173 6351 7347 6354
rect 7166 6348 7347 6351
rect 7375 6371 7439 6372
rect 6969 6328 6988 6330
rect 7003 6328 7037 6330
rect 6969 6312 7049 6328
rect 6969 6306 6988 6312
rect 6685 6280 6788 6290
rect 6639 6278 6788 6280
rect 6809 6278 6844 6290
rect 6478 6276 6640 6278
rect 6490 6256 6509 6276
rect 6524 6274 6554 6276
rect 6373 6248 6414 6256
rect 6496 6252 6509 6256
rect 6561 6260 6640 6276
rect 6672 6276 6844 6278
rect 6672 6260 6751 6276
rect 6758 6274 6788 6276
rect 6336 6238 6365 6248
rect 6379 6238 6408 6248
rect 6423 6238 6453 6252
rect 6496 6238 6539 6252
rect 6561 6248 6751 6260
rect 6816 6256 6822 6276
rect 6546 6238 6576 6248
rect 6577 6238 6735 6248
rect 6739 6238 6769 6248
rect 6773 6238 6803 6252
rect 6831 6238 6844 6276
rect 6916 6290 6945 6306
rect 6959 6290 6988 6306
rect 7003 6296 7033 6312
rect 7061 6290 7067 6338
rect 7070 6332 7089 6338
rect 7104 6332 7134 6340
rect 7070 6324 7134 6332
rect 7070 6308 7150 6324
rect 7166 6317 7228 6348
rect 7244 6317 7306 6348
rect 7375 6346 7424 6371
rect 7439 6346 7469 6362
rect 7338 6332 7368 6340
rect 7375 6338 7485 6346
rect 7338 6324 7383 6332
rect 7070 6306 7089 6308
rect 7104 6306 7150 6308
rect 7070 6290 7150 6306
rect 7177 6304 7212 6317
rect 7253 6314 7290 6317
rect 7253 6312 7295 6314
rect 7182 6301 7212 6304
rect 7191 6297 7198 6301
rect 7198 6296 7199 6297
rect 7157 6290 7167 6296
rect 6916 6282 6951 6290
rect 6916 6256 6917 6282
rect 6924 6256 6951 6282
rect 6859 6238 6889 6252
rect 6916 6248 6951 6256
rect 6953 6282 6994 6290
rect 6953 6256 6968 6282
rect 6975 6256 6994 6282
rect 7058 6278 7089 6290
rect 7104 6278 7207 6290
rect 7219 6280 7245 6306
rect 7260 6301 7290 6312
rect 7322 6308 7384 6324
rect 7322 6306 7368 6308
rect 7322 6290 7384 6306
rect 7396 6290 7402 6338
rect 7405 6330 7485 6338
rect 7405 6328 7424 6330
rect 7439 6328 7473 6330
rect 7405 6312 7485 6328
rect 7405 6290 7424 6312
rect 7439 6296 7469 6312
rect 7497 6306 7503 6380
rect 7506 6306 7525 6450
rect 7540 6306 7546 6450
rect 7555 6380 7568 6450
rect 7620 6446 7642 6450
rect 7613 6424 7642 6438
rect 7695 6424 7711 6438
rect 7749 6434 7755 6436
rect 7762 6434 7870 6450
rect 7877 6434 7883 6436
rect 7891 6434 7906 6450
rect 7972 6444 7991 6447
rect 7613 6422 7711 6424
rect 7738 6422 7906 6434
rect 7921 6424 7937 6438
rect 7972 6425 7994 6444
rect 8004 6438 8020 6439
rect 8003 6436 8020 6438
rect 8004 6431 8020 6436
rect 7994 6424 8000 6425
rect 8003 6424 8032 6431
rect 7921 6423 8032 6424
rect 7921 6422 8038 6423
rect 7597 6414 7648 6422
rect 7695 6414 7729 6422
rect 7597 6402 7622 6414
rect 7629 6402 7648 6414
rect 7702 6412 7729 6414
rect 7738 6412 7959 6422
rect 7994 6419 8000 6422
rect 7702 6408 7959 6412
rect 7597 6394 7648 6402
rect 7695 6394 7959 6408
rect 8003 6414 8038 6422
rect 7549 6346 7568 6380
rect 7613 6386 7642 6394
rect 7613 6380 7630 6386
rect 7613 6378 7647 6380
rect 7695 6378 7711 6394
rect 7712 6384 7920 6394
rect 7921 6384 7937 6394
rect 7985 6390 8000 6405
rect 8003 6402 8004 6414
rect 8011 6402 8038 6414
rect 8003 6394 8038 6402
rect 8003 6393 8032 6394
rect 7723 6380 7937 6384
rect 7738 6378 7937 6380
rect 7972 6380 7985 6390
rect 8003 6380 8020 6393
rect 7972 6378 8020 6380
rect 7614 6374 7647 6378
rect 7610 6372 7647 6374
rect 7610 6371 7677 6372
rect 7610 6366 7641 6371
rect 7647 6366 7677 6371
rect 7610 6362 7677 6366
rect 7583 6359 7677 6362
rect 7583 6352 7632 6359
rect 7583 6346 7613 6352
rect 7632 6347 7637 6352
rect 7549 6330 7629 6346
rect 7641 6338 7677 6359
rect 7738 6354 7927 6378
rect 7972 6377 8019 6378
rect 7985 6372 8019 6377
rect 7753 6351 7927 6354
rect 7746 6348 7927 6351
rect 7955 6371 8019 6372
rect 7549 6328 7568 6330
rect 7583 6328 7617 6330
rect 7549 6312 7629 6328
rect 7549 6306 7568 6312
rect 7265 6280 7368 6290
rect 7219 6278 7368 6280
rect 7389 6278 7424 6290
rect 7058 6276 7220 6278
rect 7070 6256 7089 6276
rect 7104 6274 7134 6276
rect 6953 6248 6994 6256
rect 7076 6252 7089 6256
rect 7141 6260 7220 6276
rect 7252 6276 7424 6278
rect 7252 6260 7331 6276
rect 7338 6274 7368 6276
rect 6916 6238 6945 6248
rect 6959 6238 6988 6248
rect 7003 6238 7033 6252
rect 7076 6238 7119 6252
rect 7141 6248 7331 6260
rect 7396 6256 7402 6276
rect 7126 6238 7156 6248
rect 7157 6238 7315 6248
rect 7319 6238 7349 6248
rect 7353 6238 7383 6252
rect 7411 6238 7424 6276
rect 7496 6290 7525 6306
rect 7539 6290 7568 6306
rect 7583 6296 7613 6312
rect 7641 6290 7647 6338
rect 7650 6332 7669 6338
rect 7684 6332 7714 6340
rect 7650 6324 7714 6332
rect 7650 6308 7730 6324
rect 7746 6317 7808 6348
rect 7824 6317 7886 6348
rect 7955 6346 8004 6371
rect 8019 6346 8049 6362
rect 7918 6332 7948 6340
rect 7955 6338 8065 6346
rect 7918 6324 7963 6332
rect 7650 6306 7669 6308
rect 7684 6306 7730 6308
rect 7650 6290 7730 6306
rect 7757 6304 7792 6317
rect 7833 6314 7870 6317
rect 7833 6312 7875 6314
rect 7762 6301 7792 6304
rect 7771 6297 7778 6301
rect 7778 6296 7779 6297
rect 7737 6290 7747 6296
rect 7496 6282 7531 6290
rect 7496 6256 7497 6282
rect 7504 6256 7531 6282
rect 7439 6238 7469 6252
rect 7496 6248 7531 6256
rect 7533 6282 7574 6290
rect 7533 6256 7548 6282
rect 7555 6256 7574 6282
rect 7638 6278 7669 6290
rect 7684 6278 7787 6290
rect 7799 6280 7825 6306
rect 7840 6301 7870 6312
rect 7902 6308 7964 6324
rect 7902 6306 7948 6308
rect 7902 6290 7964 6306
rect 7976 6290 7982 6338
rect 7985 6330 8065 6338
rect 7985 6328 8004 6330
rect 8019 6328 8053 6330
rect 7985 6312 8065 6328
rect 7985 6290 8004 6312
rect 8019 6296 8049 6312
rect 8077 6306 8083 6380
rect 8086 6306 8105 6450
rect 8120 6306 8126 6450
rect 8135 6380 8148 6450
rect 8200 6446 8222 6450
rect 8193 6424 8222 6438
rect 8275 6424 8291 6438
rect 8329 6434 8335 6436
rect 8342 6434 8450 6450
rect 8457 6434 8463 6436
rect 8471 6434 8486 6450
rect 8552 6444 8571 6447
rect 8193 6422 8291 6424
rect 8318 6422 8486 6434
rect 8501 6424 8517 6438
rect 8552 6425 8574 6444
rect 8584 6438 8600 6439
rect 8583 6436 8600 6438
rect 8584 6431 8600 6436
rect 8574 6424 8580 6425
rect 8583 6424 8612 6431
rect 8501 6423 8612 6424
rect 8501 6422 8618 6423
rect 8177 6414 8228 6422
rect 8275 6414 8309 6422
rect 8177 6402 8202 6414
rect 8209 6402 8228 6414
rect 8282 6412 8309 6414
rect 8318 6412 8539 6422
rect 8574 6419 8580 6422
rect 8282 6408 8539 6412
rect 8177 6394 8228 6402
rect 8275 6394 8539 6408
rect 8583 6414 8618 6422
rect 8129 6346 8148 6380
rect 8193 6386 8222 6394
rect 8193 6380 8210 6386
rect 8193 6378 8227 6380
rect 8275 6378 8291 6394
rect 8292 6384 8500 6394
rect 8501 6384 8517 6394
rect 8565 6390 8580 6405
rect 8583 6402 8584 6414
rect 8591 6402 8618 6414
rect 8583 6394 8618 6402
rect 8583 6393 8612 6394
rect 8303 6380 8517 6384
rect 8318 6378 8517 6380
rect 8552 6380 8565 6390
rect 8583 6380 8600 6393
rect 8552 6378 8600 6380
rect 8194 6374 8227 6378
rect 8190 6372 8227 6374
rect 8190 6371 8257 6372
rect 8190 6366 8221 6371
rect 8227 6366 8257 6371
rect 8190 6362 8257 6366
rect 8163 6359 8257 6362
rect 8163 6352 8212 6359
rect 8163 6346 8193 6352
rect 8212 6347 8217 6352
rect 8129 6330 8209 6346
rect 8221 6338 8257 6359
rect 8318 6354 8507 6378
rect 8552 6377 8599 6378
rect 8565 6372 8599 6377
rect 8333 6351 8507 6354
rect 8326 6348 8507 6351
rect 8535 6371 8599 6372
rect 8129 6328 8148 6330
rect 8163 6328 8197 6330
rect 8129 6312 8209 6328
rect 8129 6306 8148 6312
rect 7845 6280 7948 6290
rect 7799 6278 7948 6280
rect 7969 6278 8004 6290
rect 7638 6276 7800 6278
rect 7650 6256 7669 6276
rect 7684 6274 7714 6276
rect 7533 6248 7574 6256
rect 7656 6252 7669 6256
rect 7721 6260 7800 6276
rect 7832 6276 8004 6278
rect 7832 6260 7911 6276
rect 7918 6274 7948 6276
rect 7496 6238 7525 6248
rect 7539 6238 7568 6248
rect 7583 6238 7613 6252
rect 7656 6238 7699 6252
rect 7721 6248 7911 6260
rect 7976 6256 7982 6276
rect 7706 6238 7736 6248
rect 7737 6238 7895 6248
rect 7899 6238 7929 6248
rect 7933 6238 7963 6252
rect 7991 6238 8004 6276
rect 8076 6290 8105 6306
rect 8119 6290 8148 6306
rect 8163 6296 8193 6312
rect 8221 6290 8227 6338
rect 8230 6332 8249 6338
rect 8264 6332 8294 6340
rect 8230 6324 8294 6332
rect 8230 6308 8310 6324
rect 8326 6317 8388 6348
rect 8404 6317 8466 6348
rect 8535 6346 8584 6371
rect 8599 6346 8629 6362
rect 8498 6332 8528 6340
rect 8535 6338 8645 6346
rect 8498 6324 8543 6332
rect 8230 6306 8249 6308
rect 8264 6306 8310 6308
rect 8230 6290 8310 6306
rect 8337 6304 8372 6317
rect 8413 6314 8450 6317
rect 8413 6312 8455 6314
rect 8342 6301 8372 6304
rect 8351 6297 8358 6301
rect 8358 6296 8359 6297
rect 8317 6290 8327 6296
rect 8076 6282 8111 6290
rect 8076 6256 8077 6282
rect 8084 6256 8111 6282
rect 8019 6238 8049 6252
rect 8076 6248 8111 6256
rect 8113 6282 8154 6290
rect 8113 6256 8128 6282
rect 8135 6256 8154 6282
rect 8218 6278 8249 6290
rect 8264 6278 8367 6290
rect 8379 6280 8405 6306
rect 8420 6301 8450 6312
rect 8482 6308 8544 6324
rect 8482 6306 8528 6308
rect 8482 6290 8544 6306
rect 8556 6290 8562 6338
rect 8565 6330 8645 6338
rect 8565 6328 8584 6330
rect 8599 6328 8633 6330
rect 8565 6312 8645 6328
rect 8565 6290 8584 6312
rect 8599 6296 8629 6312
rect 8657 6306 8663 6380
rect 8666 6306 8685 6450
rect 8700 6306 8706 6450
rect 8715 6380 8728 6450
rect 8780 6446 8802 6450
rect 8773 6424 8802 6438
rect 8855 6424 8871 6438
rect 8909 6434 8915 6436
rect 8922 6434 9030 6450
rect 9037 6434 9043 6436
rect 9051 6434 9066 6450
rect 9132 6444 9151 6447
rect 8773 6422 8871 6424
rect 8898 6422 9066 6434
rect 9081 6424 9097 6438
rect 9132 6425 9154 6444
rect 9164 6438 9180 6439
rect 9163 6436 9180 6438
rect 9164 6431 9180 6436
rect 9154 6424 9160 6425
rect 9163 6424 9192 6431
rect 9081 6423 9192 6424
rect 9081 6422 9198 6423
rect 8757 6414 8808 6422
rect 8855 6414 8889 6422
rect 8757 6402 8782 6414
rect 8789 6402 8808 6414
rect 8862 6412 8889 6414
rect 8898 6412 9119 6422
rect 9154 6419 9160 6422
rect 8862 6408 9119 6412
rect 8757 6394 8808 6402
rect 8855 6394 9119 6408
rect 9163 6414 9198 6422
rect 8709 6346 8728 6380
rect 8773 6386 8802 6394
rect 8773 6380 8790 6386
rect 8773 6378 8807 6380
rect 8855 6378 8871 6394
rect 8872 6384 9080 6394
rect 9081 6384 9097 6394
rect 9145 6390 9160 6405
rect 9163 6402 9164 6414
rect 9171 6402 9198 6414
rect 9163 6394 9198 6402
rect 9163 6393 9192 6394
rect 8883 6380 9097 6384
rect 8898 6378 9097 6380
rect 9132 6380 9145 6390
rect 9163 6380 9180 6393
rect 9132 6378 9180 6380
rect 8774 6374 8807 6378
rect 8770 6372 8807 6374
rect 8770 6371 8837 6372
rect 8770 6366 8801 6371
rect 8807 6366 8837 6371
rect 8770 6362 8837 6366
rect 8743 6359 8837 6362
rect 8743 6352 8792 6359
rect 8743 6346 8773 6352
rect 8792 6347 8797 6352
rect 8709 6330 8789 6346
rect 8801 6338 8837 6359
rect 8898 6354 9087 6378
rect 9132 6377 9179 6378
rect 9145 6372 9179 6377
rect 8913 6351 9087 6354
rect 8906 6348 9087 6351
rect 9115 6371 9179 6372
rect 8709 6328 8728 6330
rect 8743 6328 8777 6330
rect 8709 6312 8789 6328
rect 8709 6306 8728 6312
rect 8425 6280 8528 6290
rect 8379 6278 8528 6280
rect 8549 6278 8584 6290
rect 8218 6276 8380 6278
rect 8230 6256 8249 6276
rect 8264 6274 8294 6276
rect 8113 6248 8154 6256
rect 8236 6252 8249 6256
rect 8301 6260 8380 6276
rect 8412 6276 8584 6278
rect 8412 6260 8491 6276
rect 8498 6274 8528 6276
rect 8076 6238 8105 6248
rect 8119 6238 8148 6248
rect 8163 6238 8193 6252
rect 8236 6238 8279 6252
rect 8301 6248 8491 6260
rect 8556 6256 8562 6276
rect 8286 6238 8316 6248
rect 8317 6238 8475 6248
rect 8479 6238 8509 6248
rect 8513 6238 8543 6252
rect 8571 6238 8584 6276
rect 8656 6290 8685 6306
rect 8699 6290 8728 6306
rect 8743 6296 8773 6312
rect 8801 6290 8807 6338
rect 8810 6332 8829 6338
rect 8844 6332 8874 6340
rect 8810 6324 8874 6332
rect 8810 6308 8890 6324
rect 8906 6317 8968 6348
rect 8984 6317 9046 6348
rect 9115 6346 9164 6371
rect 9179 6346 9209 6362
rect 9078 6332 9108 6340
rect 9115 6338 9225 6346
rect 9078 6324 9123 6332
rect 8810 6306 8829 6308
rect 8844 6306 8890 6308
rect 8810 6290 8890 6306
rect 8917 6304 8952 6317
rect 8993 6314 9030 6317
rect 8993 6312 9035 6314
rect 8922 6301 8952 6304
rect 8931 6297 8938 6301
rect 8938 6296 8939 6297
rect 8897 6290 8907 6296
rect 8656 6282 8691 6290
rect 8656 6256 8657 6282
rect 8664 6256 8691 6282
rect 8599 6238 8629 6252
rect 8656 6248 8691 6256
rect 8693 6282 8734 6290
rect 8693 6256 8708 6282
rect 8715 6256 8734 6282
rect 8798 6278 8829 6290
rect 8844 6278 8947 6290
rect 8959 6280 8985 6306
rect 9000 6301 9030 6312
rect 9062 6308 9124 6324
rect 9062 6306 9108 6308
rect 9062 6290 9124 6306
rect 9136 6290 9142 6338
rect 9145 6330 9225 6338
rect 9145 6328 9164 6330
rect 9179 6328 9213 6330
rect 9145 6312 9225 6328
rect 9145 6290 9164 6312
rect 9179 6296 9209 6312
rect 9237 6306 9243 6380
rect 9246 6306 9265 6450
rect 9280 6306 9286 6450
rect 9295 6380 9308 6450
rect 9360 6446 9382 6450
rect 9353 6424 9382 6438
rect 9435 6424 9451 6438
rect 9489 6434 9495 6436
rect 9502 6434 9610 6450
rect 9617 6434 9623 6436
rect 9631 6434 9646 6450
rect 9712 6444 9731 6447
rect 9353 6422 9451 6424
rect 9478 6422 9646 6434
rect 9661 6424 9677 6438
rect 9712 6425 9734 6444
rect 9744 6438 9760 6439
rect 9743 6436 9760 6438
rect 9744 6431 9760 6436
rect 9734 6424 9740 6425
rect 9743 6424 9772 6431
rect 9661 6423 9772 6424
rect 9661 6422 9778 6423
rect 9337 6414 9388 6422
rect 9435 6414 9469 6422
rect 9337 6402 9362 6414
rect 9369 6402 9388 6414
rect 9442 6412 9469 6414
rect 9478 6412 9699 6422
rect 9734 6419 9740 6422
rect 9442 6408 9699 6412
rect 9337 6394 9388 6402
rect 9435 6394 9699 6408
rect 9743 6414 9778 6422
rect 9289 6346 9308 6380
rect 9353 6386 9382 6394
rect 9353 6380 9370 6386
rect 9353 6378 9387 6380
rect 9435 6378 9451 6394
rect 9452 6384 9660 6394
rect 9661 6384 9677 6394
rect 9725 6390 9740 6405
rect 9743 6402 9744 6414
rect 9751 6402 9778 6414
rect 9743 6394 9778 6402
rect 9743 6393 9772 6394
rect 9463 6380 9677 6384
rect 9478 6378 9677 6380
rect 9712 6380 9725 6390
rect 9743 6380 9760 6393
rect 9712 6378 9760 6380
rect 9354 6374 9387 6378
rect 9350 6372 9387 6374
rect 9350 6371 9417 6372
rect 9350 6366 9381 6371
rect 9387 6366 9417 6371
rect 9350 6362 9417 6366
rect 9323 6359 9417 6362
rect 9323 6352 9372 6359
rect 9323 6346 9353 6352
rect 9372 6347 9377 6352
rect 9289 6330 9369 6346
rect 9381 6338 9417 6359
rect 9478 6354 9667 6378
rect 9712 6377 9759 6378
rect 9725 6372 9759 6377
rect 9493 6351 9667 6354
rect 9486 6348 9667 6351
rect 9695 6371 9759 6372
rect 9289 6328 9308 6330
rect 9323 6328 9357 6330
rect 9289 6312 9369 6328
rect 9289 6306 9308 6312
rect 9005 6280 9108 6290
rect 8959 6278 9108 6280
rect 9129 6278 9164 6290
rect 8798 6276 8960 6278
rect 8810 6256 8829 6276
rect 8844 6274 8874 6276
rect 8693 6248 8734 6256
rect 8816 6252 8829 6256
rect 8881 6260 8960 6276
rect 8992 6276 9164 6278
rect 8992 6260 9071 6276
rect 9078 6274 9108 6276
rect 8656 6238 8685 6248
rect 8699 6238 8728 6248
rect 8743 6238 8773 6252
rect 8816 6238 8859 6252
rect 8881 6248 9071 6260
rect 9136 6256 9142 6276
rect 8866 6238 8896 6248
rect 8897 6238 9055 6248
rect 9059 6238 9089 6248
rect 9093 6238 9123 6252
rect 9151 6238 9164 6276
rect 9236 6290 9265 6306
rect 9279 6290 9308 6306
rect 9323 6296 9353 6312
rect 9381 6290 9387 6338
rect 9390 6332 9409 6338
rect 9424 6332 9454 6340
rect 9390 6324 9454 6332
rect 9390 6308 9470 6324
rect 9486 6317 9548 6348
rect 9564 6317 9626 6348
rect 9695 6346 9744 6371
rect 9759 6346 9789 6362
rect 9658 6332 9688 6340
rect 9695 6338 9805 6346
rect 9658 6324 9703 6332
rect 9390 6306 9409 6308
rect 9424 6306 9470 6308
rect 9390 6290 9470 6306
rect 9497 6304 9532 6317
rect 9573 6314 9610 6317
rect 9573 6312 9615 6314
rect 9502 6301 9532 6304
rect 9511 6297 9518 6301
rect 9518 6296 9519 6297
rect 9477 6290 9487 6296
rect 9236 6282 9271 6290
rect 9236 6256 9237 6282
rect 9244 6256 9271 6282
rect 9179 6238 9209 6252
rect 9236 6248 9271 6256
rect 9273 6282 9314 6290
rect 9273 6256 9288 6282
rect 9295 6256 9314 6282
rect 9378 6278 9409 6290
rect 9424 6278 9527 6290
rect 9539 6280 9565 6306
rect 9580 6301 9610 6312
rect 9642 6308 9704 6324
rect 9642 6306 9688 6308
rect 9642 6290 9704 6306
rect 9716 6290 9722 6338
rect 9725 6330 9805 6338
rect 9725 6328 9744 6330
rect 9759 6328 9793 6330
rect 9725 6312 9805 6328
rect 9725 6290 9744 6312
rect 9759 6296 9789 6312
rect 9817 6306 9823 6380
rect 9826 6306 9845 6450
rect 9860 6306 9866 6450
rect 9875 6380 9888 6450
rect 9940 6446 9962 6450
rect 9933 6424 9962 6438
rect 10015 6424 10031 6438
rect 10069 6434 10075 6436
rect 10082 6434 10190 6450
rect 10197 6434 10203 6436
rect 10211 6434 10226 6450
rect 10292 6444 10311 6447
rect 9933 6422 10031 6424
rect 10058 6422 10226 6434
rect 10241 6424 10257 6438
rect 10292 6425 10314 6444
rect 10324 6438 10340 6439
rect 10323 6436 10340 6438
rect 10324 6431 10340 6436
rect 10314 6424 10320 6425
rect 10323 6424 10352 6431
rect 10241 6423 10352 6424
rect 10241 6422 10358 6423
rect 9917 6414 9968 6422
rect 10015 6414 10049 6422
rect 9917 6402 9942 6414
rect 9949 6402 9968 6414
rect 10022 6412 10049 6414
rect 10058 6412 10279 6422
rect 10314 6419 10320 6422
rect 10022 6408 10279 6412
rect 9917 6394 9968 6402
rect 10015 6394 10279 6408
rect 10323 6414 10358 6422
rect 9869 6346 9888 6380
rect 9933 6386 9962 6394
rect 9933 6380 9950 6386
rect 9933 6378 9967 6380
rect 10015 6378 10031 6394
rect 10032 6384 10240 6394
rect 10241 6384 10257 6394
rect 10305 6390 10320 6405
rect 10323 6402 10324 6414
rect 10331 6402 10358 6414
rect 10323 6394 10358 6402
rect 10323 6393 10352 6394
rect 10043 6380 10257 6384
rect 10058 6378 10257 6380
rect 10292 6380 10305 6390
rect 10323 6380 10340 6393
rect 10292 6378 10340 6380
rect 9934 6374 9967 6378
rect 9930 6372 9967 6374
rect 9930 6371 9997 6372
rect 9930 6366 9961 6371
rect 9967 6366 9997 6371
rect 9930 6362 9997 6366
rect 9903 6359 9997 6362
rect 9903 6352 9952 6359
rect 9903 6346 9933 6352
rect 9952 6347 9957 6352
rect 9869 6330 9949 6346
rect 9961 6338 9997 6359
rect 10058 6354 10247 6378
rect 10292 6377 10339 6378
rect 10305 6372 10339 6377
rect 10073 6351 10247 6354
rect 10066 6348 10247 6351
rect 10275 6371 10339 6372
rect 9869 6328 9888 6330
rect 9903 6328 9937 6330
rect 9869 6312 9949 6328
rect 9869 6306 9888 6312
rect 9585 6280 9688 6290
rect 9539 6278 9688 6280
rect 9709 6278 9744 6290
rect 9378 6276 9540 6278
rect 9390 6256 9409 6276
rect 9424 6274 9454 6276
rect 9273 6248 9314 6256
rect 9396 6252 9409 6256
rect 9461 6260 9540 6276
rect 9572 6276 9744 6278
rect 9572 6260 9651 6276
rect 9658 6274 9688 6276
rect 9236 6238 9265 6248
rect 9279 6238 9308 6248
rect 9323 6238 9353 6252
rect 9396 6238 9439 6252
rect 9461 6248 9651 6260
rect 9716 6256 9722 6276
rect 9446 6238 9476 6248
rect 9477 6238 9635 6248
rect 9639 6238 9669 6248
rect 9673 6238 9703 6252
rect 9731 6238 9744 6276
rect 9816 6290 9845 6306
rect 9859 6290 9888 6306
rect 9903 6296 9933 6312
rect 9961 6290 9967 6338
rect 9970 6332 9989 6338
rect 10004 6332 10034 6340
rect 9970 6324 10034 6332
rect 9970 6308 10050 6324
rect 10066 6317 10128 6348
rect 10144 6317 10206 6348
rect 10275 6346 10324 6371
rect 10339 6346 10369 6362
rect 10238 6332 10268 6340
rect 10275 6338 10385 6346
rect 10238 6324 10283 6332
rect 9970 6306 9989 6308
rect 10004 6306 10050 6308
rect 9970 6290 10050 6306
rect 10077 6304 10112 6317
rect 10153 6314 10190 6317
rect 10153 6312 10195 6314
rect 10082 6301 10112 6304
rect 10091 6297 10098 6301
rect 10098 6296 10099 6297
rect 10057 6290 10067 6296
rect 9816 6282 9851 6290
rect 9816 6256 9817 6282
rect 9824 6256 9851 6282
rect 9759 6238 9789 6252
rect 9816 6248 9851 6256
rect 9853 6282 9894 6290
rect 9853 6256 9868 6282
rect 9875 6256 9894 6282
rect 9958 6278 9989 6290
rect 10004 6278 10107 6290
rect 10119 6280 10145 6306
rect 10160 6301 10190 6312
rect 10222 6308 10284 6324
rect 10222 6306 10268 6308
rect 10222 6290 10284 6306
rect 10296 6290 10302 6338
rect 10305 6330 10385 6338
rect 10305 6328 10324 6330
rect 10339 6328 10373 6330
rect 10305 6312 10385 6328
rect 10305 6290 10324 6312
rect 10339 6296 10369 6312
rect 10397 6306 10403 6380
rect 10406 6306 10425 6450
rect 10440 6306 10446 6450
rect 10455 6380 10468 6450
rect 10520 6446 10542 6450
rect 10513 6424 10542 6438
rect 10595 6424 10611 6438
rect 10649 6434 10655 6436
rect 10662 6434 10770 6450
rect 10777 6434 10783 6436
rect 10791 6434 10806 6450
rect 10872 6444 10891 6447
rect 10513 6422 10611 6424
rect 10638 6422 10806 6434
rect 10821 6424 10837 6438
rect 10872 6425 10894 6444
rect 10904 6438 10920 6439
rect 10903 6436 10920 6438
rect 10904 6431 10920 6436
rect 10894 6424 10900 6425
rect 10903 6424 10932 6431
rect 10821 6423 10932 6424
rect 10821 6422 10938 6423
rect 10497 6414 10548 6422
rect 10595 6414 10629 6422
rect 10497 6402 10522 6414
rect 10529 6402 10548 6414
rect 10602 6412 10629 6414
rect 10638 6412 10859 6422
rect 10894 6419 10900 6422
rect 10602 6408 10859 6412
rect 10497 6394 10548 6402
rect 10595 6394 10859 6408
rect 10903 6414 10938 6422
rect 10449 6346 10468 6380
rect 10513 6386 10542 6394
rect 10513 6380 10530 6386
rect 10513 6378 10547 6380
rect 10595 6378 10611 6394
rect 10612 6384 10820 6394
rect 10821 6384 10837 6394
rect 10885 6390 10900 6405
rect 10903 6402 10904 6414
rect 10911 6402 10938 6414
rect 10903 6394 10938 6402
rect 10903 6393 10932 6394
rect 10623 6380 10837 6384
rect 10638 6378 10837 6380
rect 10872 6380 10885 6390
rect 10903 6380 10920 6393
rect 10872 6378 10920 6380
rect 10514 6374 10547 6378
rect 10510 6372 10547 6374
rect 10510 6371 10577 6372
rect 10510 6366 10541 6371
rect 10547 6366 10577 6371
rect 10510 6362 10577 6366
rect 10483 6359 10577 6362
rect 10483 6352 10532 6359
rect 10483 6346 10513 6352
rect 10532 6347 10537 6352
rect 10449 6330 10529 6346
rect 10541 6338 10577 6359
rect 10638 6354 10827 6378
rect 10872 6377 10919 6378
rect 10885 6372 10919 6377
rect 10653 6351 10827 6354
rect 10646 6348 10827 6351
rect 10855 6371 10919 6372
rect 10449 6328 10468 6330
rect 10483 6328 10517 6330
rect 10449 6312 10529 6328
rect 10449 6306 10468 6312
rect 10165 6280 10268 6290
rect 10119 6278 10268 6280
rect 10289 6278 10324 6290
rect 9958 6276 10120 6278
rect 9970 6256 9989 6276
rect 10004 6274 10034 6276
rect 9853 6248 9894 6256
rect 9976 6252 9989 6256
rect 10041 6260 10120 6276
rect 10152 6276 10324 6278
rect 10152 6260 10231 6276
rect 10238 6274 10268 6276
rect 9816 6238 9845 6248
rect 9859 6238 9888 6248
rect 9903 6238 9933 6252
rect 9976 6238 10019 6252
rect 10041 6248 10231 6260
rect 10296 6256 10302 6276
rect 10026 6238 10056 6248
rect 10057 6238 10215 6248
rect 10219 6238 10249 6248
rect 10253 6238 10283 6252
rect 10311 6238 10324 6276
rect 10396 6290 10425 6306
rect 10439 6290 10468 6306
rect 10483 6296 10513 6312
rect 10541 6290 10547 6338
rect 10550 6332 10569 6338
rect 10584 6332 10614 6340
rect 10550 6324 10614 6332
rect 10550 6308 10630 6324
rect 10646 6317 10708 6348
rect 10724 6317 10786 6348
rect 10855 6346 10904 6371
rect 10919 6346 10949 6362
rect 10818 6332 10848 6340
rect 10855 6338 10965 6346
rect 10818 6324 10863 6332
rect 10550 6306 10569 6308
rect 10584 6306 10630 6308
rect 10550 6290 10630 6306
rect 10657 6304 10692 6317
rect 10733 6314 10770 6317
rect 10733 6312 10775 6314
rect 10662 6301 10692 6304
rect 10671 6297 10678 6301
rect 10678 6296 10679 6297
rect 10637 6290 10647 6296
rect 10396 6282 10431 6290
rect 10396 6256 10397 6282
rect 10404 6256 10431 6282
rect 10339 6238 10369 6252
rect 10396 6248 10431 6256
rect 10433 6282 10474 6290
rect 10433 6256 10448 6282
rect 10455 6256 10474 6282
rect 10538 6278 10569 6290
rect 10584 6278 10687 6290
rect 10699 6280 10725 6306
rect 10740 6301 10770 6312
rect 10802 6308 10864 6324
rect 10802 6306 10848 6308
rect 10802 6290 10864 6306
rect 10876 6290 10882 6338
rect 10885 6330 10965 6338
rect 10885 6328 10904 6330
rect 10919 6328 10953 6330
rect 10885 6312 10965 6328
rect 10885 6290 10904 6312
rect 10919 6296 10949 6312
rect 10977 6306 10983 6380
rect 10986 6306 11005 6450
rect 11020 6306 11026 6450
rect 11035 6380 11048 6450
rect 11100 6446 11122 6450
rect 11093 6424 11122 6438
rect 11175 6424 11191 6438
rect 11229 6434 11235 6436
rect 11242 6434 11350 6450
rect 11357 6434 11363 6436
rect 11371 6434 11386 6450
rect 11452 6444 11471 6447
rect 11093 6422 11191 6424
rect 11218 6422 11386 6434
rect 11401 6424 11417 6438
rect 11452 6425 11474 6444
rect 11484 6438 11500 6439
rect 11483 6436 11500 6438
rect 11484 6431 11500 6436
rect 11474 6424 11480 6425
rect 11483 6424 11512 6431
rect 11401 6423 11512 6424
rect 11401 6422 11518 6423
rect 11077 6414 11128 6422
rect 11175 6414 11209 6422
rect 11077 6402 11102 6414
rect 11109 6402 11128 6414
rect 11182 6412 11209 6414
rect 11218 6412 11439 6422
rect 11474 6419 11480 6422
rect 11182 6408 11439 6412
rect 11077 6394 11128 6402
rect 11175 6394 11439 6408
rect 11483 6414 11518 6422
rect 11029 6346 11048 6380
rect 11093 6386 11122 6394
rect 11093 6380 11110 6386
rect 11093 6378 11127 6380
rect 11175 6378 11191 6394
rect 11192 6384 11400 6394
rect 11401 6384 11417 6394
rect 11465 6390 11480 6405
rect 11483 6402 11484 6414
rect 11491 6402 11518 6414
rect 11483 6394 11518 6402
rect 11483 6393 11512 6394
rect 11203 6380 11417 6384
rect 11218 6378 11417 6380
rect 11452 6380 11465 6390
rect 11483 6380 11500 6393
rect 11452 6378 11500 6380
rect 11094 6374 11127 6378
rect 11090 6372 11127 6374
rect 11090 6371 11157 6372
rect 11090 6366 11121 6371
rect 11127 6366 11157 6371
rect 11090 6362 11157 6366
rect 11063 6359 11157 6362
rect 11063 6352 11112 6359
rect 11063 6346 11093 6352
rect 11112 6347 11117 6352
rect 11029 6330 11109 6346
rect 11121 6338 11157 6359
rect 11218 6354 11407 6378
rect 11452 6377 11499 6378
rect 11465 6372 11499 6377
rect 11233 6351 11407 6354
rect 11226 6348 11407 6351
rect 11435 6371 11499 6372
rect 11029 6328 11048 6330
rect 11063 6328 11097 6330
rect 11029 6312 11109 6328
rect 11029 6306 11048 6312
rect 10745 6280 10848 6290
rect 10699 6278 10848 6280
rect 10869 6278 10904 6290
rect 10538 6276 10700 6278
rect 10550 6256 10569 6276
rect 10584 6274 10614 6276
rect 10433 6248 10474 6256
rect 10556 6252 10569 6256
rect 10621 6260 10700 6276
rect 10732 6276 10904 6278
rect 10732 6260 10811 6276
rect 10818 6274 10848 6276
rect 10396 6238 10425 6248
rect 10439 6238 10468 6248
rect 10483 6238 10513 6252
rect 10556 6238 10599 6252
rect 10621 6248 10811 6260
rect 10876 6256 10882 6276
rect 10606 6238 10636 6248
rect 10637 6238 10795 6248
rect 10799 6238 10829 6248
rect 10833 6238 10863 6252
rect 10891 6238 10904 6276
rect 10976 6290 11005 6306
rect 11019 6290 11048 6306
rect 11063 6296 11093 6312
rect 11121 6290 11127 6338
rect 11130 6332 11149 6338
rect 11164 6332 11194 6340
rect 11130 6324 11194 6332
rect 11130 6308 11210 6324
rect 11226 6317 11288 6348
rect 11304 6317 11366 6348
rect 11435 6346 11484 6371
rect 11499 6346 11529 6362
rect 11398 6332 11428 6340
rect 11435 6338 11545 6346
rect 11398 6324 11443 6332
rect 11130 6306 11149 6308
rect 11164 6306 11210 6308
rect 11130 6290 11210 6306
rect 11237 6304 11272 6317
rect 11313 6314 11350 6317
rect 11313 6312 11355 6314
rect 11242 6301 11272 6304
rect 11251 6297 11258 6301
rect 11258 6296 11259 6297
rect 11217 6290 11227 6296
rect 10976 6282 11011 6290
rect 10976 6256 10977 6282
rect 10984 6256 11011 6282
rect 10919 6238 10949 6252
rect 10976 6248 11011 6256
rect 11013 6282 11054 6290
rect 11013 6256 11028 6282
rect 11035 6256 11054 6282
rect 11118 6278 11149 6290
rect 11164 6278 11267 6290
rect 11279 6280 11305 6306
rect 11320 6301 11350 6312
rect 11382 6308 11444 6324
rect 11382 6306 11428 6308
rect 11382 6290 11444 6306
rect 11456 6290 11462 6338
rect 11465 6330 11545 6338
rect 11465 6328 11484 6330
rect 11499 6328 11533 6330
rect 11465 6312 11545 6328
rect 11465 6290 11484 6312
rect 11499 6296 11529 6312
rect 11557 6306 11563 6380
rect 11566 6306 11585 6450
rect 11600 6306 11606 6450
rect 11615 6380 11628 6450
rect 11680 6446 11702 6450
rect 11673 6424 11702 6438
rect 11755 6424 11771 6438
rect 11809 6434 11815 6436
rect 11822 6434 11930 6450
rect 11937 6434 11943 6436
rect 11951 6434 11966 6450
rect 12032 6444 12051 6447
rect 11673 6422 11771 6424
rect 11798 6422 11966 6434
rect 11981 6424 11997 6438
rect 12032 6425 12054 6444
rect 12064 6438 12080 6439
rect 12063 6436 12080 6438
rect 12064 6431 12080 6436
rect 12054 6424 12060 6425
rect 12063 6424 12092 6431
rect 11981 6423 12092 6424
rect 11981 6422 12098 6423
rect 11657 6414 11708 6422
rect 11755 6414 11789 6422
rect 11657 6402 11682 6414
rect 11689 6402 11708 6414
rect 11762 6412 11789 6414
rect 11798 6412 12019 6422
rect 12054 6419 12060 6422
rect 11762 6408 12019 6412
rect 11657 6394 11708 6402
rect 11755 6394 12019 6408
rect 12063 6414 12098 6422
rect 11609 6346 11628 6380
rect 11673 6386 11702 6394
rect 11673 6380 11690 6386
rect 11673 6378 11707 6380
rect 11755 6378 11771 6394
rect 11772 6384 11980 6394
rect 11981 6384 11997 6394
rect 12045 6390 12060 6405
rect 12063 6402 12064 6414
rect 12071 6402 12098 6414
rect 12063 6394 12098 6402
rect 12063 6393 12092 6394
rect 11783 6380 11997 6384
rect 11798 6378 11997 6380
rect 12032 6380 12045 6390
rect 12063 6380 12080 6393
rect 12032 6378 12080 6380
rect 11674 6374 11707 6378
rect 11670 6372 11707 6374
rect 11670 6371 11737 6372
rect 11670 6366 11701 6371
rect 11707 6366 11737 6371
rect 11670 6362 11737 6366
rect 11643 6359 11737 6362
rect 11643 6352 11692 6359
rect 11643 6346 11673 6352
rect 11692 6347 11697 6352
rect 11609 6330 11689 6346
rect 11701 6338 11737 6359
rect 11798 6354 11987 6378
rect 12032 6377 12079 6378
rect 12045 6372 12079 6377
rect 11813 6351 11987 6354
rect 11806 6348 11987 6351
rect 12015 6371 12079 6372
rect 11609 6328 11628 6330
rect 11643 6328 11677 6330
rect 11609 6312 11689 6328
rect 11609 6306 11628 6312
rect 11325 6280 11428 6290
rect 11279 6278 11428 6280
rect 11449 6278 11484 6290
rect 11118 6276 11280 6278
rect 11130 6256 11149 6276
rect 11164 6274 11194 6276
rect 11013 6248 11054 6256
rect 11136 6252 11149 6256
rect 11201 6260 11280 6276
rect 11312 6276 11484 6278
rect 11312 6260 11391 6276
rect 11398 6274 11428 6276
rect 10976 6238 11005 6248
rect 11019 6238 11048 6248
rect 11063 6238 11093 6252
rect 11136 6238 11179 6252
rect 11201 6248 11391 6260
rect 11456 6256 11462 6276
rect 11186 6238 11216 6248
rect 11217 6238 11375 6248
rect 11379 6238 11409 6248
rect 11413 6238 11443 6252
rect 11471 6238 11484 6276
rect 11556 6290 11585 6306
rect 11599 6290 11628 6306
rect 11643 6296 11673 6312
rect 11701 6290 11707 6338
rect 11710 6332 11729 6338
rect 11744 6332 11774 6340
rect 11710 6324 11774 6332
rect 11710 6308 11790 6324
rect 11806 6317 11868 6348
rect 11884 6317 11946 6348
rect 12015 6346 12064 6371
rect 12079 6346 12109 6362
rect 11978 6332 12008 6340
rect 12015 6338 12125 6346
rect 11978 6324 12023 6332
rect 11710 6306 11729 6308
rect 11744 6306 11790 6308
rect 11710 6290 11790 6306
rect 11817 6304 11852 6317
rect 11893 6314 11930 6317
rect 11893 6312 11935 6314
rect 11822 6301 11852 6304
rect 11831 6297 11838 6301
rect 11838 6296 11839 6297
rect 11797 6290 11807 6296
rect 11556 6282 11591 6290
rect 11556 6256 11557 6282
rect 11564 6256 11591 6282
rect 11499 6238 11529 6252
rect 11556 6248 11591 6256
rect 11593 6282 11634 6290
rect 11593 6256 11608 6282
rect 11615 6256 11634 6282
rect 11698 6278 11729 6290
rect 11744 6278 11847 6290
rect 11859 6280 11885 6306
rect 11900 6301 11930 6312
rect 11962 6308 12024 6324
rect 11962 6306 12008 6308
rect 11962 6290 12024 6306
rect 12036 6290 12042 6338
rect 12045 6330 12125 6338
rect 12045 6328 12064 6330
rect 12079 6328 12113 6330
rect 12045 6312 12125 6328
rect 12045 6290 12064 6312
rect 12079 6296 12109 6312
rect 12137 6306 12143 6380
rect 12146 6306 12165 6450
rect 12180 6306 12186 6450
rect 12195 6380 12208 6450
rect 12260 6446 12282 6450
rect 12253 6424 12282 6438
rect 12335 6424 12351 6438
rect 12389 6434 12395 6436
rect 12402 6434 12510 6450
rect 12517 6434 12523 6436
rect 12531 6434 12546 6450
rect 12612 6444 12631 6447
rect 12253 6422 12351 6424
rect 12378 6422 12546 6434
rect 12561 6424 12577 6438
rect 12612 6425 12634 6444
rect 12644 6438 12660 6439
rect 12643 6436 12660 6438
rect 12644 6431 12660 6436
rect 12634 6424 12640 6425
rect 12643 6424 12672 6431
rect 12561 6423 12672 6424
rect 12561 6422 12678 6423
rect 12237 6414 12288 6422
rect 12335 6414 12369 6422
rect 12237 6402 12262 6414
rect 12269 6402 12288 6414
rect 12342 6412 12369 6414
rect 12378 6412 12599 6422
rect 12634 6419 12640 6422
rect 12342 6408 12599 6412
rect 12237 6394 12288 6402
rect 12335 6394 12599 6408
rect 12643 6414 12678 6422
rect 12189 6346 12208 6380
rect 12253 6386 12282 6394
rect 12253 6380 12270 6386
rect 12253 6378 12287 6380
rect 12335 6378 12351 6394
rect 12352 6384 12560 6394
rect 12561 6384 12577 6394
rect 12625 6390 12640 6405
rect 12643 6402 12644 6414
rect 12651 6402 12678 6414
rect 12643 6394 12678 6402
rect 12643 6393 12672 6394
rect 12363 6380 12577 6384
rect 12378 6378 12577 6380
rect 12612 6380 12625 6390
rect 12643 6380 12660 6393
rect 12612 6378 12660 6380
rect 12254 6374 12287 6378
rect 12250 6372 12287 6374
rect 12250 6371 12317 6372
rect 12250 6366 12281 6371
rect 12287 6366 12317 6371
rect 12250 6362 12317 6366
rect 12223 6359 12317 6362
rect 12223 6352 12272 6359
rect 12223 6346 12253 6352
rect 12272 6347 12277 6352
rect 12189 6330 12269 6346
rect 12281 6338 12317 6359
rect 12378 6354 12567 6378
rect 12612 6377 12659 6378
rect 12625 6372 12659 6377
rect 12393 6351 12567 6354
rect 12386 6348 12567 6351
rect 12595 6371 12659 6372
rect 12189 6328 12208 6330
rect 12223 6328 12257 6330
rect 12189 6312 12269 6328
rect 12189 6306 12208 6312
rect 11905 6280 12008 6290
rect 11859 6278 12008 6280
rect 12029 6278 12064 6290
rect 11698 6276 11860 6278
rect 11710 6256 11729 6276
rect 11744 6274 11774 6276
rect 11593 6248 11634 6256
rect 11716 6252 11729 6256
rect 11781 6260 11860 6276
rect 11892 6276 12064 6278
rect 11892 6260 11971 6276
rect 11978 6274 12008 6276
rect 11556 6238 11585 6248
rect 11599 6238 11628 6248
rect 11643 6238 11673 6252
rect 11716 6238 11759 6252
rect 11781 6248 11971 6260
rect 12036 6256 12042 6276
rect 11766 6238 11796 6248
rect 11797 6238 11955 6248
rect 11959 6238 11989 6248
rect 11993 6238 12023 6252
rect 12051 6238 12064 6276
rect 12136 6290 12165 6306
rect 12179 6290 12208 6306
rect 12223 6296 12253 6312
rect 12281 6290 12287 6338
rect 12290 6332 12309 6338
rect 12324 6332 12354 6340
rect 12290 6324 12354 6332
rect 12290 6308 12370 6324
rect 12386 6317 12448 6348
rect 12464 6317 12526 6348
rect 12595 6346 12644 6371
rect 12659 6346 12689 6362
rect 12558 6332 12588 6340
rect 12595 6338 12705 6346
rect 12558 6324 12603 6332
rect 12290 6306 12309 6308
rect 12324 6306 12370 6308
rect 12290 6290 12370 6306
rect 12397 6304 12432 6317
rect 12473 6314 12510 6317
rect 12473 6312 12515 6314
rect 12402 6301 12432 6304
rect 12411 6297 12418 6301
rect 12418 6296 12419 6297
rect 12377 6290 12387 6296
rect 12136 6282 12171 6290
rect 12136 6256 12137 6282
rect 12144 6256 12171 6282
rect 12079 6238 12109 6252
rect 12136 6248 12171 6256
rect 12173 6282 12214 6290
rect 12173 6256 12188 6282
rect 12195 6256 12214 6282
rect 12278 6278 12309 6290
rect 12324 6278 12427 6290
rect 12439 6280 12465 6306
rect 12480 6301 12510 6312
rect 12542 6308 12604 6324
rect 12542 6306 12588 6308
rect 12542 6290 12604 6306
rect 12616 6290 12622 6338
rect 12625 6330 12705 6338
rect 12625 6328 12644 6330
rect 12659 6328 12693 6330
rect 12625 6312 12705 6328
rect 12625 6290 12644 6312
rect 12659 6296 12689 6312
rect 12717 6306 12723 6380
rect 12726 6306 12745 6450
rect 12760 6306 12766 6450
rect 12775 6380 12788 6450
rect 12840 6446 12862 6450
rect 12833 6424 12862 6438
rect 12915 6424 12931 6438
rect 12969 6434 12975 6436
rect 12982 6434 13090 6450
rect 13097 6434 13103 6436
rect 13111 6434 13126 6450
rect 13192 6444 13211 6447
rect 12833 6422 12931 6424
rect 12958 6422 13126 6434
rect 13141 6424 13157 6438
rect 13192 6425 13214 6444
rect 13224 6438 13240 6439
rect 13223 6436 13240 6438
rect 13224 6431 13240 6436
rect 13214 6424 13220 6425
rect 13223 6424 13252 6431
rect 13141 6423 13252 6424
rect 13141 6422 13258 6423
rect 12817 6414 12868 6422
rect 12915 6414 12949 6422
rect 12817 6402 12842 6414
rect 12849 6402 12868 6414
rect 12922 6412 12949 6414
rect 12958 6412 13179 6422
rect 13214 6419 13220 6422
rect 12922 6408 13179 6412
rect 12817 6394 12868 6402
rect 12915 6394 13179 6408
rect 13223 6414 13258 6422
rect 12769 6346 12788 6380
rect 12833 6386 12862 6394
rect 12833 6380 12850 6386
rect 12833 6378 12867 6380
rect 12915 6378 12931 6394
rect 12932 6384 13140 6394
rect 13141 6384 13157 6394
rect 13205 6390 13220 6405
rect 13223 6402 13224 6414
rect 13231 6402 13258 6414
rect 13223 6394 13258 6402
rect 13223 6393 13252 6394
rect 12943 6380 13157 6384
rect 12958 6378 13157 6380
rect 13192 6380 13205 6390
rect 13223 6380 13240 6393
rect 13192 6378 13240 6380
rect 12834 6374 12867 6378
rect 12830 6372 12867 6374
rect 12830 6371 12897 6372
rect 12830 6366 12861 6371
rect 12867 6366 12897 6371
rect 12830 6362 12897 6366
rect 12803 6359 12897 6362
rect 12803 6352 12852 6359
rect 12803 6346 12833 6352
rect 12852 6347 12857 6352
rect 12769 6330 12849 6346
rect 12861 6338 12897 6359
rect 12958 6354 13147 6378
rect 13192 6377 13239 6378
rect 13205 6372 13239 6377
rect 12973 6351 13147 6354
rect 12966 6348 13147 6351
rect 13175 6371 13239 6372
rect 12769 6328 12788 6330
rect 12803 6328 12837 6330
rect 12769 6312 12849 6328
rect 12769 6306 12788 6312
rect 12485 6280 12588 6290
rect 12439 6278 12588 6280
rect 12609 6278 12644 6290
rect 12278 6276 12440 6278
rect 12290 6256 12309 6276
rect 12324 6274 12354 6276
rect 12173 6248 12214 6256
rect 12296 6252 12309 6256
rect 12361 6260 12440 6276
rect 12472 6276 12644 6278
rect 12472 6260 12551 6276
rect 12558 6274 12588 6276
rect 12136 6238 12165 6248
rect 12179 6238 12208 6248
rect 12223 6238 12253 6252
rect 12296 6238 12339 6252
rect 12361 6248 12551 6260
rect 12616 6256 12622 6276
rect 12346 6238 12376 6248
rect 12377 6238 12535 6248
rect 12539 6238 12569 6248
rect 12573 6238 12603 6252
rect 12631 6238 12644 6276
rect 12716 6290 12745 6306
rect 12759 6290 12788 6306
rect 12803 6296 12833 6312
rect 12861 6290 12867 6338
rect 12870 6332 12889 6338
rect 12904 6332 12934 6340
rect 12870 6324 12934 6332
rect 12870 6308 12950 6324
rect 12966 6317 13028 6348
rect 13044 6317 13106 6348
rect 13175 6346 13224 6371
rect 13239 6346 13269 6362
rect 13138 6332 13168 6340
rect 13175 6338 13285 6346
rect 13138 6324 13183 6332
rect 12870 6306 12889 6308
rect 12904 6306 12950 6308
rect 12870 6290 12950 6306
rect 12977 6304 13012 6317
rect 13053 6314 13090 6317
rect 13053 6312 13095 6314
rect 12982 6301 13012 6304
rect 12991 6297 12998 6301
rect 12998 6296 12999 6297
rect 12957 6290 12967 6296
rect 12716 6282 12751 6290
rect 12716 6256 12717 6282
rect 12724 6256 12751 6282
rect 12659 6238 12689 6252
rect 12716 6248 12751 6256
rect 12753 6282 12794 6290
rect 12753 6256 12768 6282
rect 12775 6256 12794 6282
rect 12858 6278 12889 6290
rect 12904 6278 13007 6290
rect 13019 6280 13045 6306
rect 13060 6301 13090 6312
rect 13122 6308 13184 6324
rect 13122 6306 13168 6308
rect 13122 6290 13184 6306
rect 13196 6290 13202 6338
rect 13205 6330 13285 6338
rect 13205 6328 13224 6330
rect 13239 6328 13273 6330
rect 13205 6312 13285 6328
rect 13205 6290 13224 6312
rect 13239 6296 13269 6312
rect 13297 6306 13303 6380
rect 13306 6306 13325 6450
rect 13340 6306 13346 6450
rect 13355 6380 13368 6450
rect 13420 6446 13442 6450
rect 13413 6424 13442 6438
rect 13495 6424 13511 6438
rect 13549 6434 13555 6436
rect 13562 6434 13670 6450
rect 13677 6434 13683 6436
rect 13691 6434 13706 6450
rect 13772 6444 13791 6447
rect 13413 6422 13511 6424
rect 13538 6422 13706 6434
rect 13721 6424 13737 6438
rect 13772 6425 13794 6444
rect 13804 6438 13820 6439
rect 13803 6436 13820 6438
rect 13804 6431 13820 6436
rect 13794 6424 13800 6425
rect 13803 6424 13832 6431
rect 13721 6423 13832 6424
rect 13721 6422 13838 6423
rect 13397 6414 13448 6422
rect 13495 6414 13529 6422
rect 13397 6402 13422 6414
rect 13429 6402 13448 6414
rect 13502 6412 13529 6414
rect 13538 6412 13759 6422
rect 13794 6419 13800 6422
rect 13502 6408 13759 6412
rect 13397 6394 13448 6402
rect 13495 6394 13759 6408
rect 13803 6414 13838 6422
rect 13349 6346 13368 6380
rect 13413 6386 13442 6394
rect 13413 6380 13430 6386
rect 13413 6378 13447 6380
rect 13495 6378 13511 6394
rect 13512 6384 13720 6394
rect 13721 6384 13737 6394
rect 13785 6390 13800 6405
rect 13803 6402 13804 6414
rect 13811 6402 13838 6414
rect 13803 6394 13838 6402
rect 13803 6393 13832 6394
rect 13523 6380 13737 6384
rect 13538 6378 13737 6380
rect 13772 6380 13785 6390
rect 13803 6380 13820 6393
rect 13772 6378 13820 6380
rect 13414 6374 13447 6378
rect 13410 6372 13447 6374
rect 13410 6371 13477 6372
rect 13410 6366 13441 6371
rect 13447 6366 13477 6371
rect 13410 6362 13477 6366
rect 13383 6359 13477 6362
rect 13383 6352 13432 6359
rect 13383 6346 13413 6352
rect 13432 6347 13437 6352
rect 13349 6330 13429 6346
rect 13441 6338 13477 6359
rect 13538 6354 13727 6378
rect 13772 6377 13819 6378
rect 13785 6372 13819 6377
rect 13553 6351 13727 6354
rect 13546 6348 13727 6351
rect 13755 6371 13819 6372
rect 13349 6328 13368 6330
rect 13383 6328 13417 6330
rect 13349 6312 13429 6328
rect 13349 6306 13368 6312
rect 13065 6280 13168 6290
rect 13019 6278 13168 6280
rect 13189 6278 13224 6290
rect 12858 6276 13020 6278
rect 12870 6256 12889 6276
rect 12904 6274 12934 6276
rect 12753 6248 12794 6256
rect 12876 6252 12889 6256
rect 12941 6260 13020 6276
rect 13052 6276 13224 6278
rect 13052 6260 13131 6276
rect 13138 6274 13168 6276
rect 12716 6238 12745 6248
rect 12759 6238 12788 6248
rect 12803 6238 12833 6252
rect 12876 6238 12919 6252
rect 12941 6248 13131 6260
rect 13196 6256 13202 6276
rect 12926 6238 12956 6248
rect 12957 6238 13115 6248
rect 13119 6238 13149 6248
rect 13153 6238 13183 6252
rect 13211 6238 13224 6276
rect 13296 6290 13325 6306
rect 13339 6290 13368 6306
rect 13383 6296 13413 6312
rect 13441 6290 13447 6338
rect 13450 6332 13469 6338
rect 13484 6332 13514 6340
rect 13450 6324 13514 6332
rect 13450 6308 13530 6324
rect 13546 6317 13608 6348
rect 13624 6317 13686 6348
rect 13755 6346 13804 6371
rect 13819 6346 13849 6362
rect 13718 6332 13748 6340
rect 13755 6338 13865 6346
rect 13718 6324 13763 6332
rect 13450 6306 13469 6308
rect 13484 6306 13530 6308
rect 13450 6290 13530 6306
rect 13557 6304 13592 6317
rect 13633 6314 13670 6317
rect 13633 6312 13675 6314
rect 13562 6301 13592 6304
rect 13571 6297 13578 6301
rect 13578 6296 13579 6297
rect 13537 6290 13547 6296
rect 13296 6282 13331 6290
rect 13296 6256 13297 6282
rect 13304 6256 13331 6282
rect 13239 6238 13269 6252
rect 13296 6248 13331 6256
rect 13333 6282 13374 6290
rect 13333 6256 13348 6282
rect 13355 6256 13374 6282
rect 13438 6278 13469 6290
rect 13484 6278 13587 6290
rect 13599 6280 13625 6306
rect 13640 6301 13670 6312
rect 13702 6308 13764 6324
rect 13702 6306 13748 6308
rect 13702 6290 13764 6306
rect 13776 6290 13782 6338
rect 13785 6330 13865 6338
rect 13785 6328 13804 6330
rect 13819 6328 13853 6330
rect 13785 6312 13865 6328
rect 13785 6290 13804 6312
rect 13819 6296 13849 6312
rect 13877 6306 13883 6380
rect 13886 6306 13905 6450
rect 13920 6306 13926 6450
rect 13935 6380 13948 6450
rect 14000 6446 14022 6450
rect 13993 6424 14022 6438
rect 14075 6424 14091 6438
rect 14129 6434 14135 6436
rect 14142 6434 14250 6450
rect 14257 6434 14263 6436
rect 14271 6434 14286 6450
rect 14352 6444 14371 6447
rect 13993 6422 14091 6424
rect 14118 6422 14286 6434
rect 14301 6424 14317 6438
rect 14352 6425 14374 6444
rect 14384 6438 14400 6439
rect 14383 6436 14400 6438
rect 14384 6431 14400 6436
rect 14374 6424 14380 6425
rect 14383 6424 14412 6431
rect 14301 6423 14412 6424
rect 14301 6422 14418 6423
rect 13977 6414 14028 6422
rect 14075 6414 14109 6422
rect 13977 6402 14002 6414
rect 14009 6402 14028 6414
rect 14082 6412 14109 6414
rect 14118 6412 14339 6422
rect 14374 6419 14380 6422
rect 14082 6408 14339 6412
rect 13977 6394 14028 6402
rect 14075 6394 14339 6408
rect 14383 6414 14418 6422
rect 13929 6346 13948 6380
rect 13993 6386 14022 6394
rect 13993 6380 14010 6386
rect 13993 6378 14027 6380
rect 14075 6378 14091 6394
rect 14092 6384 14300 6394
rect 14301 6384 14317 6394
rect 14365 6390 14380 6405
rect 14383 6402 14384 6414
rect 14391 6402 14418 6414
rect 14383 6394 14418 6402
rect 14383 6393 14412 6394
rect 14103 6380 14317 6384
rect 14118 6378 14317 6380
rect 14352 6380 14365 6390
rect 14383 6380 14400 6393
rect 14352 6378 14400 6380
rect 13994 6374 14027 6378
rect 13990 6372 14027 6374
rect 13990 6371 14057 6372
rect 13990 6366 14021 6371
rect 14027 6366 14057 6371
rect 13990 6362 14057 6366
rect 13963 6359 14057 6362
rect 13963 6352 14012 6359
rect 13963 6346 13993 6352
rect 14012 6347 14017 6352
rect 13929 6330 14009 6346
rect 14021 6338 14057 6359
rect 14118 6354 14307 6378
rect 14352 6377 14399 6378
rect 14365 6372 14399 6377
rect 14133 6351 14307 6354
rect 14126 6348 14307 6351
rect 14335 6371 14399 6372
rect 13929 6328 13948 6330
rect 13963 6328 13997 6330
rect 13929 6312 14009 6328
rect 13929 6306 13948 6312
rect 13645 6280 13748 6290
rect 13599 6278 13748 6280
rect 13769 6278 13804 6290
rect 13438 6276 13600 6278
rect 13450 6256 13469 6276
rect 13484 6274 13514 6276
rect 13333 6248 13374 6256
rect 13456 6252 13469 6256
rect 13521 6260 13600 6276
rect 13632 6276 13804 6278
rect 13632 6260 13711 6276
rect 13718 6274 13748 6276
rect 13296 6238 13325 6248
rect 13339 6238 13368 6248
rect 13383 6238 13413 6252
rect 13456 6238 13499 6252
rect 13521 6248 13711 6260
rect 13776 6256 13782 6276
rect 13506 6238 13536 6248
rect 13537 6238 13695 6248
rect 13699 6238 13729 6248
rect 13733 6238 13763 6252
rect 13791 6238 13804 6276
rect 13876 6290 13905 6306
rect 13919 6290 13948 6306
rect 13963 6296 13993 6312
rect 14021 6290 14027 6338
rect 14030 6332 14049 6338
rect 14064 6332 14094 6340
rect 14030 6324 14094 6332
rect 14030 6308 14110 6324
rect 14126 6317 14188 6348
rect 14204 6317 14266 6348
rect 14335 6346 14384 6371
rect 14399 6346 14429 6362
rect 14298 6332 14328 6340
rect 14335 6338 14445 6346
rect 14298 6324 14343 6332
rect 14030 6306 14049 6308
rect 14064 6306 14110 6308
rect 14030 6290 14110 6306
rect 14137 6304 14172 6317
rect 14213 6314 14250 6317
rect 14213 6312 14255 6314
rect 14142 6301 14172 6304
rect 14151 6297 14158 6301
rect 14158 6296 14159 6297
rect 14117 6290 14127 6296
rect 13876 6282 13911 6290
rect 13876 6256 13877 6282
rect 13884 6256 13911 6282
rect 13819 6238 13849 6252
rect 13876 6248 13911 6256
rect 13913 6282 13954 6290
rect 13913 6256 13928 6282
rect 13935 6256 13954 6282
rect 14018 6278 14049 6290
rect 14064 6278 14167 6290
rect 14179 6280 14205 6306
rect 14220 6301 14250 6312
rect 14282 6308 14344 6324
rect 14282 6306 14328 6308
rect 14282 6290 14344 6306
rect 14356 6290 14362 6338
rect 14365 6330 14445 6338
rect 14365 6328 14384 6330
rect 14399 6328 14433 6330
rect 14365 6312 14445 6328
rect 14365 6290 14384 6312
rect 14399 6296 14429 6312
rect 14457 6306 14463 6380
rect 14466 6306 14485 6450
rect 14500 6306 14506 6450
rect 14515 6380 14528 6450
rect 14580 6446 14602 6450
rect 14573 6424 14602 6438
rect 14655 6424 14671 6438
rect 14709 6434 14715 6436
rect 14722 6434 14830 6450
rect 14837 6434 14843 6436
rect 14851 6434 14866 6450
rect 14932 6444 14951 6447
rect 14573 6422 14671 6424
rect 14698 6422 14866 6434
rect 14881 6424 14897 6438
rect 14932 6425 14954 6444
rect 14964 6438 14980 6439
rect 14963 6436 14980 6438
rect 14964 6431 14980 6436
rect 14954 6424 14960 6425
rect 14963 6424 14992 6431
rect 14881 6423 14992 6424
rect 14881 6422 14998 6423
rect 14557 6414 14608 6422
rect 14655 6414 14689 6422
rect 14557 6402 14582 6414
rect 14589 6402 14608 6414
rect 14662 6412 14689 6414
rect 14698 6412 14919 6422
rect 14954 6419 14960 6422
rect 14662 6408 14919 6412
rect 14557 6394 14608 6402
rect 14655 6394 14919 6408
rect 14963 6414 14998 6422
rect 14509 6346 14528 6380
rect 14573 6386 14602 6394
rect 14573 6380 14590 6386
rect 14573 6378 14607 6380
rect 14655 6378 14671 6394
rect 14672 6384 14880 6394
rect 14881 6384 14897 6394
rect 14945 6390 14960 6405
rect 14963 6402 14964 6414
rect 14971 6402 14998 6414
rect 14963 6394 14998 6402
rect 14963 6393 14992 6394
rect 14683 6380 14897 6384
rect 14698 6378 14897 6380
rect 14932 6380 14945 6390
rect 14963 6380 14980 6393
rect 14932 6378 14980 6380
rect 14574 6374 14607 6378
rect 14570 6372 14607 6374
rect 14570 6371 14637 6372
rect 14570 6366 14601 6371
rect 14607 6366 14637 6371
rect 14570 6362 14637 6366
rect 14543 6359 14637 6362
rect 14543 6352 14592 6359
rect 14543 6346 14573 6352
rect 14592 6347 14597 6352
rect 14509 6330 14589 6346
rect 14601 6338 14637 6359
rect 14698 6354 14887 6378
rect 14932 6377 14979 6378
rect 14945 6372 14979 6377
rect 14713 6351 14887 6354
rect 14706 6348 14887 6351
rect 14915 6371 14979 6372
rect 14509 6328 14528 6330
rect 14543 6328 14577 6330
rect 14509 6312 14589 6328
rect 14509 6306 14528 6312
rect 14225 6280 14328 6290
rect 14179 6278 14328 6280
rect 14349 6278 14384 6290
rect 14018 6276 14180 6278
rect 14030 6256 14049 6276
rect 14064 6274 14094 6276
rect 13913 6248 13954 6256
rect 14036 6252 14049 6256
rect 14101 6260 14180 6276
rect 14212 6276 14384 6278
rect 14212 6260 14291 6276
rect 14298 6274 14328 6276
rect 13876 6238 13905 6248
rect 13919 6238 13948 6248
rect 13963 6238 13993 6252
rect 14036 6238 14079 6252
rect 14101 6248 14291 6260
rect 14356 6256 14362 6276
rect 14086 6238 14116 6248
rect 14117 6238 14275 6248
rect 14279 6238 14309 6248
rect 14313 6238 14343 6252
rect 14371 6238 14384 6276
rect 14456 6290 14485 6306
rect 14499 6290 14528 6306
rect 14543 6296 14573 6312
rect 14601 6290 14607 6338
rect 14610 6332 14629 6338
rect 14644 6332 14674 6340
rect 14610 6324 14674 6332
rect 14610 6308 14690 6324
rect 14706 6317 14768 6348
rect 14784 6317 14846 6348
rect 14915 6346 14964 6371
rect 14979 6346 15009 6362
rect 14878 6332 14908 6340
rect 14915 6338 15025 6346
rect 14878 6324 14923 6332
rect 14610 6306 14629 6308
rect 14644 6306 14690 6308
rect 14610 6290 14690 6306
rect 14717 6304 14752 6317
rect 14793 6314 14830 6317
rect 14793 6312 14835 6314
rect 14722 6301 14752 6304
rect 14731 6297 14738 6301
rect 14738 6296 14739 6297
rect 14697 6290 14707 6296
rect 14456 6282 14491 6290
rect 14456 6256 14457 6282
rect 14464 6256 14491 6282
rect 14399 6238 14429 6252
rect 14456 6248 14491 6256
rect 14493 6282 14534 6290
rect 14493 6256 14508 6282
rect 14515 6256 14534 6282
rect 14598 6278 14629 6290
rect 14644 6278 14747 6290
rect 14759 6280 14785 6306
rect 14800 6301 14830 6312
rect 14862 6308 14924 6324
rect 14862 6306 14908 6308
rect 14862 6290 14924 6306
rect 14936 6290 14942 6338
rect 14945 6330 15025 6338
rect 14945 6328 14964 6330
rect 14979 6328 15013 6330
rect 14945 6312 15025 6328
rect 14945 6290 14964 6312
rect 14979 6296 15009 6312
rect 15037 6306 15043 6380
rect 15046 6306 15065 6450
rect 15080 6306 15086 6450
rect 15095 6380 15108 6450
rect 15160 6446 15182 6450
rect 15153 6424 15182 6438
rect 15235 6424 15251 6438
rect 15289 6434 15295 6436
rect 15302 6434 15410 6450
rect 15417 6434 15423 6436
rect 15431 6434 15446 6450
rect 15512 6444 15531 6447
rect 15153 6422 15251 6424
rect 15278 6422 15446 6434
rect 15461 6424 15477 6438
rect 15512 6425 15534 6444
rect 15544 6438 15560 6439
rect 15543 6436 15560 6438
rect 15544 6431 15560 6436
rect 15534 6424 15540 6425
rect 15543 6424 15572 6431
rect 15461 6423 15572 6424
rect 15461 6422 15578 6423
rect 15137 6414 15188 6422
rect 15235 6414 15269 6422
rect 15137 6402 15162 6414
rect 15169 6402 15188 6414
rect 15242 6412 15269 6414
rect 15278 6412 15499 6422
rect 15534 6419 15540 6422
rect 15242 6408 15499 6412
rect 15137 6394 15188 6402
rect 15235 6394 15499 6408
rect 15543 6414 15578 6422
rect 15089 6346 15108 6380
rect 15153 6386 15182 6394
rect 15153 6380 15170 6386
rect 15153 6378 15187 6380
rect 15235 6378 15251 6394
rect 15252 6384 15460 6394
rect 15461 6384 15477 6394
rect 15525 6390 15540 6405
rect 15543 6402 15544 6414
rect 15551 6402 15578 6414
rect 15543 6394 15578 6402
rect 15543 6393 15572 6394
rect 15263 6380 15477 6384
rect 15278 6378 15477 6380
rect 15512 6380 15525 6390
rect 15543 6380 15560 6393
rect 15512 6378 15560 6380
rect 15154 6374 15187 6378
rect 15150 6372 15187 6374
rect 15150 6371 15217 6372
rect 15150 6366 15181 6371
rect 15187 6366 15217 6371
rect 15150 6362 15217 6366
rect 15123 6359 15217 6362
rect 15123 6352 15172 6359
rect 15123 6346 15153 6352
rect 15172 6347 15177 6352
rect 15089 6330 15169 6346
rect 15181 6338 15217 6359
rect 15278 6354 15467 6378
rect 15512 6377 15559 6378
rect 15525 6372 15559 6377
rect 15293 6351 15467 6354
rect 15286 6348 15467 6351
rect 15495 6371 15559 6372
rect 15089 6328 15108 6330
rect 15123 6328 15157 6330
rect 15089 6312 15169 6328
rect 15089 6306 15108 6312
rect 14805 6280 14908 6290
rect 14759 6278 14908 6280
rect 14929 6278 14964 6290
rect 14598 6276 14760 6278
rect 14610 6256 14629 6276
rect 14644 6274 14674 6276
rect 14493 6248 14534 6256
rect 14616 6252 14629 6256
rect 14681 6260 14760 6276
rect 14792 6276 14964 6278
rect 14792 6260 14871 6276
rect 14878 6274 14908 6276
rect 14456 6238 14485 6248
rect 14499 6238 14528 6248
rect 14543 6238 14573 6252
rect 14616 6238 14659 6252
rect 14681 6248 14871 6260
rect 14936 6256 14942 6276
rect 14666 6238 14696 6248
rect 14697 6238 14855 6248
rect 14859 6238 14889 6248
rect 14893 6238 14923 6252
rect 14951 6238 14964 6276
rect 15036 6290 15065 6306
rect 15079 6290 15108 6306
rect 15123 6296 15153 6312
rect 15181 6290 15187 6338
rect 15190 6332 15209 6338
rect 15224 6332 15254 6340
rect 15190 6324 15254 6332
rect 15190 6308 15270 6324
rect 15286 6317 15348 6348
rect 15364 6317 15426 6348
rect 15495 6346 15544 6371
rect 15559 6346 15589 6362
rect 15458 6332 15488 6340
rect 15495 6338 15605 6346
rect 15458 6324 15503 6332
rect 15190 6306 15209 6308
rect 15224 6306 15270 6308
rect 15190 6290 15270 6306
rect 15297 6304 15332 6317
rect 15373 6314 15410 6317
rect 15373 6312 15415 6314
rect 15302 6301 15332 6304
rect 15311 6297 15318 6301
rect 15318 6296 15319 6297
rect 15277 6290 15287 6296
rect 15036 6282 15071 6290
rect 15036 6256 15037 6282
rect 15044 6256 15071 6282
rect 14979 6238 15009 6252
rect 15036 6248 15071 6256
rect 15073 6282 15114 6290
rect 15073 6256 15088 6282
rect 15095 6256 15114 6282
rect 15178 6278 15209 6290
rect 15224 6278 15327 6290
rect 15339 6280 15365 6306
rect 15380 6301 15410 6312
rect 15442 6308 15504 6324
rect 15442 6306 15488 6308
rect 15442 6290 15504 6306
rect 15516 6290 15522 6338
rect 15525 6330 15605 6338
rect 15525 6328 15544 6330
rect 15559 6328 15593 6330
rect 15525 6312 15605 6328
rect 15525 6290 15544 6312
rect 15559 6296 15589 6312
rect 15617 6306 15623 6380
rect 15626 6306 15645 6450
rect 15660 6306 15666 6450
rect 15675 6380 15688 6450
rect 15740 6446 15762 6450
rect 15733 6424 15762 6438
rect 15815 6424 15831 6438
rect 15869 6434 15875 6436
rect 15882 6434 15990 6450
rect 15997 6434 16003 6436
rect 16011 6434 16026 6450
rect 16092 6444 16111 6447
rect 15733 6422 15831 6424
rect 15858 6422 16026 6434
rect 16041 6424 16057 6438
rect 16092 6425 16114 6444
rect 16124 6438 16140 6439
rect 16123 6436 16140 6438
rect 16124 6431 16140 6436
rect 16114 6424 16120 6425
rect 16123 6424 16152 6431
rect 16041 6423 16152 6424
rect 16041 6422 16158 6423
rect 15717 6414 15768 6422
rect 15815 6414 15849 6422
rect 15717 6402 15742 6414
rect 15749 6402 15768 6414
rect 15822 6412 15849 6414
rect 15858 6412 16079 6422
rect 16114 6419 16120 6422
rect 15822 6408 16079 6412
rect 15717 6394 15768 6402
rect 15815 6394 16079 6408
rect 16123 6414 16158 6422
rect 15669 6346 15688 6380
rect 15733 6386 15762 6394
rect 15733 6380 15750 6386
rect 15733 6378 15767 6380
rect 15815 6378 15831 6394
rect 15832 6384 16040 6394
rect 16041 6384 16057 6394
rect 16105 6390 16120 6405
rect 16123 6402 16124 6414
rect 16131 6402 16158 6414
rect 16123 6394 16158 6402
rect 16123 6393 16152 6394
rect 15843 6380 16057 6384
rect 15858 6378 16057 6380
rect 16092 6380 16105 6390
rect 16123 6380 16140 6393
rect 16092 6378 16140 6380
rect 15734 6374 15767 6378
rect 15730 6372 15767 6374
rect 15730 6371 15797 6372
rect 15730 6366 15761 6371
rect 15767 6366 15797 6371
rect 15730 6362 15797 6366
rect 15703 6359 15797 6362
rect 15703 6352 15752 6359
rect 15703 6346 15733 6352
rect 15752 6347 15757 6352
rect 15669 6330 15749 6346
rect 15761 6338 15797 6359
rect 15858 6354 16047 6378
rect 16092 6377 16139 6378
rect 16105 6372 16139 6377
rect 15873 6351 16047 6354
rect 15866 6348 16047 6351
rect 16075 6371 16139 6372
rect 15669 6328 15688 6330
rect 15703 6328 15737 6330
rect 15669 6312 15749 6328
rect 15669 6306 15688 6312
rect 15385 6280 15488 6290
rect 15339 6278 15488 6280
rect 15509 6278 15544 6290
rect 15178 6276 15340 6278
rect 15190 6256 15209 6276
rect 15224 6274 15254 6276
rect 15073 6248 15114 6256
rect 15196 6252 15209 6256
rect 15261 6260 15340 6276
rect 15372 6276 15544 6278
rect 15372 6260 15451 6276
rect 15458 6274 15488 6276
rect 15036 6238 15065 6248
rect 15079 6238 15108 6248
rect 15123 6238 15153 6252
rect 15196 6238 15239 6252
rect 15261 6248 15451 6260
rect 15516 6256 15522 6276
rect 15246 6238 15276 6248
rect 15277 6238 15435 6248
rect 15439 6238 15469 6248
rect 15473 6238 15503 6252
rect 15531 6238 15544 6276
rect 15616 6290 15645 6306
rect 15659 6290 15688 6306
rect 15703 6296 15733 6312
rect 15761 6290 15767 6338
rect 15770 6332 15789 6338
rect 15804 6332 15834 6340
rect 15770 6324 15834 6332
rect 15770 6308 15850 6324
rect 15866 6317 15928 6348
rect 15944 6317 16006 6348
rect 16075 6346 16124 6371
rect 16139 6346 16169 6362
rect 16038 6332 16068 6340
rect 16075 6338 16185 6346
rect 16038 6324 16083 6332
rect 15770 6306 15789 6308
rect 15804 6306 15850 6308
rect 15770 6290 15850 6306
rect 15877 6304 15912 6317
rect 15953 6314 15990 6317
rect 15953 6312 15995 6314
rect 15882 6301 15912 6304
rect 15891 6297 15898 6301
rect 15898 6296 15899 6297
rect 15857 6290 15867 6296
rect 15616 6282 15651 6290
rect 15616 6256 15617 6282
rect 15624 6256 15651 6282
rect 15559 6238 15589 6252
rect 15616 6248 15651 6256
rect 15653 6282 15694 6290
rect 15653 6256 15668 6282
rect 15675 6256 15694 6282
rect 15758 6278 15789 6290
rect 15804 6278 15907 6290
rect 15919 6280 15945 6306
rect 15960 6301 15990 6312
rect 16022 6308 16084 6324
rect 16022 6306 16068 6308
rect 16022 6290 16084 6306
rect 16096 6290 16102 6338
rect 16105 6330 16185 6338
rect 16105 6328 16124 6330
rect 16139 6328 16173 6330
rect 16105 6312 16185 6328
rect 16105 6290 16124 6312
rect 16139 6296 16169 6312
rect 16197 6306 16203 6380
rect 16206 6306 16225 6450
rect 16240 6306 16246 6450
rect 16255 6380 16268 6450
rect 16320 6446 16342 6450
rect 16313 6424 16342 6438
rect 16395 6424 16411 6438
rect 16449 6434 16455 6436
rect 16462 6434 16570 6450
rect 16577 6434 16583 6436
rect 16591 6434 16606 6450
rect 16672 6444 16691 6447
rect 16313 6422 16411 6424
rect 16438 6422 16606 6434
rect 16621 6424 16637 6438
rect 16672 6425 16694 6444
rect 16704 6438 16720 6439
rect 16703 6436 16720 6438
rect 16704 6431 16720 6436
rect 16694 6424 16700 6425
rect 16703 6424 16732 6431
rect 16621 6423 16732 6424
rect 16621 6422 16738 6423
rect 16297 6414 16348 6422
rect 16395 6414 16429 6422
rect 16297 6402 16322 6414
rect 16329 6402 16348 6414
rect 16402 6412 16429 6414
rect 16438 6412 16659 6422
rect 16694 6419 16700 6422
rect 16402 6408 16659 6412
rect 16297 6394 16348 6402
rect 16395 6394 16659 6408
rect 16703 6414 16738 6422
rect 16249 6346 16268 6380
rect 16313 6386 16342 6394
rect 16313 6380 16330 6386
rect 16313 6378 16347 6380
rect 16395 6378 16411 6394
rect 16412 6384 16620 6394
rect 16621 6384 16637 6394
rect 16685 6390 16700 6405
rect 16703 6402 16704 6414
rect 16711 6402 16738 6414
rect 16703 6394 16738 6402
rect 16703 6393 16732 6394
rect 16423 6380 16637 6384
rect 16438 6378 16637 6380
rect 16672 6380 16685 6390
rect 16703 6380 16720 6393
rect 16672 6378 16720 6380
rect 16314 6374 16347 6378
rect 16310 6372 16347 6374
rect 16310 6371 16377 6372
rect 16310 6366 16341 6371
rect 16347 6366 16377 6371
rect 16310 6362 16377 6366
rect 16283 6359 16377 6362
rect 16283 6352 16332 6359
rect 16283 6346 16313 6352
rect 16332 6347 16337 6352
rect 16249 6330 16329 6346
rect 16341 6338 16377 6359
rect 16438 6354 16627 6378
rect 16672 6377 16719 6378
rect 16685 6372 16719 6377
rect 16453 6351 16627 6354
rect 16446 6348 16627 6351
rect 16655 6371 16719 6372
rect 16249 6328 16268 6330
rect 16283 6328 16317 6330
rect 16249 6312 16329 6328
rect 16249 6306 16268 6312
rect 15965 6280 16068 6290
rect 15919 6278 16068 6280
rect 16089 6278 16124 6290
rect 15758 6276 15920 6278
rect 15770 6256 15789 6276
rect 15804 6274 15834 6276
rect 15653 6248 15694 6256
rect 15776 6252 15789 6256
rect 15841 6260 15920 6276
rect 15952 6276 16124 6278
rect 15952 6260 16031 6276
rect 16038 6274 16068 6276
rect 15616 6238 15645 6248
rect 15659 6238 15688 6248
rect 15703 6238 15733 6252
rect 15776 6238 15819 6252
rect 15841 6248 16031 6260
rect 16096 6256 16102 6276
rect 15826 6238 15856 6248
rect 15857 6238 16015 6248
rect 16019 6238 16049 6248
rect 16053 6238 16083 6252
rect 16111 6238 16124 6276
rect 16196 6290 16225 6306
rect 16239 6290 16268 6306
rect 16283 6296 16313 6312
rect 16341 6290 16347 6338
rect 16350 6332 16369 6338
rect 16384 6332 16414 6340
rect 16350 6324 16414 6332
rect 16350 6308 16430 6324
rect 16446 6317 16508 6348
rect 16524 6317 16586 6348
rect 16655 6346 16704 6371
rect 16719 6346 16749 6362
rect 16618 6332 16648 6340
rect 16655 6338 16765 6346
rect 16618 6324 16663 6332
rect 16350 6306 16369 6308
rect 16384 6306 16430 6308
rect 16350 6290 16430 6306
rect 16457 6304 16492 6317
rect 16533 6314 16570 6317
rect 16533 6312 16575 6314
rect 16462 6301 16492 6304
rect 16471 6297 16478 6301
rect 16478 6296 16479 6297
rect 16437 6290 16447 6296
rect 16196 6282 16231 6290
rect 16196 6256 16197 6282
rect 16204 6256 16231 6282
rect 16139 6238 16169 6252
rect 16196 6248 16231 6256
rect 16233 6282 16274 6290
rect 16233 6256 16248 6282
rect 16255 6256 16274 6282
rect 16338 6278 16369 6290
rect 16384 6278 16487 6290
rect 16499 6280 16525 6306
rect 16540 6301 16570 6312
rect 16602 6308 16664 6324
rect 16602 6306 16648 6308
rect 16602 6290 16664 6306
rect 16676 6290 16682 6338
rect 16685 6330 16765 6338
rect 16685 6328 16704 6330
rect 16719 6328 16753 6330
rect 16685 6312 16765 6328
rect 16685 6290 16704 6312
rect 16719 6296 16749 6312
rect 16777 6306 16783 6380
rect 16786 6306 16805 6450
rect 16820 6306 16826 6450
rect 16835 6380 16848 6450
rect 16900 6446 16922 6450
rect 16893 6424 16922 6438
rect 16975 6424 16991 6438
rect 17029 6434 17035 6436
rect 17042 6434 17150 6450
rect 17157 6434 17163 6436
rect 17171 6434 17186 6450
rect 17252 6444 17271 6447
rect 16893 6422 16991 6424
rect 17018 6422 17186 6434
rect 17201 6424 17217 6438
rect 17252 6425 17274 6444
rect 17284 6438 17300 6439
rect 17283 6436 17300 6438
rect 17284 6431 17300 6436
rect 17274 6424 17280 6425
rect 17283 6424 17312 6431
rect 17201 6423 17312 6424
rect 17201 6422 17318 6423
rect 16877 6414 16928 6422
rect 16975 6414 17009 6422
rect 16877 6402 16902 6414
rect 16909 6402 16928 6414
rect 16982 6412 17009 6414
rect 17018 6412 17239 6422
rect 17274 6419 17280 6422
rect 16982 6408 17239 6412
rect 16877 6394 16928 6402
rect 16975 6394 17239 6408
rect 17283 6414 17318 6422
rect 16829 6346 16848 6380
rect 16893 6386 16922 6394
rect 16893 6380 16910 6386
rect 16893 6378 16927 6380
rect 16975 6378 16991 6394
rect 16992 6384 17200 6394
rect 17201 6384 17217 6394
rect 17265 6390 17280 6405
rect 17283 6402 17284 6414
rect 17291 6402 17318 6414
rect 17283 6394 17318 6402
rect 17283 6393 17312 6394
rect 17003 6380 17217 6384
rect 17018 6378 17217 6380
rect 17252 6380 17265 6390
rect 17283 6380 17300 6393
rect 17252 6378 17300 6380
rect 16894 6374 16927 6378
rect 16890 6372 16927 6374
rect 16890 6371 16957 6372
rect 16890 6366 16921 6371
rect 16927 6366 16957 6371
rect 16890 6362 16957 6366
rect 16863 6359 16957 6362
rect 16863 6352 16912 6359
rect 16863 6346 16893 6352
rect 16912 6347 16917 6352
rect 16829 6330 16909 6346
rect 16921 6338 16957 6359
rect 17018 6354 17207 6378
rect 17252 6377 17299 6378
rect 17265 6372 17299 6377
rect 17033 6351 17207 6354
rect 17026 6348 17207 6351
rect 17235 6371 17299 6372
rect 16829 6328 16848 6330
rect 16863 6328 16897 6330
rect 16829 6312 16909 6328
rect 16829 6306 16848 6312
rect 16545 6280 16648 6290
rect 16499 6278 16648 6280
rect 16669 6278 16704 6290
rect 16338 6276 16500 6278
rect 16350 6256 16369 6276
rect 16384 6274 16414 6276
rect 16233 6248 16274 6256
rect 16356 6252 16369 6256
rect 16421 6260 16500 6276
rect 16532 6276 16704 6278
rect 16532 6260 16611 6276
rect 16618 6274 16648 6276
rect 16196 6238 16225 6248
rect 16239 6238 16268 6248
rect 16283 6238 16313 6252
rect 16356 6238 16399 6252
rect 16421 6248 16611 6260
rect 16676 6256 16682 6276
rect 16406 6238 16436 6248
rect 16437 6238 16595 6248
rect 16599 6238 16629 6248
rect 16633 6238 16663 6252
rect 16691 6238 16704 6276
rect 16776 6290 16805 6306
rect 16819 6290 16848 6306
rect 16863 6296 16893 6312
rect 16921 6290 16927 6338
rect 16930 6332 16949 6338
rect 16964 6332 16994 6340
rect 16930 6324 16994 6332
rect 16930 6308 17010 6324
rect 17026 6317 17088 6348
rect 17104 6317 17166 6348
rect 17235 6346 17284 6371
rect 17299 6346 17329 6362
rect 17198 6332 17228 6340
rect 17235 6338 17345 6346
rect 17198 6324 17243 6332
rect 16930 6306 16949 6308
rect 16964 6306 17010 6308
rect 16930 6290 17010 6306
rect 17037 6304 17072 6317
rect 17113 6314 17150 6317
rect 17113 6312 17155 6314
rect 17042 6301 17072 6304
rect 17051 6297 17058 6301
rect 17058 6296 17059 6297
rect 17017 6290 17027 6296
rect 16776 6282 16811 6290
rect 16776 6256 16777 6282
rect 16784 6256 16811 6282
rect 16719 6238 16749 6252
rect 16776 6248 16811 6256
rect 16813 6282 16854 6290
rect 16813 6256 16828 6282
rect 16835 6256 16854 6282
rect 16918 6278 16949 6290
rect 16964 6278 17067 6290
rect 17079 6280 17105 6306
rect 17120 6301 17150 6312
rect 17182 6308 17244 6324
rect 17182 6306 17228 6308
rect 17182 6290 17244 6306
rect 17256 6290 17262 6338
rect 17265 6330 17345 6338
rect 17265 6328 17284 6330
rect 17299 6328 17333 6330
rect 17265 6312 17345 6328
rect 17265 6290 17284 6312
rect 17299 6296 17329 6312
rect 17357 6306 17363 6380
rect 17366 6306 17385 6450
rect 17400 6306 17406 6450
rect 17415 6380 17428 6450
rect 17480 6446 17502 6450
rect 17473 6424 17502 6438
rect 17555 6424 17571 6438
rect 17609 6434 17615 6436
rect 17622 6434 17730 6450
rect 17737 6434 17743 6436
rect 17751 6434 17766 6450
rect 17832 6444 17851 6447
rect 17473 6422 17571 6424
rect 17598 6422 17766 6434
rect 17781 6424 17797 6438
rect 17832 6425 17854 6444
rect 17864 6438 17880 6439
rect 17863 6436 17880 6438
rect 17864 6431 17880 6436
rect 17854 6424 17860 6425
rect 17863 6424 17892 6431
rect 17781 6423 17892 6424
rect 17781 6422 17898 6423
rect 17457 6414 17508 6422
rect 17555 6414 17589 6422
rect 17457 6402 17482 6414
rect 17489 6402 17508 6414
rect 17562 6412 17589 6414
rect 17598 6412 17819 6422
rect 17854 6419 17860 6422
rect 17562 6408 17819 6412
rect 17457 6394 17508 6402
rect 17555 6394 17819 6408
rect 17863 6414 17898 6422
rect 17409 6346 17428 6380
rect 17473 6386 17502 6394
rect 17473 6380 17490 6386
rect 17473 6378 17507 6380
rect 17555 6378 17571 6394
rect 17572 6384 17780 6394
rect 17781 6384 17797 6394
rect 17845 6390 17860 6405
rect 17863 6402 17864 6414
rect 17871 6402 17898 6414
rect 17863 6394 17898 6402
rect 17863 6393 17892 6394
rect 17583 6380 17797 6384
rect 17598 6378 17797 6380
rect 17832 6380 17845 6390
rect 17863 6380 17880 6393
rect 17832 6378 17880 6380
rect 17474 6374 17507 6378
rect 17470 6372 17507 6374
rect 17470 6371 17537 6372
rect 17470 6366 17501 6371
rect 17507 6366 17537 6371
rect 17470 6362 17537 6366
rect 17443 6359 17537 6362
rect 17443 6352 17492 6359
rect 17443 6346 17473 6352
rect 17492 6347 17497 6352
rect 17409 6330 17489 6346
rect 17501 6338 17537 6359
rect 17598 6354 17787 6378
rect 17832 6377 17879 6378
rect 17845 6372 17879 6377
rect 17613 6351 17787 6354
rect 17606 6348 17787 6351
rect 17815 6371 17879 6372
rect 17409 6328 17428 6330
rect 17443 6328 17477 6330
rect 17409 6312 17489 6328
rect 17409 6306 17428 6312
rect 17125 6280 17228 6290
rect 17079 6278 17228 6280
rect 17249 6278 17284 6290
rect 16918 6276 17080 6278
rect 16930 6256 16949 6276
rect 16964 6274 16994 6276
rect 16813 6248 16854 6256
rect 16936 6252 16949 6256
rect 17001 6260 17080 6276
rect 17112 6276 17284 6278
rect 17112 6260 17191 6276
rect 17198 6274 17228 6276
rect 16776 6238 16805 6248
rect 16819 6238 16848 6248
rect 16863 6238 16893 6252
rect 16936 6238 16979 6252
rect 17001 6248 17191 6260
rect 17256 6256 17262 6276
rect 16986 6238 17016 6248
rect 17017 6238 17175 6248
rect 17179 6238 17209 6248
rect 17213 6238 17243 6252
rect 17271 6238 17284 6276
rect 17356 6290 17385 6306
rect 17399 6290 17428 6306
rect 17443 6296 17473 6312
rect 17501 6290 17507 6338
rect 17510 6332 17529 6338
rect 17544 6332 17574 6340
rect 17510 6324 17574 6332
rect 17510 6308 17590 6324
rect 17606 6317 17668 6348
rect 17684 6317 17746 6348
rect 17815 6346 17864 6371
rect 17879 6346 17909 6362
rect 17778 6332 17808 6340
rect 17815 6338 17925 6346
rect 17778 6324 17823 6332
rect 17510 6306 17529 6308
rect 17544 6306 17590 6308
rect 17510 6290 17590 6306
rect 17617 6304 17652 6317
rect 17693 6314 17730 6317
rect 17693 6312 17735 6314
rect 17622 6301 17652 6304
rect 17631 6297 17638 6301
rect 17638 6296 17639 6297
rect 17597 6290 17607 6296
rect 17356 6282 17391 6290
rect 17356 6256 17357 6282
rect 17364 6256 17391 6282
rect 17299 6238 17329 6252
rect 17356 6248 17391 6256
rect 17393 6282 17434 6290
rect 17393 6256 17408 6282
rect 17415 6256 17434 6282
rect 17498 6278 17529 6290
rect 17544 6278 17647 6290
rect 17659 6280 17685 6306
rect 17700 6301 17730 6312
rect 17762 6308 17824 6324
rect 17762 6306 17808 6308
rect 17762 6290 17824 6306
rect 17836 6290 17842 6338
rect 17845 6330 17925 6338
rect 17845 6328 17864 6330
rect 17879 6328 17913 6330
rect 17845 6312 17925 6328
rect 17845 6290 17864 6312
rect 17879 6296 17909 6312
rect 17937 6306 17943 6380
rect 17946 6306 17965 6450
rect 17980 6306 17986 6450
rect 17995 6380 18008 6450
rect 18060 6446 18082 6450
rect 18053 6424 18082 6438
rect 18135 6424 18151 6438
rect 18189 6434 18195 6436
rect 18202 6434 18310 6450
rect 18317 6434 18323 6436
rect 18331 6434 18346 6450
rect 18412 6444 18431 6447
rect 18053 6422 18151 6424
rect 18178 6422 18346 6434
rect 18361 6424 18377 6438
rect 18412 6425 18434 6444
rect 18444 6438 18460 6439
rect 18443 6436 18460 6438
rect 18444 6431 18460 6436
rect 18434 6424 18440 6425
rect 18443 6424 18472 6431
rect 18361 6423 18472 6424
rect 18361 6422 18478 6423
rect 18037 6414 18088 6422
rect 18135 6414 18169 6422
rect 18037 6402 18062 6414
rect 18069 6402 18088 6414
rect 18142 6412 18169 6414
rect 18178 6412 18399 6422
rect 18434 6419 18440 6422
rect 18142 6408 18399 6412
rect 18037 6394 18088 6402
rect 18135 6394 18399 6408
rect 18443 6414 18478 6422
rect 17989 6346 18008 6380
rect 18053 6386 18082 6394
rect 18053 6380 18070 6386
rect 18053 6378 18087 6380
rect 18135 6378 18151 6394
rect 18152 6384 18360 6394
rect 18361 6384 18377 6394
rect 18425 6390 18440 6405
rect 18443 6402 18444 6414
rect 18451 6402 18478 6414
rect 18443 6394 18478 6402
rect 18443 6393 18472 6394
rect 18163 6380 18377 6384
rect 18178 6378 18377 6380
rect 18412 6380 18425 6390
rect 18443 6380 18460 6393
rect 18412 6378 18460 6380
rect 18054 6374 18087 6378
rect 18050 6372 18087 6374
rect 18050 6371 18117 6372
rect 18050 6366 18081 6371
rect 18087 6366 18117 6371
rect 18050 6362 18117 6366
rect 18023 6359 18117 6362
rect 18023 6352 18072 6359
rect 18023 6346 18053 6352
rect 18072 6347 18077 6352
rect 17989 6330 18069 6346
rect 18081 6338 18117 6359
rect 18178 6354 18367 6378
rect 18412 6377 18459 6378
rect 18425 6372 18459 6377
rect 18193 6351 18367 6354
rect 18186 6348 18367 6351
rect 18395 6371 18459 6372
rect 17989 6328 18008 6330
rect 18023 6328 18057 6330
rect 17989 6312 18069 6328
rect 17989 6306 18008 6312
rect 17705 6280 17808 6290
rect 17659 6278 17808 6280
rect 17829 6278 17864 6290
rect 17498 6276 17660 6278
rect 17510 6256 17529 6276
rect 17544 6274 17574 6276
rect 17393 6248 17434 6256
rect 17516 6252 17529 6256
rect 17581 6260 17660 6276
rect 17692 6276 17864 6278
rect 17692 6260 17771 6276
rect 17778 6274 17808 6276
rect 17356 6238 17385 6248
rect 17399 6238 17428 6248
rect 17443 6238 17473 6252
rect 17516 6238 17559 6252
rect 17581 6248 17771 6260
rect 17836 6256 17842 6276
rect 17566 6238 17596 6248
rect 17597 6238 17755 6248
rect 17759 6238 17789 6248
rect 17793 6238 17823 6252
rect 17851 6238 17864 6276
rect 17936 6290 17965 6306
rect 17979 6290 18008 6306
rect 18023 6296 18053 6312
rect 18081 6290 18087 6338
rect 18090 6332 18109 6338
rect 18124 6332 18154 6340
rect 18090 6324 18154 6332
rect 18090 6308 18170 6324
rect 18186 6317 18248 6348
rect 18264 6317 18326 6348
rect 18395 6346 18444 6371
rect 18459 6346 18489 6362
rect 18358 6332 18388 6340
rect 18395 6338 18505 6346
rect 18358 6324 18403 6332
rect 18090 6306 18109 6308
rect 18124 6306 18170 6308
rect 18090 6290 18170 6306
rect 18197 6304 18232 6317
rect 18273 6314 18310 6317
rect 18273 6312 18315 6314
rect 18202 6301 18232 6304
rect 18211 6297 18218 6301
rect 18218 6296 18219 6297
rect 18177 6290 18187 6296
rect 17936 6282 17971 6290
rect 17936 6256 17937 6282
rect 17944 6256 17971 6282
rect 17879 6238 17909 6252
rect 17936 6248 17971 6256
rect 17973 6282 18014 6290
rect 17973 6256 17988 6282
rect 17995 6256 18014 6282
rect 18078 6278 18109 6290
rect 18124 6278 18227 6290
rect 18239 6280 18265 6306
rect 18280 6301 18310 6312
rect 18342 6308 18404 6324
rect 18342 6306 18388 6308
rect 18342 6290 18404 6306
rect 18416 6290 18422 6338
rect 18425 6330 18505 6338
rect 18425 6328 18444 6330
rect 18459 6328 18493 6330
rect 18425 6312 18505 6328
rect 18425 6290 18444 6312
rect 18459 6296 18489 6312
rect 18517 6306 18523 6380
rect 18532 6306 18545 6450
rect 18285 6280 18388 6290
rect 18239 6278 18388 6280
rect 18409 6278 18444 6290
rect 18078 6276 18240 6278
rect 18090 6256 18109 6276
rect 18124 6274 18154 6276
rect 17973 6248 18014 6256
rect 18096 6252 18109 6256
rect 18161 6260 18240 6276
rect 18272 6276 18444 6278
rect 18272 6260 18351 6276
rect 18358 6274 18388 6276
rect 17936 6238 17965 6248
rect 17979 6238 18008 6248
rect 18023 6238 18053 6252
rect 18096 6238 18139 6252
rect 18161 6248 18351 6260
rect 18416 6256 18422 6276
rect 18146 6238 18176 6248
rect 18177 6238 18335 6248
rect 18339 6238 18369 6248
rect 18373 6238 18403 6252
rect 18431 6238 18444 6276
rect 18516 6290 18545 6306
rect 18516 6282 18551 6290
rect 18516 6256 18517 6282
rect 18524 6256 18551 6282
rect 18459 6238 18489 6252
rect 18516 6248 18551 6256
rect 18516 6238 18545 6248
rect -1 6232 18545 6238
rect 0 6224 18545 6232
rect 15 6194 28 6224
rect 43 6210 73 6224
rect 116 6210 159 6224
rect 166 6210 386 6224
rect 393 6210 423 6224
rect 83 6196 98 6208
rect 117 6196 130 6210
rect 198 6206 351 6210
rect 80 6194 102 6196
rect 180 6194 372 6206
rect 451 6194 464 6224
rect 479 6210 509 6224
rect 546 6194 565 6224
rect 580 6194 586 6224
rect 595 6194 608 6224
rect 623 6210 653 6224
rect 696 6210 739 6224
rect 746 6210 966 6224
rect 973 6210 1003 6224
rect 663 6196 678 6208
rect 697 6196 710 6210
rect 778 6206 931 6210
rect 660 6194 682 6196
rect 760 6194 952 6206
rect 1031 6194 1044 6224
rect 1059 6210 1089 6224
rect 1126 6194 1145 6224
rect 1160 6194 1166 6224
rect 1175 6194 1188 6224
rect 1203 6210 1233 6224
rect 1276 6210 1319 6224
rect 1326 6210 1546 6224
rect 1553 6210 1583 6224
rect 1243 6196 1258 6208
rect 1277 6196 1290 6210
rect 1358 6206 1511 6210
rect 1240 6194 1262 6196
rect 1340 6194 1532 6206
rect 1611 6194 1624 6224
rect 1639 6210 1669 6224
rect 1706 6194 1725 6224
rect 1740 6194 1746 6224
rect 1755 6194 1768 6224
rect 1783 6210 1813 6224
rect 1856 6210 1899 6224
rect 1906 6210 2126 6224
rect 2133 6210 2163 6224
rect 1823 6196 1838 6208
rect 1857 6196 1870 6210
rect 1938 6206 2091 6210
rect 1820 6194 1842 6196
rect 1920 6194 2112 6206
rect 2191 6194 2204 6224
rect 2219 6210 2249 6224
rect 2286 6194 2305 6224
rect 2320 6194 2326 6224
rect 2335 6194 2348 6224
rect 2363 6210 2393 6224
rect 2436 6210 2479 6224
rect 2486 6210 2706 6224
rect 2713 6210 2743 6224
rect 2403 6196 2418 6208
rect 2437 6196 2450 6210
rect 2518 6206 2671 6210
rect 2400 6194 2422 6196
rect 2500 6194 2692 6206
rect 2771 6194 2784 6224
rect 2799 6210 2829 6224
rect 2866 6194 2885 6224
rect 2900 6194 2906 6224
rect 2915 6194 2928 6224
rect 2943 6210 2973 6224
rect 3016 6210 3059 6224
rect 3066 6210 3286 6224
rect 3293 6210 3323 6224
rect 2983 6196 2998 6208
rect 3017 6196 3030 6210
rect 3098 6206 3251 6210
rect 2980 6194 3002 6196
rect 3080 6194 3272 6206
rect 3351 6194 3364 6224
rect 3379 6210 3409 6224
rect 3446 6194 3465 6224
rect 3480 6194 3486 6224
rect 3495 6194 3508 6224
rect 3523 6210 3553 6224
rect 3596 6210 3639 6224
rect 3646 6210 3866 6224
rect 3873 6210 3903 6224
rect 3563 6196 3578 6208
rect 3597 6196 3610 6210
rect 3678 6206 3831 6210
rect 3560 6194 3582 6196
rect 3660 6194 3852 6206
rect 3931 6194 3944 6224
rect 3959 6210 3989 6224
rect 4026 6194 4045 6224
rect 4060 6194 4066 6224
rect 4075 6194 4088 6224
rect 4103 6210 4133 6224
rect 4176 6210 4219 6224
rect 4226 6210 4446 6224
rect 4453 6210 4483 6224
rect 4143 6196 4158 6208
rect 4177 6196 4190 6210
rect 4258 6206 4411 6210
rect 4140 6194 4162 6196
rect 4240 6194 4432 6206
rect 4511 6194 4524 6224
rect 4539 6210 4569 6224
rect 4606 6194 4625 6224
rect 4640 6194 4646 6224
rect 4655 6194 4668 6224
rect 4683 6210 4713 6224
rect 4756 6210 4799 6224
rect 4806 6210 5026 6224
rect 5033 6210 5063 6224
rect 4723 6196 4738 6208
rect 4757 6196 4770 6210
rect 4838 6206 4991 6210
rect 4720 6194 4742 6196
rect 4820 6194 5012 6206
rect 5091 6194 5104 6224
rect 5119 6210 5149 6224
rect 5186 6194 5205 6224
rect 5220 6194 5226 6224
rect 5235 6194 5248 6224
rect 5263 6210 5293 6224
rect 5336 6210 5379 6224
rect 5386 6210 5606 6224
rect 5613 6210 5643 6224
rect 5303 6196 5318 6208
rect 5337 6196 5350 6210
rect 5418 6206 5571 6210
rect 5300 6194 5322 6196
rect 5400 6194 5592 6206
rect 5671 6194 5684 6224
rect 5699 6210 5729 6224
rect 5766 6194 5785 6224
rect 5800 6194 5806 6224
rect 5815 6194 5828 6224
rect 5843 6210 5873 6224
rect 5916 6210 5959 6224
rect 5966 6210 6186 6224
rect 6193 6210 6223 6224
rect 5883 6196 5898 6208
rect 5917 6196 5930 6210
rect 5998 6206 6151 6210
rect 5880 6194 5902 6196
rect 5980 6194 6172 6206
rect 6251 6194 6264 6224
rect 6279 6210 6309 6224
rect 6346 6194 6365 6224
rect 6380 6194 6386 6224
rect 6395 6194 6408 6224
rect 6423 6210 6453 6224
rect 6496 6210 6539 6224
rect 6546 6210 6766 6224
rect 6773 6210 6803 6224
rect 6463 6196 6478 6208
rect 6497 6196 6510 6210
rect 6578 6206 6731 6210
rect 6460 6194 6482 6196
rect 6560 6194 6752 6206
rect 6831 6194 6844 6224
rect 6859 6210 6889 6224
rect 6926 6194 6945 6224
rect 6960 6194 6966 6224
rect 6975 6194 6988 6224
rect 7003 6210 7033 6224
rect 7076 6210 7119 6224
rect 7126 6210 7346 6224
rect 7353 6210 7383 6224
rect 7043 6196 7058 6208
rect 7077 6196 7090 6210
rect 7158 6206 7311 6210
rect 7040 6194 7062 6196
rect 7140 6194 7332 6206
rect 7411 6194 7424 6224
rect 7439 6210 7469 6224
rect 7506 6194 7525 6224
rect 7540 6194 7546 6224
rect 7555 6194 7568 6224
rect 7583 6210 7613 6224
rect 7656 6210 7699 6224
rect 7706 6210 7926 6224
rect 7933 6210 7963 6224
rect 7623 6196 7638 6208
rect 7657 6196 7670 6210
rect 7738 6206 7891 6210
rect 7620 6194 7642 6196
rect 7720 6194 7912 6206
rect 7991 6194 8004 6224
rect 8019 6210 8049 6224
rect 8086 6194 8105 6224
rect 8120 6194 8126 6224
rect 8135 6194 8148 6224
rect 8163 6210 8193 6224
rect 8236 6210 8279 6224
rect 8286 6210 8506 6224
rect 8513 6210 8543 6224
rect 8203 6196 8218 6208
rect 8237 6196 8250 6210
rect 8318 6206 8471 6210
rect 8200 6194 8222 6196
rect 8300 6194 8492 6206
rect 8571 6194 8584 6224
rect 8599 6210 8629 6224
rect 8666 6194 8685 6224
rect 8700 6194 8706 6224
rect 8715 6194 8728 6224
rect 8743 6210 8773 6224
rect 8816 6210 8859 6224
rect 8866 6210 9086 6224
rect 9093 6210 9123 6224
rect 8783 6196 8798 6208
rect 8817 6196 8830 6210
rect 8898 6206 9051 6210
rect 8780 6194 8802 6196
rect 8880 6194 9072 6206
rect 9151 6194 9164 6224
rect 9179 6210 9209 6224
rect 9246 6194 9265 6224
rect 9280 6194 9286 6224
rect 9295 6194 9308 6224
rect 9323 6210 9353 6224
rect 9396 6210 9439 6224
rect 9446 6210 9666 6224
rect 9673 6210 9703 6224
rect 9363 6196 9378 6208
rect 9397 6196 9410 6210
rect 9478 6206 9631 6210
rect 9360 6194 9382 6196
rect 9460 6194 9652 6206
rect 9731 6194 9744 6224
rect 9759 6210 9789 6224
rect 9826 6194 9845 6224
rect 9860 6194 9866 6224
rect 9875 6194 9888 6224
rect 9903 6210 9933 6224
rect 9976 6210 10019 6224
rect 10026 6210 10246 6224
rect 10253 6210 10283 6224
rect 9943 6196 9958 6208
rect 9977 6196 9990 6210
rect 10058 6206 10211 6210
rect 9940 6194 9962 6196
rect 10040 6194 10232 6206
rect 10311 6194 10324 6224
rect 10339 6210 10369 6224
rect 10406 6194 10425 6224
rect 10440 6194 10446 6224
rect 10455 6194 10468 6224
rect 10483 6210 10513 6224
rect 10556 6210 10599 6224
rect 10606 6210 10826 6224
rect 10833 6210 10863 6224
rect 10523 6196 10538 6208
rect 10557 6196 10570 6210
rect 10638 6206 10791 6210
rect 10520 6194 10542 6196
rect 10620 6194 10812 6206
rect 10891 6194 10904 6224
rect 10919 6210 10949 6224
rect 10986 6194 11005 6224
rect 11020 6194 11026 6224
rect 11035 6194 11048 6224
rect 11063 6210 11093 6224
rect 11136 6210 11179 6224
rect 11186 6210 11406 6224
rect 11413 6210 11443 6224
rect 11103 6196 11118 6208
rect 11137 6196 11150 6210
rect 11218 6206 11371 6210
rect 11100 6194 11122 6196
rect 11200 6194 11392 6206
rect 11471 6194 11484 6224
rect 11499 6210 11529 6224
rect 11566 6194 11585 6224
rect 11600 6194 11606 6224
rect 11615 6194 11628 6224
rect 11643 6210 11673 6224
rect 11716 6210 11759 6224
rect 11766 6210 11986 6224
rect 11993 6210 12023 6224
rect 11683 6196 11698 6208
rect 11717 6196 11730 6210
rect 11798 6206 11951 6210
rect 11680 6194 11702 6196
rect 11780 6194 11972 6206
rect 12051 6194 12064 6224
rect 12079 6210 12109 6224
rect 12146 6194 12165 6224
rect 12180 6194 12186 6224
rect 12195 6194 12208 6224
rect 12223 6210 12253 6224
rect 12296 6210 12339 6224
rect 12346 6210 12566 6224
rect 12573 6210 12603 6224
rect 12263 6196 12278 6208
rect 12297 6196 12310 6210
rect 12378 6206 12531 6210
rect 12260 6194 12282 6196
rect 12360 6194 12552 6206
rect 12631 6194 12644 6224
rect 12659 6210 12689 6224
rect 12726 6194 12745 6224
rect 12760 6194 12766 6224
rect 12775 6194 12788 6224
rect 12803 6210 12833 6224
rect 12876 6210 12919 6224
rect 12926 6210 13146 6224
rect 13153 6210 13183 6224
rect 12843 6196 12858 6208
rect 12877 6196 12890 6210
rect 12958 6206 13111 6210
rect 12840 6194 12862 6196
rect 12940 6194 13132 6206
rect 13211 6194 13224 6224
rect 13239 6210 13269 6224
rect 13306 6194 13325 6224
rect 13340 6194 13346 6224
rect 13355 6194 13368 6224
rect 13383 6210 13413 6224
rect 13456 6210 13499 6224
rect 13506 6210 13726 6224
rect 13733 6210 13763 6224
rect 13423 6196 13438 6208
rect 13457 6196 13470 6210
rect 13538 6206 13691 6210
rect 13420 6194 13442 6196
rect 13520 6194 13712 6206
rect 13791 6194 13804 6224
rect 13819 6210 13849 6224
rect 13886 6194 13905 6224
rect 13920 6194 13926 6224
rect 13935 6194 13948 6224
rect 13963 6210 13993 6224
rect 14036 6210 14079 6224
rect 14086 6210 14306 6224
rect 14313 6210 14343 6224
rect 14003 6196 14018 6208
rect 14037 6196 14050 6210
rect 14118 6206 14271 6210
rect 14000 6194 14022 6196
rect 14100 6194 14292 6206
rect 14371 6194 14384 6224
rect 14399 6210 14429 6224
rect 14466 6194 14485 6224
rect 14500 6194 14506 6224
rect 14515 6194 14528 6224
rect 14543 6210 14573 6224
rect 14616 6210 14659 6224
rect 14666 6210 14886 6224
rect 14893 6210 14923 6224
rect 14583 6196 14598 6208
rect 14617 6196 14630 6210
rect 14698 6206 14851 6210
rect 14580 6194 14602 6196
rect 14680 6194 14872 6206
rect 14951 6194 14964 6224
rect 14979 6210 15009 6224
rect 15046 6194 15065 6224
rect 15080 6194 15086 6224
rect 15095 6194 15108 6224
rect 15123 6210 15153 6224
rect 15196 6210 15239 6224
rect 15246 6210 15466 6224
rect 15473 6210 15503 6224
rect 15163 6196 15178 6208
rect 15197 6196 15210 6210
rect 15278 6206 15431 6210
rect 15160 6194 15182 6196
rect 15260 6194 15452 6206
rect 15531 6194 15544 6224
rect 15559 6210 15589 6224
rect 15626 6194 15645 6224
rect 15660 6194 15666 6224
rect 15675 6194 15688 6224
rect 15703 6210 15733 6224
rect 15776 6210 15819 6224
rect 15826 6210 16046 6224
rect 16053 6210 16083 6224
rect 15743 6196 15758 6208
rect 15777 6196 15790 6210
rect 15858 6206 16011 6210
rect 15740 6194 15762 6196
rect 15840 6194 16032 6206
rect 16111 6194 16124 6224
rect 16139 6210 16169 6224
rect 16206 6194 16225 6224
rect 16240 6194 16246 6224
rect 16255 6194 16268 6224
rect 16283 6210 16313 6224
rect 16356 6210 16399 6224
rect 16406 6210 16626 6224
rect 16633 6210 16663 6224
rect 16323 6196 16338 6208
rect 16357 6196 16370 6210
rect 16438 6206 16591 6210
rect 16320 6194 16342 6196
rect 16420 6194 16612 6206
rect 16691 6194 16704 6224
rect 16719 6210 16749 6224
rect 16786 6194 16805 6224
rect 16820 6194 16826 6224
rect 16835 6194 16848 6224
rect 16863 6210 16893 6224
rect 16936 6210 16979 6224
rect 16986 6210 17206 6224
rect 17213 6210 17243 6224
rect 16903 6196 16918 6208
rect 16937 6196 16950 6210
rect 17018 6206 17171 6210
rect 16900 6194 16922 6196
rect 17000 6194 17192 6206
rect 17271 6194 17284 6224
rect 17299 6210 17329 6224
rect 17366 6194 17385 6224
rect 17400 6194 17406 6224
rect 17415 6194 17428 6224
rect 17443 6210 17473 6224
rect 17516 6210 17559 6224
rect 17566 6210 17786 6224
rect 17793 6210 17823 6224
rect 17483 6196 17498 6208
rect 17517 6196 17530 6210
rect 17598 6206 17751 6210
rect 17480 6194 17502 6196
rect 17580 6194 17772 6206
rect 17851 6194 17864 6224
rect 17879 6210 17909 6224
rect 17946 6194 17965 6224
rect 17980 6194 17986 6224
rect 17995 6194 18008 6224
rect 18023 6210 18053 6224
rect 18096 6210 18139 6224
rect 18146 6210 18366 6224
rect 18373 6210 18403 6224
rect 18063 6196 18078 6208
rect 18097 6196 18110 6210
rect 18178 6206 18331 6210
rect 18060 6194 18082 6196
rect 18160 6194 18352 6206
rect 18431 6194 18444 6224
rect 18459 6210 18489 6224
rect 18532 6194 18545 6224
rect 0 6180 18545 6194
rect 15 6110 28 6180
rect 80 6176 102 6180
rect 73 6154 102 6168
rect 155 6154 171 6168
rect 209 6164 215 6166
rect 222 6164 330 6180
rect 337 6164 343 6166
rect 351 6164 366 6180
rect 432 6174 451 6177
rect 73 6152 171 6154
rect 198 6152 366 6164
rect 381 6154 397 6168
rect 432 6155 454 6174
rect 464 6168 480 6169
rect 463 6166 480 6168
rect 464 6161 480 6166
rect 454 6154 460 6155
rect 463 6154 492 6161
rect 381 6153 492 6154
rect 381 6152 498 6153
rect 57 6144 108 6152
rect 155 6144 189 6152
rect 57 6132 82 6144
rect 89 6132 108 6144
rect 162 6142 189 6144
rect 198 6142 419 6152
rect 454 6149 460 6152
rect 162 6138 419 6142
rect 57 6124 108 6132
rect 155 6124 419 6138
rect 463 6144 498 6152
rect 9 6076 28 6110
rect 73 6116 102 6124
rect 73 6110 90 6116
rect 73 6108 107 6110
rect 155 6108 171 6124
rect 172 6114 380 6124
rect 381 6114 397 6124
rect 445 6120 460 6135
rect 463 6132 464 6144
rect 471 6132 498 6144
rect 463 6124 498 6132
rect 463 6123 492 6124
rect 183 6110 397 6114
rect 198 6108 397 6110
rect 432 6110 445 6120
rect 463 6110 480 6123
rect 432 6108 480 6110
rect 74 6104 107 6108
rect 70 6102 107 6104
rect 70 6101 137 6102
rect 70 6096 101 6101
rect 107 6096 137 6101
rect 70 6092 137 6096
rect 43 6089 137 6092
rect 43 6082 92 6089
rect 43 6076 73 6082
rect 92 6077 97 6082
rect 9 6060 89 6076
rect 101 6068 137 6089
rect 198 6084 387 6108
rect 432 6107 479 6108
rect 445 6102 479 6107
rect 213 6081 387 6084
rect 206 6078 387 6081
rect 415 6101 479 6102
rect 9 6058 28 6060
rect 43 6058 77 6060
rect 9 6042 89 6058
rect 9 6036 28 6042
rect -1 6020 28 6036
rect 43 6026 73 6042
rect 101 6020 107 6068
rect 110 6062 129 6068
rect 144 6062 174 6070
rect 110 6054 174 6062
rect 110 6038 190 6054
rect 206 6047 268 6078
rect 284 6047 346 6078
rect 415 6076 464 6101
rect 479 6076 509 6092
rect 378 6062 408 6070
rect 415 6068 525 6076
rect 378 6054 423 6062
rect 110 6036 129 6038
rect 144 6036 190 6038
rect 110 6020 190 6036
rect 217 6034 252 6047
rect 293 6044 330 6047
rect 293 6042 335 6044
rect 222 6031 252 6034
rect 231 6027 238 6031
rect 238 6026 239 6027
rect 197 6020 207 6026
rect -7 6012 34 6020
rect -7 5986 8 6012
rect 15 5986 34 6012
rect 98 6008 129 6020
rect 144 6008 247 6020
rect 259 6010 285 6036
rect 300 6031 330 6042
rect 362 6038 424 6054
rect 362 6036 408 6038
rect 362 6020 424 6036
rect 436 6020 442 6068
rect 445 6060 525 6068
rect 445 6058 464 6060
rect 479 6058 513 6060
rect 445 6042 525 6058
rect 445 6020 464 6042
rect 479 6026 509 6042
rect 537 6036 543 6110
rect 546 6036 565 6180
rect 580 6036 586 6180
rect 595 6110 608 6180
rect 660 6176 682 6180
rect 653 6154 682 6168
rect 735 6154 751 6168
rect 789 6164 795 6166
rect 802 6164 910 6180
rect 917 6164 923 6166
rect 931 6164 946 6180
rect 1012 6174 1031 6177
rect 653 6152 751 6154
rect 778 6152 946 6164
rect 961 6154 977 6168
rect 1012 6155 1034 6174
rect 1044 6168 1060 6169
rect 1043 6166 1060 6168
rect 1044 6161 1060 6166
rect 1034 6154 1040 6155
rect 1043 6154 1072 6161
rect 961 6153 1072 6154
rect 961 6152 1078 6153
rect 637 6144 688 6152
rect 735 6144 769 6152
rect 637 6132 662 6144
rect 669 6132 688 6144
rect 742 6142 769 6144
rect 778 6142 999 6152
rect 1034 6149 1040 6152
rect 742 6138 999 6142
rect 637 6124 688 6132
rect 735 6124 999 6138
rect 1043 6144 1078 6152
rect 589 6076 608 6110
rect 653 6116 682 6124
rect 653 6110 670 6116
rect 653 6108 687 6110
rect 735 6108 751 6124
rect 752 6114 960 6124
rect 961 6114 977 6124
rect 1025 6120 1040 6135
rect 1043 6132 1044 6144
rect 1051 6132 1078 6144
rect 1043 6124 1078 6132
rect 1043 6123 1072 6124
rect 763 6110 977 6114
rect 778 6108 977 6110
rect 1012 6110 1025 6120
rect 1043 6110 1060 6123
rect 1012 6108 1060 6110
rect 654 6104 687 6108
rect 650 6102 687 6104
rect 650 6101 717 6102
rect 650 6096 681 6101
rect 687 6096 717 6101
rect 650 6092 717 6096
rect 623 6089 717 6092
rect 623 6082 672 6089
rect 623 6076 653 6082
rect 672 6077 677 6082
rect 589 6060 669 6076
rect 681 6068 717 6089
rect 778 6084 967 6108
rect 1012 6107 1059 6108
rect 1025 6102 1059 6107
rect 793 6081 967 6084
rect 786 6078 967 6081
rect 995 6101 1059 6102
rect 589 6058 608 6060
rect 623 6058 657 6060
rect 589 6042 669 6058
rect 589 6036 608 6042
rect 305 6010 408 6020
rect 259 6008 408 6010
rect 429 6008 464 6020
rect 98 6006 260 6008
rect 110 5986 129 6006
rect 144 6004 174 6006
rect -7 5978 34 5986
rect 116 5982 129 5986
rect 181 5990 260 6006
rect 292 6006 464 6008
rect 292 5990 371 6006
rect 378 6004 408 6006
rect -1 5968 28 5978
rect 43 5968 73 5982
rect 116 5968 159 5982
rect 181 5978 371 5990
rect 436 5986 442 6006
rect 166 5968 196 5978
rect 197 5968 355 5978
rect 359 5968 389 5978
rect 393 5968 423 5982
rect 451 5968 464 6006
rect 536 6020 565 6036
rect 579 6020 608 6036
rect 623 6026 653 6042
rect 681 6020 687 6068
rect 690 6062 709 6068
rect 724 6062 754 6070
rect 690 6054 754 6062
rect 690 6038 770 6054
rect 786 6047 848 6078
rect 864 6047 926 6078
rect 995 6076 1044 6101
rect 1059 6076 1089 6092
rect 958 6062 988 6070
rect 995 6068 1105 6076
rect 958 6054 1003 6062
rect 690 6036 709 6038
rect 724 6036 770 6038
rect 690 6020 770 6036
rect 797 6034 832 6047
rect 873 6044 910 6047
rect 873 6042 915 6044
rect 802 6031 832 6034
rect 811 6027 818 6031
rect 818 6026 819 6027
rect 777 6020 787 6026
rect 536 6012 571 6020
rect 536 5986 537 6012
rect 544 5986 571 6012
rect 479 5968 509 5982
rect 536 5978 571 5986
rect 573 6012 614 6020
rect 573 5986 588 6012
rect 595 5986 614 6012
rect 678 6008 709 6020
rect 724 6008 827 6020
rect 839 6010 865 6036
rect 880 6031 910 6042
rect 942 6038 1004 6054
rect 942 6036 988 6038
rect 942 6020 1004 6036
rect 1016 6020 1022 6068
rect 1025 6060 1105 6068
rect 1025 6058 1044 6060
rect 1059 6058 1093 6060
rect 1025 6042 1105 6058
rect 1025 6020 1044 6042
rect 1059 6026 1089 6042
rect 1117 6036 1123 6110
rect 1126 6036 1145 6180
rect 1160 6036 1166 6180
rect 1175 6110 1188 6180
rect 1240 6176 1262 6180
rect 1233 6154 1262 6168
rect 1315 6154 1331 6168
rect 1369 6164 1375 6166
rect 1382 6164 1490 6180
rect 1497 6164 1503 6166
rect 1511 6164 1526 6180
rect 1592 6174 1611 6177
rect 1233 6152 1331 6154
rect 1358 6152 1526 6164
rect 1541 6154 1557 6168
rect 1592 6155 1614 6174
rect 1624 6168 1640 6169
rect 1623 6166 1640 6168
rect 1624 6161 1640 6166
rect 1614 6154 1620 6155
rect 1623 6154 1652 6161
rect 1541 6153 1652 6154
rect 1541 6152 1658 6153
rect 1217 6144 1268 6152
rect 1315 6144 1349 6152
rect 1217 6132 1242 6144
rect 1249 6132 1268 6144
rect 1322 6142 1349 6144
rect 1358 6142 1579 6152
rect 1614 6149 1620 6152
rect 1322 6138 1579 6142
rect 1217 6124 1268 6132
rect 1315 6124 1579 6138
rect 1623 6144 1658 6152
rect 1169 6076 1188 6110
rect 1233 6116 1262 6124
rect 1233 6110 1250 6116
rect 1233 6108 1267 6110
rect 1315 6108 1331 6124
rect 1332 6114 1540 6124
rect 1541 6114 1557 6124
rect 1605 6120 1620 6135
rect 1623 6132 1624 6144
rect 1631 6132 1658 6144
rect 1623 6124 1658 6132
rect 1623 6123 1652 6124
rect 1343 6110 1557 6114
rect 1358 6108 1557 6110
rect 1592 6110 1605 6120
rect 1623 6110 1640 6123
rect 1592 6108 1640 6110
rect 1234 6104 1267 6108
rect 1230 6102 1267 6104
rect 1230 6101 1297 6102
rect 1230 6096 1261 6101
rect 1267 6096 1297 6101
rect 1230 6092 1297 6096
rect 1203 6089 1297 6092
rect 1203 6082 1252 6089
rect 1203 6076 1233 6082
rect 1252 6077 1257 6082
rect 1169 6060 1249 6076
rect 1261 6068 1297 6089
rect 1358 6084 1547 6108
rect 1592 6107 1639 6108
rect 1605 6102 1639 6107
rect 1373 6081 1547 6084
rect 1366 6078 1547 6081
rect 1575 6101 1639 6102
rect 1169 6058 1188 6060
rect 1203 6058 1237 6060
rect 1169 6042 1249 6058
rect 1169 6036 1188 6042
rect 885 6010 988 6020
rect 839 6008 988 6010
rect 1009 6008 1044 6020
rect 678 6006 840 6008
rect 690 5986 709 6006
rect 724 6004 754 6006
rect 573 5978 614 5986
rect 696 5982 709 5986
rect 761 5990 840 6006
rect 872 6006 1044 6008
rect 872 5990 951 6006
rect 958 6004 988 6006
rect 536 5968 565 5978
rect 579 5968 608 5978
rect 623 5968 653 5982
rect 696 5968 739 5982
rect 761 5978 951 5990
rect 1016 5986 1022 6006
rect 746 5968 776 5978
rect 777 5968 935 5978
rect 939 5968 969 5978
rect 973 5968 1003 5982
rect 1031 5968 1044 6006
rect 1116 6020 1145 6036
rect 1159 6020 1188 6036
rect 1203 6026 1233 6042
rect 1261 6020 1267 6068
rect 1270 6062 1289 6068
rect 1304 6062 1334 6070
rect 1270 6054 1334 6062
rect 1270 6038 1350 6054
rect 1366 6047 1428 6078
rect 1444 6047 1506 6078
rect 1575 6076 1624 6101
rect 1639 6076 1669 6092
rect 1538 6062 1568 6070
rect 1575 6068 1685 6076
rect 1538 6054 1583 6062
rect 1270 6036 1289 6038
rect 1304 6036 1350 6038
rect 1270 6020 1350 6036
rect 1377 6034 1412 6047
rect 1453 6044 1490 6047
rect 1453 6042 1495 6044
rect 1382 6031 1412 6034
rect 1391 6027 1398 6031
rect 1398 6026 1399 6027
rect 1357 6020 1367 6026
rect 1116 6012 1151 6020
rect 1116 5986 1117 6012
rect 1124 5986 1151 6012
rect 1059 5968 1089 5982
rect 1116 5978 1151 5986
rect 1153 6012 1194 6020
rect 1153 5986 1168 6012
rect 1175 5986 1194 6012
rect 1258 6008 1289 6020
rect 1304 6008 1407 6020
rect 1419 6010 1445 6036
rect 1460 6031 1490 6042
rect 1522 6038 1584 6054
rect 1522 6036 1568 6038
rect 1522 6020 1584 6036
rect 1596 6020 1602 6068
rect 1605 6060 1685 6068
rect 1605 6058 1624 6060
rect 1639 6058 1673 6060
rect 1605 6042 1685 6058
rect 1605 6020 1624 6042
rect 1639 6026 1669 6042
rect 1697 6036 1703 6110
rect 1706 6036 1725 6180
rect 1740 6036 1746 6180
rect 1755 6110 1768 6180
rect 1820 6176 1842 6180
rect 1813 6154 1842 6168
rect 1895 6154 1911 6168
rect 1949 6164 1955 6166
rect 1962 6164 2070 6180
rect 2077 6164 2083 6166
rect 2091 6164 2106 6180
rect 2172 6174 2191 6177
rect 1813 6152 1911 6154
rect 1938 6152 2106 6164
rect 2121 6154 2137 6168
rect 2172 6155 2194 6174
rect 2204 6168 2220 6169
rect 2203 6166 2220 6168
rect 2204 6161 2220 6166
rect 2194 6154 2200 6155
rect 2203 6154 2232 6161
rect 2121 6153 2232 6154
rect 2121 6152 2238 6153
rect 1797 6144 1848 6152
rect 1895 6144 1929 6152
rect 1797 6132 1822 6144
rect 1829 6132 1848 6144
rect 1902 6142 1929 6144
rect 1938 6142 2159 6152
rect 2194 6149 2200 6152
rect 1902 6138 2159 6142
rect 1797 6124 1848 6132
rect 1895 6124 2159 6138
rect 2203 6144 2238 6152
rect 1749 6076 1768 6110
rect 1813 6116 1842 6124
rect 1813 6110 1830 6116
rect 1813 6108 1847 6110
rect 1895 6108 1911 6124
rect 1912 6114 2120 6124
rect 2121 6114 2137 6124
rect 2185 6120 2200 6135
rect 2203 6132 2204 6144
rect 2211 6132 2238 6144
rect 2203 6124 2238 6132
rect 2203 6123 2232 6124
rect 1923 6110 2137 6114
rect 1938 6108 2137 6110
rect 2172 6110 2185 6120
rect 2203 6110 2220 6123
rect 2172 6108 2220 6110
rect 1814 6104 1847 6108
rect 1810 6102 1847 6104
rect 1810 6101 1877 6102
rect 1810 6096 1841 6101
rect 1847 6096 1877 6101
rect 1810 6092 1877 6096
rect 1783 6089 1877 6092
rect 1783 6082 1832 6089
rect 1783 6076 1813 6082
rect 1832 6077 1837 6082
rect 1749 6060 1829 6076
rect 1841 6068 1877 6089
rect 1938 6084 2127 6108
rect 2172 6107 2219 6108
rect 2185 6102 2219 6107
rect 1953 6081 2127 6084
rect 1946 6078 2127 6081
rect 2155 6101 2219 6102
rect 1749 6058 1768 6060
rect 1783 6058 1817 6060
rect 1749 6042 1829 6058
rect 1749 6036 1768 6042
rect 1465 6010 1568 6020
rect 1419 6008 1568 6010
rect 1589 6008 1624 6020
rect 1258 6006 1420 6008
rect 1270 5986 1289 6006
rect 1304 6004 1334 6006
rect 1153 5978 1194 5986
rect 1276 5982 1289 5986
rect 1341 5990 1420 6006
rect 1452 6006 1624 6008
rect 1452 5990 1531 6006
rect 1538 6004 1568 6006
rect 1116 5968 1145 5978
rect 1159 5968 1188 5978
rect 1203 5968 1233 5982
rect 1276 5968 1319 5982
rect 1341 5978 1531 5990
rect 1596 5986 1602 6006
rect 1326 5968 1356 5978
rect 1357 5968 1515 5978
rect 1519 5968 1549 5978
rect 1553 5968 1583 5982
rect 1611 5968 1624 6006
rect 1696 6020 1725 6036
rect 1739 6020 1768 6036
rect 1783 6026 1813 6042
rect 1841 6020 1847 6068
rect 1850 6062 1869 6068
rect 1884 6062 1914 6070
rect 1850 6054 1914 6062
rect 1850 6038 1930 6054
rect 1946 6047 2008 6078
rect 2024 6047 2086 6078
rect 2155 6076 2204 6101
rect 2219 6076 2249 6092
rect 2118 6062 2148 6070
rect 2155 6068 2265 6076
rect 2118 6054 2163 6062
rect 1850 6036 1869 6038
rect 1884 6036 1930 6038
rect 1850 6020 1930 6036
rect 1957 6034 1992 6047
rect 2033 6044 2070 6047
rect 2033 6042 2075 6044
rect 1962 6031 1992 6034
rect 1971 6027 1978 6031
rect 1978 6026 1979 6027
rect 1937 6020 1947 6026
rect 1696 6012 1731 6020
rect 1696 5986 1697 6012
rect 1704 5986 1731 6012
rect 1639 5968 1669 5982
rect 1696 5978 1731 5986
rect 1733 6012 1774 6020
rect 1733 5986 1748 6012
rect 1755 5986 1774 6012
rect 1838 6008 1869 6020
rect 1884 6008 1987 6020
rect 1999 6010 2025 6036
rect 2040 6031 2070 6042
rect 2102 6038 2164 6054
rect 2102 6036 2148 6038
rect 2102 6020 2164 6036
rect 2176 6020 2182 6068
rect 2185 6060 2265 6068
rect 2185 6058 2204 6060
rect 2219 6058 2253 6060
rect 2185 6042 2265 6058
rect 2185 6020 2204 6042
rect 2219 6026 2249 6042
rect 2277 6036 2283 6110
rect 2286 6036 2305 6180
rect 2320 6036 2326 6180
rect 2335 6110 2348 6180
rect 2400 6176 2422 6180
rect 2393 6154 2422 6168
rect 2475 6154 2491 6168
rect 2529 6164 2535 6166
rect 2542 6164 2650 6180
rect 2657 6164 2663 6166
rect 2671 6164 2686 6180
rect 2752 6174 2771 6177
rect 2393 6152 2491 6154
rect 2518 6152 2686 6164
rect 2701 6154 2717 6168
rect 2752 6155 2774 6174
rect 2784 6168 2800 6169
rect 2783 6166 2800 6168
rect 2784 6161 2800 6166
rect 2774 6154 2780 6155
rect 2783 6154 2812 6161
rect 2701 6153 2812 6154
rect 2701 6152 2818 6153
rect 2377 6144 2428 6152
rect 2475 6144 2509 6152
rect 2377 6132 2402 6144
rect 2409 6132 2428 6144
rect 2482 6142 2509 6144
rect 2518 6142 2739 6152
rect 2774 6149 2780 6152
rect 2482 6138 2739 6142
rect 2377 6124 2428 6132
rect 2475 6124 2739 6138
rect 2783 6144 2818 6152
rect 2329 6076 2348 6110
rect 2393 6116 2422 6124
rect 2393 6110 2410 6116
rect 2393 6108 2427 6110
rect 2475 6108 2491 6124
rect 2492 6114 2700 6124
rect 2701 6114 2717 6124
rect 2765 6120 2780 6135
rect 2783 6132 2784 6144
rect 2791 6132 2818 6144
rect 2783 6124 2818 6132
rect 2783 6123 2812 6124
rect 2503 6110 2717 6114
rect 2518 6108 2717 6110
rect 2752 6110 2765 6120
rect 2783 6110 2800 6123
rect 2752 6108 2800 6110
rect 2394 6104 2427 6108
rect 2390 6102 2427 6104
rect 2390 6101 2457 6102
rect 2390 6096 2421 6101
rect 2427 6096 2457 6101
rect 2390 6092 2457 6096
rect 2363 6089 2457 6092
rect 2363 6082 2412 6089
rect 2363 6076 2393 6082
rect 2412 6077 2417 6082
rect 2329 6060 2409 6076
rect 2421 6068 2457 6089
rect 2518 6084 2707 6108
rect 2752 6107 2799 6108
rect 2765 6102 2799 6107
rect 2533 6081 2707 6084
rect 2526 6078 2707 6081
rect 2735 6101 2799 6102
rect 2329 6058 2348 6060
rect 2363 6058 2397 6060
rect 2329 6042 2409 6058
rect 2329 6036 2348 6042
rect 2045 6010 2148 6020
rect 1999 6008 2148 6010
rect 2169 6008 2204 6020
rect 1838 6006 2000 6008
rect 1850 5986 1869 6006
rect 1884 6004 1914 6006
rect 1733 5978 1774 5986
rect 1856 5982 1869 5986
rect 1921 5990 2000 6006
rect 2032 6006 2204 6008
rect 2032 5990 2111 6006
rect 2118 6004 2148 6006
rect 1696 5968 1725 5978
rect 1739 5968 1768 5978
rect 1783 5968 1813 5982
rect 1856 5968 1899 5982
rect 1921 5978 2111 5990
rect 2176 5986 2182 6006
rect 1906 5968 1936 5978
rect 1937 5968 2095 5978
rect 2099 5968 2129 5978
rect 2133 5968 2163 5982
rect 2191 5968 2204 6006
rect 2276 6020 2305 6036
rect 2319 6020 2348 6036
rect 2363 6026 2393 6042
rect 2421 6020 2427 6068
rect 2430 6062 2449 6068
rect 2464 6062 2494 6070
rect 2430 6054 2494 6062
rect 2430 6038 2510 6054
rect 2526 6047 2588 6078
rect 2604 6047 2666 6078
rect 2735 6076 2784 6101
rect 2799 6076 2829 6092
rect 2698 6062 2728 6070
rect 2735 6068 2845 6076
rect 2698 6054 2743 6062
rect 2430 6036 2449 6038
rect 2464 6036 2510 6038
rect 2430 6020 2510 6036
rect 2537 6034 2572 6047
rect 2613 6044 2650 6047
rect 2613 6042 2655 6044
rect 2542 6031 2572 6034
rect 2551 6027 2558 6031
rect 2558 6026 2559 6027
rect 2517 6020 2527 6026
rect 2276 6012 2311 6020
rect 2276 5986 2277 6012
rect 2284 5986 2311 6012
rect 2219 5968 2249 5982
rect 2276 5978 2311 5986
rect 2313 6012 2354 6020
rect 2313 5986 2328 6012
rect 2335 5986 2354 6012
rect 2418 6008 2449 6020
rect 2464 6008 2567 6020
rect 2579 6010 2605 6036
rect 2620 6031 2650 6042
rect 2682 6038 2744 6054
rect 2682 6036 2728 6038
rect 2682 6020 2744 6036
rect 2756 6020 2762 6068
rect 2765 6060 2845 6068
rect 2765 6058 2784 6060
rect 2799 6058 2833 6060
rect 2765 6042 2845 6058
rect 2765 6020 2784 6042
rect 2799 6026 2829 6042
rect 2857 6036 2863 6110
rect 2866 6036 2885 6180
rect 2900 6036 2906 6180
rect 2915 6110 2928 6180
rect 2980 6176 3002 6180
rect 2973 6154 3002 6168
rect 3055 6154 3071 6168
rect 3109 6164 3115 6166
rect 3122 6164 3230 6180
rect 3237 6164 3243 6166
rect 3251 6164 3266 6180
rect 3332 6174 3351 6177
rect 2973 6152 3071 6154
rect 3098 6152 3266 6164
rect 3281 6154 3297 6168
rect 3332 6155 3354 6174
rect 3364 6168 3380 6169
rect 3363 6166 3380 6168
rect 3364 6161 3380 6166
rect 3354 6154 3360 6155
rect 3363 6154 3392 6161
rect 3281 6153 3392 6154
rect 3281 6152 3398 6153
rect 2957 6144 3008 6152
rect 3055 6144 3089 6152
rect 2957 6132 2982 6144
rect 2989 6132 3008 6144
rect 3062 6142 3089 6144
rect 3098 6142 3319 6152
rect 3354 6149 3360 6152
rect 3062 6138 3319 6142
rect 2957 6124 3008 6132
rect 3055 6124 3319 6138
rect 3363 6144 3398 6152
rect 2909 6076 2928 6110
rect 2973 6116 3002 6124
rect 2973 6110 2990 6116
rect 2973 6108 3007 6110
rect 3055 6108 3071 6124
rect 3072 6114 3280 6124
rect 3281 6114 3297 6124
rect 3345 6120 3360 6135
rect 3363 6132 3364 6144
rect 3371 6132 3398 6144
rect 3363 6124 3398 6132
rect 3363 6123 3392 6124
rect 3083 6110 3297 6114
rect 3098 6108 3297 6110
rect 3332 6110 3345 6120
rect 3363 6110 3380 6123
rect 3332 6108 3380 6110
rect 2974 6104 3007 6108
rect 2970 6102 3007 6104
rect 2970 6101 3037 6102
rect 2970 6096 3001 6101
rect 3007 6096 3037 6101
rect 2970 6092 3037 6096
rect 2943 6089 3037 6092
rect 2943 6082 2992 6089
rect 2943 6076 2973 6082
rect 2992 6077 2997 6082
rect 2909 6060 2989 6076
rect 3001 6068 3037 6089
rect 3098 6084 3287 6108
rect 3332 6107 3379 6108
rect 3345 6102 3379 6107
rect 3113 6081 3287 6084
rect 3106 6078 3287 6081
rect 3315 6101 3379 6102
rect 2909 6058 2928 6060
rect 2943 6058 2977 6060
rect 2909 6042 2989 6058
rect 2909 6036 2928 6042
rect 2625 6010 2728 6020
rect 2579 6008 2728 6010
rect 2749 6008 2784 6020
rect 2418 6006 2580 6008
rect 2430 5986 2449 6006
rect 2464 6004 2494 6006
rect 2313 5978 2354 5986
rect 2436 5982 2449 5986
rect 2501 5990 2580 6006
rect 2612 6006 2784 6008
rect 2612 5990 2691 6006
rect 2698 6004 2728 6006
rect 2276 5968 2305 5978
rect 2319 5968 2348 5978
rect 2363 5968 2393 5982
rect 2436 5968 2479 5982
rect 2501 5978 2691 5990
rect 2756 5986 2762 6006
rect 2486 5968 2516 5978
rect 2517 5968 2675 5978
rect 2679 5968 2709 5978
rect 2713 5968 2743 5982
rect 2771 5968 2784 6006
rect 2856 6020 2885 6036
rect 2899 6020 2928 6036
rect 2943 6026 2973 6042
rect 3001 6020 3007 6068
rect 3010 6062 3029 6068
rect 3044 6062 3074 6070
rect 3010 6054 3074 6062
rect 3010 6038 3090 6054
rect 3106 6047 3168 6078
rect 3184 6047 3246 6078
rect 3315 6076 3364 6101
rect 3379 6076 3409 6092
rect 3278 6062 3308 6070
rect 3315 6068 3425 6076
rect 3278 6054 3323 6062
rect 3010 6036 3029 6038
rect 3044 6036 3090 6038
rect 3010 6020 3090 6036
rect 3117 6034 3152 6047
rect 3193 6044 3230 6047
rect 3193 6042 3235 6044
rect 3122 6031 3152 6034
rect 3131 6027 3138 6031
rect 3138 6026 3139 6027
rect 3097 6020 3107 6026
rect 2856 6012 2891 6020
rect 2856 5986 2857 6012
rect 2864 5986 2891 6012
rect 2799 5968 2829 5982
rect 2856 5978 2891 5986
rect 2893 6012 2934 6020
rect 2893 5986 2908 6012
rect 2915 5986 2934 6012
rect 2998 6008 3029 6020
rect 3044 6008 3147 6020
rect 3159 6010 3185 6036
rect 3200 6031 3230 6042
rect 3262 6038 3324 6054
rect 3262 6036 3308 6038
rect 3262 6020 3324 6036
rect 3336 6020 3342 6068
rect 3345 6060 3425 6068
rect 3345 6058 3364 6060
rect 3379 6058 3413 6060
rect 3345 6042 3425 6058
rect 3345 6020 3364 6042
rect 3379 6026 3409 6042
rect 3437 6036 3443 6110
rect 3446 6036 3465 6180
rect 3480 6036 3486 6180
rect 3495 6110 3508 6180
rect 3560 6176 3582 6180
rect 3553 6154 3582 6168
rect 3635 6154 3651 6168
rect 3689 6164 3695 6166
rect 3702 6164 3810 6180
rect 3817 6164 3823 6166
rect 3831 6164 3846 6180
rect 3912 6174 3931 6177
rect 3553 6152 3651 6154
rect 3678 6152 3846 6164
rect 3861 6154 3877 6168
rect 3912 6155 3934 6174
rect 3944 6168 3960 6169
rect 3943 6166 3960 6168
rect 3944 6161 3960 6166
rect 3934 6154 3940 6155
rect 3943 6154 3972 6161
rect 3861 6153 3972 6154
rect 3861 6152 3978 6153
rect 3537 6144 3588 6152
rect 3635 6144 3669 6152
rect 3537 6132 3562 6144
rect 3569 6132 3588 6144
rect 3642 6142 3669 6144
rect 3678 6142 3899 6152
rect 3934 6149 3940 6152
rect 3642 6138 3899 6142
rect 3537 6124 3588 6132
rect 3635 6124 3899 6138
rect 3943 6144 3978 6152
rect 3489 6076 3508 6110
rect 3553 6116 3582 6124
rect 3553 6110 3570 6116
rect 3553 6108 3587 6110
rect 3635 6108 3651 6124
rect 3652 6114 3860 6124
rect 3861 6114 3877 6124
rect 3925 6120 3940 6135
rect 3943 6132 3944 6144
rect 3951 6132 3978 6144
rect 3943 6124 3978 6132
rect 3943 6123 3972 6124
rect 3663 6110 3877 6114
rect 3678 6108 3877 6110
rect 3912 6110 3925 6120
rect 3943 6110 3960 6123
rect 3912 6108 3960 6110
rect 3554 6104 3587 6108
rect 3550 6102 3587 6104
rect 3550 6101 3617 6102
rect 3550 6096 3581 6101
rect 3587 6096 3617 6101
rect 3550 6092 3617 6096
rect 3523 6089 3617 6092
rect 3523 6082 3572 6089
rect 3523 6076 3553 6082
rect 3572 6077 3577 6082
rect 3489 6060 3569 6076
rect 3581 6068 3617 6089
rect 3678 6084 3867 6108
rect 3912 6107 3959 6108
rect 3925 6102 3959 6107
rect 3693 6081 3867 6084
rect 3686 6078 3867 6081
rect 3895 6101 3959 6102
rect 3489 6058 3508 6060
rect 3523 6058 3557 6060
rect 3489 6042 3569 6058
rect 3489 6036 3508 6042
rect 3205 6010 3308 6020
rect 3159 6008 3308 6010
rect 3329 6008 3364 6020
rect 2998 6006 3160 6008
rect 3010 5986 3029 6006
rect 3044 6004 3074 6006
rect 2893 5978 2934 5986
rect 3016 5982 3029 5986
rect 3081 5990 3160 6006
rect 3192 6006 3364 6008
rect 3192 5990 3271 6006
rect 3278 6004 3308 6006
rect 2856 5968 2885 5978
rect 2899 5968 2928 5978
rect 2943 5968 2973 5982
rect 3016 5968 3059 5982
rect 3081 5978 3271 5990
rect 3336 5986 3342 6006
rect 3066 5968 3096 5978
rect 3097 5968 3255 5978
rect 3259 5968 3289 5978
rect 3293 5968 3323 5982
rect 3351 5968 3364 6006
rect 3436 6020 3465 6036
rect 3479 6020 3508 6036
rect 3523 6026 3553 6042
rect 3581 6020 3587 6068
rect 3590 6062 3609 6068
rect 3624 6062 3654 6070
rect 3590 6054 3654 6062
rect 3590 6038 3670 6054
rect 3686 6047 3748 6078
rect 3764 6047 3826 6078
rect 3895 6076 3944 6101
rect 3959 6076 3989 6092
rect 3858 6062 3888 6070
rect 3895 6068 4005 6076
rect 3858 6054 3903 6062
rect 3590 6036 3609 6038
rect 3624 6036 3670 6038
rect 3590 6020 3670 6036
rect 3697 6034 3732 6047
rect 3773 6044 3810 6047
rect 3773 6042 3815 6044
rect 3702 6031 3732 6034
rect 3711 6027 3718 6031
rect 3718 6026 3719 6027
rect 3677 6020 3687 6026
rect 3436 6012 3471 6020
rect 3436 5986 3437 6012
rect 3444 5986 3471 6012
rect 3379 5968 3409 5982
rect 3436 5978 3471 5986
rect 3473 6012 3514 6020
rect 3473 5986 3488 6012
rect 3495 5986 3514 6012
rect 3578 6008 3609 6020
rect 3624 6008 3727 6020
rect 3739 6010 3765 6036
rect 3780 6031 3810 6042
rect 3842 6038 3904 6054
rect 3842 6036 3888 6038
rect 3842 6020 3904 6036
rect 3916 6020 3922 6068
rect 3925 6060 4005 6068
rect 3925 6058 3944 6060
rect 3959 6058 3993 6060
rect 3925 6042 4005 6058
rect 3925 6020 3944 6042
rect 3959 6026 3989 6042
rect 4017 6036 4023 6110
rect 4026 6036 4045 6180
rect 4060 6036 4066 6180
rect 4075 6110 4088 6180
rect 4140 6176 4162 6180
rect 4133 6154 4162 6168
rect 4215 6154 4231 6168
rect 4269 6164 4275 6166
rect 4282 6164 4390 6180
rect 4397 6164 4403 6166
rect 4411 6164 4426 6180
rect 4492 6174 4511 6177
rect 4133 6152 4231 6154
rect 4258 6152 4426 6164
rect 4441 6154 4457 6168
rect 4492 6155 4514 6174
rect 4524 6168 4540 6169
rect 4523 6166 4540 6168
rect 4524 6161 4540 6166
rect 4514 6154 4520 6155
rect 4523 6154 4552 6161
rect 4441 6153 4552 6154
rect 4441 6152 4558 6153
rect 4117 6144 4168 6152
rect 4215 6144 4249 6152
rect 4117 6132 4142 6144
rect 4149 6132 4168 6144
rect 4222 6142 4249 6144
rect 4258 6142 4479 6152
rect 4514 6149 4520 6152
rect 4222 6138 4479 6142
rect 4117 6124 4168 6132
rect 4215 6124 4479 6138
rect 4523 6144 4558 6152
rect 4069 6076 4088 6110
rect 4133 6116 4162 6124
rect 4133 6110 4150 6116
rect 4133 6108 4167 6110
rect 4215 6108 4231 6124
rect 4232 6114 4440 6124
rect 4441 6114 4457 6124
rect 4505 6120 4520 6135
rect 4523 6132 4524 6144
rect 4531 6132 4558 6144
rect 4523 6124 4558 6132
rect 4523 6123 4552 6124
rect 4243 6110 4457 6114
rect 4258 6108 4457 6110
rect 4492 6110 4505 6120
rect 4523 6110 4540 6123
rect 4492 6108 4540 6110
rect 4134 6104 4167 6108
rect 4130 6102 4167 6104
rect 4130 6101 4197 6102
rect 4130 6096 4161 6101
rect 4167 6096 4197 6101
rect 4130 6092 4197 6096
rect 4103 6089 4197 6092
rect 4103 6082 4152 6089
rect 4103 6076 4133 6082
rect 4152 6077 4157 6082
rect 4069 6060 4149 6076
rect 4161 6068 4197 6089
rect 4258 6084 4447 6108
rect 4492 6107 4539 6108
rect 4505 6102 4539 6107
rect 4273 6081 4447 6084
rect 4266 6078 4447 6081
rect 4475 6101 4539 6102
rect 4069 6058 4088 6060
rect 4103 6058 4137 6060
rect 4069 6042 4149 6058
rect 4069 6036 4088 6042
rect 3785 6010 3888 6020
rect 3739 6008 3888 6010
rect 3909 6008 3944 6020
rect 3578 6006 3740 6008
rect 3590 5986 3609 6006
rect 3624 6004 3654 6006
rect 3473 5978 3514 5986
rect 3596 5982 3609 5986
rect 3661 5990 3740 6006
rect 3772 6006 3944 6008
rect 3772 5990 3851 6006
rect 3858 6004 3888 6006
rect 3436 5968 3465 5978
rect 3479 5968 3508 5978
rect 3523 5968 3553 5982
rect 3596 5968 3639 5982
rect 3661 5978 3851 5990
rect 3916 5986 3922 6006
rect 3646 5968 3676 5978
rect 3677 5968 3835 5978
rect 3839 5968 3869 5978
rect 3873 5968 3903 5982
rect 3931 5968 3944 6006
rect 4016 6020 4045 6036
rect 4059 6020 4088 6036
rect 4103 6026 4133 6042
rect 4161 6020 4167 6068
rect 4170 6062 4189 6068
rect 4204 6062 4234 6070
rect 4170 6054 4234 6062
rect 4170 6038 4250 6054
rect 4266 6047 4328 6078
rect 4344 6047 4406 6078
rect 4475 6076 4524 6101
rect 4539 6076 4569 6092
rect 4438 6062 4468 6070
rect 4475 6068 4585 6076
rect 4438 6054 4483 6062
rect 4170 6036 4189 6038
rect 4204 6036 4250 6038
rect 4170 6020 4250 6036
rect 4277 6034 4312 6047
rect 4353 6044 4390 6047
rect 4353 6042 4395 6044
rect 4282 6031 4312 6034
rect 4291 6027 4298 6031
rect 4298 6026 4299 6027
rect 4257 6020 4267 6026
rect 4016 6012 4051 6020
rect 4016 5986 4017 6012
rect 4024 5986 4051 6012
rect 3959 5968 3989 5982
rect 4016 5978 4051 5986
rect 4053 6012 4094 6020
rect 4053 5986 4068 6012
rect 4075 5986 4094 6012
rect 4158 6008 4189 6020
rect 4204 6008 4307 6020
rect 4319 6010 4345 6036
rect 4360 6031 4390 6042
rect 4422 6038 4484 6054
rect 4422 6036 4468 6038
rect 4422 6020 4484 6036
rect 4496 6020 4502 6068
rect 4505 6060 4585 6068
rect 4505 6058 4524 6060
rect 4539 6058 4573 6060
rect 4505 6042 4585 6058
rect 4505 6020 4524 6042
rect 4539 6026 4569 6042
rect 4597 6036 4603 6110
rect 4606 6036 4625 6180
rect 4640 6036 4646 6180
rect 4655 6110 4668 6180
rect 4720 6176 4742 6180
rect 4713 6154 4742 6168
rect 4795 6154 4811 6168
rect 4849 6164 4855 6166
rect 4862 6164 4970 6180
rect 4977 6164 4983 6166
rect 4991 6164 5006 6180
rect 5072 6174 5091 6177
rect 4713 6152 4811 6154
rect 4838 6152 5006 6164
rect 5021 6154 5037 6168
rect 5072 6155 5094 6174
rect 5104 6168 5120 6169
rect 5103 6166 5120 6168
rect 5104 6161 5120 6166
rect 5094 6154 5100 6155
rect 5103 6154 5132 6161
rect 5021 6153 5132 6154
rect 5021 6152 5138 6153
rect 4697 6144 4748 6152
rect 4795 6144 4829 6152
rect 4697 6132 4722 6144
rect 4729 6132 4748 6144
rect 4802 6142 4829 6144
rect 4838 6142 5059 6152
rect 5094 6149 5100 6152
rect 4802 6138 5059 6142
rect 4697 6124 4748 6132
rect 4795 6124 5059 6138
rect 5103 6144 5138 6152
rect 4649 6076 4668 6110
rect 4713 6116 4742 6124
rect 4713 6110 4730 6116
rect 4713 6108 4747 6110
rect 4795 6108 4811 6124
rect 4812 6114 5020 6124
rect 5021 6114 5037 6124
rect 5085 6120 5100 6135
rect 5103 6132 5104 6144
rect 5111 6132 5138 6144
rect 5103 6124 5138 6132
rect 5103 6123 5132 6124
rect 4823 6110 5037 6114
rect 4838 6108 5037 6110
rect 5072 6110 5085 6120
rect 5103 6110 5120 6123
rect 5072 6108 5120 6110
rect 4714 6104 4747 6108
rect 4710 6102 4747 6104
rect 4710 6101 4777 6102
rect 4710 6096 4741 6101
rect 4747 6096 4777 6101
rect 4710 6092 4777 6096
rect 4683 6089 4777 6092
rect 4683 6082 4732 6089
rect 4683 6076 4713 6082
rect 4732 6077 4737 6082
rect 4649 6060 4729 6076
rect 4741 6068 4777 6089
rect 4838 6084 5027 6108
rect 5072 6107 5119 6108
rect 5085 6102 5119 6107
rect 4853 6081 5027 6084
rect 4846 6078 5027 6081
rect 5055 6101 5119 6102
rect 4649 6058 4668 6060
rect 4683 6058 4717 6060
rect 4649 6042 4729 6058
rect 4649 6036 4668 6042
rect 4365 6010 4468 6020
rect 4319 6008 4468 6010
rect 4489 6008 4524 6020
rect 4158 6006 4320 6008
rect 4170 5986 4189 6006
rect 4204 6004 4234 6006
rect 4053 5978 4094 5986
rect 4176 5982 4189 5986
rect 4241 5990 4320 6006
rect 4352 6006 4524 6008
rect 4352 5990 4431 6006
rect 4438 6004 4468 6006
rect 4016 5968 4045 5978
rect 4059 5968 4088 5978
rect 4103 5968 4133 5982
rect 4176 5968 4219 5982
rect 4241 5978 4431 5990
rect 4496 5986 4502 6006
rect 4226 5968 4256 5978
rect 4257 5968 4415 5978
rect 4419 5968 4449 5978
rect 4453 5968 4483 5982
rect 4511 5968 4524 6006
rect 4596 6020 4625 6036
rect 4639 6020 4668 6036
rect 4683 6026 4713 6042
rect 4741 6020 4747 6068
rect 4750 6062 4769 6068
rect 4784 6062 4814 6070
rect 4750 6054 4814 6062
rect 4750 6038 4830 6054
rect 4846 6047 4908 6078
rect 4924 6047 4986 6078
rect 5055 6076 5104 6101
rect 5119 6076 5149 6092
rect 5018 6062 5048 6070
rect 5055 6068 5165 6076
rect 5018 6054 5063 6062
rect 4750 6036 4769 6038
rect 4784 6036 4830 6038
rect 4750 6020 4830 6036
rect 4857 6034 4892 6047
rect 4933 6044 4970 6047
rect 4933 6042 4975 6044
rect 4862 6031 4892 6034
rect 4871 6027 4878 6031
rect 4878 6026 4879 6027
rect 4837 6020 4847 6026
rect 4596 6012 4631 6020
rect 4596 5986 4597 6012
rect 4604 5986 4631 6012
rect 4539 5968 4569 5982
rect 4596 5978 4631 5986
rect 4633 6012 4674 6020
rect 4633 5986 4648 6012
rect 4655 5986 4674 6012
rect 4738 6008 4769 6020
rect 4784 6008 4887 6020
rect 4899 6010 4925 6036
rect 4940 6031 4970 6042
rect 5002 6038 5064 6054
rect 5002 6036 5048 6038
rect 5002 6020 5064 6036
rect 5076 6020 5082 6068
rect 5085 6060 5165 6068
rect 5085 6058 5104 6060
rect 5119 6058 5153 6060
rect 5085 6042 5165 6058
rect 5085 6020 5104 6042
rect 5119 6026 5149 6042
rect 5177 6036 5183 6110
rect 5186 6036 5205 6180
rect 5220 6036 5226 6180
rect 5235 6110 5248 6180
rect 5300 6176 5322 6180
rect 5293 6154 5322 6168
rect 5375 6154 5391 6168
rect 5429 6164 5435 6166
rect 5442 6164 5550 6180
rect 5557 6164 5563 6166
rect 5571 6164 5586 6180
rect 5652 6174 5671 6177
rect 5293 6152 5391 6154
rect 5418 6152 5586 6164
rect 5601 6154 5617 6168
rect 5652 6155 5674 6174
rect 5684 6168 5700 6169
rect 5683 6166 5700 6168
rect 5684 6161 5700 6166
rect 5674 6154 5680 6155
rect 5683 6154 5712 6161
rect 5601 6153 5712 6154
rect 5601 6152 5718 6153
rect 5277 6144 5328 6152
rect 5375 6144 5409 6152
rect 5277 6132 5302 6144
rect 5309 6132 5328 6144
rect 5382 6142 5409 6144
rect 5418 6142 5639 6152
rect 5674 6149 5680 6152
rect 5382 6138 5639 6142
rect 5277 6124 5328 6132
rect 5375 6124 5639 6138
rect 5683 6144 5718 6152
rect 5229 6076 5248 6110
rect 5293 6116 5322 6124
rect 5293 6110 5310 6116
rect 5293 6108 5327 6110
rect 5375 6108 5391 6124
rect 5392 6114 5600 6124
rect 5601 6114 5617 6124
rect 5665 6120 5680 6135
rect 5683 6132 5684 6144
rect 5691 6132 5718 6144
rect 5683 6124 5718 6132
rect 5683 6123 5712 6124
rect 5403 6110 5617 6114
rect 5418 6108 5617 6110
rect 5652 6110 5665 6120
rect 5683 6110 5700 6123
rect 5652 6108 5700 6110
rect 5294 6104 5327 6108
rect 5290 6102 5327 6104
rect 5290 6101 5357 6102
rect 5290 6096 5321 6101
rect 5327 6096 5357 6101
rect 5290 6092 5357 6096
rect 5263 6089 5357 6092
rect 5263 6082 5312 6089
rect 5263 6076 5293 6082
rect 5312 6077 5317 6082
rect 5229 6060 5309 6076
rect 5321 6068 5357 6089
rect 5418 6084 5607 6108
rect 5652 6107 5699 6108
rect 5665 6102 5699 6107
rect 5433 6081 5607 6084
rect 5426 6078 5607 6081
rect 5635 6101 5699 6102
rect 5229 6058 5248 6060
rect 5263 6058 5297 6060
rect 5229 6042 5309 6058
rect 5229 6036 5248 6042
rect 4945 6010 5048 6020
rect 4899 6008 5048 6010
rect 5069 6008 5104 6020
rect 4738 6006 4900 6008
rect 4750 5986 4769 6006
rect 4784 6004 4814 6006
rect 4633 5978 4674 5986
rect 4756 5982 4769 5986
rect 4821 5990 4900 6006
rect 4932 6006 5104 6008
rect 4932 5990 5011 6006
rect 5018 6004 5048 6006
rect 4596 5968 4625 5978
rect 4639 5968 4668 5978
rect 4683 5968 4713 5982
rect 4756 5968 4799 5982
rect 4821 5978 5011 5990
rect 5076 5986 5082 6006
rect 4806 5968 4836 5978
rect 4837 5968 4995 5978
rect 4999 5968 5029 5978
rect 5033 5968 5063 5982
rect 5091 5968 5104 6006
rect 5176 6020 5205 6036
rect 5219 6020 5248 6036
rect 5263 6026 5293 6042
rect 5321 6020 5327 6068
rect 5330 6062 5349 6068
rect 5364 6062 5394 6070
rect 5330 6054 5394 6062
rect 5330 6038 5410 6054
rect 5426 6047 5488 6078
rect 5504 6047 5566 6078
rect 5635 6076 5684 6101
rect 5699 6076 5729 6092
rect 5598 6062 5628 6070
rect 5635 6068 5745 6076
rect 5598 6054 5643 6062
rect 5330 6036 5349 6038
rect 5364 6036 5410 6038
rect 5330 6020 5410 6036
rect 5437 6034 5472 6047
rect 5513 6044 5550 6047
rect 5513 6042 5555 6044
rect 5442 6031 5472 6034
rect 5451 6027 5458 6031
rect 5458 6026 5459 6027
rect 5417 6020 5427 6026
rect 5176 6012 5211 6020
rect 5176 5986 5177 6012
rect 5184 5986 5211 6012
rect 5119 5968 5149 5982
rect 5176 5978 5211 5986
rect 5213 6012 5254 6020
rect 5213 5986 5228 6012
rect 5235 5986 5254 6012
rect 5318 6008 5349 6020
rect 5364 6008 5467 6020
rect 5479 6010 5505 6036
rect 5520 6031 5550 6042
rect 5582 6038 5644 6054
rect 5582 6036 5628 6038
rect 5582 6020 5644 6036
rect 5656 6020 5662 6068
rect 5665 6060 5745 6068
rect 5665 6058 5684 6060
rect 5699 6058 5733 6060
rect 5665 6042 5745 6058
rect 5665 6020 5684 6042
rect 5699 6026 5729 6042
rect 5757 6036 5763 6110
rect 5766 6036 5785 6180
rect 5800 6036 5806 6180
rect 5815 6110 5828 6180
rect 5880 6176 5902 6180
rect 5873 6154 5902 6168
rect 5955 6154 5971 6168
rect 6009 6164 6015 6166
rect 6022 6164 6130 6180
rect 6137 6164 6143 6166
rect 6151 6164 6166 6180
rect 6232 6174 6251 6177
rect 5873 6152 5971 6154
rect 5998 6152 6166 6164
rect 6181 6154 6197 6168
rect 6232 6155 6254 6174
rect 6264 6168 6280 6169
rect 6263 6166 6280 6168
rect 6264 6161 6280 6166
rect 6254 6154 6260 6155
rect 6263 6154 6292 6161
rect 6181 6153 6292 6154
rect 6181 6152 6298 6153
rect 5857 6144 5908 6152
rect 5955 6144 5989 6152
rect 5857 6132 5882 6144
rect 5889 6132 5908 6144
rect 5962 6142 5989 6144
rect 5998 6142 6219 6152
rect 6254 6149 6260 6152
rect 5962 6138 6219 6142
rect 5857 6124 5908 6132
rect 5955 6124 6219 6138
rect 6263 6144 6298 6152
rect 5809 6076 5828 6110
rect 5873 6116 5902 6124
rect 5873 6110 5890 6116
rect 5873 6108 5907 6110
rect 5955 6108 5971 6124
rect 5972 6114 6180 6124
rect 6181 6114 6197 6124
rect 6245 6120 6260 6135
rect 6263 6132 6264 6144
rect 6271 6132 6298 6144
rect 6263 6124 6298 6132
rect 6263 6123 6292 6124
rect 5983 6110 6197 6114
rect 5998 6108 6197 6110
rect 6232 6110 6245 6120
rect 6263 6110 6280 6123
rect 6232 6108 6280 6110
rect 5874 6104 5907 6108
rect 5870 6102 5907 6104
rect 5870 6101 5937 6102
rect 5870 6096 5901 6101
rect 5907 6096 5937 6101
rect 5870 6092 5937 6096
rect 5843 6089 5937 6092
rect 5843 6082 5892 6089
rect 5843 6076 5873 6082
rect 5892 6077 5897 6082
rect 5809 6060 5889 6076
rect 5901 6068 5937 6089
rect 5998 6084 6187 6108
rect 6232 6107 6279 6108
rect 6245 6102 6279 6107
rect 6013 6081 6187 6084
rect 6006 6078 6187 6081
rect 6215 6101 6279 6102
rect 5809 6058 5828 6060
rect 5843 6058 5877 6060
rect 5809 6042 5889 6058
rect 5809 6036 5828 6042
rect 5525 6010 5628 6020
rect 5479 6008 5628 6010
rect 5649 6008 5684 6020
rect 5318 6006 5480 6008
rect 5330 5986 5349 6006
rect 5364 6004 5394 6006
rect 5213 5978 5254 5986
rect 5336 5982 5349 5986
rect 5401 5990 5480 6006
rect 5512 6006 5684 6008
rect 5512 5990 5591 6006
rect 5598 6004 5628 6006
rect 5176 5968 5205 5978
rect 5219 5968 5248 5978
rect 5263 5968 5293 5982
rect 5336 5968 5379 5982
rect 5401 5978 5591 5990
rect 5656 5986 5662 6006
rect 5386 5968 5416 5978
rect 5417 5968 5575 5978
rect 5579 5968 5609 5978
rect 5613 5968 5643 5982
rect 5671 5968 5684 6006
rect 5756 6020 5785 6036
rect 5799 6020 5828 6036
rect 5843 6026 5873 6042
rect 5901 6020 5907 6068
rect 5910 6062 5929 6068
rect 5944 6062 5974 6070
rect 5910 6054 5974 6062
rect 5910 6038 5990 6054
rect 6006 6047 6068 6078
rect 6084 6047 6146 6078
rect 6215 6076 6264 6101
rect 6279 6076 6309 6092
rect 6178 6062 6208 6070
rect 6215 6068 6325 6076
rect 6178 6054 6223 6062
rect 5910 6036 5929 6038
rect 5944 6036 5990 6038
rect 5910 6020 5990 6036
rect 6017 6034 6052 6047
rect 6093 6044 6130 6047
rect 6093 6042 6135 6044
rect 6022 6031 6052 6034
rect 6031 6027 6038 6031
rect 6038 6026 6039 6027
rect 5997 6020 6007 6026
rect 5756 6012 5791 6020
rect 5756 5986 5757 6012
rect 5764 5986 5791 6012
rect 5699 5968 5729 5982
rect 5756 5978 5791 5986
rect 5793 6012 5834 6020
rect 5793 5986 5808 6012
rect 5815 5986 5834 6012
rect 5898 6008 5929 6020
rect 5944 6008 6047 6020
rect 6059 6010 6085 6036
rect 6100 6031 6130 6042
rect 6162 6038 6224 6054
rect 6162 6036 6208 6038
rect 6162 6020 6224 6036
rect 6236 6020 6242 6068
rect 6245 6060 6325 6068
rect 6245 6058 6264 6060
rect 6279 6058 6313 6060
rect 6245 6042 6325 6058
rect 6245 6020 6264 6042
rect 6279 6026 6309 6042
rect 6337 6036 6343 6110
rect 6346 6036 6365 6180
rect 6380 6036 6386 6180
rect 6395 6110 6408 6180
rect 6460 6176 6482 6180
rect 6453 6154 6482 6168
rect 6535 6154 6551 6168
rect 6589 6164 6595 6166
rect 6602 6164 6710 6180
rect 6717 6164 6723 6166
rect 6731 6164 6746 6180
rect 6812 6174 6831 6177
rect 6453 6152 6551 6154
rect 6578 6152 6746 6164
rect 6761 6154 6777 6168
rect 6812 6155 6834 6174
rect 6844 6168 6860 6169
rect 6843 6166 6860 6168
rect 6844 6161 6860 6166
rect 6834 6154 6840 6155
rect 6843 6154 6872 6161
rect 6761 6153 6872 6154
rect 6761 6152 6878 6153
rect 6437 6144 6488 6152
rect 6535 6144 6569 6152
rect 6437 6132 6462 6144
rect 6469 6132 6488 6144
rect 6542 6142 6569 6144
rect 6578 6142 6799 6152
rect 6834 6149 6840 6152
rect 6542 6138 6799 6142
rect 6437 6124 6488 6132
rect 6535 6124 6799 6138
rect 6843 6144 6878 6152
rect 6389 6076 6408 6110
rect 6453 6116 6482 6124
rect 6453 6110 6470 6116
rect 6453 6108 6487 6110
rect 6535 6108 6551 6124
rect 6552 6114 6760 6124
rect 6761 6114 6777 6124
rect 6825 6120 6840 6135
rect 6843 6132 6844 6144
rect 6851 6132 6878 6144
rect 6843 6124 6878 6132
rect 6843 6123 6872 6124
rect 6563 6110 6777 6114
rect 6578 6108 6777 6110
rect 6812 6110 6825 6120
rect 6843 6110 6860 6123
rect 6812 6108 6860 6110
rect 6454 6104 6487 6108
rect 6450 6102 6487 6104
rect 6450 6101 6517 6102
rect 6450 6096 6481 6101
rect 6487 6096 6517 6101
rect 6450 6092 6517 6096
rect 6423 6089 6517 6092
rect 6423 6082 6472 6089
rect 6423 6076 6453 6082
rect 6472 6077 6477 6082
rect 6389 6060 6469 6076
rect 6481 6068 6517 6089
rect 6578 6084 6767 6108
rect 6812 6107 6859 6108
rect 6825 6102 6859 6107
rect 6593 6081 6767 6084
rect 6586 6078 6767 6081
rect 6795 6101 6859 6102
rect 6389 6058 6408 6060
rect 6423 6058 6457 6060
rect 6389 6042 6469 6058
rect 6389 6036 6408 6042
rect 6105 6010 6208 6020
rect 6059 6008 6208 6010
rect 6229 6008 6264 6020
rect 5898 6006 6060 6008
rect 5910 5986 5929 6006
rect 5944 6004 5974 6006
rect 5793 5978 5834 5986
rect 5916 5982 5929 5986
rect 5981 5990 6060 6006
rect 6092 6006 6264 6008
rect 6092 5990 6171 6006
rect 6178 6004 6208 6006
rect 5756 5968 5785 5978
rect 5799 5968 5828 5978
rect 5843 5968 5873 5982
rect 5916 5968 5959 5982
rect 5981 5978 6171 5990
rect 6236 5986 6242 6006
rect 5966 5968 5996 5978
rect 5997 5968 6155 5978
rect 6159 5968 6189 5978
rect 6193 5968 6223 5982
rect 6251 5968 6264 6006
rect 6336 6020 6365 6036
rect 6379 6020 6408 6036
rect 6423 6026 6453 6042
rect 6481 6020 6487 6068
rect 6490 6062 6509 6068
rect 6524 6062 6554 6070
rect 6490 6054 6554 6062
rect 6490 6038 6570 6054
rect 6586 6047 6648 6078
rect 6664 6047 6726 6078
rect 6795 6076 6844 6101
rect 6859 6076 6889 6092
rect 6758 6062 6788 6070
rect 6795 6068 6905 6076
rect 6758 6054 6803 6062
rect 6490 6036 6509 6038
rect 6524 6036 6570 6038
rect 6490 6020 6570 6036
rect 6597 6034 6632 6047
rect 6673 6044 6710 6047
rect 6673 6042 6715 6044
rect 6602 6031 6632 6034
rect 6611 6027 6618 6031
rect 6618 6026 6619 6027
rect 6577 6020 6587 6026
rect 6336 6012 6371 6020
rect 6336 5986 6337 6012
rect 6344 5986 6371 6012
rect 6279 5968 6309 5982
rect 6336 5978 6371 5986
rect 6373 6012 6414 6020
rect 6373 5986 6388 6012
rect 6395 5986 6414 6012
rect 6478 6008 6509 6020
rect 6524 6008 6627 6020
rect 6639 6010 6665 6036
rect 6680 6031 6710 6042
rect 6742 6038 6804 6054
rect 6742 6036 6788 6038
rect 6742 6020 6804 6036
rect 6816 6020 6822 6068
rect 6825 6060 6905 6068
rect 6825 6058 6844 6060
rect 6859 6058 6893 6060
rect 6825 6042 6905 6058
rect 6825 6020 6844 6042
rect 6859 6026 6889 6042
rect 6917 6036 6923 6110
rect 6926 6036 6945 6180
rect 6960 6036 6966 6180
rect 6975 6110 6988 6180
rect 7040 6176 7062 6180
rect 7033 6154 7062 6168
rect 7115 6154 7131 6168
rect 7169 6164 7175 6166
rect 7182 6164 7290 6180
rect 7297 6164 7303 6166
rect 7311 6164 7326 6180
rect 7392 6174 7411 6177
rect 7033 6152 7131 6154
rect 7158 6152 7326 6164
rect 7341 6154 7357 6168
rect 7392 6155 7414 6174
rect 7424 6168 7440 6169
rect 7423 6166 7440 6168
rect 7424 6161 7440 6166
rect 7414 6154 7420 6155
rect 7423 6154 7452 6161
rect 7341 6153 7452 6154
rect 7341 6152 7458 6153
rect 7017 6144 7068 6152
rect 7115 6144 7149 6152
rect 7017 6132 7042 6144
rect 7049 6132 7068 6144
rect 7122 6142 7149 6144
rect 7158 6142 7379 6152
rect 7414 6149 7420 6152
rect 7122 6138 7379 6142
rect 7017 6124 7068 6132
rect 7115 6124 7379 6138
rect 7423 6144 7458 6152
rect 6969 6076 6988 6110
rect 7033 6116 7062 6124
rect 7033 6110 7050 6116
rect 7033 6108 7067 6110
rect 7115 6108 7131 6124
rect 7132 6114 7340 6124
rect 7341 6114 7357 6124
rect 7405 6120 7420 6135
rect 7423 6132 7424 6144
rect 7431 6132 7458 6144
rect 7423 6124 7458 6132
rect 7423 6123 7452 6124
rect 7143 6110 7357 6114
rect 7158 6108 7357 6110
rect 7392 6110 7405 6120
rect 7423 6110 7440 6123
rect 7392 6108 7440 6110
rect 7034 6104 7067 6108
rect 7030 6102 7067 6104
rect 7030 6101 7097 6102
rect 7030 6096 7061 6101
rect 7067 6096 7097 6101
rect 7030 6092 7097 6096
rect 7003 6089 7097 6092
rect 7003 6082 7052 6089
rect 7003 6076 7033 6082
rect 7052 6077 7057 6082
rect 6969 6060 7049 6076
rect 7061 6068 7097 6089
rect 7158 6084 7347 6108
rect 7392 6107 7439 6108
rect 7405 6102 7439 6107
rect 7173 6081 7347 6084
rect 7166 6078 7347 6081
rect 7375 6101 7439 6102
rect 6969 6058 6988 6060
rect 7003 6058 7037 6060
rect 6969 6042 7049 6058
rect 6969 6036 6988 6042
rect 6685 6010 6788 6020
rect 6639 6008 6788 6010
rect 6809 6008 6844 6020
rect 6478 6006 6640 6008
rect 6490 5986 6509 6006
rect 6524 6004 6554 6006
rect 6373 5978 6414 5986
rect 6496 5982 6509 5986
rect 6561 5990 6640 6006
rect 6672 6006 6844 6008
rect 6672 5990 6751 6006
rect 6758 6004 6788 6006
rect 6336 5968 6365 5978
rect 6379 5968 6408 5978
rect 6423 5968 6453 5982
rect 6496 5968 6539 5982
rect 6561 5978 6751 5990
rect 6816 5986 6822 6006
rect 6546 5968 6576 5978
rect 6577 5968 6735 5978
rect 6739 5968 6769 5978
rect 6773 5968 6803 5982
rect 6831 5968 6844 6006
rect 6916 6020 6945 6036
rect 6959 6020 6988 6036
rect 7003 6026 7033 6042
rect 7061 6020 7067 6068
rect 7070 6062 7089 6068
rect 7104 6062 7134 6070
rect 7070 6054 7134 6062
rect 7070 6038 7150 6054
rect 7166 6047 7228 6078
rect 7244 6047 7306 6078
rect 7375 6076 7424 6101
rect 7439 6076 7469 6092
rect 7338 6062 7368 6070
rect 7375 6068 7485 6076
rect 7338 6054 7383 6062
rect 7070 6036 7089 6038
rect 7104 6036 7150 6038
rect 7070 6020 7150 6036
rect 7177 6034 7212 6047
rect 7253 6044 7290 6047
rect 7253 6042 7295 6044
rect 7182 6031 7212 6034
rect 7191 6027 7198 6031
rect 7198 6026 7199 6027
rect 7157 6020 7167 6026
rect 6916 6012 6951 6020
rect 6916 5986 6917 6012
rect 6924 5986 6951 6012
rect 6859 5968 6889 5982
rect 6916 5978 6951 5986
rect 6953 6012 6994 6020
rect 6953 5986 6968 6012
rect 6975 5986 6994 6012
rect 7058 6008 7089 6020
rect 7104 6008 7207 6020
rect 7219 6010 7245 6036
rect 7260 6031 7290 6042
rect 7322 6038 7384 6054
rect 7322 6036 7368 6038
rect 7322 6020 7384 6036
rect 7396 6020 7402 6068
rect 7405 6060 7485 6068
rect 7405 6058 7424 6060
rect 7439 6058 7473 6060
rect 7405 6042 7485 6058
rect 7405 6020 7424 6042
rect 7439 6026 7469 6042
rect 7497 6036 7503 6110
rect 7506 6036 7525 6180
rect 7540 6036 7546 6180
rect 7555 6110 7568 6180
rect 7620 6176 7642 6180
rect 7613 6154 7642 6168
rect 7695 6154 7711 6168
rect 7749 6164 7755 6166
rect 7762 6164 7870 6180
rect 7877 6164 7883 6166
rect 7891 6164 7906 6180
rect 7972 6174 7991 6177
rect 7613 6152 7711 6154
rect 7738 6152 7906 6164
rect 7921 6154 7937 6168
rect 7972 6155 7994 6174
rect 8004 6168 8020 6169
rect 8003 6166 8020 6168
rect 8004 6161 8020 6166
rect 7994 6154 8000 6155
rect 8003 6154 8032 6161
rect 7921 6153 8032 6154
rect 7921 6152 8038 6153
rect 7597 6144 7648 6152
rect 7695 6144 7729 6152
rect 7597 6132 7622 6144
rect 7629 6132 7648 6144
rect 7702 6142 7729 6144
rect 7738 6142 7959 6152
rect 7994 6149 8000 6152
rect 7702 6138 7959 6142
rect 7597 6124 7648 6132
rect 7695 6124 7959 6138
rect 8003 6144 8038 6152
rect 7549 6076 7568 6110
rect 7613 6116 7642 6124
rect 7613 6110 7630 6116
rect 7613 6108 7647 6110
rect 7695 6108 7711 6124
rect 7712 6114 7920 6124
rect 7921 6114 7937 6124
rect 7985 6120 8000 6135
rect 8003 6132 8004 6144
rect 8011 6132 8038 6144
rect 8003 6124 8038 6132
rect 8003 6123 8032 6124
rect 7723 6110 7937 6114
rect 7738 6108 7937 6110
rect 7972 6110 7985 6120
rect 8003 6110 8020 6123
rect 7972 6108 8020 6110
rect 7614 6104 7647 6108
rect 7610 6102 7647 6104
rect 7610 6101 7677 6102
rect 7610 6096 7641 6101
rect 7647 6096 7677 6101
rect 7610 6092 7677 6096
rect 7583 6089 7677 6092
rect 7583 6082 7632 6089
rect 7583 6076 7613 6082
rect 7632 6077 7637 6082
rect 7549 6060 7629 6076
rect 7641 6068 7677 6089
rect 7738 6084 7927 6108
rect 7972 6107 8019 6108
rect 7985 6102 8019 6107
rect 7753 6081 7927 6084
rect 7746 6078 7927 6081
rect 7955 6101 8019 6102
rect 7549 6058 7568 6060
rect 7583 6058 7617 6060
rect 7549 6042 7629 6058
rect 7549 6036 7568 6042
rect 7265 6010 7368 6020
rect 7219 6008 7368 6010
rect 7389 6008 7424 6020
rect 7058 6006 7220 6008
rect 7070 5986 7089 6006
rect 7104 6004 7134 6006
rect 6953 5978 6994 5986
rect 7076 5982 7089 5986
rect 7141 5990 7220 6006
rect 7252 6006 7424 6008
rect 7252 5990 7331 6006
rect 7338 6004 7368 6006
rect 6916 5968 6945 5978
rect 6959 5968 6988 5978
rect 7003 5968 7033 5982
rect 7076 5968 7119 5982
rect 7141 5978 7331 5990
rect 7396 5986 7402 6006
rect 7126 5968 7156 5978
rect 7157 5968 7315 5978
rect 7319 5968 7349 5978
rect 7353 5968 7383 5982
rect 7411 5968 7424 6006
rect 7496 6020 7525 6036
rect 7539 6020 7568 6036
rect 7583 6026 7613 6042
rect 7641 6020 7647 6068
rect 7650 6062 7669 6068
rect 7684 6062 7714 6070
rect 7650 6054 7714 6062
rect 7650 6038 7730 6054
rect 7746 6047 7808 6078
rect 7824 6047 7886 6078
rect 7955 6076 8004 6101
rect 8019 6076 8049 6092
rect 7918 6062 7948 6070
rect 7955 6068 8065 6076
rect 7918 6054 7963 6062
rect 7650 6036 7669 6038
rect 7684 6036 7730 6038
rect 7650 6020 7730 6036
rect 7757 6034 7792 6047
rect 7833 6044 7870 6047
rect 7833 6042 7875 6044
rect 7762 6031 7792 6034
rect 7771 6027 7778 6031
rect 7778 6026 7779 6027
rect 7737 6020 7747 6026
rect 7496 6012 7531 6020
rect 7496 5986 7497 6012
rect 7504 5986 7531 6012
rect 7439 5968 7469 5982
rect 7496 5978 7531 5986
rect 7533 6012 7574 6020
rect 7533 5986 7548 6012
rect 7555 5986 7574 6012
rect 7638 6008 7669 6020
rect 7684 6008 7787 6020
rect 7799 6010 7825 6036
rect 7840 6031 7870 6042
rect 7902 6038 7964 6054
rect 7902 6036 7948 6038
rect 7902 6020 7964 6036
rect 7976 6020 7982 6068
rect 7985 6060 8065 6068
rect 7985 6058 8004 6060
rect 8019 6058 8053 6060
rect 7985 6042 8065 6058
rect 7985 6020 8004 6042
rect 8019 6026 8049 6042
rect 8077 6036 8083 6110
rect 8086 6036 8105 6180
rect 8120 6036 8126 6180
rect 8135 6110 8148 6180
rect 8200 6176 8222 6180
rect 8193 6154 8222 6168
rect 8275 6154 8291 6168
rect 8329 6164 8335 6166
rect 8342 6164 8450 6180
rect 8457 6164 8463 6166
rect 8471 6164 8486 6180
rect 8552 6174 8571 6177
rect 8193 6152 8291 6154
rect 8318 6152 8486 6164
rect 8501 6154 8517 6168
rect 8552 6155 8574 6174
rect 8584 6168 8600 6169
rect 8583 6166 8600 6168
rect 8584 6161 8600 6166
rect 8574 6154 8580 6155
rect 8583 6154 8612 6161
rect 8501 6153 8612 6154
rect 8501 6152 8618 6153
rect 8177 6144 8228 6152
rect 8275 6144 8309 6152
rect 8177 6132 8202 6144
rect 8209 6132 8228 6144
rect 8282 6142 8309 6144
rect 8318 6142 8539 6152
rect 8574 6149 8580 6152
rect 8282 6138 8539 6142
rect 8177 6124 8228 6132
rect 8275 6124 8539 6138
rect 8583 6144 8618 6152
rect 8129 6076 8148 6110
rect 8193 6116 8222 6124
rect 8193 6110 8210 6116
rect 8193 6108 8227 6110
rect 8275 6108 8291 6124
rect 8292 6114 8500 6124
rect 8501 6114 8517 6124
rect 8565 6120 8580 6135
rect 8583 6132 8584 6144
rect 8591 6132 8618 6144
rect 8583 6124 8618 6132
rect 8583 6123 8612 6124
rect 8303 6110 8517 6114
rect 8318 6108 8517 6110
rect 8552 6110 8565 6120
rect 8583 6110 8600 6123
rect 8552 6108 8600 6110
rect 8194 6104 8227 6108
rect 8190 6102 8227 6104
rect 8190 6101 8257 6102
rect 8190 6096 8221 6101
rect 8227 6096 8257 6101
rect 8190 6092 8257 6096
rect 8163 6089 8257 6092
rect 8163 6082 8212 6089
rect 8163 6076 8193 6082
rect 8212 6077 8217 6082
rect 8129 6060 8209 6076
rect 8221 6068 8257 6089
rect 8318 6084 8507 6108
rect 8552 6107 8599 6108
rect 8565 6102 8599 6107
rect 8333 6081 8507 6084
rect 8326 6078 8507 6081
rect 8535 6101 8599 6102
rect 8129 6058 8148 6060
rect 8163 6058 8197 6060
rect 8129 6042 8209 6058
rect 8129 6036 8148 6042
rect 7845 6010 7948 6020
rect 7799 6008 7948 6010
rect 7969 6008 8004 6020
rect 7638 6006 7800 6008
rect 7650 5986 7669 6006
rect 7684 6004 7714 6006
rect 7533 5978 7574 5986
rect 7656 5982 7669 5986
rect 7721 5990 7800 6006
rect 7832 6006 8004 6008
rect 7832 5990 7911 6006
rect 7918 6004 7948 6006
rect 7496 5968 7525 5978
rect 7539 5968 7568 5978
rect 7583 5968 7613 5982
rect 7656 5968 7699 5982
rect 7721 5978 7911 5990
rect 7976 5986 7982 6006
rect 7706 5968 7736 5978
rect 7737 5968 7895 5978
rect 7899 5968 7929 5978
rect 7933 5968 7963 5982
rect 7991 5968 8004 6006
rect 8076 6020 8105 6036
rect 8119 6020 8148 6036
rect 8163 6026 8193 6042
rect 8221 6020 8227 6068
rect 8230 6062 8249 6068
rect 8264 6062 8294 6070
rect 8230 6054 8294 6062
rect 8230 6038 8310 6054
rect 8326 6047 8388 6078
rect 8404 6047 8466 6078
rect 8535 6076 8584 6101
rect 8599 6076 8629 6092
rect 8498 6062 8528 6070
rect 8535 6068 8645 6076
rect 8498 6054 8543 6062
rect 8230 6036 8249 6038
rect 8264 6036 8310 6038
rect 8230 6020 8310 6036
rect 8337 6034 8372 6047
rect 8413 6044 8450 6047
rect 8413 6042 8455 6044
rect 8342 6031 8372 6034
rect 8351 6027 8358 6031
rect 8358 6026 8359 6027
rect 8317 6020 8327 6026
rect 8076 6012 8111 6020
rect 8076 5986 8077 6012
rect 8084 5986 8111 6012
rect 8019 5968 8049 5982
rect 8076 5978 8111 5986
rect 8113 6012 8154 6020
rect 8113 5986 8128 6012
rect 8135 5986 8154 6012
rect 8218 6008 8249 6020
rect 8264 6008 8367 6020
rect 8379 6010 8405 6036
rect 8420 6031 8450 6042
rect 8482 6038 8544 6054
rect 8482 6036 8528 6038
rect 8482 6020 8544 6036
rect 8556 6020 8562 6068
rect 8565 6060 8645 6068
rect 8565 6058 8584 6060
rect 8599 6058 8633 6060
rect 8565 6042 8645 6058
rect 8565 6020 8584 6042
rect 8599 6026 8629 6042
rect 8657 6036 8663 6110
rect 8666 6036 8685 6180
rect 8700 6036 8706 6180
rect 8715 6110 8728 6180
rect 8780 6176 8802 6180
rect 8773 6154 8802 6168
rect 8855 6154 8871 6168
rect 8909 6164 8915 6166
rect 8922 6164 9030 6180
rect 9037 6164 9043 6166
rect 9051 6164 9066 6180
rect 9132 6174 9151 6177
rect 8773 6152 8871 6154
rect 8898 6152 9066 6164
rect 9081 6154 9097 6168
rect 9132 6155 9154 6174
rect 9164 6168 9180 6169
rect 9163 6166 9180 6168
rect 9164 6161 9180 6166
rect 9154 6154 9160 6155
rect 9163 6154 9192 6161
rect 9081 6153 9192 6154
rect 9081 6152 9198 6153
rect 8757 6144 8808 6152
rect 8855 6144 8889 6152
rect 8757 6132 8782 6144
rect 8789 6132 8808 6144
rect 8862 6142 8889 6144
rect 8898 6142 9119 6152
rect 9154 6149 9160 6152
rect 8862 6138 9119 6142
rect 8757 6124 8808 6132
rect 8855 6124 9119 6138
rect 9163 6144 9198 6152
rect 8709 6076 8728 6110
rect 8773 6116 8802 6124
rect 8773 6110 8790 6116
rect 8773 6108 8807 6110
rect 8855 6108 8871 6124
rect 8872 6114 9080 6124
rect 9081 6114 9097 6124
rect 9145 6120 9160 6135
rect 9163 6132 9164 6144
rect 9171 6132 9198 6144
rect 9163 6124 9198 6132
rect 9163 6123 9192 6124
rect 8883 6110 9097 6114
rect 8898 6108 9097 6110
rect 9132 6110 9145 6120
rect 9163 6110 9180 6123
rect 9132 6108 9180 6110
rect 8774 6104 8807 6108
rect 8770 6102 8807 6104
rect 8770 6101 8837 6102
rect 8770 6096 8801 6101
rect 8807 6096 8837 6101
rect 8770 6092 8837 6096
rect 8743 6089 8837 6092
rect 8743 6082 8792 6089
rect 8743 6076 8773 6082
rect 8792 6077 8797 6082
rect 8709 6060 8789 6076
rect 8801 6068 8837 6089
rect 8898 6084 9087 6108
rect 9132 6107 9179 6108
rect 9145 6102 9179 6107
rect 8913 6081 9087 6084
rect 8906 6078 9087 6081
rect 9115 6101 9179 6102
rect 8709 6058 8728 6060
rect 8743 6058 8777 6060
rect 8709 6042 8789 6058
rect 8709 6036 8728 6042
rect 8425 6010 8528 6020
rect 8379 6008 8528 6010
rect 8549 6008 8584 6020
rect 8218 6006 8380 6008
rect 8230 5986 8249 6006
rect 8264 6004 8294 6006
rect 8113 5978 8154 5986
rect 8236 5982 8249 5986
rect 8301 5990 8380 6006
rect 8412 6006 8584 6008
rect 8412 5990 8491 6006
rect 8498 6004 8528 6006
rect 8076 5968 8105 5978
rect 8119 5968 8148 5978
rect 8163 5968 8193 5982
rect 8236 5968 8279 5982
rect 8301 5978 8491 5990
rect 8556 5986 8562 6006
rect 8286 5968 8316 5978
rect 8317 5968 8475 5978
rect 8479 5968 8509 5978
rect 8513 5968 8543 5982
rect 8571 5968 8584 6006
rect 8656 6020 8685 6036
rect 8699 6020 8728 6036
rect 8743 6026 8773 6042
rect 8801 6020 8807 6068
rect 8810 6062 8829 6068
rect 8844 6062 8874 6070
rect 8810 6054 8874 6062
rect 8810 6038 8890 6054
rect 8906 6047 8968 6078
rect 8984 6047 9046 6078
rect 9115 6076 9164 6101
rect 9179 6076 9209 6092
rect 9078 6062 9108 6070
rect 9115 6068 9225 6076
rect 9078 6054 9123 6062
rect 8810 6036 8829 6038
rect 8844 6036 8890 6038
rect 8810 6020 8890 6036
rect 8917 6034 8952 6047
rect 8993 6044 9030 6047
rect 8993 6042 9035 6044
rect 8922 6031 8952 6034
rect 8931 6027 8938 6031
rect 8938 6026 8939 6027
rect 8897 6020 8907 6026
rect 8656 6012 8691 6020
rect 8656 5986 8657 6012
rect 8664 5986 8691 6012
rect 8599 5968 8629 5982
rect 8656 5978 8691 5986
rect 8693 6012 8734 6020
rect 8693 5986 8708 6012
rect 8715 5986 8734 6012
rect 8798 6008 8829 6020
rect 8844 6008 8947 6020
rect 8959 6010 8985 6036
rect 9000 6031 9030 6042
rect 9062 6038 9124 6054
rect 9062 6036 9108 6038
rect 9062 6020 9124 6036
rect 9136 6020 9142 6068
rect 9145 6060 9225 6068
rect 9145 6058 9164 6060
rect 9179 6058 9213 6060
rect 9145 6042 9225 6058
rect 9145 6020 9164 6042
rect 9179 6026 9209 6042
rect 9237 6036 9243 6110
rect 9246 6036 9265 6180
rect 9280 6036 9286 6180
rect 9295 6110 9308 6180
rect 9360 6176 9382 6180
rect 9353 6154 9382 6168
rect 9435 6154 9451 6168
rect 9489 6164 9495 6166
rect 9502 6164 9610 6180
rect 9617 6164 9623 6166
rect 9631 6164 9646 6180
rect 9712 6174 9731 6177
rect 9353 6152 9451 6154
rect 9478 6152 9646 6164
rect 9661 6154 9677 6168
rect 9712 6155 9734 6174
rect 9744 6168 9760 6169
rect 9743 6166 9760 6168
rect 9744 6161 9760 6166
rect 9734 6154 9740 6155
rect 9743 6154 9772 6161
rect 9661 6153 9772 6154
rect 9661 6152 9778 6153
rect 9337 6144 9388 6152
rect 9435 6144 9469 6152
rect 9337 6132 9362 6144
rect 9369 6132 9388 6144
rect 9442 6142 9469 6144
rect 9478 6142 9699 6152
rect 9734 6149 9740 6152
rect 9442 6138 9699 6142
rect 9337 6124 9388 6132
rect 9435 6124 9699 6138
rect 9743 6144 9778 6152
rect 9289 6076 9308 6110
rect 9353 6116 9382 6124
rect 9353 6110 9370 6116
rect 9353 6108 9387 6110
rect 9435 6108 9451 6124
rect 9452 6114 9660 6124
rect 9661 6114 9677 6124
rect 9725 6120 9740 6135
rect 9743 6132 9744 6144
rect 9751 6132 9778 6144
rect 9743 6124 9778 6132
rect 9743 6123 9772 6124
rect 9463 6110 9677 6114
rect 9478 6108 9677 6110
rect 9712 6110 9725 6120
rect 9743 6110 9760 6123
rect 9712 6108 9760 6110
rect 9354 6104 9387 6108
rect 9350 6102 9387 6104
rect 9350 6101 9417 6102
rect 9350 6096 9381 6101
rect 9387 6096 9417 6101
rect 9350 6092 9417 6096
rect 9323 6089 9417 6092
rect 9323 6082 9372 6089
rect 9323 6076 9353 6082
rect 9372 6077 9377 6082
rect 9289 6060 9369 6076
rect 9381 6068 9417 6089
rect 9478 6084 9667 6108
rect 9712 6107 9759 6108
rect 9725 6102 9759 6107
rect 9493 6081 9667 6084
rect 9486 6078 9667 6081
rect 9695 6101 9759 6102
rect 9289 6058 9308 6060
rect 9323 6058 9357 6060
rect 9289 6042 9369 6058
rect 9289 6036 9308 6042
rect 9005 6010 9108 6020
rect 8959 6008 9108 6010
rect 9129 6008 9164 6020
rect 8798 6006 8960 6008
rect 8810 5986 8829 6006
rect 8844 6004 8874 6006
rect 8693 5978 8734 5986
rect 8816 5982 8829 5986
rect 8881 5990 8960 6006
rect 8992 6006 9164 6008
rect 8992 5990 9071 6006
rect 9078 6004 9108 6006
rect 8656 5968 8685 5978
rect 8699 5968 8728 5978
rect 8743 5968 8773 5982
rect 8816 5968 8859 5982
rect 8881 5978 9071 5990
rect 9136 5986 9142 6006
rect 8866 5968 8896 5978
rect 8897 5968 9055 5978
rect 9059 5968 9089 5978
rect 9093 5968 9123 5982
rect 9151 5968 9164 6006
rect 9236 6020 9265 6036
rect 9279 6020 9308 6036
rect 9323 6026 9353 6042
rect 9381 6020 9387 6068
rect 9390 6062 9409 6068
rect 9424 6062 9454 6070
rect 9390 6054 9454 6062
rect 9390 6038 9470 6054
rect 9486 6047 9548 6078
rect 9564 6047 9626 6078
rect 9695 6076 9744 6101
rect 9759 6076 9789 6092
rect 9658 6062 9688 6070
rect 9695 6068 9805 6076
rect 9658 6054 9703 6062
rect 9390 6036 9409 6038
rect 9424 6036 9470 6038
rect 9390 6020 9470 6036
rect 9497 6034 9532 6047
rect 9573 6044 9610 6047
rect 9573 6042 9615 6044
rect 9502 6031 9532 6034
rect 9511 6027 9518 6031
rect 9518 6026 9519 6027
rect 9477 6020 9487 6026
rect 9236 6012 9271 6020
rect 9236 5986 9237 6012
rect 9244 5986 9271 6012
rect 9179 5968 9209 5982
rect 9236 5978 9271 5986
rect 9273 6012 9314 6020
rect 9273 5986 9288 6012
rect 9295 5986 9314 6012
rect 9378 6008 9409 6020
rect 9424 6008 9527 6020
rect 9539 6010 9565 6036
rect 9580 6031 9610 6042
rect 9642 6038 9704 6054
rect 9642 6036 9688 6038
rect 9642 6020 9704 6036
rect 9716 6020 9722 6068
rect 9725 6060 9805 6068
rect 9725 6058 9744 6060
rect 9759 6058 9793 6060
rect 9725 6042 9805 6058
rect 9725 6020 9744 6042
rect 9759 6026 9789 6042
rect 9817 6036 9823 6110
rect 9826 6036 9845 6180
rect 9860 6036 9866 6180
rect 9875 6110 9888 6180
rect 9940 6176 9962 6180
rect 9933 6154 9962 6168
rect 10015 6154 10031 6168
rect 10069 6164 10075 6166
rect 10082 6164 10190 6180
rect 10197 6164 10203 6166
rect 10211 6164 10226 6180
rect 10292 6174 10311 6177
rect 9933 6152 10031 6154
rect 10058 6152 10226 6164
rect 10241 6154 10257 6168
rect 10292 6155 10314 6174
rect 10324 6168 10340 6169
rect 10323 6166 10340 6168
rect 10324 6161 10340 6166
rect 10314 6154 10320 6155
rect 10323 6154 10352 6161
rect 10241 6153 10352 6154
rect 10241 6152 10358 6153
rect 9917 6144 9968 6152
rect 10015 6144 10049 6152
rect 9917 6132 9942 6144
rect 9949 6132 9968 6144
rect 10022 6142 10049 6144
rect 10058 6142 10279 6152
rect 10314 6149 10320 6152
rect 10022 6138 10279 6142
rect 9917 6124 9968 6132
rect 10015 6124 10279 6138
rect 10323 6144 10358 6152
rect 9869 6076 9888 6110
rect 9933 6116 9962 6124
rect 9933 6110 9950 6116
rect 9933 6108 9967 6110
rect 10015 6108 10031 6124
rect 10032 6114 10240 6124
rect 10241 6114 10257 6124
rect 10305 6120 10320 6135
rect 10323 6132 10324 6144
rect 10331 6132 10358 6144
rect 10323 6124 10358 6132
rect 10323 6123 10352 6124
rect 10043 6110 10257 6114
rect 10058 6108 10257 6110
rect 10292 6110 10305 6120
rect 10323 6110 10340 6123
rect 10292 6108 10340 6110
rect 9934 6104 9967 6108
rect 9930 6102 9967 6104
rect 9930 6101 9997 6102
rect 9930 6096 9961 6101
rect 9967 6096 9997 6101
rect 9930 6092 9997 6096
rect 9903 6089 9997 6092
rect 9903 6082 9952 6089
rect 9903 6076 9933 6082
rect 9952 6077 9957 6082
rect 9869 6060 9949 6076
rect 9961 6068 9997 6089
rect 10058 6084 10247 6108
rect 10292 6107 10339 6108
rect 10305 6102 10339 6107
rect 10073 6081 10247 6084
rect 10066 6078 10247 6081
rect 10275 6101 10339 6102
rect 9869 6058 9888 6060
rect 9903 6058 9937 6060
rect 9869 6042 9949 6058
rect 9869 6036 9888 6042
rect 9585 6010 9688 6020
rect 9539 6008 9688 6010
rect 9709 6008 9744 6020
rect 9378 6006 9540 6008
rect 9390 5986 9409 6006
rect 9424 6004 9454 6006
rect 9273 5978 9314 5986
rect 9396 5982 9409 5986
rect 9461 5990 9540 6006
rect 9572 6006 9744 6008
rect 9572 5990 9651 6006
rect 9658 6004 9688 6006
rect 9236 5968 9265 5978
rect 9279 5968 9308 5978
rect 9323 5968 9353 5982
rect 9396 5968 9439 5982
rect 9461 5978 9651 5990
rect 9716 5986 9722 6006
rect 9446 5968 9476 5978
rect 9477 5968 9635 5978
rect 9639 5968 9669 5978
rect 9673 5968 9703 5982
rect 9731 5968 9744 6006
rect 9816 6020 9845 6036
rect 9859 6020 9888 6036
rect 9903 6026 9933 6042
rect 9961 6020 9967 6068
rect 9970 6062 9989 6068
rect 10004 6062 10034 6070
rect 9970 6054 10034 6062
rect 9970 6038 10050 6054
rect 10066 6047 10128 6078
rect 10144 6047 10206 6078
rect 10275 6076 10324 6101
rect 10339 6076 10369 6092
rect 10238 6062 10268 6070
rect 10275 6068 10385 6076
rect 10238 6054 10283 6062
rect 9970 6036 9989 6038
rect 10004 6036 10050 6038
rect 9970 6020 10050 6036
rect 10077 6034 10112 6047
rect 10153 6044 10190 6047
rect 10153 6042 10195 6044
rect 10082 6031 10112 6034
rect 10091 6027 10098 6031
rect 10098 6026 10099 6027
rect 10057 6020 10067 6026
rect 9816 6012 9851 6020
rect 9816 5986 9817 6012
rect 9824 5986 9851 6012
rect 9759 5968 9789 5982
rect 9816 5978 9851 5986
rect 9853 6012 9894 6020
rect 9853 5986 9868 6012
rect 9875 5986 9894 6012
rect 9958 6008 9989 6020
rect 10004 6008 10107 6020
rect 10119 6010 10145 6036
rect 10160 6031 10190 6042
rect 10222 6038 10284 6054
rect 10222 6036 10268 6038
rect 10222 6020 10284 6036
rect 10296 6020 10302 6068
rect 10305 6060 10385 6068
rect 10305 6058 10324 6060
rect 10339 6058 10373 6060
rect 10305 6042 10385 6058
rect 10305 6020 10324 6042
rect 10339 6026 10369 6042
rect 10397 6036 10403 6110
rect 10406 6036 10425 6180
rect 10440 6036 10446 6180
rect 10455 6110 10468 6180
rect 10520 6176 10542 6180
rect 10513 6154 10542 6168
rect 10595 6154 10611 6168
rect 10649 6164 10655 6166
rect 10662 6164 10770 6180
rect 10777 6164 10783 6166
rect 10791 6164 10806 6180
rect 10872 6174 10891 6177
rect 10513 6152 10611 6154
rect 10638 6152 10806 6164
rect 10821 6154 10837 6168
rect 10872 6155 10894 6174
rect 10904 6168 10920 6169
rect 10903 6166 10920 6168
rect 10904 6161 10920 6166
rect 10894 6154 10900 6155
rect 10903 6154 10932 6161
rect 10821 6153 10932 6154
rect 10821 6152 10938 6153
rect 10497 6144 10548 6152
rect 10595 6144 10629 6152
rect 10497 6132 10522 6144
rect 10529 6132 10548 6144
rect 10602 6142 10629 6144
rect 10638 6142 10859 6152
rect 10894 6149 10900 6152
rect 10602 6138 10859 6142
rect 10497 6124 10548 6132
rect 10595 6124 10859 6138
rect 10903 6144 10938 6152
rect 10449 6076 10468 6110
rect 10513 6116 10542 6124
rect 10513 6110 10530 6116
rect 10513 6108 10547 6110
rect 10595 6108 10611 6124
rect 10612 6114 10820 6124
rect 10821 6114 10837 6124
rect 10885 6120 10900 6135
rect 10903 6132 10904 6144
rect 10911 6132 10938 6144
rect 10903 6124 10938 6132
rect 10903 6123 10932 6124
rect 10623 6110 10837 6114
rect 10638 6108 10837 6110
rect 10872 6110 10885 6120
rect 10903 6110 10920 6123
rect 10872 6108 10920 6110
rect 10514 6104 10547 6108
rect 10510 6102 10547 6104
rect 10510 6101 10577 6102
rect 10510 6096 10541 6101
rect 10547 6096 10577 6101
rect 10510 6092 10577 6096
rect 10483 6089 10577 6092
rect 10483 6082 10532 6089
rect 10483 6076 10513 6082
rect 10532 6077 10537 6082
rect 10449 6060 10529 6076
rect 10541 6068 10577 6089
rect 10638 6084 10827 6108
rect 10872 6107 10919 6108
rect 10885 6102 10919 6107
rect 10653 6081 10827 6084
rect 10646 6078 10827 6081
rect 10855 6101 10919 6102
rect 10449 6058 10468 6060
rect 10483 6058 10517 6060
rect 10449 6042 10529 6058
rect 10449 6036 10468 6042
rect 10165 6010 10268 6020
rect 10119 6008 10268 6010
rect 10289 6008 10324 6020
rect 9958 6006 10120 6008
rect 9970 5986 9989 6006
rect 10004 6004 10034 6006
rect 9853 5978 9894 5986
rect 9976 5982 9989 5986
rect 10041 5990 10120 6006
rect 10152 6006 10324 6008
rect 10152 5990 10231 6006
rect 10238 6004 10268 6006
rect 9816 5968 9845 5978
rect 9859 5968 9888 5978
rect 9903 5968 9933 5982
rect 9976 5968 10019 5982
rect 10041 5978 10231 5990
rect 10296 5986 10302 6006
rect 10026 5968 10056 5978
rect 10057 5968 10215 5978
rect 10219 5968 10249 5978
rect 10253 5968 10283 5982
rect 10311 5968 10324 6006
rect 10396 6020 10425 6036
rect 10439 6020 10468 6036
rect 10483 6026 10513 6042
rect 10541 6020 10547 6068
rect 10550 6062 10569 6068
rect 10584 6062 10614 6070
rect 10550 6054 10614 6062
rect 10550 6038 10630 6054
rect 10646 6047 10708 6078
rect 10724 6047 10786 6078
rect 10855 6076 10904 6101
rect 10919 6076 10949 6092
rect 10818 6062 10848 6070
rect 10855 6068 10965 6076
rect 10818 6054 10863 6062
rect 10550 6036 10569 6038
rect 10584 6036 10630 6038
rect 10550 6020 10630 6036
rect 10657 6034 10692 6047
rect 10733 6044 10770 6047
rect 10733 6042 10775 6044
rect 10662 6031 10692 6034
rect 10671 6027 10678 6031
rect 10678 6026 10679 6027
rect 10637 6020 10647 6026
rect 10396 6012 10431 6020
rect 10396 5986 10397 6012
rect 10404 5986 10431 6012
rect 10339 5968 10369 5982
rect 10396 5978 10431 5986
rect 10433 6012 10474 6020
rect 10433 5986 10448 6012
rect 10455 5986 10474 6012
rect 10538 6008 10569 6020
rect 10584 6008 10687 6020
rect 10699 6010 10725 6036
rect 10740 6031 10770 6042
rect 10802 6038 10864 6054
rect 10802 6036 10848 6038
rect 10802 6020 10864 6036
rect 10876 6020 10882 6068
rect 10885 6060 10965 6068
rect 10885 6058 10904 6060
rect 10919 6058 10953 6060
rect 10885 6042 10965 6058
rect 10885 6020 10904 6042
rect 10919 6026 10949 6042
rect 10977 6036 10983 6110
rect 10986 6036 11005 6180
rect 11020 6036 11026 6180
rect 11035 6110 11048 6180
rect 11100 6176 11122 6180
rect 11093 6154 11122 6168
rect 11175 6154 11191 6168
rect 11229 6164 11235 6166
rect 11242 6164 11350 6180
rect 11357 6164 11363 6166
rect 11371 6164 11386 6180
rect 11452 6174 11471 6177
rect 11093 6152 11191 6154
rect 11218 6152 11386 6164
rect 11401 6154 11417 6168
rect 11452 6155 11474 6174
rect 11484 6168 11500 6169
rect 11483 6166 11500 6168
rect 11484 6161 11500 6166
rect 11474 6154 11480 6155
rect 11483 6154 11512 6161
rect 11401 6153 11512 6154
rect 11401 6152 11518 6153
rect 11077 6144 11128 6152
rect 11175 6144 11209 6152
rect 11077 6132 11102 6144
rect 11109 6132 11128 6144
rect 11182 6142 11209 6144
rect 11218 6142 11439 6152
rect 11474 6149 11480 6152
rect 11182 6138 11439 6142
rect 11077 6124 11128 6132
rect 11175 6124 11439 6138
rect 11483 6144 11518 6152
rect 11029 6076 11048 6110
rect 11093 6116 11122 6124
rect 11093 6110 11110 6116
rect 11093 6108 11127 6110
rect 11175 6108 11191 6124
rect 11192 6114 11400 6124
rect 11401 6114 11417 6124
rect 11465 6120 11480 6135
rect 11483 6132 11484 6144
rect 11491 6132 11518 6144
rect 11483 6124 11518 6132
rect 11483 6123 11512 6124
rect 11203 6110 11417 6114
rect 11218 6108 11417 6110
rect 11452 6110 11465 6120
rect 11483 6110 11500 6123
rect 11452 6108 11500 6110
rect 11094 6104 11127 6108
rect 11090 6102 11127 6104
rect 11090 6101 11157 6102
rect 11090 6096 11121 6101
rect 11127 6096 11157 6101
rect 11090 6092 11157 6096
rect 11063 6089 11157 6092
rect 11063 6082 11112 6089
rect 11063 6076 11093 6082
rect 11112 6077 11117 6082
rect 11029 6060 11109 6076
rect 11121 6068 11157 6089
rect 11218 6084 11407 6108
rect 11452 6107 11499 6108
rect 11465 6102 11499 6107
rect 11233 6081 11407 6084
rect 11226 6078 11407 6081
rect 11435 6101 11499 6102
rect 11029 6058 11048 6060
rect 11063 6058 11097 6060
rect 11029 6042 11109 6058
rect 11029 6036 11048 6042
rect 10745 6010 10848 6020
rect 10699 6008 10848 6010
rect 10869 6008 10904 6020
rect 10538 6006 10700 6008
rect 10550 5986 10569 6006
rect 10584 6004 10614 6006
rect 10433 5978 10474 5986
rect 10556 5982 10569 5986
rect 10621 5990 10700 6006
rect 10732 6006 10904 6008
rect 10732 5990 10811 6006
rect 10818 6004 10848 6006
rect 10396 5968 10425 5978
rect 10439 5968 10468 5978
rect 10483 5968 10513 5982
rect 10556 5968 10599 5982
rect 10621 5978 10811 5990
rect 10876 5986 10882 6006
rect 10606 5968 10636 5978
rect 10637 5968 10795 5978
rect 10799 5968 10829 5978
rect 10833 5968 10863 5982
rect 10891 5968 10904 6006
rect 10976 6020 11005 6036
rect 11019 6020 11048 6036
rect 11063 6026 11093 6042
rect 11121 6020 11127 6068
rect 11130 6062 11149 6068
rect 11164 6062 11194 6070
rect 11130 6054 11194 6062
rect 11130 6038 11210 6054
rect 11226 6047 11288 6078
rect 11304 6047 11366 6078
rect 11435 6076 11484 6101
rect 11499 6076 11529 6092
rect 11398 6062 11428 6070
rect 11435 6068 11545 6076
rect 11398 6054 11443 6062
rect 11130 6036 11149 6038
rect 11164 6036 11210 6038
rect 11130 6020 11210 6036
rect 11237 6034 11272 6047
rect 11313 6044 11350 6047
rect 11313 6042 11355 6044
rect 11242 6031 11272 6034
rect 11251 6027 11258 6031
rect 11258 6026 11259 6027
rect 11217 6020 11227 6026
rect 10976 6012 11011 6020
rect 10976 5986 10977 6012
rect 10984 5986 11011 6012
rect 10919 5968 10949 5982
rect 10976 5978 11011 5986
rect 11013 6012 11054 6020
rect 11013 5986 11028 6012
rect 11035 5986 11054 6012
rect 11118 6008 11149 6020
rect 11164 6008 11267 6020
rect 11279 6010 11305 6036
rect 11320 6031 11350 6042
rect 11382 6038 11444 6054
rect 11382 6036 11428 6038
rect 11382 6020 11444 6036
rect 11456 6020 11462 6068
rect 11465 6060 11545 6068
rect 11465 6058 11484 6060
rect 11499 6058 11533 6060
rect 11465 6042 11545 6058
rect 11465 6020 11484 6042
rect 11499 6026 11529 6042
rect 11557 6036 11563 6110
rect 11566 6036 11585 6180
rect 11600 6036 11606 6180
rect 11615 6110 11628 6180
rect 11680 6176 11702 6180
rect 11673 6154 11702 6168
rect 11755 6154 11771 6168
rect 11809 6164 11815 6166
rect 11822 6164 11930 6180
rect 11937 6164 11943 6166
rect 11951 6164 11966 6180
rect 12032 6174 12051 6177
rect 11673 6152 11771 6154
rect 11798 6152 11966 6164
rect 11981 6154 11997 6168
rect 12032 6155 12054 6174
rect 12064 6168 12080 6169
rect 12063 6166 12080 6168
rect 12064 6161 12080 6166
rect 12054 6154 12060 6155
rect 12063 6154 12092 6161
rect 11981 6153 12092 6154
rect 11981 6152 12098 6153
rect 11657 6144 11708 6152
rect 11755 6144 11789 6152
rect 11657 6132 11682 6144
rect 11689 6132 11708 6144
rect 11762 6142 11789 6144
rect 11798 6142 12019 6152
rect 12054 6149 12060 6152
rect 11762 6138 12019 6142
rect 11657 6124 11708 6132
rect 11755 6124 12019 6138
rect 12063 6144 12098 6152
rect 11609 6076 11628 6110
rect 11673 6116 11702 6124
rect 11673 6110 11690 6116
rect 11673 6108 11707 6110
rect 11755 6108 11771 6124
rect 11772 6114 11980 6124
rect 11981 6114 11997 6124
rect 12045 6120 12060 6135
rect 12063 6132 12064 6144
rect 12071 6132 12098 6144
rect 12063 6124 12098 6132
rect 12063 6123 12092 6124
rect 11783 6110 11997 6114
rect 11798 6108 11997 6110
rect 12032 6110 12045 6120
rect 12063 6110 12080 6123
rect 12032 6108 12080 6110
rect 11674 6104 11707 6108
rect 11670 6102 11707 6104
rect 11670 6101 11737 6102
rect 11670 6096 11701 6101
rect 11707 6096 11737 6101
rect 11670 6092 11737 6096
rect 11643 6089 11737 6092
rect 11643 6082 11692 6089
rect 11643 6076 11673 6082
rect 11692 6077 11697 6082
rect 11609 6060 11689 6076
rect 11701 6068 11737 6089
rect 11798 6084 11987 6108
rect 12032 6107 12079 6108
rect 12045 6102 12079 6107
rect 11813 6081 11987 6084
rect 11806 6078 11987 6081
rect 12015 6101 12079 6102
rect 11609 6058 11628 6060
rect 11643 6058 11677 6060
rect 11609 6042 11689 6058
rect 11609 6036 11628 6042
rect 11325 6010 11428 6020
rect 11279 6008 11428 6010
rect 11449 6008 11484 6020
rect 11118 6006 11280 6008
rect 11130 5986 11149 6006
rect 11164 6004 11194 6006
rect 11013 5978 11054 5986
rect 11136 5982 11149 5986
rect 11201 5990 11280 6006
rect 11312 6006 11484 6008
rect 11312 5990 11391 6006
rect 11398 6004 11428 6006
rect 10976 5968 11005 5978
rect 11019 5968 11048 5978
rect 11063 5968 11093 5982
rect 11136 5968 11179 5982
rect 11201 5978 11391 5990
rect 11456 5986 11462 6006
rect 11186 5968 11216 5978
rect 11217 5968 11375 5978
rect 11379 5968 11409 5978
rect 11413 5968 11443 5982
rect 11471 5968 11484 6006
rect 11556 6020 11585 6036
rect 11599 6020 11628 6036
rect 11643 6026 11673 6042
rect 11701 6020 11707 6068
rect 11710 6062 11729 6068
rect 11744 6062 11774 6070
rect 11710 6054 11774 6062
rect 11710 6038 11790 6054
rect 11806 6047 11868 6078
rect 11884 6047 11946 6078
rect 12015 6076 12064 6101
rect 12079 6076 12109 6092
rect 11978 6062 12008 6070
rect 12015 6068 12125 6076
rect 11978 6054 12023 6062
rect 11710 6036 11729 6038
rect 11744 6036 11790 6038
rect 11710 6020 11790 6036
rect 11817 6034 11852 6047
rect 11893 6044 11930 6047
rect 11893 6042 11935 6044
rect 11822 6031 11852 6034
rect 11831 6027 11838 6031
rect 11838 6026 11839 6027
rect 11797 6020 11807 6026
rect 11556 6012 11591 6020
rect 11556 5986 11557 6012
rect 11564 5986 11591 6012
rect 11499 5968 11529 5982
rect 11556 5978 11591 5986
rect 11593 6012 11634 6020
rect 11593 5986 11608 6012
rect 11615 5986 11634 6012
rect 11698 6008 11729 6020
rect 11744 6008 11847 6020
rect 11859 6010 11885 6036
rect 11900 6031 11930 6042
rect 11962 6038 12024 6054
rect 11962 6036 12008 6038
rect 11962 6020 12024 6036
rect 12036 6020 12042 6068
rect 12045 6060 12125 6068
rect 12045 6058 12064 6060
rect 12079 6058 12113 6060
rect 12045 6042 12125 6058
rect 12045 6020 12064 6042
rect 12079 6026 12109 6042
rect 12137 6036 12143 6110
rect 12146 6036 12165 6180
rect 12180 6036 12186 6180
rect 12195 6110 12208 6180
rect 12260 6176 12282 6180
rect 12253 6154 12282 6168
rect 12335 6154 12351 6168
rect 12389 6164 12395 6166
rect 12402 6164 12510 6180
rect 12517 6164 12523 6166
rect 12531 6164 12546 6180
rect 12612 6174 12631 6177
rect 12253 6152 12351 6154
rect 12378 6152 12546 6164
rect 12561 6154 12577 6168
rect 12612 6155 12634 6174
rect 12644 6168 12660 6169
rect 12643 6166 12660 6168
rect 12644 6161 12660 6166
rect 12634 6154 12640 6155
rect 12643 6154 12672 6161
rect 12561 6153 12672 6154
rect 12561 6152 12678 6153
rect 12237 6144 12288 6152
rect 12335 6144 12369 6152
rect 12237 6132 12262 6144
rect 12269 6132 12288 6144
rect 12342 6142 12369 6144
rect 12378 6142 12599 6152
rect 12634 6149 12640 6152
rect 12342 6138 12599 6142
rect 12237 6124 12288 6132
rect 12335 6124 12599 6138
rect 12643 6144 12678 6152
rect 12189 6076 12208 6110
rect 12253 6116 12282 6124
rect 12253 6110 12270 6116
rect 12253 6108 12287 6110
rect 12335 6108 12351 6124
rect 12352 6114 12560 6124
rect 12561 6114 12577 6124
rect 12625 6120 12640 6135
rect 12643 6132 12644 6144
rect 12651 6132 12678 6144
rect 12643 6124 12678 6132
rect 12643 6123 12672 6124
rect 12363 6110 12577 6114
rect 12378 6108 12577 6110
rect 12612 6110 12625 6120
rect 12643 6110 12660 6123
rect 12612 6108 12660 6110
rect 12254 6104 12287 6108
rect 12250 6102 12287 6104
rect 12250 6101 12317 6102
rect 12250 6096 12281 6101
rect 12287 6096 12317 6101
rect 12250 6092 12317 6096
rect 12223 6089 12317 6092
rect 12223 6082 12272 6089
rect 12223 6076 12253 6082
rect 12272 6077 12277 6082
rect 12189 6060 12269 6076
rect 12281 6068 12317 6089
rect 12378 6084 12567 6108
rect 12612 6107 12659 6108
rect 12625 6102 12659 6107
rect 12393 6081 12567 6084
rect 12386 6078 12567 6081
rect 12595 6101 12659 6102
rect 12189 6058 12208 6060
rect 12223 6058 12257 6060
rect 12189 6042 12269 6058
rect 12189 6036 12208 6042
rect 11905 6010 12008 6020
rect 11859 6008 12008 6010
rect 12029 6008 12064 6020
rect 11698 6006 11860 6008
rect 11710 5986 11729 6006
rect 11744 6004 11774 6006
rect 11593 5978 11634 5986
rect 11716 5982 11729 5986
rect 11781 5990 11860 6006
rect 11892 6006 12064 6008
rect 11892 5990 11971 6006
rect 11978 6004 12008 6006
rect 11556 5968 11585 5978
rect 11599 5968 11628 5978
rect 11643 5968 11673 5982
rect 11716 5968 11759 5982
rect 11781 5978 11971 5990
rect 12036 5986 12042 6006
rect 11766 5968 11796 5978
rect 11797 5968 11955 5978
rect 11959 5968 11989 5978
rect 11993 5968 12023 5982
rect 12051 5968 12064 6006
rect 12136 6020 12165 6036
rect 12179 6020 12208 6036
rect 12223 6026 12253 6042
rect 12281 6020 12287 6068
rect 12290 6062 12309 6068
rect 12324 6062 12354 6070
rect 12290 6054 12354 6062
rect 12290 6038 12370 6054
rect 12386 6047 12448 6078
rect 12464 6047 12526 6078
rect 12595 6076 12644 6101
rect 12659 6076 12689 6092
rect 12558 6062 12588 6070
rect 12595 6068 12705 6076
rect 12558 6054 12603 6062
rect 12290 6036 12309 6038
rect 12324 6036 12370 6038
rect 12290 6020 12370 6036
rect 12397 6034 12432 6047
rect 12473 6044 12510 6047
rect 12473 6042 12515 6044
rect 12402 6031 12432 6034
rect 12411 6027 12418 6031
rect 12418 6026 12419 6027
rect 12377 6020 12387 6026
rect 12136 6012 12171 6020
rect 12136 5986 12137 6012
rect 12144 5986 12171 6012
rect 12079 5968 12109 5982
rect 12136 5978 12171 5986
rect 12173 6012 12214 6020
rect 12173 5986 12188 6012
rect 12195 5986 12214 6012
rect 12278 6008 12309 6020
rect 12324 6008 12427 6020
rect 12439 6010 12465 6036
rect 12480 6031 12510 6042
rect 12542 6038 12604 6054
rect 12542 6036 12588 6038
rect 12542 6020 12604 6036
rect 12616 6020 12622 6068
rect 12625 6060 12705 6068
rect 12625 6058 12644 6060
rect 12659 6058 12693 6060
rect 12625 6042 12705 6058
rect 12625 6020 12644 6042
rect 12659 6026 12689 6042
rect 12717 6036 12723 6110
rect 12726 6036 12745 6180
rect 12760 6036 12766 6180
rect 12775 6110 12788 6180
rect 12840 6176 12862 6180
rect 12833 6154 12862 6168
rect 12915 6154 12931 6168
rect 12969 6164 12975 6166
rect 12982 6164 13090 6180
rect 13097 6164 13103 6166
rect 13111 6164 13126 6180
rect 13192 6174 13211 6177
rect 12833 6152 12931 6154
rect 12958 6152 13126 6164
rect 13141 6154 13157 6168
rect 13192 6155 13214 6174
rect 13224 6168 13240 6169
rect 13223 6166 13240 6168
rect 13224 6161 13240 6166
rect 13214 6154 13220 6155
rect 13223 6154 13252 6161
rect 13141 6153 13252 6154
rect 13141 6152 13258 6153
rect 12817 6144 12868 6152
rect 12915 6144 12949 6152
rect 12817 6132 12842 6144
rect 12849 6132 12868 6144
rect 12922 6142 12949 6144
rect 12958 6142 13179 6152
rect 13214 6149 13220 6152
rect 12922 6138 13179 6142
rect 12817 6124 12868 6132
rect 12915 6124 13179 6138
rect 13223 6144 13258 6152
rect 12769 6076 12788 6110
rect 12833 6116 12862 6124
rect 12833 6110 12850 6116
rect 12833 6108 12867 6110
rect 12915 6108 12931 6124
rect 12932 6114 13140 6124
rect 13141 6114 13157 6124
rect 13205 6120 13220 6135
rect 13223 6132 13224 6144
rect 13231 6132 13258 6144
rect 13223 6124 13258 6132
rect 13223 6123 13252 6124
rect 12943 6110 13157 6114
rect 12958 6108 13157 6110
rect 13192 6110 13205 6120
rect 13223 6110 13240 6123
rect 13192 6108 13240 6110
rect 12834 6104 12867 6108
rect 12830 6102 12867 6104
rect 12830 6101 12897 6102
rect 12830 6096 12861 6101
rect 12867 6096 12897 6101
rect 12830 6092 12897 6096
rect 12803 6089 12897 6092
rect 12803 6082 12852 6089
rect 12803 6076 12833 6082
rect 12852 6077 12857 6082
rect 12769 6060 12849 6076
rect 12861 6068 12897 6089
rect 12958 6084 13147 6108
rect 13192 6107 13239 6108
rect 13205 6102 13239 6107
rect 12973 6081 13147 6084
rect 12966 6078 13147 6081
rect 13175 6101 13239 6102
rect 12769 6058 12788 6060
rect 12803 6058 12837 6060
rect 12769 6042 12849 6058
rect 12769 6036 12788 6042
rect 12485 6010 12588 6020
rect 12439 6008 12588 6010
rect 12609 6008 12644 6020
rect 12278 6006 12440 6008
rect 12290 5986 12309 6006
rect 12324 6004 12354 6006
rect 12173 5978 12214 5986
rect 12296 5982 12309 5986
rect 12361 5990 12440 6006
rect 12472 6006 12644 6008
rect 12472 5990 12551 6006
rect 12558 6004 12588 6006
rect 12136 5968 12165 5978
rect 12179 5968 12208 5978
rect 12223 5968 12253 5982
rect 12296 5968 12339 5982
rect 12361 5978 12551 5990
rect 12616 5986 12622 6006
rect 12346 5968 12376 5978
rect 12377 5968 12535 5978
rect 12539 5968 12569 5978
rect 12573 5968 12603 5982
rect 12631 5968 12644 6006
rect 12716 6020 12745 6036
rect 12759 6020 12788 6036
rect 12803 6026 12833 6042
rect 12861 6020 12867 6068
rect 12870 6062 12889 6068
rect 12904 6062 12934 6070
rect 12870 6054 12934 6062
rect 12870 6038 12950 6054
rect 12966 6047 13028 6078
rect 13044 6047 13106 6078
rect 13175 6076 13224 6101
rect 13239 6076 13269 6092
rect 13138 6062 13168 6070
rect 13175 6068 13285 6076
rect 13138 6054 13183 6062
rect 12870 6036 12889 6038
rect 12904 6036 12950 6038
rect 12870 6020 12950 6036
rect 12977 6034 13012 6047
rect 13053 6044 13090 6047
rect 13053 6042 13095 6044
rect 12982 6031 13012 6034
rect 12991 6027 12998 6031
rect 12998 6026 12999 6027
rect 12957 6020 12967 6026
rect 12716 6012 12751 6020
rect 12716 5986 12717 6012
rect 12724 5986 12751 6012
rect 12659 5968 12689 5982
rect 12716 5978 12751 5986
rect 12753 6012 12794 6020
rect 12753 5986 12768 6012
rect 12775 5986 12794 6012
rect 12858 6008 12889 6020
rect 12904 6008 13007 6020
rect 13019 6010 13045 6036
rect 13060 6031 13090 6042
rect 13122 6038 13184 6054
rect 13122 6036 13168 6038
rect 13122 6020 13184 6036
rect 13196 6020 13202 6068
rect 13205 6060 13285 6068
rect 13205 6058 13224 6060
rect 13239 6058 13273 6060
rect 13205 6042 13285 6058
rect 13205 6020 13224 6042
rect 13239 6026 13269 6042
rect 13297 6036 13303 6110
rect 13306 6036 13325 6180
rect 13340 6036 13346 6180
rect 13355 6110 13368 6180
rect 13420 6176 13442 6180
rect 13413 6154 13442 6168
rect 13495 6154 13511 6168
rect 13549 6164 13555 6166
rect 13562 6164 13670 6180
rect 13677 6164 13683 6166
rect 13691 6164 13706 6180
rect 13772 6174 13791 6177
rect 13413 6152 13511 6154
rect 13538 6152 13706 6164
rect 13721 6154 13737 6168
rect 13772 6155 13794 6174
rect 13804 6168 13820 6169
rect 13803 6166 13820 6168
rect 13804 6161 13820 6166
rect 13794 6154 13800 6155
rect 13803 6154 13832 6161
rect 13721 6153 13832 6154
rect 13721 6152 13838 6153
rect 13397 6144 13448 6152
rect 13495 6144 13529 6152
rect 13397 6132 13422 6144
rect 13429 6132 13448 6144
rect 13502 6142 13529 6144
rect 13538 6142 13759 6152
rect 13794 6149 13800 6152
rect 13502 6138 13759 6142
rect 13397 6124 13448 6132
rect 13495 6124 13759 6138
rect 13803 6144 13838 6152
rect 13349 6076 13368 6110
rect 13413 6116 13442 6124
rect 13413 6110 13430 6116
rect 13413 6108 13447 6110
rect 13495 6108 13511 6124
rect 13512 6114 13720 6124
rect 13721 6114 13737 6124
rect 13785 6120 13800 6135
rect 13803 6132 13804 6144
rect 13811 6132 13838 6144
rect 13803 6124 13838 6132
rect 13803 6123 13832 6124
rect 13523 6110 13737 6114
rect 13538 6108 13737 6110
rect 13772 6110 13785 6120
rect 13803 6110 13820 6123
rect 13772 6108 13820 6110
rect 13414 6104 13447 6108
rect 13410 6102 13447 6104
rect 13410 6101 13477 6102
rect 13410 6096 13441 6101
rect 13447 6096 13477 6101
rect 13410 6092 13477 6096
rect 13383 6089 13477 6092
rect 13383 6082 13432 6089
rect 13383 6076 13413 6082
rect 13432 6077 13437 6082
rect 13349 6060 13429 6076
rect 13441 6068 13477 6089
rect 13538 6084 13727 6108
rect 13772 6107 13819 6108
rect 13785 6102 13819 6107
rect 13553 6081 13727 6084
rect 13546 6078 13727 6081
rect 13755 6101 13819 6102
rect 13349 6058 13368 6060
rect 13383 6058 13417 6060
rect 13349 6042 13429 6058
rect 13349 6036 13368 6042
rect 13065 6010 13168 6020
rect 13019 6008 13168 6010
rect 13189 6008 13224 6020
rect 12858 6006 13020 6008
rect 12870 5986 12889 6006
rect 12904 6004 12934 6006
rect 12753 5978 12794 5986
rect 12876 5982 12889 5986
rect 12941 5990 13020 6006
rect 13052 6006 13224 6008
rect 13052 5990 13131 6006
rect 13138 6004 13168 6006
rect 12716 5968 12745 5978
rect 12759 5968 12788 5978
rect 12803 5968 12833 5982
rect 12876 5968 12919 5982
rect 12941 5978 13131 5990
rect 13196 5986 13202 6006
rect 12926 5968 12956 5978
rect 12957 5968 13115 5978
rect 13119 5968 13149 5978
rect 13153 5968 13183 5982
rect 13211 5968 13224 6006
rect 13296 6020 13325 6036
rect 13339 6020 13368 6036
rect 13383 6026 13413 6042
rect 13441 6020 13447 6068
rect 13450 6062 13469 6068
rect 13484 6062 13514 6070
rect 13450 6054 13514 6062
rect 13450 6038 13530 6054
rect 13546 6047 13608 6078
rect 13624 6047 13686 6078
rect 13755 6076 13804 6101
rect 13819 6076 13849 6092
rect 13718 6062 13748 6070
rect 13755 6068 13865 6076
rect 13718 6054 13763 6062
rect 13450 6036 13469 6038
rect 13484 6036 13530 6038
rect 13450 6020 13530 6036
rect 13557 6034 13592 6047
rect 13633 6044 13670 6047
rect 13633 6042 13675 6044
rect 13562 6031 13592 6034
rect 13571 6027 13578 6031
rect 13578 6026 13579 6027
rect 13537 6020 13547 6026
rect 13296 6012 13331 6020
rect 13296 5986 13297 6012
rect 13304 5986 13331 6012
rect 13239 5968 13269 5982
rect 13296 5978 13331 5986
rect 13333 6012 13374 6020
rect 13333 5986 13348 6012
rect 13355 5986 13374 6012
rect 13438 6008 13469 6020
rect 13484 6008 13587 6020
rect 13599 6010 13625 6036
rect 13640 6031 13670 6042
rect 13702 6038 13764 6054
rect 13702 6036 13748 6038
rect 13702 6020 13764 6036
rect 13776 6020 13782 6068
rect 13785 6060 13865 6068
rect 13785 6058 13804 6060
rect 13819 6058 13853 6060
rect 13785 6042 13865 6058
rect 13785 6020 13804 6042
rect 13819 6026 13849 6042
rect 13877 6036 13883 6110
rect 13886 6036 13905 6180
rect 13920 6036 13926 6180
rect 13935 6110 13948 6180
rect 14000 6176 14022 6180
rect 13993 6154 14022 6168
rect 14075 6154 14091 6168
rect 14129 6164 14135 6166
rect 14142 6164 14250 6180
rect 14257 6164 14263 6166
rect 14271 6164 14286 6180
rect 14352 6174 14371 6177
rect 13993 6152 14091 6154
rect 14118 6152 14286 6164
rect 14301 6154 14317 6168
rect 14352 6155 14374 6174
rect 14384 6168 14400 6169
rect 14383 6166 14400 6168
rect 14384 6161 14400 6166
rect 14374 6154 14380 6155
rect 14383 6154 14412 6161
rect 14301 6153 14412 6154
rect 14301 6152 14418 6153
rect 13977 6144 14028 6152
rect 14075 6144 14109 6152
rect 13977 6132 14002 6144
rect 14009 6132 14028 6144
rect 14082 6142 14109 6144
rect 14118 6142 14339 6152
rect 14374 6149 14380 6152
rect 14082 6138 14339 6142
rect 13977 6124 14028 6132
rect 14075 6124 14339 6138
rect 14383 6144 14418 6152
rect 13929 6076 13948 6110
rect 13993 6116 14022 6124
rect 13993 6110 14010 6116
rect 13993 6108 14027 6110
rect 14075 6108 14091 6124
rect 14092 6114 14300 6124
rect 14301 6114 14317 6124
rect 14365 6120 14380 6135
rect 14383 6132 14384 6144
rect 14391 6132 14418 6144
rect 14383 6124 14418 6132
rect 14383 6123 14412 6124
rect 14103 6110 14317 6114
rect 14118 6108 14317 6110
rect 14352 6110 14365 6120
rect 14383 6110 14400 6123
rect 14352 6108 14400 6110
rect 13994 6104 14027 6108
rect 13990 6102 14027 6104
rect 13990 6101 14057 6102
rect 13990 6096 14021 6101
rect 14027 6096 14057 6101
rect 13990 6092 14057 6096
rect 13963 6089 14057 6092
rect 13963 6082 14012 6089
rect 13963 6076 13993 6082
rect 14012 6077 14017 6082
rect 13929 6060 14009 6076
rect 14021 6068 14057 6089
rect 14118 6084 14307 6108
rect 14352 6107 14399 6108
rect 14365 6102 14399 6107
rect 14133 6081 14307 6084
rect 14126 6078 14307 6081
rect 14335 6101 14399 6102
rect 13929 6058 13948 6060
rect 13963 6058 13997 6060
rect 13929 6042 14009 6058
rect 13929 6036 13948 6042
rect 13645 6010 13748 6020
rect 13599 6008 13748 6010
rect 13769 6008 13804 6020
rect 13438 6006 13600 6008
rect 13450 5986 13469 6006
rect 13484 6004 13514 6006
rect 13333 5978 13374 5986
rect 13456 5982 13469 5986
rect 13521 5990 13600 6006
rect 13632 6006 13804 6008
rect 13632 5990 13711 6006
rect 13718 6004 13748 6006
rect 13296 5968 13325 5978
rect 13339 5968 13368 5978
rect 13383 5968 13413 5982
rect 13456 5968 13499 5982
rect 13521 5978 13711 5990
rect 13776 5986 13782 6006
rect 13506 5968 13536 5978
rect 13537 5968 13695 5978
rect 13699 5968 13729 5978
rect 13733 5968 13763 5982
rect 13791 5968 13804 6006
rect 13876 6020 13905 6036
rect 13919 6020 13948 6036
rect 13963 6026 13993 6042
rect 14021 6020 14027 6068
rect 14030 6062 14049 6068
rect 14064 6062 14094 6070
rect 14030 6054 14094 6062
rect 14030 6038 14110 6054
rect 14126 6047 14188 6078
rect 14204 6047 14266 6078
rect 14335 6076 14384 6101
rect 14399 6076 14429 6092
rect 14298 6062 14328 6070
rect 14335 6068 14445 6076
rect 14298 6054 14343 6062
rect 14030 6036 14049 6038
rect 14064 6036 14110 6038
rect 14030 6020 14110 6036
rect 14137 6034 14172 6047
rect 14213 6044 14250 6047
rect 14213 6042 14255 6044
rect 14142 6031 14172 6034
rect 14151 6027 14158 6031
rect 14158 6026 14159 6027
rect 14117 6020 14127 6026
rect 13876 6012 13911 6020
rect 13876 5986 13877 6012
rect 13884 5986 13911 6012
rect 13819 5968 13849 5982
rect 13876 5978 13911 5986
rect 13913 6012 13954 6020
rect 13913 5986 13928 6012
rect 13935 5986 13954 6012
rect 14018 6008 14049 6020
rect 14064 6008 14167 6020
rect 14179 6010 14205 6036
rect 14220 6031 14250 6042
rect 14282 6038 14344 6054
rect 14282 6036 14328 6038
rect 14282 6020 14344 6036
rect 14356 6020 14362 6068
rect 14365 6060 14445 6068
rect 14365 6058 14384 6060
rect 14399 6058 14433 6060
rect 14365 6042 14445 6058
rect 14365 6020 14384 6042
rect 14399 6026 14429 6042
rect 14457 6036 14463 6110
rect 14466 6036 14485 6180
rect 14500 6036 14506 6180
rect 14515 6110 14528 6180
rect 14580 6176 14602 6180
rect 14573 6154 14602 6168
rect 14655 6154 14671 6168
rect 14709 6164 14715 6166
rect 14722 6164 14830 6180
rect 14837 6164 14843 6166
rect 14851 6164 14866 6180
rect 14932 6174 14951 6177
rect 14573 6152 14671 6154
rect 14698 6152 14866 6164
rect 14881 6154 14897 6168
rect 14932 6155 14954 6174
rect 14964 6168 14980 6169
rect 14963 6166 14980 6168
rect 14964 6161 14980 6166
rect 14954 6154 14960 6155
rect 14963 6154 14992 6161
rect 14881 6153 14992 6154
rect 14881 6152 14998 6153
rect 14557 6144 14608 6152
rect 14655 6144 14689 6152
rect 14557 6132 14582 6144
rect 14589 6132 14608 6144
rect 14662 6142 14689 6144
rect 14698 6142 14919 6152
rect 14954 6149 14960 6152
rect 14662 6138 14919 6142
rect 14557 6124 14608 6132
rect 14655 6124 14919 6138
rect 14963 6144 14998 6152
rect 14509 6076 14528 6110
rect 14573 6116 14602 6124
rect 14573 6110 14590 6116
rect 14573 6108 14607 6110
rect 14655 6108 14671 6124
rect 14672 6114 14880 6124
rect 14881 6114 14897 6124
rect 14945 6120 14960 6135
rect 14963 6132 14964 6144
rect 14971 6132 14998 6144
rect 14963 6124 14998 6132
rect 14963 6123 14992 6124
rect 14683 6110 14897 6114
rect 14698 6108 14897 6110
rect 14932 6110 14945 6120
rect 14963 6110 14980 6123
rect 14932 6108 14980 6110
rect 14574 6104 14607 6108
rect 14570 6102 14607 6104
rect 14570 6101 14637 6102
rect 14570 6096 14601 6101
rect 14607 6096 14637 6101
rect 14570 6092 14637 6096
rect 14543 6089 14637 6092
rect 14543 6082 14592 6089
rect 14543 6076 14573 6082
rect 14592 6077 14597 6082
rect 14509 6060 14589 6076
rect 14601 6068 14637 6089
rect 14698 6084 14887 6108
rect 14932 6107 14979 6108
rect 14945 6102 14979 6107
rect 14713 6081 14887 6084
rect 14706 6078 14887 6081
rect 14915 6101 14979 6102
rect 14509 6058 14528 6060
rect 14543 6058 14577 6060
rect 14509 6042 14589 6058
rect 14509 6036 14528 6042
rect 14225 6010 14328 6020
rect 14179 6008 14328 6010
rect 14349 6008 14384 6020
rect 14018 6006 14180 6008
rect 14030 5986 14049 6006
rect 14064 6004 14094 6006
rect 13913 5978 13954 5986
rect 14036 5982 14049 5986
rect 14101 5990 14180 6006
rect 14212 6006 14384 6008
rect 14212 5990 14291 6006
rect 14298 6004 14328 6006
rect 13876 5968 13905 5978
rect 13919 5968 13948 5978
rect 13963 5968 13993 5982
rect 14036 5968 14079 5982
rect 14101 5978 14291 5990
rect 14356 5986 14362 6006
rect 14086 5968 14116 5978
rect 14117 5968 14275 5978
rect 14279 5968 14309 5978
rect 14313 5968 14343 5982
rect 14371 5968 14384 6006
rect 14456 6020 14485 6036
rect 14499 6020 14528 6036
rect 14543 6026 14573 6042
rect 14601 6020 14607 6068
rect 14610 6062 14629 6068
rect 14644 6062 14674 6070
rect 14610 6054 14674 6062
rect 14610 6038 14690 6054
rect 14706 6047 14768 6078
rect 14784 6047 14846 6078
rect 14915 6076 14964 6101
rect 14979 6076 15009 6092
rect 14878 6062 14908 6070
rect 14915 6068 15025 6076
rect 14878 6054 14923 6062
rect 14610 6036 14629 6038
rect 14644 6036 14690 6038
rect 14610 6020 14690 6036
rect 14717 6034 14752 6047
rect 14793 6044 14830 6047
rect 14793 6042 14835 6044
rect 14722 6031 14752 6034
rect 14731 6027 14738 6031
rect 14738 6026 14739 6027
rect 14697 6020 14707 6026
rect 14456 6012 14491 6020
rect 14456 5986 14457 6012
rect 14464 5986 14491 6012
rect 14399 5968 14429 5982
rect 14456 5978 14491 5986
rect 14493 6012 14534 6020
rect 14493 5986 14508 6012
rect 14515 5986 14534 6012
rect 14598 6008 14629 6020
rect 14644 6008 14747 6020
rect 14759 6010 14785 6036
rect 14800 6031 14830 6042
rect 14862 6038 14924 6054
rect 14862 6036 14908 6038
rect 14862 6020 14924 6036
rect 14936 6020 14942 6068
rect 14945 6060 15025 6068
rect 14945 6058 14964 6060
rect 14979 6058 15013 6060
rect 14945 6042 15025 6058
rect 14945 6020 14964 6042
rect 14979 6026 15009 6042
rect 15037 6036 15043 6110
rect 15046 6036 15065 6180
rect 15080 6036 15086 6180
rect 15095 6110 15108 6180
rect 15160 6176 15182 6180
rect 15153 6154 15182 6168
rect 15235 6154 15251 6168
rect 15289 6164 15295 6166
rect 15302 6164 15410 6180
rect 15417 6164 15423 6166
rect 15431 6164 15446 6180
rect 15512 6174 15531 6177
rect 15153 6152 15251 6154
rect 15278 6152 15446 6164
rect 15461 6154 15477 6168
rect 15512 6155 15534 6174
rect 15544 6168 15560 6169
rect 15543 6166 15560 6168
rect 15544 6161 15560 6166
rect 15534 6154 15540 6155
rect 15543 6154 15572 6161
rect 15461 6153 15572 6154
rect 15461 6152 15578 6153
rect 15137 6144 15188 6152
rect 15235 6144 15269 6152
rect 15137 6132 15162 6144
rect 15169 6132 15188 6144
rect 15242 6142 15269 6144
rect 15278 6142 15499 6152
rect 15534 6149 15540 6152
rect 15242 6138 15499 6142
rect 15137 6124 15188 6132
rect 15235 6124 15499 6138
rect 15543 6144 15578 6152
rect 15089 6076 15108 6110
rect 15153 6116 15182 6124
rect 15153 6110 15170 6116
rect 15153 6108 15187 6110
rect 15235 6108 15251 6124
rect 15252 6114 15460 6124
rect 15461 6114 15477 6124
rect 15525 6120 15540 6135
rect 15543 6132 15544 6144
rect 15551 6132 15578 6144
rect 15543 6124 15578 6132
rect 15543 6123 15572 6124
rect 15263 6110 15477 6114
rect 15278 6108 15477 6110
rect 15512 6110 15525 6120
rect 15543 6110 15560 6123
rect 15512 6108 15560 6110
rect 15154 6104 15187 6108
rect 15150 6102 15187 6104
rect 15150 6101 15217 6102
rect 15150 6096 15181 6101
rect 15187 6096 15217 6101
rect 15150 6092 15217 6096
rect 15123 6089 15217 6092
rect 15123 6082 15172 6089
rect 15123 6076 15153 6082
rect 15172 6077 15177 6082
rect 15089 6060 15169 6076
rect 15181 6068 15217 6089
rect 15278 6084 15467 6108
rect 15512 6107 15559 6108
rect 15525 6102 15559 6107
rect 15293 6081 15467 6084
rect 15286 6078 15467 6081
rect 15495 6101 15559 6102
rect 15089 6058 15108 6060
rect 15123 6058 15157 6060
rect 15089 6042 15169 6058
rect 15089 6036 15108 6042
rect 14805 6010 14908 6020
rect 14759 6008 14908 6010
rect 14929 6008 14964 6020
rect 14598 6006 14760 6008
rect 14610 5986 14629 6006
rect 14644 6004 14674 6006
rect 14493 5978 14534 5986
rect 14616 5982 14629 5986
rect 14681 5990 14760 6006
rect 14792 6006 14964 6008
rect 14792 5990 14871 6006
rect 14878 6004 14908 6006
rect 14456 5968 14485 5978
rect 14499 5968 14528 5978
rect 14543 5968 14573 5982
rect 14616 5968 14659 5982
rect 14681 5978 14871 5990
rect 14936 5986 14942 6006
rect 14666 5968 14696 5978
rect 14697 5968 14855 5978
rect 14859 5968 14889 5978
rect 14893 5968 14923 5982
rect 14951 5968 14964 6006
rect 15036 6020 15065 6036
rect 15079 6020 15108 6036
rect 15123 6026 15153 6042
rect 15181 6020 15187 6068
rect 15190 6062 15209 6068
rect 15224 6062 15254 6070
rect 15190 6054 15254 6062
rect 15190 6038 15270 6054
rect 15286 6047 15348 6078
rect 15364 6047 15426 6078
rect 15495 6076 15544 6101
rect 15559 6076 15589 6092
rect 15458 6062 15488 6070
rect 15495 6068 15605 6076
rect 15458 6054 15503 6062
rect 15190 6036 15209 6038
rect 15224 6036 15270 6038
rect 15190 6020 15270 6036
rect 15297 6034 15332 6047
rect 15373 6044 15410 6047
rect 15373 6042 15415 6044
rect 15302 6031 15332 6034
rect 15311 6027 15318 6031
rect 15318 6026 15319 6027
rect 15277 6020 15287 6026
rect 15036 6012 15071 6020
rect 15036 5986 15037 6012
rect 15044 5986 15071 6012
rect 14979 5968 15009 5982
rect 15036 5978 15071 5986
rect 15073 6012 15114 6020
rect 15073 5986 15088 6012
rect 15095 5986 15114 6012
rect 15178 6008 15209 6020
rect 15224 6008 15327 6020
rect 15339 6010 15365 6036
rect 15380 6031 15410 6042
rect 15442 6038 15504 6054
rect 15442 6036 15488 6038
rect 15442 6020 15504 6036
rect 15516 6020 15522 6068
rect 15525 6060 15605 6068
rect 15525 6058 15544 6060
rect 15559 6058 15593 6060
rect 15525 6042 15605 6058
rect 15525 6020 15544 6042
rect 15559 6026 15589 6042
rect 15617 6036 15623 6110
rect 15626 6036 15645 6180
rect 15660 6036 15666 6180
rect 15675 6110 15688 6180
rect 15740 6176 15762 6180
rect 15733 6154 15762 6168
rect 15815 6154 15831 6168
rect 15869 6164 15875 6166
rect 15882 6164 15990 6180
rect 15997 6164 16003 6166
rect 16011 6164 16026 6180
rect 16092 6174 16111 6177
rect 15733 6152 15831 6154
rect 15858 6152 16026 6164
rect 16041 6154 16057 6168
rect 16092 6155 16114 6174
rect 16124 6168 16140 6169
rect 16123 6166 16140 6168
rect 16124 6161 16140 6166
rect 16114 6154 16120 6155
rect 16123 6154 16152 6161
rect 16041 6153 16152 6154
rect 16041 6152 16158 6153
rect 15717 6144 15768 6152
rect 15815 6144 15849 6152
rect 15717 6132 15742 6144
rect 15749 6132 15768 6144
rect 15822 6142 15849 6144
rect 15858 6142 16079 6152
rect 16114 6149 16120 6152
rect 15822 6138 16079 6142
rect 15717 6124 15768 6132
rect 15815 6124 16079 6138
rect 16123 6144 16158 6152
rect 15669 6076 15688 6110
rect 15733 6116 15762 6124
rect 15733 6110 15750 6116
rect 15733 6108 15767 6110
rect 15815 6108 15831 6124
rect 15832 6114 16040 6124
rect 16041 6114 16057 6124
rect 16105 6120 16120 6135
rect 16123 6132 16124 6144
rect 16131 6132 16158 6144
rect 16123 6124 16158 6132
rect 16123 6123 16152 6124
rect 15843 6110 16057 6114
rect 15858 6108 16057 6110
rect 16092 6110 16105 6120
rect 16123 6110 16140 6123
rect 16092 6108 16140 6110
rect 15734 6104 15767 6108
rect 15730 6102 15767 6104
rect 15730 6101 15797 6102
rect 15730 6096 15761 6101
rect 15767 6096 15797 6101
rect 15730 6092 15797 6096
rect 15703 6089 15797 6092
rect 15703 6082 15752 6089
rect 15703 6076 15733 6082
rect 15752 6077 15757 6082
rect 15669 6060 15749 6076
rect 15761 6068 15797 6089
rect 15858 6084 16047 6108
rect 16092 6107 16139 6108
rect 16105 6102 16139 6107
rect 15873 6081 16047 6084
rect 15866 6078 16047 6081
rect 16075 6101 16139 6102
rect 15669 6058 15688 6060
rect 15703 6058 15737 6060
rect 15669 6042 15749 6058
rect 15669 6036 15688 6042
rect 15385 6010 15488 6020
rect 15339 6008 15488 6010
rect 15509 6008 15544 6020
rect 15178 6006 15340 6008
rect 15190 5986 15209 6006
rect 15224 6004 15254 6006
rect 15073 5978 15114 5986
rect 15196 5982 15209 5986
rect 15261 5990 15340 6006
rect 15372 6006 15544 6008
rect 15372 5990 15451 6006
rect 15458 6004 15488 6006
rect 15036 5968 15065 5978
rect 15079 5968 15108 5978
rect 15123 5968 15153 5982
rect 15196 5968 15239 5982
rect 15261 5978 15451 5990
rect 15516 5986 15522 6006
rect 15246 5968 15276 5978
rect 15277 5968 15435 5978
rect 15439 5968 15469 5978
rect 15473 5968 15503 5982
rect 15531 5968 15544 6006
rect 15616 6020 15645 6036
rect 15659 6020 15688 6036
rect 15703 6026 15733 6042
rect 15761 6020 15767 6068
rect 15770 6062 15789 6068
rect 15804 6062 15834 6070
rect 15770 6054 15834 6062
rect 15770 6038 15850 6054
rect 15866 6047 15928 6078
rect 15944 6047 16006 6078
rect 16075 6076 16124 6101
rect 16139 6076 16169 6092
rect 16038 6062 16068 6070
rect 16075 6068 16185 6076
rect 16038 6054 16083 6062
rect 15770 6036 15789 6038
rect 15804 6036 15850 6038
rect 15770 6020 15850 6036
rect 15877 6034 15912 6047
rect 15953 6044 15990 6047
rect 15953 6042 15995 6044
rect 15882 6031 15912 6034
rect 15891 6027 15898 6031
rect 15898 6026 15899 6027
rect 15857 6020 15867 6026
rect 15616 6012 15651 6020
rect 15616 5986 15617 6012
rect 15624 5986 15651 6012
rect 15559 5968 15589 5982
rect 15616 5978 15651 5986
rect 15653 6012 15694 6020
rect 15653 5986 15668 6012
rect 15675 5986 15694 6012
rect 15758 6008 15789 6020
rect 15804 6008 15907 6020
rect 15919 6010 15945 6036
rect 15960 6031 15990 6042
rect 16022 6038 16084 6054
rect 16022 6036 16068 6038
rect 16022 6020 16084 6036
rect 16096 6020 16102 6068
rect 16105 6060 16185 6068
rect 16105 6058 16124 6060
rect 16139 6058 16173 6060
rect 16105 6042 16185 6058
rect 16105 6020 16124 6042
rect 16139 6026 16169 6042
rect 16197 6036 16203 6110
rect 16206 6036 16225 6180
rect 16240 6036 16246 6180
rect 16255 6110 16268 6180
rect 16320 6176 16342 6180
rect 16313 6154 16342 6168
rect 16395 6154 16411 6168
rect 16449 6164 16455 6166
rect 16462 6164 16570 6180
rect 16577 6164 16583 6166
rect 16591 6164 16606 6180
rect 16672 6174 16691 6177
rect 16313 6152 16411 6154
rect 16438 6152 16606 6164
rect 16621 6154 16637 6168
rect 16672 6155 16694 6174
rect 16704 6168 16720 6169
rect 16703 6166 16720 6168
rect 16704 6161 16720 6166
rect 16694 6154 16700 6155
rect 16703 6154 16732 6161
rect 16621 6153 16732 6154
rect 16621 6152 16738 6153
rect 16297 6144 16348 6152
rect 16395 6144 16429 6152
rect 16297 6132 16322 6144
rect 16329 6132 16348 6144
rect 16402 6142 16429 6144
rect 16438 6142 16659 6152
rect 16694 6149 16700 6152
rect 16402 6138 16659 6142
rect 16297 6124 16348 6132
rect 16395 6124 16659 6138
rect 16703 6144 16738 6152
rect 16249 6076 16268 6110
rect 16313 6116 16342 6124
rect 16313 6110 16330 6116
rect 16313 6108 16347 6110
rect 16395 6108 16411 6124
rect 16412 6114 16620 6124
rect 16621 6114 16637 6124
rect 16685 6120 16700 6135
rect 16703 6132 16704 6144
rect 16711 6132 16738 6144
rect 16703 6124 16738 6132
rect 16703 6123 16732 6124
rect 16423 6110 16637 6114
rect 16438 6108 16637 6110
rect 16672 6110 16685 6120
rect 16703 6110 16720 6123
rect 16672 6108 16720 6110
rect 16314 6104 16347 6108
rect 16310 6102 16347 6104
rect 16310 6101 16377 6102
rect 16310 6096 16341 6101
rect 16347 6096 16377 6101
rect 16310 6092 16377 6096
rect 16283 6089 16377 6092
rect 16283 6082 16332 6089
rect 16283 6076 16313 6082
rect 16332 6077 16337 6082
rect 16249 6060 16329 6076
rect 16341 6068 16377 6089
rect 16438 6084 16627 6108
rect 16672 6107 16719 6108
rect 16685 6102 16719 6107
rect 16453 6081 16627 6084
rect 16446 6078 16627 6081
rect 16655 6101 16719 6102
rect 16249 6058 16268 6060
rect 16283 6058 16317 6060
rect 16249 6042 16329 6058
rect 16249 6036 16268 6042
rect 15965 6010 16068 6020
rect 15919 6008 16068 6010
rect 16089 6008 16124 6020
rect 15758 6006 15920 6008
rect 15770 5986 15789 6006
rect 15804 6004 15834 6006
rect 15653 5978 15694 5986
rect 15776 5982 15789 5986
rect 15841 5990 15920 6006
rect 15952 6006 16124 6008
rect 15952 5990 16031 6006
rect 16038 6004 16068 6006
rect 15616 5968 15645 5978
rect 15659 5968 15688 5978
rect 15703 5968 15733 5982
rect 15776 5968 15819 5982
rect 15841 5978 16031 5990
rect 16096 5986 16102 6006
rect 15826 5968 15856 5978
rect 15857 5968 16015 5978
rect 16019 5968 16049 5978
rect 16053 5968 16083 5982
rect 16111 5968 16124 6006
rect 16196 6020 16225 6036
rect 16239 6020 16268 6036
rect 16283 6026 16313 6042
rect 16341 6020 16347 6068
rect 16350 6062 16369 6068
rect 16384 6062 16414 6070
rect 16350 6054 16414 6062
rect 16350 6038 16430 6054
rect 16446 6047 16508 6078
rect 16524 6047 16586 6078
rect 16655 6076 16704 6101
rect 16719 6076 16749 6092
rect 16618 6062 16648 6070
rect 16655 6068 16765 6076
rect 16618 6054 16663 6062
rect 16350 6036 16369 6038
rect 16384 6036 16430 6038
rect 16350 6020 16430 6036
rect 16457 6034 16492 6047
rect 16533 6044 16570 6047
rect 16533 6042 16575 6044
rect 16462 6031 16492 6034
rect 16471 6027 16478 6031
rect 16478 6026 16479 6027
rect 16437 6020 16447 6026
rect 16196 6012 16231 6020
rect 16196 5986 16197 6012
rect 16204 5986 16231 6012
rect 16139 5968 16169 5982
rect 16196 5978 16231 5986
rect 16233 6012 16274 6020
rect 16233 5986 16248 6012
rect 16255 5986 16274 6012
rect 16338 6008 16369 6020
rect 16384 6008 16487 6020
rect 16499 6010 16525 6036
rect 16540 6031 16570 6042
rect 16602 6038 16664 6054
rect 16602 6036 16648 6038
rect 16602 6020 16664 6036
rect 16676 6020 16682 6068
rect 16685 6060 16765 6068
rect 16685 6058 16704 6060
rect 16719 6058 16753 6060
rect 16685 6042 16765 6058
rect 16685 6020 16704 6042
rect 16719 6026 16749 6042
rect 16777 6036 16783 6110
rect 16786 6036 16805 6180
rect 16820 6036 16826 6180
rect 16835 6110 16848 6180
rect 16900 6176 16922 6180
rect 16893 6154 16922 6168
rect 16975 6154 16991 6168
rect 17029 6164 17035 6166
rect 17042 6164 17150 6180
rect 17157 6164 17163 6166
rect 17171 6164 17186 6180
rect 17252 6174 17271 6177
rect 16893 6152 16991 6154
rect 17018 6152 17186 6164
rect 17201 6154 17217 6168
rect 17252 6155 17274 6174
rect 17284 6168 17300 6169
rect 17283 6166 17300 6168
rect 17284 6161 17300 6166
rect 17274 6154 17280 6155
rect 17283 6154 17312 6161
rect 17201 6153 17312 6154
rect 17201 6152 17318 6153
rect 16877 6144 16928 6152
rect 16975 6144 17009 6152
rect 16877 6132 16902 6144
rect 16909 6132 16928 6144
rect 16982 6142 17009 6144
rect 17018 6142 17239 6152
rect 17274 6149 17280 6152
rect 16982 6138 17239 6142
rect 16877 6124 16928 6132
rect 16975 6124 17239 6138
rect 17283 6144 17318 6152
rect 16829 6076 16848 6110
rect 16893 6116 16922 6124
rect 16893 6110 16910 6116
rect 16893 6108 16927 6110
rect 16975 6108 16991 6124
rect 16992 6114 17200 6124
rect 17201 6114 17217 6124
rect 17265 6120 17280 6135
rect 17283 6132 17284 6144
rect 17291 6132 17318 6144
rect 17283 6124 17318 6132
rect 17283 6123 17312 6124
rect 17003 6110 17217 6114
rect 17018 6108 17217 6110
rect 17252 6110 17265 6120
rect 17283 6110 17300 6123
rect 17252 6108 17300 6110
rect 16894 6104 16927 6108
rect 16890 6102 16927 6104
rect 16890 6101 16957 6102
rect 16890 6096 16921 6101
rect 16927 6096 16957 6101
rect 16890 6092 16957 6096
rect 16863 6089 16957 6092
rect 16863 6082 16912 6089
rect 16863 6076 16893 6082
rect 16912 6077 16917 6082
rect 16829 6060 16909 6076
rect 16921 6068 16957 6089
rect 17018 6084 17207 6108
rect 17252 6107 17299 6108
rect 17265 6102 17299 6107
rect 17033 6081 17207 6084
rect 17026 6078 17207 6081
rect 17235 6101 17299 6102
rect 16829 6058 16848 6060
rect 16863 6058 16897 6060
rect 16829 6042 16909 6058
rect 16829 6036 16848 6042
rect 16545 6010 16648 6020
rect 16499 6008 16648 6010
rect 16669 6008 16704 6020
rect 16338 6006 16500 6008
rect 16350 5986 16369 6006
rect 16384 6004 16414 6006
rect 16233 5978 16274 5986
rect 16356 5982 16369 5986
rect 16421 5990 16500 6006
rect 16532 6006 16704 6008
rect 16532 5990 16611 6006
rect 16618 6004 16648 6006
rect 16196 5968 16225 5978
rect 16239 5968 16268 5978
rect 16283 5968 16313 5982
rect 16356 5968 16399 5982
rect 16421 5978 16611 5990
rect 16676 5986 16682 6006
rect 16406 5968 16436 5978
rect 16437 5968 16595 5978
rect 16599 5968 16629 5978
rect 16633 5968 16663 5982
rect 16691 5968 16704 6006
rect 16776 6020 16805 6036
rect 16819 6020 16848 6036
rect 16863 6026 16893 6042
rect 16921 6020 16927 6068
rect 16930 6062 16949 6068
rect 16964 6062 16994 6070
rect 16930 6054 16994 6062
rect 16930 6038 17010 6054
rect 17026 6047 17088 6078
rect 17104 6047 17166 6078
rect 17235 6076 17284 6101
rect 17299 6076 17329 6092
rect 17198 6062 17228 6070
rect 17235 6068 17345 6076
rect 17198 6054 17243 6062
rect 16930 6036 16949 6038
rect 16964 6036 17010 6038
rect 16930 6020 17010 6036
rect 17037 6034 17072 6047
rect 17113 6044 17150 6047
rect 17113 6042 17155 6044
rect 17042 6031 17072 6034
rect 17051 6027 17058 6031
rect 17058 6026 17059 6027
rect 17017 6020 17027 6026
rect 16776 6012 16811 6020
rect 16776 5986 16777 6012
rect 16784 5986 16811 6012
rect 16719 5968 16749 5982
rect 16776 5978 16811 5986
rect 16813 6012 16854 6020
rect 16813 5986 16828 6012
rect 16835 5986 16854 6012
rect 16918 6008 16949 6020
rect 16964 6008 17067 6020
rect 17079 6010 17105 6036
rect 17120 6031 17150 6042
rect 17182 6038 17244 6054
rect 17182 6036 17228 6038
rect 17182 6020 17244 6036
rect 17256 6020 17262 6068
rect 17265 6060 17345 6068
rect 17265 6058 17284 6060
rect 17299 6058 17333 6060
rect 17265 6042 17345 6058
rect 17265 6020 17284 6042
rect 17299 6026 17329 6042
rect 17357 6036 17363 6110
rect 17366 6036 17385 6180
rect 17400 6036 17406 6180
rect 17415 6110 17428 6180
rect 17480 6176 17502 6180
rect 17473 6154 17502 6168
rect 17555 6154 17571 6168
rect 17609 6164 17615 6166
rect 17622 6164 17730 6180
rect 17737 6164 17743 6166
rect 17751 6164 17766 6180
rect 17832 6174 17851 6177
rect 17473 6152 17571 6154
rect 17598 6152 17766 6164
rect 17781 6154 17797 6168
rect 17832 6155 17854 6174
rect 17864 6168 17880 6169
rect 17863 6166 17880 6168
rect 17864 6161 17880 6166
rect 17854 6154 17860 6155
rect 17863 6154 17892 6161
rect 17781 6153 17892 6154
rect 17781 6152 17898 6153
rect 17457 6144 17508 6152
rect 17555 6144 17589 6152
rect 17457 6132 17482 6144
rect 17489 6132 17508 6144
rect 17562 6142 17589 6144
rect 17598 6142 17819 6152
rect 17854 6149 17860 6152
rect 17562 6138 17819 6142
rect 17457 6124 17508 6132
rect 17555 6124 17819 6138
rect 17863 6144 17898 6152
rect 17409 6076 17428 6110
rect 17473 6116 17502 6124
rect 17473 6110 17490 6116
rect 17473 6108 17507 6110
rect 17555 6108 17571 6124
rect 17572 6114 17780 6124
rect 17781 6114 17797 6124
rect 17845 6120 17860 6135
rect 17863 6132 17864 6144
rect 17871 6132 17898 6144
rect 17863 6124 17898 6132
rect 17863 6123 17892 6124
rect 17583 6110 17797 6114
rect 17598 6108 17797 6110
rect 17832 6110 17845 6120
rect 17863 6110 17880 6123
rect 17832 6108 17880 6110
rect 17474 6104 17507 6108
rect 17470 6102 17507 6104
rect 17470 6101 17537 6102
rect 17470 6096 17501 6101
rect 17507 6096 17537 6101
rect 17470 6092 17537 6096
rect 17443 6089 17537 6092
rect 17443 6082 17492 6089
rect 17443 6076 17473 6082
rect 17492 6077 17497 6082
rect 17409 6060 17489 6076
rect 17501 6068 17537 6089
rect 17598 6084 17787 6108
rect 17832 6107 17879 6108
rect 17845 6102 17879 6107
rect 17613 6081 17787 6084
rect 17606 6078 17787 6081
rect 17815 6101 17879 6102
rect 17409 6058 17428 6060
rect 17443 6058 17477 6060
rect 17409 6042 17489 6058
rect 17409 6036 17428 6042
rect 17125 6010 17228 6020
rect 17079 6008 17228 6010
rect 17249 6008 17284 6020
rect 16918 6006 17080 6008
rect 16930 5986 16949 6006
rect 16964 6004 16994 6006
rect 16813 5978 16854 5986
rect 16936 5982 16949 5986
rect 17001 5990 17080 6006
rect 17112 6006 17284 6008
rect 17112 5990 17191 6006
rect 17198 6004 17228 6006
rect 16776 5968 16805 5978
rect 16819 5968 16848 5978
rect 16863 5968 16893 5982
rect 16936 5968 16979 5982
rect 17001 5978 17191 5990
rect 17256 5986 17262 6006
rect 16986 5968 17016 5978
rect 17017 5968 17175 5978
rect 17179 5968 17209 5978
rect 17213 5968 17243 5982
rect 17271 5968 17284 6006
rect 17356 6020 17385 6036
rect 17399 6020 17428 6036
rect 17443 6026 17473 6042
rect 17501 6020 17507 6068
rect 17510 6062 17529 6068
rect 17544 6062 17574 6070
rect 17510 6054 17574 6062
rect 17510 6038 17590 6054
rect 17606 6047 17668 6078
rect 17684 6047 17746 6078
rect 17815 6076 17864 6101
rect 17879 6076 17909 6092
rect 17778 6062 17808 6070
rect 17815 6068 17925 6076
rect 17778 6054 17823 6062
rect 17510 6036 17529 6038
rect 17544 6036 17590 6038
rect 17510 6020 17590 6036
rect 17617 6034 17652 6047
rect 17693 6044 17730 6047
rect 17693 6042 17735 6044
rect 17622 6031 17652 6034
rect 17631 6027 17638 6031
rect 17638 6026 17639 6027
rect 17597 6020 17607 6026
rect 17356 6012 17391 6020
rect 17356 5986 17357 6012
rect 17364 5986 17391 6012
rect 17299 5968 17329 5982
rect 17356 5978 17391 5986
rect 17393 6012 17434 6020
rect 17393 5986 17408 6012
rect 17415 5986 17434 6012
rect 17498 6008 17529 6020
rect 17544 6008 17647 6020
rect 17659 6010 17685 6036
rect 17700 6031 17730 6042
rect 17762 6038 17824 6054
rect 17762 6036 17808 6038
rect 17762 6020 17824 6036
rect 17836 6020 17842 6068
rect 17845 6060 17925 6068
rect 17845 6058 17864 6060
rect 17879 6058 17913 6060
rect 17845 6042 17925 6058
rect 17845 6020 17864 6042
rect 17879 6026 17909 6042
rect 17937 6036 17943 6110
rect 17946 6036 17965 6180
rect 17980 6036 17986 6180
rect 17995 6110 18008 6180
rect 18060 6176 18082 6180
rect 18053 6154 18082 6168
rect 18135 6154 18151 6168
rect 18189 6164 18195 6166
rect 18202 6164 18310 6180
rect 18317 6164 18323 6166
rect 18331 6164 18346 6180
rect 18412 6174 18431 6177
rect 18053 6152 18151 6154
rect 18178 6152 18346 6164
rect 18361 6154 18377 6168
rect 18412 6155 18434 6174
rect 18444 6168 18460 6169
rect 18443 6166 18460 6168
rect 18444 6161 18460 6166
rect 18434 6154 18440 6155
rect 18443 6154 18472 6161
rect 18361 6153 18472 6154
rect 18361 6152 18478 6153
rect 18037 6144 18088 6152
rect 18135 6144 18169 6152
rect 18037 6132 18062 6144
rect 18069 6132 18088 6144
rect 18142 6142 18169 6144
rect 18178 6142 18399 6152
rect 18434 6149 18440 6152
rect 18142 6138 18399 6142
rect 18037 6124 18088 6132
rect 18135 6124 18399 6138
rect 18443 6144 18478 6152
rect 17989 6076 18008 6110
rect 18053 6116 18082 6124
rect 18053 6110 18070 6116
rect 18053 6108 18087 6110
rect 18135 6108 18151 6124
rect 18152 6114 18360 6124
rect 18361 6114 18377 6124
rect 18425 6120 18440 6135
rect 18443 6132 18444 6144
rect 18451 6132 18478 6144
rect 18443 6124 18478 6132
rect 18443 6123 18472 6124
rect 18163 6110 18377 6114
rect 18178 6108 18377 6110
rect 18412 6110 18425 6120
rect 18443 6110 18460 6123
rect 18412 6108 18460 6110
rect 18054 6104 18087 6108
rect 18050 6102 18087 6104
rect 18050 6101 18117 6102
rect 18050 6096 18081 6101
rect 18087 6096 18117 6101
rect 18050 6092 18117 6096
rect 18023 6089 18117 6092
rect 18023 6082 18072 6089
rect 18023 6076 18053 6082
rect 18072 6077 18077 6082
rect 17989 6060 18069 6076
rect 18081 6068 18117 6089
rect 18178 6084 18367 6108
rect 18412 6107 18459 6108
rect 18425 6102 18459 6107
rect 18193 6081 18367 6084
rect 18186 6078 18367 6081
rect 18395 6101 18459 6102
rect 17989 6058 18008 6060
rect 18023 6058 18057 6060
rect 17989 6042 18069 6058
rect 17989 6036 18008 6042
rect 17705 6010 17808 6020
rect 17659 6008 17808 6010
rect 17829 6008 17864 6020
rect 17498 6006 17660 6008
rect 17510 5986 17529 6006
rect 17544 6004 17574 6006
rect 17393 5978 17434 5986
rect 17516 5982 17529 5986
rect 17581 5990 17660 6006
rect 17692 6006 17864 6008
rect 17692 5990 17771 6006
rect 17778 6004 17808 6006
rect 17356 5968 17385 5978
rect 17399 5968 17428 5978
rect 17443 5968 17473 5982
rect 17516 5968 17559 5982
rect 17581 5978 17771 5990
rect 17836 5986 17842 6006
rect 17566 5968 17596 5978
rect 17597 5968 17755 5978
rect 17759 5968 17789 5978
rect 17793 5968 17823 5982
rect 17851 5968 17864 6006
rect 17936 6020 17965 6036
rect 17979 6020 18008 6036
rect 18023 6026 18053 6042
rect 18081 6020 18087 6068
rect 18090 6062 18109 6068
rect 18124 6062 18154 6070
rect 18090 6054 18154 6062
rect 18090 6038 18170 6054
rect 18186 6047 18248 6078
rect 18264 6047 18326 6078
rect 18395 6076 18444 6101
rect 18459 6076 18489 6092
rect 18358 6062 18388 6070
rect 18395 6068 18505 6076
rect 18358 6054 18403 6062
rect 18090 6036 18109 6038
rect 18124 6036 18170 6038
rect 18090 6020 18170 6036
rect 18197 6034 18232 6047
rect 18273 6044 18310 6047
rect 18273 6042 18315 6044
rect 18202 6031 18232 6034
rect 18211 6027 18218 6031
rect 18218 6026 18219 6027
rect 18177 6020 18187 6026
rect 17936 6012 17971 6020
rect 17936 5986 17937 6012
rect 17944 5986 17971 6012
rect 17879 5968 17909 5982
rect 17936 5978 17971 5986
rect 17973 6012 18014 6020
rect 17973 5986 17988 6012
rect 17995 5986 18014 6012
rect 18078 6008 18109 6020
rect 18124 6008 18227 6020
rect 18239 6010 18265 6036
rect 18280 6031 18310 6042
rect 18342 6038 18404 6054
rect 18342 6036 18388 6038
rect 18342 6020 18404 6036
rect 18416 6020 18422 6068
rect 18425 6060 18505 6068
rect 18425 6058 18444 6060
rect 18459 6058 18493 6060
rect 18425 6042 18505 6058
rect 18425 6020 18444 6042
rect 18459 6026 18489 6042
rect 18517 6036 18523 6110
rect 18532 6036 18545 6180
rect 18285 6010 18388 6020
rect 18239 6008 18388 6010
rect 18409 6008 18444 6020
rect 18078 6006 18240 6008
rect 18090 5986 18109 6006
rect 18124 6004 18154 6006
rect 17973 5978 18014 5986
rect 18096 5982 18109 5986
rect 18161 5990 18240 6006
rect 18272 6006 18444 6008
rect 18272 5990 18351 6006
rect 18358 6004 18388 6006
rect 17936 5968 17965 5978
rect 17979 5968 18008 5978
rect 18023 5968 18053 5982
rect 18096 5968 18139 5982
rect 18161 5978 18351 5990
rect 18416 5986 18422 6006
rect 18146 5968 18176 5978
rect 18177 5968 18335 5978
rect 18339 5968 18369 5978
rect 18373 5968 18403 5982
rect 18431 5968 18444 6006
rect 18516 6020 18545 6036
rect 18516 6012 18551 6020
rect 18516 5986 18517 6012
rect 18524 5986 18551 6012
rect 18459 5968 18489 5982
rect 18516 5978 18551 5986
rect 18516 5968 18545 5978
rect -1 5962 18545 5968
rect 0 5954 18545 5962
rect 15 5924 28 5954
rect 43 5940 73 5954
rect 116 5940 159 5954
rect 166 5940 386 5954
rect 393 5940 423 5954
rect 83 5926 98 5938
rect 117 5926 130 5940
rect 198 5936 351 5940
rect 80 5924 102 5926
rect 180 5924 372 5936
rect 451 5924 464 5954
rect 479 5940 509 5954
rect 546 5924 565 5954
rect 580 5924 586 5954
rect 595 5924 608 5954
rect 623 5940 653 5954
rect 696 5940 739 5954
rect 746 5940 966 5954
rect 973 5940 1003 5954
rect 663 5926 678 5938
rect 697 5926 710 5940
rect 778 5936 931 5940
rect 660 5924 682 5926
rect 760 5924 952 5936
rect 1031 5924 1044 5954
rect 1059 5940 1089 5954
rect 1126 5924 1145 5954
rect 1160 5924 1166 5954
rect 1175 5924 1188 5954
rect 1203 5940 1233 5954
rect 1276 5940 1319 5954
rect 1326 5940 1546 5954
rect 1553 5940 1583 5954
rect 1243 5926 1258 5938
rect 1277 5926 1290 5940
rect 1358 5936 1511 5940
rect 1240 5924 1262 5926
rect 1340 5924 1532 5936
rect 1611 5924 1624 5954
rect 1639 5940 1669 5954
rect 1706 5924 1725 5954
rect 1740 5924 1746 5954
rect 1755 5924 1768 5954
rect 1783 5940 1813 5954
rect 1856 5940 1899 5954
rect 1906 5940 2126 5954
rect 2133 5940 2163 5954
rect 1823 5926 1838 5938
rect 1857 5926 1870 5940
rect 1938 5936 2091 5940
rect 1820 5924 1842 5926
rect 1920 5924 2112 5936
rect 2191 5924 2204 5954
rect 2219 5940 2249 5954
rect 2286 5924 2305 5954
rect 2320 5924 2326 5954
rect 2335 5924 2348 5954
rect 2363 5940 2393 5954
rect 2436 5940 2479 5954
rect 2486 5940 2706 5954
rect 2713 5940 2743 5954
rect 2403 5926 2418 5938
rect 2437 5926 2450 5940
rect 2518 5936 2671 5940
rect 2400 5924 2422 5926
rect 2500 5924 2692 5936
rect 2771 5924 2784 5954
rect 2799 5940 2829 5954
rect 2866 5924 2885 5954
rect 2900 5924 2906 5954
rect 2915 5924 2928 5954
rect 2943 5940 2973 5954
rect 3016 5940 3059 5954
rect 3066 5940 3286 5954
rect 3293 5940 3323 5954
rect 2983 5926 2998 5938
rect 3017 5926 3030 5940
rect 3098 5936 3251 5940
rect 2980 5924 3002 5926
rect 3080 5924 3272 5936
rect 3351 5924 3364 5954
rect 3379 5940 3409 5954
rect 3446 5924 3465 5954
rect 3480 5924 3486 5954
rect 3495 5924 3508 5954
rect 3523 5940 3553 5954
rect 3596 5940 3639 5954
rect 3646 5940 3866 5954
rect 3873 5940 3903 5954
rect 3563 5926 3578 5938
rect 3597 5926 3610 5940
rect 3678 5936 3831 5940
rect 3560 5924 3582 5926
rect 3660 5924 3852 5936
rect 3931 5924 3944 5954
rect 3959 5940 3989 5954
rect 4026 5924 4045 5954
rect 4060 5924 4066 5954
rect 4075 5924 4088 5954
rect 4103 5940 4133 5954
rect 4176 5940 4219 5954
rect 4226 5940 4446 5954
rect 4453 5940 4483 5954
rect 4143 5926 4158 5938
rect 4177 5926 4190 5940
rect 4258 5936 4411 5940
rect 4140 5924 4162 5926
rect 4240 5924 4432 5936
rect 4511 5924 4524 5954
rect 4539 5940 4569 5954
rect 4606 5924 4625 5954
rect 4640 5924 4646 5954
rect 4655 5924 4668 5954
rect 4683 5940 4713 5954
rect 4756 5940 4799 5954
rect 4806 5940 5026 5954
rect 5033 5940 5063 5954
rect 4723 5926 4738 5938
rect 4757 5926 4770 5940
rect 4838 5936 4991 5940
rect 4720 5924 4742 5926
rect 4820 5924 5012 5936
rect 5091 5924 5104 5954
rect 5119 5940 5149 5954
rect 5186 5924 5205 5954
rect 5220 5924 5226 5954
rect 5235 5924 5248 5954
rect 5263 5940 5293 5954
rect 5336 5940 5379 5954
rect 5386 5940 5606 5954
rect 5613 5940 5643 5954
rect 5303 5926 5318 5938
rect 5337 5926 5350 5940
rect 5418 5936 5571 5940
rect 5300 5924 5322 5926
rect 5400 5924 5592 5936
rect 5671 5924 5684 5954
rect 5699 5940 5729 5954
rect 5766 5924 5785 5954
rect 5800 5924 5806 5954
rect 5815 5924 5828 5954
rect 5843 5940 5873 5954
rect 5916 5940 5959 5954
rect 5966 5940 6186 5954
rect 6193 5940 6223 5954
rect 5883 5926 5898 5938
rect 5917 5926 5930 5940
rect 5998 5936 6151 5940
rect 5880 5924 5902 5926
rect 5980 5924 6172 5936
rect 6251 5924 6264 5954
rect 6279 5940 6309 5954
rect 6346 5924 6365 5954
rect 6380 5924 6386 5954
rect 6395 5924 6408 5954
rect 6423 5940 6453 5954
rect 6496 5940 6539 5954
rect 6546 5940 6766 5954
rect 6773 5940 6803 5954
rect 6463 5926 6478 5938
rect 6497 5926 6510 5940
rect 6578 5936 6731 5940
rect 6460 5924 6482 5926
rect 6560 5924 6752 5936
rect 6831 5924 6844 5954
rect 6859 5940 6889 5954
rect 6926 5924 6945 5954
rect 6960 5924 6966 5954
rect 6975 5924 6988 5954
rect 7003 5940 7033 5954
rect 7076 5940 7119 5954
rect 7126 5940 7346 5954
rect 7353 5940 7383 5954
rect 7043 5926 7058 5938
rect 7077 5926 7090 5940
rect 7158 5936 7311 5940
rect 7040 5924 7062 5926
rect 7140 5924 7332 5936
rect 7411 5924 7424 5954
rect 7439 5940 7469 5954
rect 7506 5924 7525 5954
rect 7540 5924 7546 5954
rect 7555 5924 7568 5954
rect 7583 5940 7613 5954
rect 7656 5940 7699 5954
rect 7706 5940 7926 5954
rect 7933 5940 7963 5954
rect 7623 5926 7638 5938
rect 7657 5926 7670 5940
rect 7738 5936 7891 5940
rect 7620 5924 7642 5926
rect 7720 5924 7912 5936
rect 7991 5924 8004 5954
rect 8019 5940 8049 5954
rect 8086 5924 8105 5954
rect 8120 5924 8126 5954
rect 8135 5924 8148 5954
rect 8163 5940 8193 5954
rect 8236 5940 8279 5954
rect 8286 5940 8506 5954
rect 8513 5940 8543 5954
rect 8203 5926 8218 5938
rect 8237 5926 8250 5940
rect 8318 5936 8471 5940
rect 8200 5924 8222 5926
rect 8300 5924 8492 5936
rect 8571 5924 8584 5954
rect 8599 5940 8629 5954
rect 8666 5924 8685 5954
rect 8700 5924 8706 5954
rect 8715 5924 8728 5954
rect 8743 5940 8773 5954
rect 8816 5940 8859 5954
rect 8866 5940 9086 5954
rect 9093 5940 9123 5954
rect 8783 5926 8798 5938
rect 8817 5926 8830 5940
rect 8898 5936 9051 5940
rect 8780 5924 8802 5926
rect 8880 5924 9072 5936
rect 9151 5924 9164 5954
rect 9179 5940 9209 5954
rect 9246 5924 9265 5954
rect 9280 5924 9286 5954
rect 9295 5924 9308 5954
rect 9323 5940 9353 5954
rect 9396 5940 9439 5954
rect 9446 5940 9666 5954
rect 9673 5940 9703 5954
rect 9363 5926 9378 5938
rect 9397 5926 9410 5940
rect 9478 5936 9631 5940
rect 9360 5924 9382 5926
rect 9460 5924 9652 5936
rect 9731 5924 9744 5954
rect 9759 5940 9789 5954
rect 9826 5924 9845 5954
rect 9860 5924 9866 5954
rect 9875 5924 9888 5954
rect 9903 5940 9933 5954
rect 9976 5940 10019 5954
rect 10026 5940 10246 5954
rect 10253 5940 10283 5954
rect 9943 5926 9958 5938
rect 9977 5926 9990 5940
rect 10058 5936 10211 5940
rect 9940 5924 9962 5926
rect 10040 5924 10232 5936
rect 10311 5924 10324 5954
rect 10339 5940 10369 5954
rect 10406 5924 10425 5954
rect 10440 5924 10446 5954
rect 10455 5924 10468 5954
rect 10483 5940 10513 5954
rect 10556 5940 10599 5954
rect 10606 5940 10826 5954
rect 10833 5940 10863 5954
rect 10523 5926 10538 5938
rect 10557 5926 10570 5940
rect 10638 5936 10791 5940
rect 10520 5924 10542 5926
rect 10620 5924 10812 5936
rect 10891 5924 10904 5954
rect 10919 5940 10949 5954
rect 10986 5924 11005 5954
rect 11020 5924 11026 5954
rect 11035 5924 11048 5954
rect 11063 5940 11093 5954
rect 11136 5940 11179 5954
rect 11186 5940 11406 5954
rect 11413 5940 11443 5954
rect 11103 5926 11118 5938
rect 11137 5926 11150 5940
rect 11218 5936 11371 5940
rect 11100 5924 11122 5926
rect 11200 5924 11392 5936
rect 11471 5924 11484 5954
rect 11499 5940 11529 5954
rect 11566 5924 11585 5954
rect 11600 5924 11606 5954
rect 11615 5924 11628 5954
rect 11643 5940 11673 5954
rect 11716 5940 11759 5954
rect 11766 5940 11986 5954
rect 11993 5940 12023 5954
rect 11683 5926 11698 5938
rect 11717 5926 11730 5940
rect 11798 5936 11951 5940
rect 11680 5924 11702 5926
rect 11780 5924 11972 5936
rect 12051 5924 12064 5954
rect 12079 5940 12109 5954
rect 12146 5924 12165 5954
rect 12180 5924 12186 5954
rect 12195 5924 12208 5954
rect 12223 5940 12253 5954
rect 12296 5940 12339 5954
rect 12346 5940 12566 5954
rect 12573 5940 12603 5954
rect 12263 5926 12278 5938
rect 12297 5926 12310 5940
rect 12378 5936 12531 5940
rect 12260 5924 12282 5926
rect 12360 5924 12552 5936
rect 12631 5924 12644 5954
rect 12659 5940 12689 5954
rect 12726 5924 12745 5954
rect 12760 5924 12766 5954
rect 12775 5924 12788 5954
rect 12803 5940 12833 5954
rect 12876 5940 12919 5954
rect 12926 5940 13146 5954
rect 13153 5940 13183 5954
rect 12843 5926 12858 5938
rect 12877 5926 12890 5940
rect 12958 5936 13111 5940
rect 12840 5924 12862 5926
rect 12940 5924 13132 5936
rect 13211 5924 13224 5954
rect 13239 5940 13269 5954
rect 13306 5924 13325 5954
rect 13340 5924 13346 5954
rect 13355 5924 13368 5954
rect 13383 5940 13413 5954
rect 13456 5940 13499 5954
rect 13506 5940 13726 5954
rect 13733 5940 13763 5954
rect 13423 5926 13438 5938
rect 13457 5926 13470 5940
rect 13538 5936 13691 5940
rect 13420 5924 13442 5926
rect 13520 5924 13712 5936
rect 13791 5924 13804 5954
rect 13819 5940 13849 5954
rect 13886 5924 13905 5954
rect 13920 5924 13926 5954
rect 13935 5924 13948 5954
rect 13963 5940 13993 5954
rect 14036 5940 14079 5954
rect 14086 5940 14306 5954
rect 14313 5940 14343 5954
rect 14003 5926 14018 5938
rect 14037 5926 14050 5940
rect 14118 5936 14271 5940
rect 14000 5924 14022 5926
rect 14100 5924 14292 5936
rect 14371 5924 14384 5954
rect 14399 5940 14429 5954
rect 14466 5924 14485 5954
rect 14500 5924 14506 5954
rect 14515 5924 14528 5954
rect 14543 5940 14573 5954
rect 14616 5940 14659 5954
rect 14666 5940 14886 5954
rect 14893 5940 14923 5954
rect 14583 5926 14598 5938
rect 14617 5926 14630 5940
rect 14698 5936 14851 5940
rect 14580 5924 14602 5926
rect 14680 5924 14872 5936
rect 14951 5924 14964 5954
rect 14979 5940 15009 5954
rect 15046 5924 15065 5954
rect 15080 5924 15086 5954
rect 15095 5924 15108 5954
rect 15123 5940 15153 5954
rect 15196 5940 15239 5954
rect 15246 5940 15466 5954
rect 15473 5940 15503 5954
rect 15163 5926 15178 5938
rect 15197 5926 15210 5940
rect 15278 5936 15431 5940
rect 15160 5924 15182 5926
rect 15260 5924 15452 5936
rect 15531 5924 15544 5954
rect 15559 5940 15589 5954
rect 15626 5924 15645 5954
rect 15660 5924 15666 5954
rect 15675 5924 15688 5954
rect 15703 5940 15733 5954
rect 15776 5940 15819 5954
rect 15826 5940 16046 5954
rect 16053 5940 16083 5954
rect 15743 5926 15758 5938
rect 15777 5926 15790 5940
rect 15858 5936 16011 5940
rect 15740 5924 15762 5926
rect 15840 5924 16032 5936
rect 16111 5924 16124 5954
rect 16139 5940 16169 5954
rect 16206 5924 16225 5954
rect 16240 5924 16246 5954
rect 16255 5924 16268 5954
rect 16283 5940 16313 5954
rect 16356 5940 16399 5954
rect 16406 5940 16626 5954
rect 16633 5940 16663 5954
rect 16323 5926 16338 5938
rect 16357 5926 16370 5940
rect 16438 5936 16591 5940
rect 16320 5924 16342 5926
rect 16420 5924 16612 5936
rect 16691 5924 16704 5954
rect 16719 5940 16749 5954
rect 16786 5924 16805 5954
rect 16820 5924 16826 5954
rect 16835 5924 16848 5954
rect 16863 5940 16893 5954
rect 16936 5940 16979 5954
rect 16986 5940 17206 5954
rect 17213 5940 17243 5954
rect 16903 5926 16918 5938
rect 16937 5926 16950 5940
rect 17018 5936 17171 5940
rect 16900 5924 16922 5926
rect 17000 5924 17192 5936
rect 17271 5924 17284 5954
rect 17299 5940 17329 5954
rect 17366 5924 17385 5954
rect 17400 5924 17406 5954
rect 17415 5924 17428 5954
rect 17443 5940 17473 5954
rect 17516 5940 17559 5954
rect 17566 5940 17786 5954
rect 17793 5940 17823 5954
rect 17483 5926 17498 5938
rect 17517 5926 17530 5940
rect 17598 5936 17751 5940
rect 17480 5924 17502 5926
rect 17580 5924 17772 5936
rect 17851 5924 17864 5954
rect 17879 5940 17909 5954
rect 17946 5924 17965 5954
rect 17980 5924 17986 5954
rect 17995 5924 18008 5954
rect 18023 5940 18053 5954
rect 18096 5940 18139 5954
rect 18146 5940 18366 5954
rect 18373 5940 18403 5954
rect 18063 5926 18078 5938
rect 18097 5926 18110 5940
rect 18178 5936 18331 5940
rect 18060 5924 18082 5926
rect 18160 5924 18352 5936
rect 18431 5924 18444 5954
rect 18459 5940 18489 5954
rect 18532 5924 18545 5954
rect 0 5910 18545 5924
rect 15 5840 28 5910
rect 80 5906 102 5910
rect 73 5884 102 5898
rect 155 5884 171 5898
rect 209 5894 215 5896
rect 222 5894 330 5910
rect 337 5894 343 5896
rect 351 5894 366 5910
rect 432 5904 451 5907
rect 73 5882 171 5884
rect 198 5882 366 5894
rect 381 5884 397 5898
rect 432 5885 454 5904
rect 464 5898 480 5899
rect 463 5896 480 5898
rect 464 5891 480 5896
rect 454 5884 460 5885
rect 463 5884 492 5891
rect 381 5883 492 5884
rect 381 5882 498 5883
rect 57 5874 108 5882
rect 155 5874 189 5882
rect 57 5862 82 5874
rect 89 5862 108 5874
rect 162 5872 189 5874
rect 198 5872 419 5882
rect 454 5879 460 5882
rect 162 5868 419 5872
rect 57 5854 108 5862
rect 155 5854 419 5868
rect 463 5874 498 5882
rect 9 5806 28 5840
rect 73 5846 102 5854
rect 73 5840 90 5846
rect 73 5838 107 5840
rect 155 5838 171 5854
rect 172 5844 380 5854
rect 381 5844 397 5854
rect 445 5850 460 5865
rect 463 5862 464 5874
rect 471 5862 498 5874
rect 463 5854 498 5862
rect 463 5853 492 5854
rect 183 5840 397 5844
rect 198 5838 397 5840
rect 432 5840 445 5850
rect 463 5840 480 5853
rect 432 5838 480 5840
rect 74 5834 107 5838
rect 70 5832 107 5834
rect 70 5831 137 5832
rect 70 5826 101 5831
rect 107 5826 137 5831
rect 70 5822 137 5826
rect 43 5819 137 5822
rect 43 5812 92 5819
rect 43 5806 73 5812
rect 92 5807 97 5812
rect 9 5790 89 5806
rect 101 5798 137 5819
rect 198 5814 387 5838
rect 432 5837 479 5838
rect 445 5832 479 5837
rect 213 5811 387 5814
rect 206 5808 387 5811
rect 415 5831 479 5832
rect 9 5788 28 5790
rect 43 5788 77 5790
rect 9 5772 89 5788
rect 9 5766 28 5772
rect -1 5750 28 5766
rect 43 5756 73 5772
rect 101 5750 107 5798
rect 110 5792 129 5798
rect 144 5792 174 5800
rect 110 5784 174 5792
rect 110 5768 190 5784
rect 206 5777 268 5808
rect 284 5777 346 5808
rect 415 5806 464 5831
rect 479 5806 509 5822
rect 378 5792 408 5800
rect 415 5798 525 5806
rect 378 5784 423 5792
rect 110 5766 129 5768
rect 144 5766 190 5768
rect 110 5750 190 5766
rect 217 5764 252 5777
rect 293 5774 330 5777
rect 293 5772 335 5774
rect 222 5761 252 5764
rect 231 5757 238 5761
rect 238 5756 239 5757
rect 197 5750 207 5756
rect -7 5742 34 5750
rect -7 5716 8 5742
rect 15 5716 34 5742
rect 98 5738 129 5750
rect 144 5738 247 5750
rect 259 5740 285 5766
rect 300 5761 330 5772
rect 362 5768 424 5784
rect 362 5766 408 5768
rect 362 5750 424 5766
rect 436 5750 442 5798
rect 445 5790 525 5798
rect 445 5788 464 5790
rect 479 5788 513 5790
rect 445 5772 525 5788
rect 445 5750 464 5772
rect 479 5756 509 5772
rect 537 5766 543 5840
rect 546 5766 565 5910
rect 580 5766 586 5910
rect 595 5840 608 5910
rect 660 5906 682 5910
rect 653 5884 682 5898
rect 735 5884 751 5898
rect 789 5894 795 5896
rect 802 5894 910 5910
rect 917 5894 923 5896
rect 931 5894 946 5910
rect 1012 5904 1031 5907
rect 653 5882 751 5884
rect 778 5882 946 5894
rect 961 5884 977 5898
rect 1012 5885 1034 5904
rect 1044 5898 1060 5899
rect 1043 5896 1060 5898
rect 1044 5891 1060 5896
rect 1034 5884 1040 5885
rect 1043 5884 1072 5891
rect 961 5883 1072 5884
rect 961 5882 1078 5883
rect 637 5874 688 5882
rect 735 5874 769 5882
rect 637 5862 662 5874
rect 669 5862 688 5874
rect 742 5872 769 5874
rect 778 5872 999 5882
rect 1034 5879 1040 5882
rect 742 5868 999 5872
rect 637 5854 688 5862
rect 735 5854 999 5868
rect 1043 5874 1078 5882
rect 589 5806 608 5840
rect 653 5846 682 5854
rect 653 5840 670 5846
rect 653 5838 687 5840
rect 735 5838 751 5854
rect 752 5844 960 5854
rect 961 5844 977 5854
rect 1025 5850 1040 5865
rect 1043 5862 1044 5874
rect 1051 5862 1078 5874
rect 1043 5854 1078 5862
rect 1043 5853 1072 5854
rect 763 5840 977 5844
rect 778 5838 977 5840
rect 1012 5840 1025 5850
rect 1043 5840 1060 5853
rect 1012 5838 1060 5840
rect 654 5834 687 5838
rect 650 5832 687 5834
rect 650 5831 717 5832
rect 650 5826 681 5831
rect 687 5826 717 5831
rect 650 5822 717 5826
rect 623 5819 717 5822
rect 623 5812 672 5819
rect 623 5806 653 5812
rect 672 5807 677 5812
rect 589 5790 669 5806
rect 681 5798 717 5819
rect 778 5814 967 5838
rect 1012 5837 1059 5838
rect 1025 5832 1059 5837
rect 793 5811 967 5814
rect 786 5808 967 5811
rect 995 5831 1059 5832
rect 589 5788 608 5790
rect 623 5788 657 5790
rect 589 5772 669 5788
rect 589 5766 608 5772
rect 305 5740 408 5750
rect 259 5738 408 5740
rect 429 5738 464 5750
rect 98 5736 260 5738
rect 110 5716 129 5736
rect 144 5734 174 5736
rect -7 5708 34 5716
rect 116 5712 129 5716
rect 181 5720 260 5736
rect 292 5736 464 5738
rect 292 5720 371 5736
rect 378 5734 408 5736
rect -1 5698 28 5708
rect 43 5698 73 5712
rect 116 5698 159 5712
rect 181 5708 371 5720
rect 436 5716 442 5736
rect 166 5698 196 5708
rect 197 5698 355 5708
rect 359 5698 389 5708
rect 393 5698 423 5712
rect 451 5698 464 5736
rect 536 5750 565 5766
rect 579 5750 608 5766
rect 623 5756 653 5772
rect 681 5750 687 5798
rect 690 5792 709 5798
rect 724 5792 754 5800
rect 690 5784 754 5792
rect 690 5768 770 5784
rect 786 5777 848 5808
rect 864 5777 926 5808
rect 995 5806 1044 5831
rect 1059 5806 1089 5822
rect 958 5792 988 5800
rect 995 5798 1105 5806
rect 958 5784 1003 5792
rect 690 5766 709 5768
rect 724 5766 770 5768
rect 690 5750 770 5766
rect 797 5764 832 5777
rect 873 5774 910 5777
rect 873 5772 915 5774
rect 802 5761 832 5764
rect 811 5757 818 5761
rect 818 5756 819 5757
rect 777 5750 787 5756
rect 536 5742 571 5750
rect 536 5716 537 5742
rect 544 5716 571 5742
rect 479 5698 509 5712
rect 536 5708 571 5716
rect 573 5742 614 5750
rect 573 5716 588 5742
rect 595 5716 614 5742
rect 678 5738 709 5750
rect 724 5738 827 5750
rect 839 5740 865 5766
rect 880 5761 910 5772
rect 942 5768 1004 5784
rect 942 5766 988 5768
rect 942 5750 1004 5766
rect 1016 5750 1022 5798
rect 1025 5790 1105 5798
rect 1025 5788 1044 5790
rect 1059 5788 1093 5790
rect 1025 5772 1105 5788
rect 1025 5750 1044 5772
rect 1059 5756 1089 5772
rect 1117 5766 1123 5840
rect 1126 5766 1145 5910
rect 1160 5766 1166 5910
rect 1175 5840 1188 5910
rect 1240 5906 1262 5910
rect 1233 5884 1262 5898
rect 1315 5884 1331 5898
rect 1369 5894 1375 5896
rect 1382 5894 1490 5910
rect 1497 5894 1503 5896
rect 1511 5894 1526 5910
rect 1592 5904 1611 5907
rect 1233 5882 1331 5884
rect 1358 5882 1526 5894
rect 1541 5884 1557 5898
rect 1592 5885 1614 5904
rect 1624 5898 1640 5899
rect 1623 5896 1640 5898
rect 1624 5891 1640 5896
rect 1614 5884 1620 5885
rect 1623 5884 1652 5891
rect 1541 5883 1652 5884
rect 1541 5882 1658 5883
rect 1217 5874 1268 5882
rect 1315 5874 1349 5882
rect 1217 5862 1242 5874
rect 1249 5862 1268 5874
rect 1322 5872 1349 5874
rect 1358 5872 1579 5882
rect 1614 5879 1620 5882
rect 1322 5868 1579 5872
rect 1217 5854 1268 5862
rect 1315 5854 1579 5868
rect 1623 5874 1658 5882
rect 1169 5806 1188 5840
rect 1233 5846 1262 5854
rect 1233 5840 1250 5846
rect 1233 5838 1267 5840
rect 1315 5838 1331 5854
rect 1332 5844 1540 5854
rect 1541 5844 1557 5854
rect 1605 5850 1620 5865
rect 1623 5862 1624 5874
rect 1631 5862 1658 5874
rect 1623 5854 1658 5862
rect 1623 5853 1652 5854
rect 1343 5840 1557 5844
rect 1358 5838 1557 5840
rect 1592 5840 1605 5850
rect 1623 5840 1640 5853
rect 1592 5838 1640 5840
rect 1234 5834 1267 5838
rect 1230 5832 1267 5834
rect 1230 5831 1297 5832
rect 1230 5826 1261 5831
rect 1267 5826 1297 5831
rect 1230 5822 1297 5826
rect 1203 5819 1297 5822
rect 1203 5812 1252 5819
rect 1203 5806 1233 5812
rect 1252 5807 1257 5812
rect 1169 5790 1249 5806
rect 1261 5798 1297 5819
rect 1358 5814 1547 5838
rect 1592 5837 1639 5838
rect 1605 5832 1639 5837
rect 1373 5811 1547 5814
rect 1366 5808 1547 5811
rect 1575 5831 1639 5832
rect 1169 5788 1188 5790
rect 1203 5788 1237 5790
rect 1169 5772 1249 5788
rect 1169 5766 1188 5772
rect 885 5740 988 5750
rect 839 5738 988 5740
rect 1009 5738 1044 5750
rect 678 5736 840 5738
rect 690 5716 709 5736
rect 724 5734 754 5736
rect 573 5708 614 5716
rect 696 5712 709 5716
rect 761 5720 840 5736
rect 872 5736 1044 5738
rect 872 5720 951 5736
rect 958 5734 988 5736
rect 536 5698 565 5708
rect 579 5698 608 5708
rect 623 5698 653 5712
rect 696 5698 739 5712
rect 761 5708 951 5720
rect 1016 5716 1022 5736
rect 746 5698 776 5708
rect 777 5698 935 5708
rect 939 5698 969 5708
rect 973 5698 1003 5712
rect 1031 5698 1044 5736
rect 1116 5750 1145 5766
rect 1159 5750 1188 5766
rect 1203 5756 1233 5772
rect 1261 5750 1267 5798
rect 1270 5792 1289 5798
rect 1304 5792 1334 5800
rect 1270 5784 1334 5792
rect 1270 5768 1350 5784
rect 1366 5777 1428 5808
rect 1444 5777 1506 5808
rect 1575 5806 1624 5831
rect 1639 5806 1669 5822
rect 1538 5792 1568 5800
rect 1575 5798 1685 5806
rect 1538 5784 1583 5792
rect 1270 5766 1289 5768
rect 1304 5766 1350 5768
rect 1270 5750 1350 5766
rect 1377 5764 1412 5777
rect 1453 5774 1490 5777
rect 1453 5772 1495 5774
rect 1382 5761 1412 5764
rect 1391 5757 1398 5761
rect 1398 5756 1399 5757
rect 1357 5750 1367 5756
rect 1116 5742 1151 5750
rect 1116 5716 1117 5742
rect 1124 5716 1151 5742
rect 1059 5698 1089 5712
rect 1116 5708 1151 5716
rect 1153 5742 1194 5750
rect 1153 5716 1168 5742
rect 1175 5716 1194 5742
rect 1258 5738 1289 5750
rect 1304 5738 1407 5750
rect 1419 5740 1445 5766
rect 1460 5761 1490 5772
rect 1522 5768 1584 5784
rect 1522 5766 1568 5768
rect 1522 5750 1584 5766
rect 1596 5750 1602 5798
rect 1605 5790 1685 5798
rect 1605 5788 1624 5790
rect 1639 5788 1673 5790
rect 1605 5772 1685 5788
rect 1605 5750 1624 5772
rect 1639 5756 1669 5772
rect 1697 5766 1703 5840
rect 1706 5766 1725 5910
rect 1740 5766 1746 5910
rect 1755 5840 1768 5910
rect 1820 5906 1842 5910
rect 1813 5884 1842 5898
rect 1895 5884 1911 5898
rect 1949 5894 1955 5896
rect 1962 5894 2070 5910
rect 2077 5894 2083 5896
rect 2091 5894 2106 5910
rect 2172 5904 2191 5907
rect 1813 5882 1911 5884
rect 1938 5882 2106 5894
rect 2121 5884 2137 5898
rect 2172 5885 2194 5904
rect 2204 5898 2220 5899
rect 2203 5896 2220 5898
rect 2204 5891 2220 5896
rect 2194 5884 2200 5885
rect 2203 5884 2232 5891
rect 2121 5883 2232 5884
rect 2121 5882 2238 5883
rect 1797 5874 1848 5882
rect 1895 5874 1929 5882
rect 1797 5862 1822 5874
rect 1829 5862 1848 5874
rect 1902 5872 1929 5874
rect 1938 5872 2159 5882
rect 2194 5879 2200 5882
rect 1902 5868 2159 5872
rect 1797 5854 1848 5862
rect 1895 5854 2159 5868
rect 2203 5874 2238 5882
rect 1749 5806 1768 5840
rect 1813 5846 1842 5854
rect 1813 5840 1830 5846
rect 1813 5838 1847 5840
rect 1895 5838 1911 5854
rect 1912 5844 2120 5854
rect 2121 5844 2137 5854
rect 2185 5850 2200 5865
rect 2203 5862 2204 5874
rect 2211 5862 2238 5874
rect 2203 5854 2238 5862
rect 2203 5853 2232 5854
rect 1923 5840 2137 5844
rect 1938 5838 2137 5840
rect 2172 5840 2185 5850
rect 2203 5840 2220 5853
rect 2172 5838 2220 5840
rect 1814 5834 1847 5838
rect 1810 5832 1847 5834
rect 1810 5831 1877 5832
rect 1810 5826 1841 5831
rect 1847 5826 1877 5831
rect 1810 5822 1877 5826
rect 1783 5819 1877 5822
rect 1783 5812 1832 5819
rect 1783 5806 1813 5812
rect 1832 5807 1837 5812
rect 1749 5790 1829 5806
rect 1841 5798 1877 5819
rect 1938 5814 2127 5838
rect 2172 5837 2219 5838
rect 2185 5832 2219 5837
rect 1953 5811 2127 5814
rect 1946 5808 2127 5811
rect 2155 5831 2219 5832
rect 1749 5788 1768 5790
rect 1783 5788 1817 5790
rect 1749 5772 1829 5788
rect 1749 5766 1768 5772
rect 1465 5740 1568 5750
rect 1419 5738 1568 5740
rect 1589 5738 1624 5750
rect 1258 5736 1420 5738
rect 1270 5716 1289 5736
rect 1304 5734 1334 5736
rect 1153 5708 1194 5716
rect 1276 5712 1289 5716
rect 1341 5720 1420 5736
rect 1452 5736 1624 5738
rect 1452 5720 1531 5736
rect 1538 5734 1568 5736
rect 1116 5698 1145 5708
rect 1159 5698 1188 5708
rect 1203 5698 1233 5712
rect 1276 5698 1319 5712
rect 1341 5708 1531 5720
rect 1596 5716 1602 5736
rect 1326 5698 1356 5708
rect 1357 5698 1515 5708
rect 1519 5698 1549 5708
rect 1553 5698 1583 5712
rect 1611 5698 1624 5736
rect 1696 5750 1725 5766
rect 1739 5750 1768 5766
rect 1783 5756 1813 5772
rect 1841 5750 1847 5798
rect 1850 5792 1869 5798
rect 1884 5792 1914 5800
rect 1850 5784 1914 5792
rect 1850 5768 1930 5784
rect 1946 5777 2008 5808
rect 2024 5777 2086 5808
rect 2155 5806 2204 5831
rect 2219 5806 2249 5822
rect 2118 5792 2148 5800
rect 2155 5798 2265 5806
rect 2118 5784 2163 5792
rect 1850 5766 1869 5768
rect 1884 5766 1930 5768
rect 1850 5750 1930 5766
rect 1957 5764 1992 5777
rect 2033 5774 2070 5777
rect 2033 5772 2075 5774
rect 1962 5761 1992 5764
rect 1971 5757 1978 5761
rect 1978 5756 1979 5757
rect 1937 5750 1947 5756
rect 1696 5742 1731 5750
rect 1696 5716 1697 5742
rect 1704 5716 1731 5742
rect 1639 5698 1669 5712
rect 1696 5708 1731 5716
rect 1733 5742 1774 5750
rect 1733 5716 1748 5742
rect 1755 5716 1774 5742
rect 1838 5738 1869 5750
rect 1884 5738 1987 5750
rect 1999 5740 2025 5766
rect 2040 5761 2070 5772
rect 2102 5768 2164 5784
rect 2102 5766 2148 5768
rect 2102 5750 2164 5766
rect 2176 5750 2182 5798
rect 2185 5790 2265 5798
rect 2185 5788 2204 5790
rect 2219 5788 2253 5790
rect 2185 5772 2265 5788
rect 2185 5750 2204 5772
rect 2219 5756 2249 5772
rect 2277 5766 2283 5840
rect 2286 5766 2305 5910
rect 2320 5766 2326 5910
rect 2335 5840 2348 5910
rect 2400 5906 2422 5910
rect 2393 5884 2422 5898
rect 2475 5884 2491 5898
rect 2529 5894 2535 5896
rect 2542 5894 2650 5910
rect 2657 5894 2663 5896
rect 2671 5894 2686 5910
rect 2752 5904 2771 5907
rect 2393 5882 2491 5884
rect 2518 5882 2686 5894
rect 2701 5884 2717 5898
rect 2752 5885 2774 5904
rect 2784 5898 2800 5899
rect 2783 5896 2800 5898
rect 2784 5891 2800 5896
rect 2774 5884 2780 5885
rect 2783 5884 2812 5891
rect 2701 5883 2812 5884
rect 2701 5882 2818 5883
rect 2377 5874 2428 5882
rect 2475 5874 2509 5882
rect 2377 5862 2402 5874
rect 2409 5862 2428 5874
rect 2482 5872 2509 5874
rect 2518 5872 2739 5882
rect 2774 5879 2780 5882
rect 2482 5868 2739 5872
rect 2377 5854 2428 5862
rect 2475 5854 2739 5868
rect 2783 5874 2818 5882
rect 2329 5806 2348 5840
rect 2393 5846 2422 5854
rect 2393 5840 2410 5846
rect 2393 5838 2427 5840
rect 2475 5838 2491 5854
rect 2492 5844 2700 5854
rect 2701 5844 2717 5854
rect 2765 5850 2780 5865
rect 2783 5862 2784 5874
rect 2791 5862 2818 5874
rect 2783 5854 2818 5862
rect 2783 5853 2812 5854
rect 2503 5840 2717 5844
rect 2518 5838 2717 5840
rect 2752 5840 2765 5850
rect 2783 5840 2800 5853
rect 2752 5838 2800 5840
rect 2394 5834 2427 5838
rect 2390 5832 2427 5834
rect 2390 5831 2457 5832
rect 2390 5826 2421 5831
rect 2427 5826 2457 5831
rect 2390 5822 2457 5826
rect 2363 5819 2457 5822
rect 2363 5812 2412 5819
rect 2363 5806 2393 5812
rect 2412 5807 2417 5812
rect 2329 5790 2409 5806
rect 2421 5798 2457 5819
rect 2518 5814 2707 5838
rect 2752 5837 2799 5838
rect 2765 5832 2799 5837
rect 2533 5811 2707 5814
rect 2526 5808 2707 5811
rect 2735 5831 2799 5832
rect 2329 5788 2348 5790
rect 2363 5788 2397 5790
rect 2329 5772 2409 5788
rect 2329 5766 2348 5772
rect 2045 5740 2148 5750
rect 1999 5738 2148 5740
rect 2169 5738 2204 5750
rect 1838 5736 2000 5738
rect 1850 5716 1869 5736
rect 1884 5734 1914 5736
rect 1733 5708 1774 5716
rect 1856 5712 1869 5716
rect 1921 5720 2000 5736
rect 2032 5736 2204 5738
rect 2032 5720 2111 5736
rect 2118 5734 2148 5736
rect 1696 5698 1725 5708
rect 1739 5698 1768 5708
rect 1783 5698 1813 5712
rect 1856 5698 1899 5712
rect 1921 5708 2111 5720
rect 2176 5716 2182 5736
rect 1906 5698 1936 5708
rect 1937 5698 2095 5708
rect 2099 5698 2129 5708
rect 2133 5698 2163 5712
rect 2191 5698 2204 5736
rect 2276 5750 2305 5766
rect 2319 5750 2348 5766
rect 2363 5756 2393 5772
rect 2421 5750 2427 5798
rect 2430 5792 2449 5798
rect 2464 5792 2494 5800
rect 2430 5784 2494 5792
rect 2430 5768 2510 5784
rect 2526 5777 2588 5808
rect 2604 5777 2666 5808
rect 2735 5806 2784 5831
rect 2799 5806 2829 5822
rect 2698 5792 2728 5800
rect 2735 5798 2845 5806
rect 2698 5784 2743 5792
rect 2430 5766 2449 5768
rect 2464 5766 2510 5768
rect 2430 5750 2510 5766
rect 2537 5764 2572 5777
rect 2613 5774 2650 5777
rect 2613 5772 2655 5774
rect 2542 5761 2572 5764
rect 2551 5757 2558 5761
rect 2558 5756 2559 5757
rect 2517 5750 2527 5756
rect 2276 5742 2311 5750
rect 2276 5716 2277 5742
rect 2284 5716 2311 5742
rect 2219 5698 2249 5712
rect 2276 5708 2311 5716
rect 2313 5742 2354 5750
rect 2313 5716 2328 5742
rect 2335 5716 2354 5742
rect 2418 5738 2449 5750
rect 2464 5738 2567 5750
rect 2579 5740 2605 5766
rect 2620 5761 2650 5772
rect 2682 5768 2744 5784
rect 2682 5766 2728 5768
rect 2682 5750 2744 5766
rect 2756 5750 2762 5798
rect 2765 5790 2845 5798
rect 2765 5788 2784 5790
rect 2799 5788 2833 5790
rect 2765 5772 2845 5788
rect 2765 5750 2784 5772
rect 2799 5756 2829 5772
rect 2857 5766 2863 5840
rect 2866 5766 2885 5910
rect 2900 5766 2906 5910
rect 2915 5840 2928 5910
rect 2980 5906 3002 5910
rect 2973 5884 3002 5898
rect 3055 5884 3071 5898
rect 3109 5894 3115 5896
rect 3122 5894 3230 5910
rect 3237 5894 3243 5896
rect 3251 5894 3266 5910
rect 3332 5904 3351 5907
rect 2973 5882 3071 5884
rect 3098 5882 3266 5894
rect 3281 5884 3297 5898
rect 3332 5885 3354 5904
rect 3364 5898 3380 5899
rect 3363 5896 3380 5898
rect 3364 5891 3380 5896
rect 3354 5884 3360 5885
rect 3363 5884 3392 5891
rect 3281 5883 3392 5884
rect 3281 5882 3398 5883
rect 2957 5874 3008 5882
rect 3055 5874 3089 5882
rect 2957 5862 2982 5874
rect 2989 5862 3008 5874
rect 3062 5872 3089 5874
rect 3098 5872 3319 5882
rect 3354 5879 3360 5882
rect 3062 5868 3319 5872
rect 2957 5854 3008 5862
rect 3055 5854 3319 5868
rect 3363 5874 3398 5882
rect 2909 5806 2928 5840
rect 2973 5846 3002 5854
rect 2973 5840 2990 5846
rect 2973 5838 3007 5840
rect 3055 5838 3071 5854
rect 3072 5844 3280 5854
rect 3281 5844 3297 5854
rect 3345 5850 3360 5865
rect 3363 5862 3364 5874
rect 3371 5862 3398 5874
rect 3363 5854 3398 5862
rect 3363 5853 3392 5854
rect 3083 5840 3297 5844
rect 3098 5838 3297 5840
rect 3332 5840 3345 5850
rect 3363 5840 3380 5853
rect 3332 5838 3380 5840
rect 2974 5834 3007 5838
rect 2970 5832 3007 5834
rect 2970 5831 3037 5832
rect 2970 5826 3001 5831
rect 3007 5826 3037 5831
rect 2970 5822 3037 5826
rect 2943 5819 3037 5822
rect 2943 5812 2992 5819
rect 2943 5806 2973 5812
rect 2992 5807 2997 5812
rect 2909 5790 2989 5806
rect 3001 5798 3037 5819
rect 3098 5814 3287 5838
rect 3332 5837 3379 5838
rect 3345 5832 3379 5837
rect 3113 5811 3287 5814
rect 3106 5808 3287 5811
rect 3315 5831 3379 5832
rect 2909 5788 2928 5790
rect 2943 5788 2977 5790
rect 2909 5772 2989 5788
rect 2909 5766 2928 5772
rect 2625 5740 2728 5750
rect 2579 5738 2728 5740
rect 2749 5738 2784 5750
rect 2418 5736 2580 5738
rect 2430 5716 2449 5736
rect 2464 5734 2494 5736
rect 2313 5708 2354 5716
rect 2436 5712 2449 5716
rect 2501 5720 2580 5736
rect 2612 5736 2784 5738
rect 2612 5720 2691 5736
rect 2698 5734 2728 5736
rect 2276 5698 2305 5708
rect 2319 5698 2348 5708
rect 2363 5698 2393 5712
rect 2436 5698 2479 5712
rect 2501 5708 2691 5720
rect 2756 5716 2762 5736
rect 2486 5698 2516 5708
rect 2517 5698 2675 5708
rect 2679 5698 2709 5708
rect 2713 5698 2743 5712
rect 2771 5698 2784 5736
rect 2856 5750 2885 5766
rect 2899 5750 2928 5766
rect 2943 5756 2973 5772
rect 3001 5750 3007 5798
rect 3010 5792 3029 5798
rect 3044 5792 3074 5800
rect 3010 5784 3074 5792
rect 3010 5768 3090 5784
rect 3106 5777 3168 5808
rect 3184 5777 3246 5808
rect 3315 5806 3364 5831
rect 3379 5806 3409 5822
rect 3278 5792 3308 5800
rect 3315 5798 3425 5806
rect 3278 5784 3323 5792
rect 3010 5766 3029 5768
rect 3044 5766 3090 5768
rect 3010 5750 3090 5766
rect 3117 5764 3152 5777
rect 3193 5774 3230 5777
rect 3193 5772 3235 5774
rect 3122 5761 3152 5764
rect 3131 5757 3138 5761
rect 3138 5756 3139 5757
rect 3097 5750 3107 5756
rect 2856 5742 2891 5750
rect 2856 5716 2857 5742
rect 2864 5716 2891 5742
rect 2799 5698 2829 5712
rect 2856 5708 2891 5716
rect 2893 5742 2934 5750
rect 2893 5716 2908 5742
rect 2915 5716 2934 5742
rect 2998 5738 3029 5750
rect 3044 5738 3147 5750
rect 3159 5740 3185 5766
rect 3200 5761 3230 5772
rect 3262 5768 3324 5784
rect 3262 5766 3308 5768
rect 3262 5750 3324 5766
rect 3336 5750 3342 5798
rect 3345 5790 3425 5798
rect 3345 5788 3364 5790
rect 3379 5788 3413 5790
rect 3345 5772 3425 5788
rect 3345 5750 3364 5772
rect 3379 5756 3409 5772
rect 3437 5766 3443 5840
rect 3446 5766 3465 5910
rect 3480 5766 3486 5910
rect 3495 5840 3508 5910
rect 3560 5906 3582 5910
rect 3553 5884 3582 5898
rect 3635 5884 3651 5898
rect 3689 5894 3695 5896
rect 3702 5894 3810 5910
rect 3817 5894 3823 5896
rect 3831 5894 3846 5910
rect 3912 5904 3931 5907
rect 3553 5882 3651 5884
rect 3678 5882 3846 5894
rect 3861 5884 3877 5898
rect 3912 5885 3934 5904
rect 3944 5898 3960 5899
rect 3943 5896 3960 5898
rect 3944 5891 3960 5896
rect 3934 5884 3940 5885
rect 3943 5884 3972 5891
rect 3861 5883 3972 5884
rect 3861 5882 3978 5883
rect 3537 5874 3588 5882
rect 3635 5874 3669 5882
rect 3537 5862 3562 5874
rect 3569 5862 3588 5874
rect 3642 5872 3669 5874
rect 3678 5872 3899 5882
rect 3934 5879 3940 5882
rect 3642 5868 3899 5872
rect 3537 5854 3588 5862
rect 3635 5854 3899 5868
rect 3943 5874 3978 5882
rect 3489 5806 3508 5840
rect 3553 5846 3582 5854
rect 3553 5840 3570 5846
rect 3553 5838 3587 5840
rect 3635 5838 3651 5854
rect 3652 5844 3860 5854
rect 3861 5844 3877 5854
rect 3925 5850 3940 5865
rect 3943 5862 3944 5874
rect 3951 5862 3978 5874
rect 3943 5854 3978 5862
rect 3943 5853 3972 5854
rect 3663 5840 3877 5844
rect 3678 5838 3877 5840
rect 3912 5840 3925 5850
rect 3943 5840 3960 5853
rect 3912 5838 3960 5840
rect 3554 5834 3587 5838
rect 3550 5832 3587 5834
rect 3550 5831 3617 5832
rect 3550 5826 3581 5831
rect 3587 5826 3617 5831
rect 3550 5822 3617 5826
rect 3523 5819 3617 5822
rect 3523 5812 3572 5819
rect 3523 5806 3553 5812
rect 3572 5807 3577 5812
rect 3489 5790 3569 5806
rect 3581 5798 3617 5819
rect 3678 5814 3867 5838
rect 3912 5837 3959 5838
rect 3925 5832 3959 5837
rect 3693 5811 3867 5814
rect 3686 5808 3867 5811
rect 3895 5831 3959 5832
rect 3489 5788 3508 5790
rect 3523 5788 3557 5790
rect 3489 5772 3569 5788
rect 3489 5766 3508 5772
rect 3205 5740 3308 5750
rect 3159 5738 3308 5740
rect 3329 5738 3364 5750
rect 2998 5736 3160 5738
rect 3010 5716 3029 5736
rect 3044 5734 3074 5736
rect 2893 5708 2934 5716
rect 3016 5712 3029 5716
rect 3081 5720 3160 5736
rect 3192 5736 3364 5738
rect 3192 5720 3271 5736
rect 3278 5734 3308 5736
rect 2856 5698 2885 5708
rect 2899 5698 2928 5708
rect 2943 5698 2973 5712
rect 3016 5698 3059 5712
rect 3081 5708 3271 5720
rect 3336 5716 3342 5736
rect 3066 5698 3096 5708
rect 3097 5698 3255 5708
rect 3259 5698 3289 5708
rect 3293 5698 3323 5712
rect 3351 5698 3364 5736
rect 3436 5750 3465 5766
rect 3479 5750 3508 5766
rect 3523 5756 3553 5772
rect 3581 5750 3587 5798
rect 3590 5792 3609 5798
rect 3624 5792 3654 5800
rect 3590 5784 3654 5792
rect 3590 5768 3670 5784
rect 3686 5777 3748 5808
rect 3764 5777 3826 5808
rect 3895 5806 3944 5831
rect 3959 5806 3989 5822
rect 3858 5792 3888 5800
rect 3895 5798 4005 5806
rect 3858 5784 3903 5792
rect 3590 5766 3609 5768
rect 3624 5766 3670 5768
rect 3590 5750 3670 5766
rect 3697 5764 3732 5777
rect 3773 5774 3810 5777
rect 3773 5772 3815 5774
rect 3702 5761 3732 5764
rect 3711 5757 3718 5761
rect 3718 5756 3719 5757
rect 3677 5750 3687 5756
rect 3436 5742 3471 5750
rect 3436 5716 3437 5742
rect 3444 5716 3471 5742
rect 3379 5698 3409 5712
rect 3436 5708 3471 5716
rect 3473 5742 3514 5750
rect 3473 5716 3488 5742
rect 3495 5716 3514 5742
rect 3578 5738 3609 5750
rect 3624 5738 3727 5750
rect 3739 5740 3765 5766
rect 3780 5761 3810 5772
rect 3842 5768 3904 5784
rect 3842 5766 3888 5768
rect 3842 5750 3904 5766
rect 3916 5750 3922 5798
rect 3925 5790 4005 5798
rect 3925 5788 3944 5790
rect 3959 5788 3993 5790
rect 3925 5772 4005 5788
rect 3925 5750 3944 5772
rect 3959 5756 3989 5772
rect 4017 5766 4023 5840
rect 4026 5766 4045 5910
rect 4060 5766 4066 5910
rect 4075 5840 4088 5910
rect 4140 5906 4162 5910
rect 4133 5884 4162 5898
rect 4215 5884 4231 5898
rect 4269 5894 4275 5896
rect 4282 5894 4390 5910
rect 4397 5894 4403 5896
rect 4411 5894 4426 5910
rect 4492 5904 4511 5907
rect 4133 5882 4231 5884
rect 4258 5882 4426 5894
rect 4441 5884 4457 5898
rect 4492 5885 4514 5904
rect 4524 5898 4540 5899
rect 4523 5896 4540 5898
rect 4524 5891 4540 5896
rect 4514 5884 4520 5885
rect 4523 5884 4552 5891
rect 4441 5883 4552 5884
rect 4441 5882 4558 5883
rect 4117 5874 4168 5882
rect 4215 5874 4249 5882
rect 4117 5862 4142 5874
rect 4149 5862 4168 5874
rect 4222 5872 4249 5874
rect 4258 5872 4479 5882
rect 4514 5879 4520 5882
rect 4222 5868 4479 5872
rect 4117 5854 4168 5862
rect 4215 5854 4479 5868
rect 4523 5874 4558 5882
rect 4069 5806 4088 5840
rect 4133 5846 4162 5854
rect 4133 5840 4150 5846
rect 4133 5838 4167 5840
rect 4215 5838 4231 5854
rect 4232 5844 4440 5854
rect 4441 5844 4457 5854
rect 4505 5850 4520 5865
rect 4523 5862 4524 5874
rect 4531 5862 4558 5874
rect 4523 5854 4558 5862
rect 4523 5853 4552 5854
rect 4243 5840 4457 5844
rect 4258 5838 4457 5840
rect 4492 5840 4505 5850
rect 4523 5840 4540 5853
rect 4492 5838 4540 5840
rect 4134 5834 4167 5838
rect 4130 5832 4167 5834
rect 4130 5831 4197 5832
rect 4130 5826 4161 5831
rect 4167 5826 4197 5831
rect 4130 5822 4197 5826
rect 4103 5819 4197 5822
rect 4103 5812 4152 5819
rect 4103 5806 4133 5812
rect 4152 5807 4157 5812
rect 4069 5790 4149 5806
rect 4161 5798 4197 5819
rect 4258 5814 4447 5838
rect 4492 5837 4539 5838
rect 4505 5832 4539 5837
rect 4273 5811 4447 5814
rect 4266 5808 4447 5811
rect 4475 5831 4539 5832
rect 4069 5788 4088 5790
rect 4103 5788 4137 5790
rect 4069 5772 4149 5788
rect 4069 5766 4088 5772
rect 3785 5740 3888 5750
rect 3739 5738 3888 5740
rect 3909 5738 3944 5750
rect 3578 5736 3740 5738
rect 3590 5716 3609 5736
rect 3624 5734 3654 5736
rect 3473 5708 3514 5716
rect 3596 5712 3609 5716
rect 3661 5720 3740 5736
rect 3772 5736 3944 5738
rect 3772 5720 3851 5736
rect 3858 5734 3888 5736
rect 3436 5698 3465 5708
rect 3479 5698 3508 5708
rect 3523 5698 3553 5712
rect 3596 5698 3639 5712
rect 3661 5708 3851 5720
rect 3916 5716 3922 5736
rect 3646 5698 3676 5708
rect 3677 5698 3835 5708
rect 3839 5698 3869 5708
rect 3873 5698 3903 5712
rect 3931 5698 3944 5736
rect 4016 5750 4045 5766
rect 4059 5750 4088 5766
rect 4103 5756 4133 5772
rect 4161 5750 4167 5798
rect 4170 5792 4189 5798
rect 4204 5792 4234 5800
rect 4170 5784 4234 5792
rect 4170 5768 4250 5784
rect 4266 5777 4328 5808
rect 4344 5777 4406 5808
rect 4475 5806 4524 5831
rect 4539 5806 4569 5822
rect 4438 5792 4468 5800
rect 4475 5798 4585 5806
rect 4438 5784 4483 5792
rect 4170 5766 4189 5768
rect 4204 5766 4250 5768
rect 4170 5750 4250 5766
rect 4277 5764 4312 5777
rect 4353 5774 4390 5777
rect 4353 5772 4395 5774
rect 4282 5761 4312 5764
rect 4291 5757 4298 5761
rect 4298 5756 4299 5757
rect 4257 5750 4267 5756
rect 4016 5742 4051 5750
rect 4016 5716 4017 5742
rect 4024 5716 4051 5742
rect 3959 5698 3989 5712
rect 4016 5708 4051 5716
rect 4053 5742 4094 5750
rect 4053 5716 4068 5742
rect 4075 5716 4094 5742
rect 4158 5738 4189 5750
rect 4204 5738 4307 5750
rect 4319 5740 4345 5766
rect 4360 5761 4390 5772
rect 4422 5768 4484 5784
rect 4422 5766 4468 5768
rect 4422 5750 4484 5766
rect 4496 5750 4502 5798
rect 4505 5790 4585 5798
rect 4505 5788 4524 5790
rect 4539 5788 4573 5790
rect 4505 5772 4585 5788
rect 4505 5750 4524 5772
rect 4539 5756 4569 5772
rect 4597 5766 4603 5840
rect 4606 5766 4625 5910
rect 4640 5766 4646 5910
rect 4655 5840 4668 5910
rect 4720 5906 4742 5910
rect 4713 5884 4742 5898
rect 4795 5884 4811 5898
rect 4849 5894 4855 5896
rect 4862 5894 4970 5910
rect 4977 5894 4983 5896
rect 4991 5894 5006 5910
rect 5072 5904 5091 5907
rect 4713 5882 4811 5884
rect 4838 5882 5006 5894
rect 5021 5884 5037 5898
rect 5072 5885 5094 5904
rect 5104 5898 5120 5899
rect 5103 5896 5120 5898
rect 5104 5891 5120 5896
rect 5094 5884 5100 5885
rect 5103 5884 5132 5891
rect 5021 5883 5132 5884
rect 5021 5882 5138 5883
rect 4697 5874 4748 5882
rect 4795 5874 4829 5882
rect 4697 5862 4722 5874
rect 4729 5862 4748 5874
rect 4802 5872 4829 5874
rect 4838 5872 5059 5882
rect 5094 5879 5100 5882
rect 4802 5868 5059 5872
rect 4697 5854 4748 5862
rect 4795 5854 5059 5868
rect 5103 5874 5138 5882
rect 4649 5806 4668 5840
rect 4713 5846 4742 5854
rect 4713 5840 4730 5846
rect 4713 5838 4747 5840
rect 4795 5838 4811 5854
rect 4812 5844 5020 5854
rect 5021 5844 5037 5854
rect 5085 5850 5100 5865
rect 5103 5862 5104 5874
rect 5111 5862 5138 5874
rect 5103 5854 5138 5862
rect 5103 5853 5132 5854
rect 4823 5840 5037 5844
rect 4838 5838 5037 5840
rect 5072 5840 5085 5850
rect 5103 5840 5120 5853
rect 5072 5838 5120 5840
rect 4714 5834 4747 5838
rect 4710 5832 4747 5834
rect 4710 5831 4777 5832
rect 4710 5826 4741 5831
rect 4747 5826 4777 5831
rect 4710 5822 4777 5826
rect 4683 5819 4777 5822
rect 4683 5812 4732 5819
rect 4683 5806 4713 5812
rect 4732 5807 4737 5812
rect 4649 5790 4729 5806
rect 4741 5798 4777 5819
rect 4838 5814 5027 5838
rect 5072 5837 5119 5838
rect 5085 5832 5119 5837
rect 4853 5811 5027 5814
rect 4846 5808 5027 5811
rect 5055 5831 5119 5832
rect 4649 5788 4668 5790
rect 4683 5788 4717 5790
rect 4649 5772 4729 5788
rect 4649 5766 4668 5772
rect 4365 5740 4468 5750
rect 4319 5738 4468 5740
rect 4489 5738 4524 5750
rect 4158 5736 4320 5738
rect 4170 5716 4189 5736
rect 4204 5734 4234 5736
rect 4053 5708 4094 5716
rect 4176 5712 4189 5716
rect 4241 5720 4320 5736
rect 4352 5736 4524 5738
rect 4352 5720 4431 5736
rect 4438 5734 4468 5736
rect 4016 5698 4045 5708
rect 4059 5698 4088 5708
rect 4103 5698 4133 5712
rect 4176 5698 4219 5712
rect 4241 5708 4431 5720
rect 4496 5716 4502 5736
rect 4226 5698 4256 5708
rect 4257 5698 4415 5708
rect 4419 5698 4449 5708
rect 4453 5698 4483 5712
rect 4511 5698 4524 5736
rect 4596 5750 4625 5766
rect 4639 5750 4668 5766
rect 4683 5756 4713 5772
rect 4741 5750 4747 5798
rect 4750 5792 4769 5798
rect 4784 5792 4814 5800
rect 4750 5784 4814 5792
rect 4750 5768 4830 5784
rect 4846 5777 4908 5808
rect 4924 5777 4986 5808
rect 5055 5806 5104 5831
rect 5119 5806 5149 5822
rect 5018 5792 5048 5800
rect 5055 5798 5165 5806
rect 5018 5784 5063 5792
rect 4750 5766 4769 5768
rect 4784 5766 4830 5768
rect 4750 5750 4830 5766
rect 4857 5764 4892 5777
rect 4933 5774 4970 5777
rect 4933 5772 4975 5774
rect 4862 5761 4892 5764
rect 4871 5757 4878 5761
rect 4878 5756 4879 5757
rect 4837 5750 4847 5756
rect 4596 5742 4631 5750
rect 4596 5716 4597 5742
rect 4604 5716 4631 5742
rect 4539 5698 4569 5712
rect 4596 5708 4631 5716
rect 4633 5742 4674 5750
rect 4633 5716 4648 5742
rect 4655 5716 4674 5742
rect 4738 5738 4769 5750
rect 4784 5738 4887 5750
rect 4899 5740 4925 5766
rect 4940 5761 4970 5772
rect 5002 5768 5064 5784
rect 5002 5766 5048 5768
rect 5002 5750 5064 5766
rect 5076 5750 5082 5798
rect 5085 5790 5165 5798
rect 5085 5788 5104 5790
rect 5119 5788 5153 5790
rect 5085 5772 5165 5788
rect 5085 5750 5104 5772
rect 5119 5756 5149 5772
rect 5177 5766 5183 5840
rect 5186 5766 5205 5910
rect 5220 5766 5226 5910
rect 5235 5840 5248 5910
rect 5300 5906 5322 5910
rect 5293 5884 5322 5898
rect 5375 5884 5391 5898
rect 5429 5894 5435 5896
rect 5442 5894 5550 5910
rect 5557 5894 5563 5896
rect 5571 5894 5586 5910
rect 5652 5904 5671 5907
rect 5293 5882 5391 5884
rect 5418 5882 5586 5894
rect 5601 5884 5617 5898
rect 5652 5885 5674 5904
rect 5684 5898 5700 5899
rect 5683 5896 5700 5898
rect 5684 5891 5700 5896
rect 5674 5884 5680 5885
rect 5683 5884 5712 5891
rect 5601 5883 5712 5884
rect 5601 5882 5718 5883
rect 5277 5874 5328 5882
rect 5375 5874 5409 5882
rect 5277 5862 5302 5874
rect 5309 5862 5328 5874
rect 5382 5872 5409 5874
rect 5418 5872 5639 5882
rect 5674 5879 5680 5882
rect 5382 5868 5639 5872
rect 5277 5854 5328 5862
rect 5375 5854 5639 5868
rect 5683 5874 5718 5882
rect 5229 5806 5248 5840
rect 5293 5846 5322 5854
rect 5293 5840 5310 5846
rect 5293 5838 5327 5840
rect 5375 5838 5391 5854
rect 5392 5844 5600 5854
rect 5601 5844 5617 5854
rect 5665 5850 5680 5865
rect 5683 5862 5684 5874
rect 5691 5862 5718 5874
rect 5683 5854 5718 5862
rect 5683 5853 5712 5854
rect 5403 5840 5617 5844
rect 5418 5838 5617 5840
rect 5652 5840 5665 5850
rect 5683 5840 5700 5853
rect 5652 5838 5700 5840
rect 5294 5834 5327 5838
rect 5290 5832 5327 5834
rect 5290 5831 5357 5832
rect 5290 5826 5321 5831
rect 5327 5826 5357 5831
rect 5290 5822 5357 5826
rect 5263 5819 5357 5822
rect 5263 5812 5312 5819
rect 5263 5806 5293 5812
rect 5312 5807 5317 5812
rect 5229 5790 5309 5806
rect 5321 5798 5357 5819
rect 5418 5814 5607 5838
rect 5652 5837 5699 5838
rect 5665 5832 5699 5837
rect 5433 5811 5607 5814
rect 5426 5808 5607 5811
rect 5635 5831 5699 5832
rect 5229 5788 5248 5790
rect 5263 5788 5297 5790
rect 5229 5772 5309 5788
rect 5229 5766 5248 5772
rect 4945 5740 5048 5750
rect 4899 5738 5048 5740
rect 5069 5738 5104 5750
rect 4738 5736 4900 5738
rect 4750 5716 4769 5736
rect 4784 5734 4814 5736
rect 4633 5708 4674 5716
rect 4756 5712 4769 5716
rect 4821 5720 4900 5736
rect 4932 5736 5104 5738
rect 4932 5720 5011 5736
rect 5018 5734 5048 5736
rect 4596 5698 4625 5708
rect 4639 5698 4668 5708
rect 4683 5698 4713 5712
rect 4756 5698 4799 5712
rect 4821 5708 5011 5720
rect 5076 5716 5082 5736
rect 4806 5698 4836 5708
rect 4837 5698 4995 5708
rect 4999 5698 5029 5708
rect 5033 5698 5063 5712
rect 5091 5698 5104 5736
rect 5176 5750 5205 5766
rect 5219 5750 5248 5766
rect 5263 5756 5293 5772
rect 5321 5750 5327 5798
rect 5330 5792 5349 5798
rect 5364 5792 5394 5800
rect 5330 5784 5394 5792
rect 5330 5768 5410 5784
rect 5426 5777 5488 5808
rect 5504 5777 5566 5808
rect 5635 5806 5684 5831
rect 5699 5806 5729 5822
rect 5598 5792 5628 5800
rect 5635 5798 5745 5806
rect 5598 5784 5643 5792
rect 5330 5766 5349 5768
rect 5364 5766 5410 5768
rect 5330 5750 5410 5766
rect 5437 5764 5472 5777
rect 5513 5774 5550 5777
rect 5513 5772 5555 5774
rect 5442 5761 5472 5764
rect 5451 5757 5458 5761
rect 5458 5756 5459 5757
rect 5417 5750 5427 5756
rect 5176 5742 5211 5750
rect 5176 5716 5177 5742
rect 5184 5716 5211 5742
rect 5119 5698 5149 5712
rect 5176 5708 5211 5716
rect 5213 5742 5254 5750
rect 5213 5716 5228 5742
rect 5235 5716 5254 5742
rect 5318 5738 5349 5750
rect 5364 5738 5467 5750
rect 5479 5740 5505 5766
rect 5520 5761 5550 5772
rect 5582 5768 5644 5784
rect 5582 5766 5628 5768
rect 5582 5750 5644 5766
rect 5656 5750 5662 5798
rect 5665 5790 5745 5798
rect 5665 5788 5684 5790
rect 5699 5788 5733 5790
rect 5665 5772 5745 5788
rect 5665 5750 5684 5772
rect 5699 5756 5729 5772
rect 5757 5766 5763 5840
rect 5766 5766 5785 5910
rect 5800 5766 5806 5910
rect 5815 5840 5828 5910
rect 5880 5906 5902 5910
rect 5873 5884 5902 5898
rect 5955 5884 5971 5898
rect 6009 5894 6015 5896
rect 6022 5894 6130 5910
rect 6137 5894 6143 5896
rect 6151 5894 6166 5910
rect 6232 5904 6251 5907
rect 5873 5882 5971 5884
rect 5998 5882 6166 5894
rect 6181 5884 6197 5898
rect 6232 5885 6254 5904
rect 6264 5898 6280 5899
rect 6263 5896 6280 5898
rect 6264 5891 6280 5896
rect 6254 5884 6260 5885
rect 6263 5884 6292 5891
rect 6181 5883 6292 5884
rect 6181 5882 6298 5883
rect 5857 5874 5908 5882
rect 5955 5874 5989 5882
rect 5857 5862 5882 5874
rect 5889 5862 5908 5874
rect 5962 5872 5989 5874
rect 5998 5872 6219 5882
rect 6254 5879 6260 5882
rect 5962 5868 6219 5872
rect 5857 5854 5908 5862
rect 5955 5854 6219 5868
rect 6263 5874 6298 5882
rect 5809 5806 5828 5840
rect 5873 5846 5902 5854
rect 5873 5840 5890 5846
rect 5873 5838 5907 5840
rect 5955 5838 5971 5854
rect 5972 5844 6180 5854
rect 6181 5844 6197 5854
rect 6245 5850 6260 5865
rect 6263 5862 6264 5874
rect 6271 5862 6298 5874
rect 6263 5854 6298 5862
rect 6263 5853 6292 5854
rect 5983 5840 6197 5844
rect 5998 5838 6197 5840
rect 6232 5840 6245 5850
rect 6263 5840 6280 5853
rect 6232 5838 6280 5840
rect 5874 5834 5907 5838
rect 5870 5832 5907 5834
rect 5870 5831 5937 5832
rect 5870 5826 5901 5831
rect 5907 5826 5937 5831
rect 5870 5822 5937 5826
rect 5843 5819 5937 5822
rect 5843 5812 5892 5819
rect 5843 5806 5873 5812
rect 5892 5807 5897 5812
rect 5809 5790 5889 5806
rect 5901 5798 5937 5819
rect 5998 5814 6187 5838
rect 6232 5837 6279 5838
rect 6245 5832 6279 5837
rect 6013 5811 6187 5814
rect 6006 5808 6187 5811
rect 6215 5831 6279 5832
rect 5809 5788 5828 5790
rect 5843 5788 5877 5790
rect 5809 5772 5889 5788
rect 5809 5766 5828 5772
rect 5525 5740 5628 5750
rect 5479 5738 5628 5740
rect 5649 5738 5684 5750
rect 5318 5736 5480 5738
rect 5330 5716 5349 5736
rect 5364 5734 5394 5736
rect 5213 5708 5254 5716
rect 5336 5712 5349 5716
rect 5401 5720 5480 5736
rect 5512 5736 5684 5738
rect 5512 5720 5591 5736
rect 5598 5734 5628 5736
rect 5176 5698 5205 5708
rect 5219 5698 5248 5708
rect 5263 5698 5293 5712
rect 5336 5698 5379 5712
rect 5401 5708 5591 5720
rect 5656 5716 5662 5736
rect 5386 5698 5416 5708
rect 5417 5698 5575 5708
rect 5579 5698 5609 5708
rect 5613 5698 5643 5712
rect 5671 5698 5684 5736
rect 5756 5750 5785 5766
rect 5799 5750 5828 5766
rect 5843 5756 5873 5772
rect 5901 5750 5907 5798
rect 5910 5792 5929 5798
rect 5944 5792 5974 5800
rect 5910 5784 5974 5792
rect 5910 5768 5990 5784
rect 6006 5777 6068 5808
rect 6084 5777 6146 5808
rect 6215 5806 6264 5831
rect 6279 5806 6309 5822
rect 6178 5792 6208 5800
rect 6215 5798 6325 5806
rect 6178 5784 6223 5792
rect 5910 5766 5929 5768
rect 5944 5766 5990 5768
rect 5910 5750 5990 5766
rect 6017 5764 6052 5777
rect 6093 5774 6130 5777
rect 6093 5772 6135 5774
rect 6022 5761 6052 5764
rect 6031 5757 6038 5761
rect 6038 5756 6039 5757
rect 5997 5750 6007 5756
rect 5756 5742 5791 5750
rect 5756 5716 5757 5742
rect 5764 5716 5791 5742
rect 5699 5698 5729 5712
rect 5756 5708 5791 5716
rect 5793 5742 5834 5750
rect 5793 5716 5808 5742
rect 5815 5716 5834 5742
rect 5898 5738 5929 5750
rect 5944 5738 6047 5750
rect 6059 5740 6085 5766
rect 6100 5761 6130 5772
rect 6162 5768 6224 5784
rect 6162 5766 6208 5768
rect 6162 5750 6224 5766
rect 6236 5750 6242 5798
rect 6245 5790 6325 5798
rect 6245 5788 6264 5790
rect 6279 5788 6313 5790
rect 6245 5772 6325 5788
rect 6245 5750 6264 5772
rect 6279 5756 6309 5772
rect 6337 5766 6343 5840
rect 6346 5766 6365 5910
rect 6380 5766 6386 5910
rect 6395 5840 6408 5910
rect 6460 5906 6482 5910
rect 6453 5884 6482 5898
rect 6535 5884 6551 5898
rect 6589 5894 6595 5896
rect 6602 5894 6710 5910
rect 6717 5894 6723 5896
rect 6731 5894 6746 5910
rect 6812 5904 6831 5907
rect 6453 5882 6551 5884
rect 6578 5882 6746 5894
rect 6761 5884 6777 5898
rect 6812 5885 6834 5904
rect 6844 5898 6860 5899
rect 6843 5896 6860 5898
rect 6844 5891 6860 5896
rect 6834 5884 6840 5885
rect 6843 5884 6872 5891
rect 6761 5883 6872 5884
rect 6761 5882 6878 5883
rect 6437 5874 6488 5882
rect 6535 5874 6569 5882
rect 6437 5862 6462 5874
rect 6469 5862 6488 5874
rect 6542 5872 6569 5874
rect 6578 5872 6799 5882
rect 6834 5879 6840 5882
rect 6542 5868 6799 5872
rect 6437 5854 6488 5862
rect 6535 5854 6799 5868
rect 6843 5874 6878 5882
rect 6389 5806 6408 5840
rect 6453 5846 6482 5854
rect 6453 5840 6470 5846
rect 6453 5838 6487 5840
rect 6535 5838 6551 5854
rect 6552 5844 6760 5854
rect 6761 5844 6777 5854
rect 6825 5850 6840 5865
rect 6843 5862 6844 5874
rect 6851 5862 6878 5874
rect 6843 5854 6878 5862
rect 6843 5853 6872 5854
rect 6563 5840 6777 5844
rect 6578 5838 6777 5840
rect 6812 5840 6825 5850
rect 6843 5840 6860 5853
rect 6812 5838 6860 5840
rect 6454 5834 6487 5838
rect 6450 5832 6487 5834
rect 6450 5831 6517 5832
rect 6450 5826 6481 5831
rect 6487 5826 6517 5831
rect 6450 5822 6517 5826
rect 6423 5819 6517 5822
rect 6423 5812 6472 5819
rect 6423 5806 6453 5812
rect 6472 5807 6477 5812
rect 6389 5790 6469 5806
rect 6481 5798 6517 5819
rect 6578 5814 6767 5838
rect 6812 5837 6859 5838
rect 6825 5832 6859 5837
rect 6593 5811 6767 5814
rect 6586 5808 6767 5811
rect 6795 5831 6859 5832
rect 6389 5788 6408 5790
rect 6423 5788 6457 5790
rect 6389 5772 6469 5788
rect 6389 5766 6408 5772
rect 6105 5740 6208 5750
rect 6059 5738 6208 5740
rect 6229 5738 6264 5750
rect 5898 5736 6060 5738
rect 5910 5716 5929 5736
rect 5944 5734 5974 5736
rect 5793 5708 5834 5716
rect 5916 5712 5929 5716
rect 5981 5720 6060 5736
rect 6092 5736 6264 5738
rect 6092 5720 6171 5736
rect 6178 5734 6208 5736
rect 5756 5698 5785 5708
rect 5799 5698 5828 5708
rect 5843 5698 5873 5712
rect 5916 5698 5959 5712
rect 5981 5708 6171 5720
rect 6236 5716 6242 5736
rect 5966 5698 5996 5708
rect 5997 5698 6155 5708
rect 6159 5698 6189 5708
rect 6193 5698 6223 5712
rect 6251 5698 6264 5736
rect 6336 5750 6365 5766
rect 6379 5750 6408 5766
rect 6423 5756 6453 5772
rect 6481 5750 6487 5798
rect 6490 5792 6509 5798
rect 6524 5792 6554 5800
rect 6490 5784 6554 5792
rect 6490 5768 6570 5784
rect 6586 5777 6648 5808
rect 6664 5777 6726 5808
rect 6795 5806 6844 5831
rect 6859 5806 6889 5822
rect 6758 5792 6788 5800
rect 6795 5798 6905 5806
rect 6758 5784 6803 5792
rect 6490 5766 6509 5768
rect 6524 5766 6570 5768
rect 6490 5750 6570 5766
rect 6597 5764 6632 5777
rect 6673 5774 6710 5777
rect 6673 5772 6715 5774
rect 6602 5761 6632 5764
rect 6611 5757 6618 5761
rect 6618 5756 6619 5757
rect 6577 5750 6587 5756
rect 6336 5742 6371 5750
rect 6336 5716 6337 5742
rect 6344 5716 6371 5742
rect 6279 5698 6309 5712
rect 6336 5708 6371 5716
rect 6373 5742 6414 5750
rect 6373 5716 6388 5742
rect 6395 5716 6414 5742
rect 6478 5738 6509 5750
rect 6524 5738 6627 5750
rect 6639 5740 6665 5766
rect 6680 5761 6710 5772
rect 6742 5768 6804 5784
rect 6742 5766 6788 5768
rect 6742 5750 6804 5766
rect 6816 5750 6822 5798
rect 6825 5790 6905 5798
rect 6825 5788 6844 5790
rect 6859 5788 6893 5790
rect 6825 5772 6905 5788
rect 6825 5750 6844 5772
rect 6859 5756 6889 5772
rect 6917 5766 6923 5840
rect 6926 5766 6945 5910
rect 6960 5766 6966 5910
rect 6975 5840 6988 5910
rect 7040 5906 7062 5910
rect 7033 5884 7062 5898
rect 7115 5884 7131 5898
rect 7169 5894 7175 5896
rect 7182 5894 7290 5910
rect 7297 5894 7303 5896
rect 7311 5894 7326 5910
rect 7392 5904 7411 5907
rect 7033 5882 7131 5884
rect 7158 5882 7326 5894
rect 7341 5884 7357 5898
rect 7392 5885 7414 5904
rect 7424 5898 7440 5899
rect 7423 5896 7440 5898
rect 7424 5891 7440 5896
rect 7414 5884 7420 5885
rect 7423 5884 7452 5891
rect 7341 5883 7452 5884
rect 7341 5882 7458 5883
rect 7017 5874 7068 5882
rect 7115 5874 7149 5882
rect 7017 5862 7042 5874
rect 7049 5862 7068 5874
rect 7122 5872 7149 5874
rect 7158 5872 7379 5882
rect 7414 5879 7420 5882
rect 7122 5868 7379 5872
rect 7017 5854 7068 5862
rect 7115 5854 7379 5868
rect 7423 5874 7458 5882
rect 6969 5806 6988 5840
rect 7033 5846 7062 5854
rect 7033 5840 7050 5846
rect 7033 5838 7067 5840
rect 7115 5838 7131 5854
rect 7132 5844 7340 5854
rect 7341 5844 7357 5854
rect 7405 5850 7420 5865
rect 7423 5862 7424 5874
rect 7431 5862 7458 5874
rect 7423 5854 7458 5862
rect 7423 5853 7452 5854
rect 7143 5840 7357 5844
rect 7158 5838 7357 5840
rect 7392 5840 7405 5850
rect 7423 5840 7440 5853
rect 7392 5838 7440 5840
rect 7034 5834 7067 5838
rect 7030 5832 7067 5834
rect 7030 5831 7097 5832
rect 7030 5826 7061 5831
rect 7067 5826 7097 5831
rect 7030 5822 7097 5826
rect 7003 5819 7097 5822
rect 7003 5812 7052 5819
rect 7003 5806 7033 5812
rect 7052 5807 7057 5812
rect 6969 5790 7049 5806
rect 7061 5798 7097 5819
rect 7158 5814 7347 5838
rect 7392 5837 7439 5838
rect 7405 5832 7439 5837
rect 7173 5811 7347 5814
rect 7166 5808 7347 5811
rect 7375 5831 7439 5832
rect 6969 5788 6988 5790
rect 7003 5788 7037 5790
rect 6969 5772 7049 5788
rect 6969 5766 6988 5772
rect 6685 5740 6788 5750
rect 6639 5738 6788 5740
rect 6809 5738 6844 5750
rect 6478 5736 6640 5738
rect 6490 5716 6509 5736
rect 6524 5734 6554 5736
rect 6373 5708 6414 5716
rect 6496 5712 6509 5716
rect 6561 5720 6640 5736
rect 6672 5736 6844 5738
rect 6672 5720 6751 5736
rect 6758 5734 6788 5736
rect 6336 5698 6365 5708
rect 6379 5698 6408 5708
rect 6423 5698 6453 5712
rect 6496 5698 6539 5712
rect 6561 5708 6751 5720
rect 6816 5716 6822 5736
rect 6546 5698 6576 5708
rect 6577 5698 6735 5708
rect 6739 5698 6769 5708
rect 6773 5698 6803 5712
rect 6831 5698 6844 5736
rect 6916 5750 6945 5766
rect 6959 5750 6988 5766
rect 7003 5756 7033 5772
rect 7061 5750 7067 5798
rect 7070 5792 7089 5798
rect 7104 5792 7134 5800
rect 7070 5784 7134 5792
rect 7070 5768 7150 5784
rect 7166 5777 7228 5808
rect 7244 5777 7306 5808
rect 7375 5806 7424 5831
rect 7439 5806 7469 5822
rect 7338 5792 7368 5800
rect 7375 5798 7485 5806
rect 7338 5784 7383 5792
rect 7070 5766 7089 5768
rect 7104 5766 7150 5768
rect 7070 5750 7150 5766
rect 7177 5764 7212 5777
rect 7253 5774 7290 5777
rect 7253 5772 7295 5774
rect 7182 5761 7212 5764
rect 7191 5757 7198 5761
rect 7198 5756 7199 5757
rect 7157 5750 7167 5756
rect 6916 5742 6951 5750
rect 6916 5716 6917 5742
rect 6924 5716 6951 5742
rect 6859 5698 6889 5712
rect 6916 5708 6951 5716
rect 6953 5742 6994 5750
rect 6953 5716 6968 5742
rect 6975 5716 6994 5742
rect 7058 5738 7089 5750
rect 7104 5738 7207 5750
rect 7219 5740 7245 5766
rect 7260 5761 7290 5772
rect 7322 5768 7384 5784
rect 7322 5766 7368 5768
rect 7322 5750 7384 5766
rect 7396 5750 7402 5798
rect 7405 5790 7485 5798
rect 7405 5788 7424 5790
rect 7439 5788 7473 5790
rect 7405 5772 7485 5788
rect 7405 5750 7424 5772
rect 7439 5756 7469 5772
rect 7497 5766 7503 5840
rect 7506 5766 7525 5910
rect 7540 5766 7546 5910
rect 7555 5840 7568 5910
rect 7620 5906 7642 5910
rect 7613 5884 7642 5898
rect 7695 5884 7711 5898
rect 7749 5894 7755 5896
rect 7762 5894 7870 5910
rect 7877 5894 7883 5896
rect 7891 5894 7906 5910
rect 7972 5904 7991 5907
rect 7613 5882 7711 5884
rect 7738 5882 7906 5894
rect 7921 5884 7937 5898
rect 7972 5885 7994 5904
rect 8004 5898 8020 5899
rect 8003 5896 8020 5898
rect 8004 5891 8020 5896
rect 7994 5884 8000 5885
rect 8003 5884 8032 5891
rect 7921 5883 8032 5884
rect 7921 5882 8038 5883
rect 7597 5874 7648 5882
rect 7695 5874 7729 5882
rect 7597 5862 7622 5874
rect 7629 5862 7648 5874
rect 7702 5872 7729 5874
rect 7738 5872 7959 5882
rect 7994 5879 8000 5882
rect 7702 5868 7959 5872
rect 7597 5854 7648 5862
rect 7695 5854 7959 5868
rect 8003 5874 8038 5882
rect 7549 5806 7568 5840
rect 7613 5846 7642 5854
rect 7613 5840 7630 5846
rect 7613 5838 7647 5840
rect 7695 5838 7711 5854
rect 7712 5844 7920 5854
rect 7921 5844 7937 5854
rect 7985 5850 8000 5865
rect 8003 5862 8004 5874
rect 8011 5862 8038 5874
rect 8003 5854 8038 5862
rect 8003 5853 8032 5854
rect 7723 5840 7937 5844
rect 7738 5838 7937 5840
rect 7972 5840 7985 5850
rect 8003 5840 8020 5853
rect 7972 5838 8020 5840
rect 7614 5834 7647 5838
rect 7610 5832 7647 5834
rect 7610 5831 7677 5832
rect 7610 5826 7641 5831
rect 7647 5826 7677 5831
rect 7610 5822 7677 5826
rect 7583 5819 7677 5822
rect 7583 5812 7632 5819
rect 7583 5806 7613 5812
rect 7632 5807 7637 5812
rect 7549 5790 7629 5806
rect 7641 5798 7677 5819
rect 7738 5814 7927 5838
rect 7972 5837 8019 5838
rect 7985 5832 8019 5837
rect 7753 5811 7927 5814
rect 7746 5808 7927 5811
rect 7955 5831 8019 5832
rect 7549 5788 7568 5790
rect 7583 5788 7617 5790
rect 7549 5772 7629 5788
rect 7549 5766 7568 5772
rect 7265 5740 7368 5750
rect 7219 5738 7368 5740
rect 7389 5738 7424 5750
rect 7058 5736 7220 5738
rect 7070 5716 7089 5736
rect 7104 5734 7134 5736
rect 6953 5708 6994 5716
rect 7076 5712 7089 5716
rect 7141 5720 7220 5736
rect 7252 5736 7424 5738
rect 7252 5720 7331 5736
rect 7338 5734 7368 5736
rect 6916 5698 6945 5708
rect 6959 5698 6988 5708
rect 7003 5698 7033 5712
rect 7076 5698 7119 5712
rect 7141 5708 7331 5720
rect 7396 5716 7402 5736
rect 7126 5698 7156 5708
rect 7157 5698 7315 5708
rect 7319 5698 7349 5708
rect 7353 5698 7383 5712
rect 7411 5698 7424 5736
rect 7496 5750 7525 5766
rect 7539 5750 7568 5766
rect 7583 5756 7613 5772
rect 7641 5750 7647 5798
rect 7650 5792 7669 5798
rect 7684 5792 7714 5800
rect 7650 5784 7714 5792
rect 7650 5768 7730 5784
rect 7746 5777 7808 5808
rect 7824 5777 7886 5808
rect 7955 5806 8004 5831
rect 8019 5806 8049 5822
rect 7918 5792 7948 5800
rect 7955 5798 8065 5806
rect 7918 5784 7963 5792
rect 7650 5766 7669 5768
rect 7684 5766 7730 5768
rect 7650 5750 7730 5766
rect 7757 5764 7792 5777
rect 7833 5774 7870 5777
rect 7833 5772 7875 5774
rect 7762 5761 7792 5764
rect 7771 5757 7778 5761
rect 7778 5756 7779 5757
rect 7737 5750 7747 5756
rect 7496 5742 7531 5750
rect 7496 5716 7497 5742
rect 7504 5716 7531 5742
rect 7439 5698 7469 5712
rect 7496 5708 7531 5716
rect 7533 5742 7574 5750
rect 7533 5716 7548 5742
rect 7555 5716 7574 5742
rect 7638 5738 7669 5750
rect 7684 5738 7787 5750
rect 7799 5740 7825 5766
rect 7840 5761 7870 5772
rect 7902 5768 7964 5784
rect 7902 5766 7948 5768
rect 7902 5750 7964 5766
rect 7976 5750 7982 5798
rect 7985 5790 8065 5798
rect 7985 5788 8004 5790
rect 8019 5788 8053 5790
rect 7985 5772 8065 5788
rect 7985 5750 8004 5772
rect 8019 5756 8049 5772
rect 8077 5766 8083 5840
rect 8086 5766 8105 5910
rect 8120 5766 8126 5910
rect 8135 5840 8148 5910
rect 8200 5906 8222 5910
rect 8193 5884 8222 5898
rect 8275 5884 8291 5898
rect 8329 5894 8335 5896
rect 8342 5894 8450 5910
rect 8457 5894 8463 5896
rect 8471 5894 8486 5910
rect 8552 5904 8571 5907
rect 8193 5882 8291 5884
rect 8318 5882 8486 5894
rect 8501 5884 8517 5898
rect 8552 5885 8574 5904
rect 8584 5898 8600 5899
rect 8583 5896 8600 5898
rect 8584 5891 8600 5896
rect 8574 5884 8580 5885
rect 8583 5884 8612 5891
rect 8501 5883 8612 5884
rect 8501 5882 8618 5883
rect 8177 5874 8228 5882
rect 8275 5874 8309 5882
rect 8177 5862 8202 5874
rect 8209 5862 8228 5874
rect 8282 5872 8309 5874
rect 8318 5872 8539 5882
rect 8574 5879 8580 5882
rect 8282 5868 8539 5872
rect 8177 5854 8228 5862
rect 8275 5854 8539 5868
rect 8583 5874 8618 5882
rect 8129 5806 8148 5840
rect 8193 5846 8222 5854
rect 8193 5840 8210 5846
rect 8193 5838 8227 5840
rect 8275 5838 8291 5854
rect 8292 5844 8500 5854
rect 8501 5844 8517 5854
rect 8565 5850 8580 5865
rect 8583 5862 8584 5874
rect 8591 5862 8618 5874
rect 8583 5854 8618 5862
rect 8583 5853 8612 5854
rect 8303 5840 8517 5844
rect 8318 5838 8517 5840
rect 8552 5840 8565 5850
rect 8583 5840 8600 5853
rect 8552 5838 8600 5840
rect 8194 5834 8227 5838
rect 8190 5832 8227 5834
rect 8190 5831 8257 5832
rect 8190 5826 8221 5831
rect 8227 5826 8257 5831
rect 8190 5822 8257 5826
rect 8163 5819 8257 5822
rect 8163 5812 8212 5819
rect 8163 5806 8193 5812
rect 8212 5807 8217 5812
rect 8129 5790 8209 5806
rect 8221 5798 8257 5819
rect 8318 5814 8507 5838
rect 8552 5837 8599 5838
rect 8565 5832 8599 5837
rect 8333 5811 8507 5814
rect 8326 5808 8507 5811
rect 8535 5831 8599 5832
rect 8129 5788 8148 5790
rect 8163 5788 8197 5790
rect 8129 5772 8209 5788
rect 8129 5766 8148 5772
rect 7845 5740 7948 5750
rect 7799 5738 7948 5740
rect 7969 5738 8004 5750
rect 7638 5736 7800 5738
rect 7650 5716 7669 5736
rect 7684 5734 7714 5736
rect 7533 5708 7574 5716
rect 7656 5712 7669 5716
rect 7721 5720 7800 5736
rect 7832 5736 8004 5738
rect 7832 5720 7911 5736
rect 7918 5734 7948 5736
rect 7496 5698 7525 5708
rect 7539 5698 7568 5708
rect 7583 5698 7613 5712
rect 7656 5698 7699 5712
rect 7721 5708 7911 5720
rect 7976 5716 7982 5736
rect 7706 5698 7736 5708
rect 7737 5698 7895 5708
rect 7899 5698 7929 5708
rect 7933 5698 7963 5712
rect 7991 5698 8004 5736
rect 8076 5750 8105 5766
rect 8119 5750 8148 5766
rect 8163 5756 8193 5772
rect 8221 5750 8227 5798
rect 8230 5792 8249 5798
rect 8264 5792 8294 5800
rect 8230 5784 8294 5792
rect 8230 5768 8310 5784
rect 8326 5777 8388 5808
rect 8404 5777 8466 5808
rect 8535 5806 8584 5831
rect 8599 5806 8629 5822
rect 8498 5792 8528 5800
rect 8535 5798 8645 5806
rect 8498 5784 8543 5792
rect 8230 5766 8249 5768
rect 8264 5766 8310 5768
rect 8230 5750 8310 5766
rect 8337 5764 8372 5777
rect 8413 5774 8450 5777
rect 8413 5772 8455 5774
rect 8342 5761 8372 5764
rect 8351 5757 8358 5761
rect 8358 5756 8359 5757
rect 8317 5750 8327 5756
rect 8076 5742 8111 5750
rect 8076 5716 8077 5742
rect 8084 5716 8111 5742
rect 8019 5698 8049 5712
rect 8076 5708 8111 5716
rect 8113 5742 8154 5750
rect 8113 5716 8128 5742
rect 8135 5716 8154 5742
rect 8218 5738 8249 5750
rect 8264 5738 8367 5750
rect 8379 5740 8405 5766
rect 8420 5761 8450 5772
rect 8482 5768 8544 5784
rect 8482 5766 8528 5768
rect 8482 5750 8544 5766
rect 8556 5750 8562 5798
rect 8565 5790 8645 5798
rect 8565 5788 8584 5790
rect 8599 5788 8633 5790
rect 8565 5772 8645 5788
rect 8565 5750 8584 5772
rect 8599 5756 8629 5772
rect 8657 5766 8663 5840
rect 8666 5766 8685 5910
rect 8700 5766 8706 5910
rect 8715 5840 8728 5910
rect 8780 5906 8802 5910
rect 8773 5884 8802 5898
rect 8855 5884 8871 5898
rect 8909 5894 8915 5896
rect 8922 5894 9030 5910
rect 9037 5894 9043 5896
rect 9051 5894 9066 5910
rect 9132 5904 9151 5907
rect 8773 5882 8871 5884
rect 8898 5882 9066 5894
rect 9081 5884 9097 5898
rect 9132 5885 9154 5904
rect 9164 5898 9180 5899
rect 9163 5896 9180 5898
rect 9164 5891 9180 5896
rect 9154 5884 9160 5885
rect 9163 5884 9192 5891
rect 9081 5883 9192 5884
rect 9081 5882 9198 5883
rect 8757 5874 8808 5882
rect 8855 5874 8889 5882
rect 8757 5862 8782 5874
rect 8789 5862 8808 5874
rect 8862 5872 8889 5874
rect 8898 5872 9119 5882
rect 9154 5879 9160 5882
rect 8862 5868 9119 5872
rect 8757 5854 8808 5862
rect 8855 5854 9119 5868
rect 9163 5874 9198 5882
rect 8709 5806 8728 5840
rect 8773 5846 8802 5854
rect 8773 5840 8790 5846
rect 8773 5838 8807 5840
rect 8855 5838 8871 5854
rect 8872 5844 9080 5854
rect 9081 5844 9097 5854
rect 9145 5850 9160 5865
rect 9163 5862 9164 5874
rect 9171 5862 9198 5874
rect 9163 5854 9198 5862
rect 9163 5853 9192 5854
rect 8883 5840 9097 5844
rect 8898 5838 9097 5840
rect 9132 5840 9145 5850
rect 9163 5840 9180 5853
rect 9132 5838 9180 5840
rect 8774 5834 8807 5838
rect 8770 5832 8807 5834
rect 8770 5831 8837 5832
rect 8770 5826 8801 5831
rect 8807 5826 8837 5831
rect 8770 5822 8837 5826
rect 8743 5819 8837 5822
rect 8743 5812 8792 5819
rect 8743 5806 8773 5812
rect 8792 5807 8797 5812
rect 8709 5790 8789 5806
rect 8801 5798 8837 5819
rect 8898 5814 9087 5838
rect 9132 5837 9179 5838
rect 9145 5832 9179 5837
rect 8913 5811 9087 5814
rect 8906 5808 9087 5811
rect 9115 5831 9179 5832
rect 8709 5788 8728 5790
rect 8743 5788 8777 5790
rect 8709 5772 8789 5788
rect 8709 5766 8728 5772
rect 8425 5740 8528 5750
rect 8379 5738 8528 5740
rect 8549 5738 8584 5750
rect 8218 5736 8380 5738
rect 8230 5716 8249 5736
rect 8264 5734 8294 5736
rect 8113 5708 8154 5716
rect 8236 5712 8249 5716
rect 8301 5720 8380 5736
rect 8412 5736 8584 5738
rect 8412 5720 8491 5736
rect 8498 5734 8528 5736
rect 8076 5698 8105 5708
rect 8119 5698 8148 5708
rect 8163 5698 8193 5712
rect 8236 5698 8279 5712
rect 8301 5708 8491 5720
rect 8556 5716 8562 5736
rect 8286 5698 8316 5708
rect 8317 5698 8475 5708
rect 8479 5698 8509 5708
rect 8513 5698 8543 5712
rect 8571 5698 8584 5736
rect 8656 5750 8685 5766
rect 8699 5750 8728 5766
rect 8743 5756 8773 5772
rect 8801 5750 8807 5798
rect 8810 5792 8829 5798
rect 8844 5792 8874 5800
rect 8810 5784 8874 5792
rect 8810 5768 8890 5784
rect 8906 5777 8968 5808
rect 8984 5777 9046 5808
rect 9115 5806 9164 5831
rect 9179 5806 9209 5822
rect 9078 5792 9108 5800
rect 9115 5798 9225 5806
rect 9078 5784 9123 5792
rect 8810 5766 8829 5768
rect 8844 5766 8890 5768
rect 8810 5750 8890 5766
rect 8917 5764 8952 5777
rect 8993 5774 9030 5777
rect 8993 5772 9035 5774
rect 8922 5761 8952 5764
rect 8931 5757 8938 5761
rect 8938 5756 8939 5757
rect 8897 5750 8907 5756
rect 8656 5742 8691 5750
rect 8656 5716 8657 5742
rect 8664 5716 8691 5742
rect 8599 5698 8629 5712
rect 8656 5708 8691 5716
rect 8693 5742 8734 5750
rect 8693 5716 8708 5742
rect 8715 5716 8734 5742
rect 8798 5738 8829 5750
rect 8844 5738 8947 5750
rect 8959 5740 8985 5766
rect 9000 5761 9030 5772
rect 9062 5768 9124 5784
rect 9062 5766 9108 5768
rect 9062 5750 9124 5766
rect 9136 5750 9142 5798
rect 9145 5790 9225 5798
rect 9145 5788 9164 5790
rect 9179 5788 9213 5790
rect 9145 5772 9225 5788
rect 9145 5750 9164 5772
rect 9179 5756 9209 5772
rect 9237 5766 9243 5840
rect 9246 5766 9265 5910
rect 9280 5766 9286 5910
rect 9295 5840 9308 5910
rect 9360 5906 9382 5910
rect 9353 5884 9382 5898
rect 9435 5884 9451 5898
rect 9489 5894 9495 5896
rect 9502 5894 9610 5910
rect 9617 5894 9623 5896
rect 9631 5894 9646 5910
rect 9712 5904 9731 5907
rect 9353 5882 9451 5884
rect 9478 5882 9646 5894
rect 9661 5884 9677 5898
rect 9712 5885 9734 5904
rect 9744 5898 9760 5899
rect 9743 5896 9760 5898
rect 9744 5891 9760 5896
rect 9734 5884 9740 5885
rect 9743 5884 9772 5891
rect 9661 5883 9772 5884
rect 9661 5882 9778 5883
rect 9337 5874 9388 5882
rect 9435 5874 9469 5882
rect 9337 5862 9362 5874
rect 9369 5862 9388 5874
rect 9442 5872 9469 5874
rect 9478 5872 9699 5882
rect 9734 5879 9740 5882
rect 9442 5868 9699 5872
rect 9337 5854 9388 5862
rect 9435 5854 9699 5868
rect 9743 5874 9778 5882
rect 9289 5806 9308 5840
rect 9353 5846 9382 5854
rect 9353 5840 9370 5846
rect 9353 5838 9387 5840
rect 9435 5838 9451 5854
rect 9452 5844 9660 5854
rect 9661 5844 9677 5854
rect 9725 5850 9740 5865
rect 9743 5862 9744 5874
rect 9751 5862 9778 5874
rect 9743 5854 9778 5862
rect 9743 5853 9772 5854
rect 9463 5840 9677 5844
rect 9478 5838 9677 5840
rect 9712 5840 9725 5850
rect 9743 5840 9760 5853
rect 9712 5838 9760 5840
rect 9354 5834 9387 5838
rect 9350 5832 9387 5834
rect 9350 5831 9417 5832
rect 9350 5826 9381 5831
rect 9387 5826 9417 5831
rect 9350 5822 9417 5826
rect 9323 5819 9417 5822
rect 9323 5812 9372 5819
rect 9323 5806 9353 5812
rect 9372 5807 9377 5812
rect 9289 5790 9369 5806
rect 9381 5798 9417 5819
rect 9478 5814 9667 5838
rect 9712 5837 9759 5838
rect 9725 5832 9759 5837
rect 9493 5811 9667 5814
rect 9486 5808 9667 5811
rect 9695 5831 9759 5832
rect 9289 5788 9308 5790
rect 9323 5788 9357 5790
rect 9289 5772 9369 5788
rect 9289 5766 9308 5772
rect 9005 5740 9108 5750
rect 8959 5738 9108 5740
rect 9129 5738 9164 5750
rect 8798 5736 8960 5738
rect 8810 5716 8829 5736
rect 8844 5734 8874 5736
rect 8693 5708 8734 5716
rect 8816 5712 8829 5716
rect 8881 5720 8960 5736
rect 8992 5736 9164 5738
rect 8992 5720 9071 5736
rect 9078 5734 9108 5736
rect 8656 5698 8685 5708
rect 8699 5698 8728 5708
rect 8743 5698 8773 5712
rect 8816 5698 8859 5712
rect 8881 5708 9071 5720
rect 9136 5716 9142 5736
rect 8866 5698 8896 5708
rect 8897 5698 9055 5708
rect 9059 5698 9089 5708
rect 9093 5698 9123 5712
rect 9151 5698 9164 5736
rect 9236 5750 9265 5766
rect 9279 5750 9308 5766
rect 9323 5756 9353 5772
rect 9381 5750 9387 5798
rect 9390 5792 9409 5798
rect 9424 5792 9454 5800
rect 9390 5784 9454 5792
rect 9390 5768 9470 5784
rect 9486 5777 9548 5808
rect 9564 5777 9626 5808
rect 9695 5806 9744 5831
rect 9759 5806 9789 5822
rect 9658 5792 9688 5800
rect 9695 5798 9805 5806
rect 9658 5784 9703 5792
rect 9390 5766 9409 5768
rect 9424 5766 9470 5768
rect 9390 5750 9470 5766
rect 9497 5764 9532 5777
rect 9573 5774 9610 5777
rect 9573 5772 9615 5774
rect 9502 5761 9532 5764
rect 9511 5757 9518 5761
rect 9518 5756 9519 5757
rect 9477 5750 9487 5756
rect 9236 5742 9271 5750
rect 9236 5716 9237 5742
rect 9244 5716 9271 5742
rect 9179 5698 9209 5712
rect 9236 5708 9271 5716
rect 9273 5742 9314 5750
rect 9273 5716 9288 5742
rect 9295 5716 9314 5742
rect 9378 5738 9409 5750
rect 9424 5738 9527 5750
rect 9539 5740 9565 5766
rect 9580 5761 9610 5772
rect 9642 5768 9704 5784
rect 9642 5766 9688 5768
rect 9642 5750 9704 5766
rect 9716 5750 9722 5798
rect 9725 5790 9805 5798
rect 9725 5788 9744 5790
rect 9759 5788 9793 5790
rect 9725 5772 9805 5788
rect 9725 5750 9744 5772
rect 9759 5756 9789 5772
rect 9817 5766 9823 5840
rect 9826 5766 9845 5910
rect 9860 5766 9866 5910
rect 9875 5840 9888 5910
rect 9940 5906 9962 5910
rect 9933 5884 9962 5898
rect 10015 5884 10031 5898
rect 10069 5894 10075 5896
rect 10082 5894 10190 5910
rect 10197 5894 10203 5896
rect 10211 5894 10226 5910
rect 10292 5904 10311 5907
rect 9933 5882 10031 5884
rect 10058 5882 10226 5894
rect 10241 5884 10257 5898
rect 10292 5885 10314 5904
rect 10324 5898 10340 5899
rect 10323 5896 10340 5898
rect 10324 5891 10340 5896
rect 10314 5884 10320 5885
rect 10323 5884 10352 5891
rect 10241 5883 10352 5884
rect 10241 5882 10358 5883
rect 9917 5874 9968 5882
rect 10015 5874 10049 5882
rect 9917 5862 9942 5874
rect 9949 5862 9968 5874
rect 10022 5872 10049 5874
rect 10058 5872 10279 5882
rect 10314 5879 10320 5882
rect 10022 5868 10279 5872
rect 9917 5854 9968 5862
rect 10015 5854 10279 5868
rect 10323 5874 10358 5882
rect 9869 5806 9888 5840
rect 9933 5846 9962 5854
rect 9933 5840 9950 5846
rect 9933 5838 9967 5840
rect 10015 5838 10031 5854
rect 10032 5844 10240 5854
rect 10241 5844 10257 5854
rect 10305 5850 10320 5865
rect 10323 5862 10324 5874
rect 10331 5862 10358 5874
rect 10323 5854 10358 5862
rect 10323 5853 10352 5854
rect 10043 5840 10257 5844
rect 10058 5838 10257 5840
rect 10292 5840 10305 5850
rect 10323 5840 10340 5853
rect 10292 5838 10340 5840
rect 9934 5834 9967 5838
rect 9930 5832 9967 5834
rect 9930 5831 9997 5832
rect 9930 5826 9961 5831
rect 9967 5826 9997 5831
rect 9930 5822 9997 5826
rect 9903 5819 9997 5822
rect 9903 5812 9952 5819
rect 9903 5806 9933 5812
rect 9952 5807 9957 5812
rect 9869 5790 9949 5806
rect 9961 5798 9997 5819
rect 10058 5814 10247 5838
rect 10292 5837 10339 5838
rect 10305 5832 10339 5837
rect 10073 5811 10247 5814
rect 10066 5808 10247 5811
rect 10275 5831 10339 5832
rect 9869 5788 9888 5790
rect 9903 5788 9937 5790
rect 9869 5772 9949 5788
rect 9869 5766 9888 5772
rect 9585 5740 9688 5750
rect 9539 5738 9688 5740
rect 9709 5738 9744 5750
rect 9378 5736 9540 5738
rect 9390 5716 9409 5736
rect 9424 5734 9454 5736
rect 9273 5708 9314 5716
rect 9396 5712 9409 5716
rect 9461 5720 9540 5736
rect 9572 5736 9744 5738
rect 9572 5720 9651 5736
rect 9658 5734 9688 5736
rect 9236 5698 9265 5708
rect 9279 5698 9308 5708
rect 9323 5698 9353 5712
rect 9396 5698 9439 5712
rect 9461 5708 9651 5720
rect 9716 5716 9722 5736
rect 9446 5698 9476 5708
rect 9477 5698 9635 5708
rect 9639 5698 9669 5708
rect 9673 5698 9703 5712
rect 9731 5698 9744 5736
rect 9816 5750 9845 5766
rect 9859 5750 9888 5766
rect 9903 5756 9933 5772
rect 9961 5750 9967 5798
rect 9970 5792 9989 5798
rect 10004 5792 10034 5800
rect 9970 5784 10034 5792
rect 9970 5768 10050 5784
rect 10066 5777 10128 5808
rect 10144 5777 10206 5808
rect 10275 5806 10324 5831
rect 10339 5806 10369 5822
rect 10238 5792 10268 5800
rect 10275 5798 10385 5806
rect 10238 5784 10283 5792
rect 9970 5766 9989 5768
rect 10004 5766 10050 5768
rect 9970 5750 10050 5766
rect 10077 5764 10112 5777
rect 10153 5774 10190 5777
rect 10153 5772 10195 5774
rect 10082 5761 10112 5764
rect 10091 5757 10098 5761
rect 10098 5756 10099 5757
rect 10057 5750 10067 5756
rect 9816 5742 9851 5750
rect 9816 5716 9817 5742
rect 9824 5716 9851 5742
rect 9759 5698 9789 5712
rect 9816 5708 9851 5716
rect 9853 5742 9894 5750
rect 9853 5716 9868 5742
rect 9875 5716 9894 5742
rect 9958 5738 9989 5750
rect 10004 5738 10107 5750
rect 10119 5740 10145 5766
rect 10160 5761 10190 5772
rect 10222 5768 10284 5784
rect 10222 5766 10268 5768
rect 10222 5750 10284 5766
rect 10296 5750 10302 5798
rect 10305 5790 10385 5798
rect 10305 5788 10324 5790
rect 10339 5788 10373 5790
rect 10305 5772 10385 5788
rect 10305 5750 10324 5772
rect 10339 5756 10369 5772
rect 10397 5766 10403 5840
rect 10406 5766 10425 5910
rect 10440 5766 10446 5910
rect 10455 5840 10468 5910
rect 10520 5906 10542 5910
rect 10513 5884 10542 5898
rect 10595 5884 10611 5898
rect 10649 5894 10655 5896
rect 10662 5894 10770 5910
rect 10777 5894 10783 5896
rect 10791 5894 10806 5910
rect 10872 5904 10891 5907
rect 10513 5882 10611 5884
rect 10638 5882 10806 5894
rect 10821 5884 10837 5898
rect 10872 5885 10894 5904
rect 10904 5898 10920 5899
rect 10903 5896 10920 5898
rect 10904 5891 10920 5896
rect 10894 5884 10900 5885
rect 10903 5884 10932 5891
rect 10821 5883 10932 5884
rect 10821 5882 10938 5883
rect 10497 5874 10548 5882
rect 10595 5874 10629 5882
rect 10497 5862 10522 5874
rect 10529 5862 10548 5874
rect 10602 5872 10629 5874
rect 10638 5872 10859 5882
rect 10894 5879 10900 5882
rect 10602 5868 10859 5872
rect 10497 5854 10548 5862
rect 10595 5854 10859 5868
rect 10903 5874 10938 5882
rect 10449 5806 10468 5840
rect 10513 5846 10542 5854
rect 10513 5840 10530 5846
rect 10513 5838 10547 5840
rect 10595 5838 10611 5854
rect 10612 5844 10820 5854
rect 10821 5844 10837 5854
rect 10885 5850 10900 5865
rect 10903 5862 10904 5874
rect 10911 5862 10938 5874
rect 10903 5854 10938 5862
rect 10903 5853 10932 5854
rect 10623 5840 10837 5844
rect 10638 5838 10837 5840
rect 10872 5840 10885 5850
rect 10903 5840 10920 5853
rect 10872 5838 10920 5840
rect 10514 5834 10547 5838
rect 10510 5832 10547 5834
rect 10510 5831 10577 5832
rect 10510 5826 10541 5831
rect 10547 5826 10577 5831
rect 10510 5822 10577 5826
rect 10483 5819 10577 5822
rect 10483 5812 10532 5819
rect 10483 5806 10513 5812
rect 10532 5807 10537 5812
rect 10449 5790 10529 5806
rect 10541 5798 10577 5819
rect 10638 5814 10827 5838
rect 10872 5837 10919 5838
rect 10885 5832 10919 5837
rect 10653 5811 10827 5814
rect 10646 5808 10827 5811
rect 10855 5831 10919 5832
rect 10449 5788 10468 5790
rect 10483 5788 10517 5790
rect 10449 5772 10529 5788
rect 10449 5766 10468 5772
rect 10165 5740 10268 5750
rect 10119 5738 10268 5740
rect 10289 5738 10324 5750
rect 9958 5736 10120 5738
rect 9970 5716 9989 5736
rect 10004 5734 10034 5736
rect 9853 5708 9894 5716
rect 9976 5712 9989 5716
rect 10041 5720 10120 5736
rect 10152 5736 10324 5738
rect 10152 5720 10231 5736
rect 10238 5734 10268 5736
rect 9816 5698 9845 5708
rect 9859 5698 9888 5708
rect 9903 5698 9933 5712
rect 9976 5698 10019 5712
rect 10041 5708 10231 5720
rect 10296 5716 10302 5736
rect 10026 5698 10056 5708
rect 10057 5698 10215 5708
rect 10219 5698 10249 5708
rect 10253 5698 10283 5712
rect 10311 5698 10324 5736
rect 10396 5750 10425 5766
rect 10439 5750 10468 5766
rect 10483 5756 10513 5772
rect 10541 5750 10547 5798
rect 10550 5792 10569 5798
rect 10584 5792 10614 5800
rect 10550 5784 10614 5792
rect 10550 5768 10630 5784
rect 10646 5777 10708 5808
rect 10724 5777 10786 5808
rect 10855 5806 10904 5831
rect 10919 5806 10949 5822
rect 10818 5792 10848 5800
rect 10855 5798 10965 5806
rect 10818 5784 10863 5792
rect 10550 5766 10569 5768
rect 10584 5766 10630 5768
rect 10550 5750 10630 5766
rect 10657 5764 10692 5777
rect 10733 5774 10770 5777
rect 10733 5772 10775 5774
rect 10662 5761 10692 5764
rect 10671 5757 10678 5761
rect 10678 5756 10679 5757
rect 10637 5750 10647 5756
rect 10396 5742 10431 5750
rect 10396 5716 10397 5742
rect 10404 5716 10431 5742
rect 10339 5698 10369 5712
rect 10396 5708 10431 5716
rect 10433 5742 10474 5750
rect 10433 5716 10448 5742
rect 10455 5716 10474 5742
rect 10538 5738 10569 5750
rect 10584 5738 10687 5750
rect 10699 5740 10725 5766
rect 10740 5761 10770 5772
rect 10802 5768 10864 5784
rect 10802 5766 10848 5768
rect 10802 5750 10864 5766
rect 10876 5750 10882 5798
rect 10885 5790 10965 5798
rect 10885 5788 10904 5790
rect 10919 5788 10953 5790
rect 10885 5772 10965 5788
rect 10885 5750 10904 5772
rect 10919 5756 10949 5772
rect 10977 5766 10983 5840
rect 10986 5766 11005 5910
rect 11020 5766 11026 5910
rect 11035 5840 11048 5910
rect 11100 5906 11122 5910
rect 11093 5884 11122 5898
rect 11175 5884 11191 5898
rect 11229 5894 11235 5896
rect 11242 5894 11350 5910
rect 11357 5894 11363 5896
rect 11371 5894 11386 5910
rect 11452 5904 11471 5907
rect 11093 5882 11191 5884
rect 11218 5882 11386 5894
rect 11401 5884 11417 5898
rect 11452 5885 11474 5904
rect 11484 5898 11500 5899
rect 11483 5896 11500 5898
rect 11484 5891 11500 5896
rect 11474 5884 11480 5885
rect 11483 5884 11512 5891
rect 11401 5883 11512 5884
rect 11401 5882 11518 5883
rect 11077 5874 11128 5882
rect 11175 5874 11209 5882
rect 11077 5862 11102 5874
rect 11109 5862 11128 5874
rect 11182 5872 11209 5874
rect 11218 5872 11439 5882
rect 11474 5879 11480 5882
rect 11182 5868 11439 5872
rect 11077 5854 11128 5862
rect 11175 5854 11439 5868
rect 11483 5874 11518 5882
rect 11029 5806 11048 5840
rect 11093 5846 11122 5854
rect 11093 5840 11110 5846
rect 11093 5838 11127 5840
rect 11175 5838 11191 5854
rect 11192 5844 11400 5854
rect 11401 5844 11417 5854
rect 11465 5850 11480 5865
rect 11483 5862 11484 5874
rect 11491 5862 11518 5874
rect 11483 5854 11518 5862
rect 11483 5853 11512 5854
rect 11203 5840 11417 5844
rect 11218 5838 11417 5840
rect 11452 5840 11465 5850
rect 11483 5840 11500 5853
rect 11452 5838 11500 5840
rect 11094 5834 11127 5838
rect 11090 5832 11127 5834
rect 11090 5831 11157 5832
rect 11090 5826 11121 5831
rect 11127 5826 11157 5831
rect 11090 5822 11157 5826
rect 11063 5819 11157 5822
rect 11063 5812 11112 5819
rect 11063 5806 11093 5812
rect 11112 5807 11117 5812
rect 11029 5790 11109 5806
rect 11121 5798 11157 5819
rect 11218 5814 11407 5838
rect 11452 5837 11499 5838
rect 11465 5832 11499 5837
rect 11233 5811 11407 5814
rect 11226 5808 11407 5811
rect 11435 5831 11499 5832
rect 11029 5788 11048 5790
rect 11063 5788 11097 5790
rect 11029 5772 11109 5788
rect 11029 5766 11048 5772
rect 10745 5740 10848 5750
rect 10699 5738 10848 5740
rect 10869 5738 10904 5750
rect 10538 5736 10700 5738
rect 10550 5716 10569 5736
rect 10584 5734 10614 5736
rect 10433 5708 10474 5716
rect 10556 5712 10569 5716
rect 10621 5720 10700 5736
rect 10732 5736 10904 5738
rect 10732 5720 10811 5736
rect 10818 5734 10848 5736
rect 10396 5698 10425 5708
rect 10439 5698 10468 5708
rect 10483 5698 10513 5712
rect 10556 5698 10599 5712
rect 10621 5708 10811 5720
rect 10876 5716 10882 5736
rect 10606 5698 10636 5708
rect 10637 5698 10795 5708
rect 10799 5698 10829 5708
rect 10833 5698 10863 5712
rect 10891 5698 10904 5736
rect 10976 5750 11005 5766
rect 11019 5750 11048 5766
rect 11063 5756 11093 5772
rect 11121 5750 11127 5798
rect 11130 5792 11149 5798
rect 11164 5792 11194 5800
rect 11130 5784 11194 5792
rect 11130 5768 11210 5784
rect 11226 5777 11288 5808
rect 11304 5777 11366 5808
rect 11435 5806 11484 5831
rect 11499 5806 11529 5822
rect 11398 5792 11428 5800
rect 11435 5798 11545 5806
rect 11398 5784 11443 5792
rect 11130 5766 11149 5768
rect 11164 5766 11210 5768
rect 11130 5750 11210 5766
rect 11237 5764 11272 5777
rect 11313 5774 11350 5777
rect 11313 5772 11355 5774
rect 11242 5761 11272 5764
rect 11251 5757 11258 5761
rect 11258 5756 11259 5757
rect 11217 5750 11227 5756
rect 10976 5742 11011 5750
rect 10976 5716 10977 5742
rect 10984 5716 11011 5742
rect 10919 5698 10949 5712
rect 10976 5708 11011 5716
rect 11013 5742 11054 5750
rect 11013 5716 11028 5742
rect 11035 5716 11054 5742
rect 11118 5738 11149 5750
rect 11164 5738 11267 5750
rect 11279 5740 11305 5766
rect 11320 5761 11350 5772
rect 11382 5768 11444 5784
rect 11382 5766 11428 5768
rect 11382 5750 11444 5766
rect 11456 5750 11462 5798
rect 11465 5790 11545 5798
rect 11465 5788 11484 5790
rect 11499 5788 11533 5790
rect 11465 5772 11545 5788
rect 11465 5750 11484 5772
rect 11499 5756 11529 5772
rect 11557 5766 11563 5840
rect 11566 5766 11585 5910
rect 11600 5766 11606 5910
rect 11615 5840 11628 5910
rect 11680 5906 11702 5910
rect 11673 5884 11702 5898
rect 11755 5884 11771 5898
rect 11809 5894 11815 5896
rect 11822 5894 11930 5910
rect 11937 5894 11943 5896
rect 11951 5894 11966 5910
rect 12032 5904 12051 5907
rect 11673 5882 11771 5884
rect 11798 5882 11966 5894
rect 11981 5884 11997 5898
rect 12032 5885 12054 5904
rect 12064 5898 12080 5899
rect 12063 5896 12080 5898
rect 12064 5891 12080 5896
rect 12054 5884 12060 5885
rect 12063 5884 12092 5891
rect 11981 5883 12092 5884
rect 11981 5882 12098 5883
rect 11657 5874 11708 5882
rect 11755 5874 11789 5882
rect 11657 5862 11682 5874
rect 11689 5862 11708 5874
rect 11762 5872 11789 5874
rect 11798 5872 12019 5882
rect 12054 5879 12060 5882
rect 11762 5868 12019 5872
rect 11657 5854 11708 5862
rect 11755 5854 12019 5868
rect 12063 5874 12098 5882
rect 11609 5806 11628 5840
rect 11673 5846 11702 5854
rect 11673 5840 11690 5846
rect 11673 5838 11707 5840
rect 11755 5838 11771 5854
rect 11772 5844 11980 5854
rect 11981 5844 11997 5854
rect 12045 5850 12060 5865
rect 12063 5862 12064 5874
rect 12071 5862 12098 5874
rect 12063 5854 12098 5862
rect 12063 5853 12092 5854
rect 11783 5840 11997 5844
rect 11798 5838 11997 5840
rect 12032 5840 12045 5850
rect 12063 5840 12080 5853
rect 12032 5838 12080 5840
rect 11674 5834 11707 5838
rect 11670 5832 11707 5834
rect 11670 5831 11737 5832
rect 11670 5826 11701 5831
rect 11707 5826 11737 5831
rect 11670 5822 11737 5826
rect 11643 5819 11737 5822
rect 11643 5812 11692 5819
rect 11643 5806 11673 5812
rect 11692 5807 11697 5812
rect 11609 5790 11689 5806
rect 11701 5798 11737 5819
rect 11798 5814 11987 5838
rect 12032 5837 12079 5838
rect 12045 5832 12079 5837
rect 11813 5811 11987 5814
rect 11806 5808 11987 5811
rect 12015 5831 12079 5832
rect 11609 5788 11628 5790
rect 11643 5788 11677 5790
rect 11609 5772 11689 5788
rect 11609 5766 11628 5772
rect 11325 5740 11428 5750
rect 11279 5738 11428 5740
rect 11449 5738 11484 5750
rect 11118 5736 11280 5738
rect 11130 5716 11149 5736
rect 11164 5734 11194 5736
rect 11013 5708 11054 5716
rect 11136 5712 11149 5716
rect 11201 5720 11280 5736
rect 11312 5736 11484 5738
rect 11312 5720 11391 5736
rect 11398 5734 11428 5736
rect 10976 5698 11005 5708
rect 11019 5698 11048 5708
rect 11063 5698 11093 5712
rect 11136 5698 11179 5712
rect 11201 5708 11391 5720
rect 11456 5716 11462 5736
rect 11186 5698 11216 5708
rect 11217 5698 11375 5708
rect 11379 5698 11409 5708
rect 11413 5698 11443 5712
rect 11471 5698 11484 5736
rect 11556 5750 11585 5766
rect 11599 5750 11628 5766
rect 11643 5756 11673 5772
rect 11701 5750 11707 5798
rect 11710 5792 11729 5798
rect 11744 5792 11774 5800
rect 11710 5784 11774 5792
rect 11710 5768 11790 5784
rect 11806 5777 11868 5808
rect 11884 5777 11946 5808
rect 12015 5806 12064 5831
rect 12079 5806 12109 5822
rect 11978 5792 12008 5800
rect 12015 5798 12125 5806
rect 11978 5784 12023 5792
rect 11710 5766 11729 5768
rect 11744 5766 11790 5768
rect 11710 5750 11790 5766
rect 11817 5764 11852 5777
rect 11893 5774 11930 5777
rect 11893 5772 11935 5774
rect 11822 5761 11852 5764
rect 11831 5757 11838 5761
rect 11838 5756 11839 5757
rect 11797 5750 11807 5756
rect 11556 5742 11591 5750
rect 11556 5716 11557 5742
rect 11564 5716 11591 5742
rect 11499 5698 11529 5712
rect 11556 5708 11591 5716
rect 11593 5742 11634 5750
rect 11593 5716 11608 5742
rect 11615 5716 11634 5742
rect 11698 5738 11729 5750
rect 11744 5738 11847 5750
rect 11859 5740 11885 5766
rect 11900 5761 11930 5772
rect 11962 5768 12024 5784
rect 11962 5766 12008 5768
rect 11962 5750 12024 5766
rect 12036 5750 12042 5798
rect 12045 5790 12125 5798
rect 12045 5788 12064 5790
rect 12079 5788 12113 5790
rect 12045 5772 12125 5788
rect 12045 5750 12064 5772
rect 12079 5756 12109 5772
rect 12137 5766 12143 5840
rect 12146 5766 12165 5910
rect 12180 5766 12186 5910
rect 12195 5840 12208 5910
rect 12260 5906 12282 5910
rect 12253 5884 12282 5898
rect 12335 5884 12351 5898
rect 12389 5894 12395 5896
rect 12402 5894 12510 5910
rect 12517 5894 12523 5896
rect 12531 5894 12546 5910
rect 12612 5904 12631 5907
rect 12253 5882 12351 5884
rect 12378 5882 12546 5894
rect 12561 5884 12577 5898
rect 12612 5885 12634 5904
rect 12644 5898 12660 5899
rect 12643 5896 12660 5898
rect 12644 5891 12660 5896
rect 12634 5884 12640 5885
rect 12643 5884 12672 5891
rect 12561 5883 12672 5884
rect 12561 5882 12678 5883
rect 12237 5874 12288 5882
rect 12335 5874 12369 5882
rect 12237 5862 12262 5874
rect 12269 5862 12288 5874
rect 12342 5872 12369 5874
rect 12378 5872 12599 5882
rect 12634 5879 12640 5882
rect 12342 5868 12599 5872
rect 12237 5854 12288 5862
rect 12335 5854 12599 5868
rect 12643 5874 12678 5882
rect 12189 5806 12208 5840
rect 12253 5846 12282 5854
rect 12253 5840 12270 5846
rect 12253 5838 12287 5840
rect 12335 5838 12351 5854
rect 12352 5844 12560 5854
rect 12561 5844 12577 5854
rect 12625 5850 12640 5865
rect 12643 5862 12644 5874
rect 12651 5862 12678 5874
rect 12643 5854 12678 5862
rect 12643 5853 12672 5854
rect 12363 5840 12577 5844
rect 12378 5838 12577 5840
rect 12612 5840 12625 5850
rect 12643 5840 12660 5853
rect 12612 5838 12660 5840
rect 12254 5834 12287 5838
rect 12250 5832 12287 5834
rect 12250 5831 12317 5832
rect 12250 5826 12281 5831
rect 12287 5826 12317 5831
rect 12250 5822 12317 5826
rect 12223 5819 12317 5822
rect 12223 5812 12272 5819
rect 12223 5806 12253 5812
rect 12272 5807 12277 5812
rect 12189 5790 12269 5806
rect 12281 5798 12317 5819
rect 12378 5814 12567 5838
rect 12612 5837 12659 5838
rect 12625 5832 12659 5837
rect 12393 5811 12567 5814
rect 12386 5808 12567 5811
rect 12595 5831 12659 5832
rect 12189 5788 12208 5790
rect 12223 5788 12257 5790
rect 12189 5772 12269 5788
rect 12189 5766 12208 5772
rect 11905 5740 12008 5750
rect 11859 5738 12008 5740
rect 12029 5738 12064 5750
rect 11698 5736 11860 5738
rect 11710 5716 11729 5736
rect 11744 5734 11774 5736
rect 11593 5708 11634 5716
rect 11716 5712 11729 5716
rect 11781 5720 11860 5736
rect 11892 5736 12064 5738
rect 11892 5720 11971 5736
rect 11978 5734 12008 5736
rect 11556 5698 11585 5708
rect 11599 5698 11628 5708
rect 11643 5698 11673 5712
rect 11716 5698 11759 5712
rect 11781 5708 11971 5720
rect 12036 5716 12042 5736
rect 11766 5698 11796 5708
rect 11797 5698 11955 5708
rect 11959 5698 11989 5708
rect 11993 5698 12023 5712
rect 12051 5698 12064 5736
rect 12136 5750 12165 5766
rect 12179 5750 12208 5766
rect 12223 5756 12253 5772
rect 12281 5750 12287 5798
rect 12290 5792 12309 5798
rect 12324 5792 12354 5800
rect 12290 5784 12354 5792
rect 12290 5768 12370 5784
rect 12386 5777 12448 5808
rect 12464 5777 12526 5808
rect 12595 5806 12644 5831
rect 12659 5806 12689 5822
rect 12558 5792 12588 5800
rect 12595 5798 12705 5806
rect 12558 5784 12603 5792
rect 12290 5766 12309 5768
rect 12324 5766 12370 5768
rect 12290 5750 12370 5766
rect 12397 5764 12432 5777
rect 12473 5774 12510 5777
rect 12473 5772 12515 5774
rect 12402 5761 12432 5764
rect 12411 5757 12418 5761
rect 12418 5756 12419 5757
rect 12377 5750 12387 5756
rect 12136 5742 12171 5750
rect 12136 5716 12137 5742
rect 12144 5716 12171 5742
rect 12079 5698 12109 5712
rect 12136 5708 12171 5716
rect 12173 5742 12214 5750
rect 12173 5716 12188 5742
rect 12195 5716 12214 5742
rect 12278 5738 12309 5750
rect 12324 5738 12427 5750
rect 12439 5740 12465 5766
rect 12480 5761 12510 5772
rect 12542 5768 12604 5784
rect 12542 5766 12588 5768
rect 12542 5750 12604 5766
rect 12616 5750 12622 5798
rect 12625 5790 12705 5798
rect 12625 5788 12644 5790
rect 12659 5788 12693 5790
rect 12625 5772 12705 5788
rect 12625 5750 12644 5772
rect 12659 5756 12689 5772
rect 12717 5766 12723 5840
rect 12726 5766 12745 5910
rect 12760 5766 12766 5910
rect 12775 5840 12788 5910
rect 12840 5906 12862 5910
rect 12833 5884 12862 5898
rect 12915 5884 12931 5898
rect 12969 5894 12975 5896
rect 12982 5894 13090 5910
rect 13097 5894 13103 5896
rect 13111 5894 13126 5910
rect 13192 5904 13211 5907
rect 12833 5882 12931 5884
rect 12958 5882 13126 5894
rect 13141 5884 13157 5898
rect 13192 5885 13214 5904
rect 13224 5898 13240 5899
rect 13223 5896 13240 5898
rect 13224 5891 13240 5896
rect 13214 5884 13220 5885
rect 13223 5884 13252 5891
rect 13141 5883 13252 5884
rect 13141 5882 13258 5883
rect 12817 5874 12868 5882
rect 12915 5874 12949 5882
rect 12817 5862 12842 5874
rect 12849 5862 12868 5874
rect 12922 5872 12949 5874
rect 12958 5872 13179 5882
rect 13214 5879 13220 5882
rect 12922 5868 13179 5872
rect 12817 5854 12868 5862
rect 12915 5854 13179 5868
rect 13223 5874 13258 5882
rect 12769 5806 12788 5840
rect 12833 5846 12862 5854
rect 12833 5840 12850 5846
rect 12833 5838 12867 5840
rect 12915 5838 12931 5854
rect 12932 5844 13140 5854
rect 13141 5844 13157 5854
rect 13205 5850 13220 5865
rect 13223 5862 13224 5874
rect 13231 5862 13258 5874
rect 13223 5854 13258 5862
rect 13223 5853 13252 5854
rect 12943 5840 13157 5844
rect 12958 5838 13157 5840
rect 13192 5840 13205 5850
rect 13223 5840 13240 5853
rect 13192 5838 13240 5840
rect 12834 5834 12867 5838
rect 12830 5832 12867 5834
rect 12830 5831 12897 5832
rect 12830 5826 12861 5831
rect 12867 5826 12897 5831
rect 12830 5822 12897 5826
rect 12803 5819 12897 5822
rect 12803 5812 12852 5819
rect 12803 5806 12833 5812
rect 12852 5807 12857 5812
rect 12769 5790 12849 5806
rect 12861 5798 12897 5819
rect 12958 5814 13147 5838
rect 13192 5837 13239 5838
rect 13205 5832 13239 5837
rect 12973 5811 13147 5814
rect 12966 5808 13147 5811
rect 13175 5831 13239 5832
rect 12769 5788 12788 5790
rect 12803 5788 12837 5790
rect 12769 5772 12849 5788
rect 12769 5766 12788 5772
rect 12485 5740 12588 5750
rect 12439 5738 12588 5740
rect 12609 5738 12644 5750
rect 12278 5736 12440 5738
rect 12290 5716 12309 5736
rect 12324 5734 12354 5736
rect 12173 5708 12214 5716
rect 12296 5712 12309 5716
rect 12361 5720 12440 5736
rect 12472 5736 12644 5738
rect 12472 5720 12551 5736
rect 12558 5734 12588 5736
rect 12136 5698 12165 5708
rect 12179 5698 12208 5708
rect 12223 5698 12253 5712
rect 12296 5698 12339 5712
rect 12361 5708 12551 5720
rect 12616 5716 12622 5736
rect 12346 5698 12376 5708
rect 12377 5698 12535 5708
rect 12539 5698 12569 5708
rect 12573 5698 12603 5712
rect 12631 5698 12644 5736
rect 12716 5750 12745 5766
rect 12759 5750 12788 5766
rect 12803 5756 12833 5772
rect 12861 5750 12867 5798
rect 12870 5792 12889 5798
rect 12904 5792 12934 5800
rect 12870 5784 12934 5792
rect 12870 5768 12950 5784
rect 12966 5777 13028 5808
rect 13044 5777 13106 5808
rect 13175 5806 13224 5831
rect 13239 5806 13269 5822
rect 13138 5792 13168 5800
rect 13175 5798 13285 5806
rect 13138 5784 13183 5792
rect 12870 5766 12889 5768
rect 12904 5766 12950 5768
rect 12870 5750 12950 5766
rect 12977 5764 13012 5777
rect 13053 5774 13090 5777
rect 13053 5772 13095 5774
rect 12982 5761 13012 5764
rect 12991 5757 12998 5761
rect 12998 5756 12999 5757
rect 12957 5750 12967 5756
rect 12716 5742 12751 5750
rect 12716 5716 12717 5742
rect 12724 5716 12751 5742
rect 12659 5698 12689 5712
rect 12716 5708 12751 5716
rect 12753 5742 12794 5750
rect 12753 5716 12768 5742
rect 12775 5716 12794 5742
rect 12858 5738 12889 5750
rect 12904 5738 13007 5750
rect 13019 5740 13045 5766
rect 13060 5761 13090 5772
rect 13122 5768 13184 5784
rect 13122 5766 13168 5768
rect 13122 5750 13184 5766
rect 13196 5750 13202 5798
rect 13205 5790 13285 5798
rect 13205 5788 13224 5790
rect 13239 5788 13273 5790
rect 13205 5772 13285 5788
rect 13205 5750 13224 5772
rect 13239 5756 13269 5772
rect 13297 5766 13303 5840
rect 13306 5766 13325 5910
rect 13340 5766 13346 5910
rect 13355 5840 13368 5910
rect 13420 5906 13442 5910
rect 13413 5884 13442 5898
rect 13495 5884 13511 5898
rect 13549 5894 13555 5896
rect 13562 5894 13670 5910
rect 13677 5894 13683 5896
rect 13691 5894 13706 5910
rect 13772 5904 13791 5907
rect 13413 5882 13511 5884
rect 13538 5882 13706 5894
rect 13721 5884 13737 5898
rect 13772 5885 13794 5904
rect 13804 5898 13820 5899
rect 13803 5896 13820 5898
rect 13804 5891 13820 5896
rect 13794 5884 13800 5885
rect 13803 5884 13832 5891
rect 13721 5883 13832 5884
rect 13721 5882 13838 5883
rect 13397 5874 13448 5882
rect 13495 5874 13529 5882
rect 13397 5862 13422 5874
rect 13429 5862 13448 5874
rect 13502 5872 13529 5874
rect 13538 5872 13759 5882
rect 13794 5879 13800 5882
rect 13502 5868 13759 5872
rect 13397 5854 13448 5862
rect 13495 5854 13759 5868
rect 13803 5874 13838 5882
rect 13349 5806 13368 5840
rect 13413 5846 13442 5854
rect 13413 5840 13430 5846
rect 13413 5838 13447 5840
rect 13495 5838 13511 5854
rect 13512 5844 13720 5854
rect 13721 5844 13737 5854
rect 13785 5850 13800 5865
rect 13803 5862 13804 5874
rect 13811 5862 13838 5874
rect 13803 5854 13838 5862
rect 13803 5853 13832 5854
rect 13523 5840 13737 5844
rect 13538 5838 13737 5840
rect 13772 5840 13785 5850
rect 13803 5840 13820 5853
rect 13772 5838 13820 5840
rect 13414 5834 13447 5838
rect 13410 5832 13447 5834
rect 13410 5831 13477 5832
rect 13410 5826 13441 5831
rect 13447 5826 13477 5831
rect 13410 5822 13477 5826
rect 13383 5819 13477 5822
rect 13383 5812 13432 5819
rect 13383 5806 13413 5812
rect 13432 5807 13437 5812
rect 13349 5790 13429 5806
rect 13441 5798 13477 5819
rect 13538 5814 13727 5838
rect 13772 5837 13819 5838
rect 13785 5832 13819 5837
rect 13553 5811 13727 5814
rect 13546 5808 13727 5811
rect 13755 5831 13819 5832
rect 13349 5788 13368 5790
rect 13383 5788 13417 5790
rect 13349 5772 13429 5788
rect 13349 5766 13368 5772
rect 13065 5740 13168 5750
rect 13019 5738 13168 5740
rect 13189 5738 13224 5750
rect 12858 5736 13020 5738
rect 12870 5716 12889 5736
rect 12904 5734 12934 5736
rect 12753 5708 12794 5716
rect 12876 5712 12889 5716
rect 12941 5720 13020 5736
rect 13052 5736 13224 5738
rect 13052 5720 13131 5736
rect 13138 5734 13168 5736
rect 12716 5698 12745 5708
rect 12759 5698 12788 5708
rect 12803 5698 12833 5712
rect 12876 5698 12919 5712
rect 12941 5708 13131 5720
rect 13196 5716 13202 5736
rect 12926 5698 12956 5708
rect 12957 5698 13115 5708
rect 13119 5698 13149 5708
rect 13153 5698 13183 5712
rect 13211 5698 13224 5736
rect 13296 5750 13325 5766
rect 13339 5750 13368 5766
rect 13383 5756 13413 5772
rect 13441 5750 13447 5798
rect 13450 5792 13469 5798
rect 13484 5792 13514 5800
rect 13450 5784 13514 5792
rect 13450 5768 13530 5784
rect 13546 5777 13608 5808
rect 13624 5777 13686 5808
rect 13755 5806 13804 5831
rect 13819 5806 13849 5822
rect 13718 5792 13748 5800
rect 13755 5798 13865 5806
rect 13718 5784 13763 5792
rect 13450 5766 13469 5768
rect 13484 5766 13530 5768
rect 13450 5750 13530 5766
rect 13557 5764 13592 5777
rect 13633 5774 13670 5777
rect 13633 5772 13675 5774
rect 13562 5761 13592 5764
rect 13571 5757 13578 5761
rect 13578 5756 13579 5757
rect 13537 5750 13547 5756
rect 13296 5742 13331 5750
rect 13296 5716 13297 5742
rect 13304 5716 13331 5742
rect 13239 5698 13269 5712
rect 13296 5708 13331 5716
rect 13333 5742 13374 5750
rect 13333 5716 13348 5742
rect 13355 5716 13374 5742
rect 13438 5738 13469 5750
rect 13484 5738 13587 5750
rect 13599 5740 13625 5766
rect 13640 5761 13670 5772
rect 13702 5768 13764 5784
rect 13702 5766 13748 5768
rect 13702 5750 13764 5766
rect 13776 5750 13782 5798
rect 13785 5790 13865 5798
rect 13785 5788 13804 5790
rect 13819 5788 13853 5790
rect 13785 5772 13865 5788
rect 13785 5750 13804 5772
rect 13819 5756 13849 5772
rect 13877 5766 13883 5840
rect 13886 5766 13905 5910
rect 13920 5766 13926 5910
rect 13935 5840 13948 5910
rect 14000 5906 14022 5910
rect 13993 5884 14022 5898
rect 14075 5884 14091 5898
rect 14129 5894 14135 5896
rect 14142 5894 14250 5910
rect 14257 5894 14263 5896
rect 14271 5894 14286 5910
rect 14352 5904 14371 5907
rect 13993 5882 14091 5884
rect 14118 5882 14286 5894
rect 14301 5884 14317 5898
rect 14352 5885 14374 5904
rect 14384 5898 14400 5899
rect 14383 5896 14400 5898
rect 14384 5891 14400 5896
rect 14374 5884 14380 5885
rect 14383 5884 14412 5891
rect 14301 5883 14412 5884
rect 14301 5882 14418 5883
rect 13977 5874 14028 5882
rect 14075 5874 14109 5882
rect 13977 5862 14002 5874
rect 14009 5862 14028 5874
rect 14082 5872 14109 5874
rect 14118 5872 14339 5882
rect 14374 5879 14380 5882
rect 14082 5868 14339 5872
rect 13977 5854 14028 5862
rect 14075 5854 14339 5868
rect 14383 5874 14418 5882
rect 13929 5806 13948 5840
rect 13993 5846 14022 5854
rect 13993 5840 14010 5846
rect 13993 5838 14027 5840
rect 14075 5838 14091 5854
rect 14092 5844 14300 5854
rect 14301 5844 14317 5854
rect 14365 5850 14380 5865
rect 14383 5862 14384 5874
rect 14391 5862 14418 5874
rect 14383 5854 14418 5862
rect 14383 5853 14412 5854
rect 14103 5840 14317 5844
rect 14118 5838 14317 5840
rect 14352 5840 14365 5850
rect 14383 5840 14400 5853
rect 14352 5838 14400 5840
rect 13994 5834 14027 5838
rect 13990 5832 14027 5834
rect 13990 5831 14057 5832
rect 13990 5826 14021 5831
rect 14027 5826 14057 5831
rect 13990 5822 14057 5826
rect 13963 5819 14057 5822
rect 13963 5812 14012 5819
rect 13963 5806 13993 5812
rect 14012 5807 14017 5812
rect 13929 5790 14009 5806
rect 14021 5798 14057 5819
rect 14118 5814 14307 5838
rect 14352 5837 14399 5838
rect 14365 5832 14399 5837
rect 14133 5811 14307 5814
rect 14126 5808 14307 5811
rect 14335 5831 14399 5832
rect 13929 5788 13948 5790
rect 13963 5788 13997 5790
rect 13929 5772 14009 5788
rect 13929 5766 13948 5772
rect 13645 5740 13748 5750
rect 13599 5738 13748 5740
rect 13769 5738 13804 5750
rect 13438 5736 13600 5738
rect 13450 5716 13469 5736
rect 13484 5734 13514 5736
rect 13333 5708 13374 5716
rect 13456 5712 13469 5716
rect 13521 5720 13600 5736
rect 13632 5736 13804 5738
rect 13632 5720 13711 5736
rect 13718 5734 13748 5736
rect 13296 5698 13325 5708
rect 13339 5698 13368 5708
rect 13383 5698 13413 5712
rect 13456 5698 13499 5712
rect 13521 5708 13711 5720
rect 13776 5716 13782 5736
rect 13506 5698 13536 5708
rect 13537 5698 13695 5708
rect 13699 5698 13729 5708
rect 13733 5698 13763 5712
rect 13791 5698 13804 5736
rect 13876 5750 13905 5766
rect 13919 5750 13948 5766
rect 13963 5756 13993 5772
rect 14021 5750 14027 5798
rect 14030 5792 14049 5798
rect 14064 5792 14094 5800
rect 14030 5784 14094 5792
rect 14030 5768 14110 5784
rect 14126 5777 14188 5808
rect 14204 5777 14266 5808
rect 14335 5806 14384 5831
rect 14399 5806 14429 5822
rect 14298 5792 14328 5800
rect 14335 5798 14445 5806
rect 14298 5784 14343 5792
rect 14030 5766 14049 5768
rect 14064 5766 14110 5768
rect 14030 5750 14110 5766
rect 14137 5764 14172 5777
rect 14213 5774 14250 5777
rect 14213 5772 14255 5774
rect 14142 5761 14172 5764
rect 14151 5757 14158 5761
rect 14158 5756 14159 5757
rect 14117 5750 14127 5756
rect 13876 5742 13911 5750
rect 13876 5716 13877 5742
rect 13884 5716 13911 5742
rect 13819 5698 13849 5712
rect 13876 5708 13911 5716
rect 13913 5742 13954 5750
rect 13913 5716 13928 5742
rect 13935 5716 13954 5742
rect 14018 5738 14049 5750
rect 14064 5738 14167 5750
rect 14179 5740 14205 5766
rect 14220 5761 14250 5772
rect 14282 5768 14344 5784
rect 14282 5766 14328 5768
rect 14282 5750 14344 5766
rect 14356 5750 14362 5798
rect 14365 5790 14445 5798
rect 14365 5788 14384 5790
rect 14399 5788 14433 5790
rect 14365 5772 14445 5788
rect 14365 5750 14384 5772
rect 14399 5756 14429 5772
rect 14457 5766 14463 5840
rect 14466 5766 14485 5910
rect 14500 5766 14506 5910
rect 14515 5840 14528 5910
rect 14580 5906 14602 5910
rect 14573 5884 14602 5898
rect 14655 5884 14671 5898
rect 14709 5894 14715 5896
rect 14722 5894 14830 5910
rect 14837 5894 14843 5896
rect 14851 5894 14866 5910
rect 14932 5904 14951 5907
rect 14573 5882 14671 5884
rect 14698 5882 14866 5894
rect 14881 5884 14897 5898
rect 14932 5885 14954 5904
rect 14964 5898 14980 5899
rect 14963 5896 14980 5898
rect 14964 5891 14980 5896
rect 14954 5884 14960 5885
rect 14963 5884 14992 5891
rect 14881 5883 14992 5884
rect 14881 5882 14998 5883
rect 14557 5874 14608 5882
rect 14655 5874 14689 5882
rect 14557 5862 14582 5874
rect 14589 5862 14608 5874
rect 14662 5872 14689 5874
rect 14698 5872 14919 5882
rect 14954 5879 14960 5882
rect 14662 5868 14919 5872
rect 14557 5854 14608 5862
rect 14655 5854 14919 5868
rect 14963 5874 14998 5882
rect 14509 5806 14528 5840
rect 14573 5846 14602 5854
rect 14573 5840 14590 5846
rect 14573 5838 14607 5840
rect 14655 5838 14671 5854
rect 14672 5844 14880 5854
rect 14881 5844 14897 5854
rect 14945 5850 14960 5865
rect 14963 5862 14964 5874
rect 14971 5862 14998 5874
rect 14963 5854 14998 5862
rect 14963 5853 14992 5854
rect 14683 5840 14897 5844
rect 14698 5838 14897 5840
rect 14932 5840 14945 5850
rect 14963 5840 14980 5853
rect 14932 5838 14980 5840
rect 14574 5834 14607 5838
rect 14570 5832 14607 5834
rect 14570 5831 14637 5832
rect 14570 5826 14601 5831
rect 14607 5826 14637 5831
rect 14570 5822 14637 5826
rect 14543 5819 14637 5822
rect 14543 5812 14592 5819
rect 14543 5806 14573 5812
rect 14592 5807 14597 5812
rect 14509 5790 14589 5806
rect 14601 5798 14637 5819
rect 14698 5814 14887 5838
rect 14932 5837 14979 5838
rect 14945 5832 14979 5837
rect 14713 5811 14887 5814
rect 14706 5808 14887 5811
rect 14915 5831 14979 5832
rect 14509 5788 14528 5790
rect 14543 5788 14577 5790
rect 14509 5772 14589 5788
rect 14509 5766 14528 5772
rect 14225 5740 14328 5750
rect 14179 5738 14328 5740
rect 14349 5738 14384 5750
rect 14018 5736 14180 5738
rect 14030 5716 14049 5736
rect 14064 5734 14094 5736
rect 13913 5708 13954 5716
rect 14036 5712 14049 5716
rect 14101 5720 14180 5736
rect 14212 5736 14384 5738
rect 14212 5720 14291 5736
rect 14298 5734 14328 5736
rect 13876 5698 13905 5708
rect 13919 5698 13948 5708
rect 13963 5698 13993 5712
rect 14036 5698 14079 5712
rect 14101 5708 14291 5720
rect 14356 5716 14362 5736
rect 14086 5698 14116 5708
rect 14117 5698 14275 5708
rect 14279 5698 14309 5708
rect 14313 5698 14343 5712
rect 14371 5698 14384 5736
rect 14456 5750 14485 5766
rect 14499 5750 14528 5766
rect 14543 5756 14573 5772
rect 14601 5750 14607 5798
rect 14610 5792 14629 5798
rect 14644 5792 14674 5800
rect 14610 5784 14674 5792
rect 14610 5768 14690 5784
rect 14706 5777 14768 5808
rect 14784 5777 14846 5808
rect 14915 5806 14964 5831
rect 14979 5806 15009 5822
rect 14878 5792 14908 5800
rect 14915 5798 15025 5806
rect 14878 5784 14923 5792
rect 14610 5766 14629 5768
rect 14644 5766 14690 5768
rect 14610 5750 14690 5766
rect 14717 5764 14752 5777
rect 14793 5774 14830 5777
rect 14793 5772 14835 5774
rect 14722 5761 14752 5764
rect 14731 5757 14738 5761
rect 14738 5756 14739 5757
rect 14697 5750 14707 5756
rect 14456 5742 14491 5750
rect 14456 5716 14457 5742
rect 14464 5716 14491 5742
rect 14399 5698 14429 5712
rect 14456 5708 14491 5716
rect 14493 5742 14534 5750
rect 14493 5716 14508 5742
rect 14515 5716 14534 5742
rect 14598 5738 14629 5750
rect 14644 5738 14747 5750
rect 14759 5740 14785 5766
rect 14800 5761 14830 5772
rect 14862 5768 14924 5784
rect 14862 5766 14908 5768
rect 14862 5750 14924 5766
rect 14936 5750 14942 5798
rect 14945 5790 15025 5798
rect 14945 5788 14964 5790
rect 14979 5788 15013 5790
rect 14945 5772 15025 5788
rect 14945 5750 14964 5772
rect 14979 5756 15009 5772
rect 15037 5766 15043 5840
rect 15046 5766 15065 5910
rect 15080 5766 15086 5910
rect 15095 5840 15108 5910
rect 15160 5906 15182 5910
rect 15153 5884 15182 5898
rect 15235 5884 15251 5898
rect 15289 5894 15295 5896
rect 15302 5894 15410 5910
rect 15417 5894 15423 5896
rect 15431 5894 15446 5910
rect 15512 5904 15531 5907
rect 15153 5882 15251 5884
rect 15278 5882 15446 5894
rect 15461 5884 15477 5898
rect 15512 5885 15534 5904
rect 15544 5898 15560 5899
rect 15543 5896 15560 5898
rect 15544 5891 15560 5896
rect 15534 5884 15540 5885
rect 15543 5884 15572 5891
rect 15461 5883 15572 5884
rect 15461 5882 15578 5883
rect 15137 5874 15188 5882
rect 15235 5874 15269 5882
rect 15137 5862 15162 5874
rect 15169 5862 15188 5874
rect 15242 5872 15269 5874
rect 15278 5872 15499 5882
rect 15534 5879 15540 5882
rect 15242 5868 15499 5872
rect 15137 5854 15188 5862
rect 15235 5854 15499 5868
rect 15543 5874 15578 5882
rect 15089 5806 15108 5840
rect 15153 5846 15182 5854
rect 15153 5840 15170 5846
rect 15153 5838 15187 5840
rect 15235 5838 15251 5854
rect 15252 5844 15460 5854
rect 15461 5844 15477 5854
rect 15525 5850 15540 5865
rect 15543 5862 15544 5874
rect 15551 5862 15578 5874
rect 15543 5854 15578 5862
rect 15543 5853 15572 5854
rect 15263 5840 15477 5844
rect 15278 5838 15477 5840
rect 15512 5840 15525 5850
rect 15543 5840 15560 5853
rect 15512 5838 15560 5840
rect 15154 5834 15187 5838
rect 15150 5832 15187 5834
rect 15150 5831 15217 5832
rect 15150 5826 15181 5831
rect 15187 5826 15217 5831
rect 15150 5822 15217 5826
rect 15123 5819 15217 5822
rect 15123 5812 15172 5819
rect 15123 5806 15153 5812
rect 15172 5807 15177 5812
rect 15089 5790 15169 5806
rect 15181 5798 15217 5819
rect 15278 5814 15467 5838
rect 15512 5837 15559 5838
rect 15525 5832 15559 5837
rect 15293 5811 15467 5814
rect 15286 5808 15467 5811
rect 15495 5831 15559 5832
rect 15089 5788 15108 5790
rect 15123 5788 15157 5790
rect 15089 5772 15169 5788
rect 15089 5766 15108 5772
rect 14805 5740 14908 5750
rect 14759 5738 14908 5740
rect 14929 5738 14964 5750
rect 14598 5736 14760 5738
rect 14610 5716 14629 5736
rect 14644 5734 14674 5736
rect 14493 5708 14534 5716
rect 14616 5712 14629 5716
rect 14681 5720 14760 5736
rect 14792 5736 14964 5738
rect 14792 5720 14871 5736
rect 14878 5734 14908 5736
rect 14456 5698 14485 5708
rect 14499 5698 14528 5708
rect 14543 5698 14573 5712
rect 14616 5698 14659 5712
rect 14681 5708 14871 5720
rect 14936 5716 14942 5736
rect 14666 5698 14696 5708
rect 14697 5698 14855 5708
rect 14859 5698 14889 5708
rect 14893 5698 14923 5712
rect 14951 5698 14964 5736
rect 15036 5750 15065 5766
rect 15079 5750 15108 5766
rect 15123 5756 15153 5772
rect 15181 5750 15187 5798
rect 15190 5792 15209 5798
rect 15224 5792 15254 5800
rect 15190 5784 15254 5792
rect 15190 5768 15270 5784
rect 15286 5777 15348 5808
rect 15364 5777 15426 5808
rect 15495 5806 15544 5831
rect 15559 5806 15589 5822
rect 15458 5792 15488 5800
rect 15495 5798 15605 5806
rect 15458 5784 15503 5792
rect 15190 5766 15209 5768
rect 15224 5766 15270 5768
rect 15190 5750 15270 5766
rect 15297 5764 15332 5777
rect 15373 5774 15410 5777
rect 15373 5772 15415 5774
rect 15302 5761 15332 5764
rect 15311 5757 15318 5761
rect 15318 5756 15319 5757
rect 15277 5750 15287 5756
rect 15036 5742 15071 5750
rect 15036 5716 15037 5742
rect 15044 5716 15071 5742
rect 14979 5698 15009 5712
rect 15036 5708 15071 5716
rect 15073 5742 15114 5750
rect 15073 5716 15088 5742
rect 15095 5716 15114 5742
rect 15178 5738 15209 5750
rect 15224 5738 15327 5750
rect 15339 5740 15365 5766
rect 15380 5761 15410 5772
rect 15442 5768 15504 5784
rect 15442 5766 15488 5768
rect 15442 5750 15504 5766
rect 15516 5750 15522 5798
rect 15525 5790 15605 5798
rect 15525 5788 15544 5790
rect 15559 5788 15593 5790
rect 15525 5772 15605 5788
rect 15525 5750 15544 5772
rect 15559 5756 15589 5772
rect 15617 5766 15623 5840
rect 15626 5766 15645 5910
rect 15660 5766 15666 5910
rect 15675 5840 15688 5910
rect 15740 5906 15762 5910
rect 15733 5884 15762 5898
rect 15815 5884 15831 5898
rect 15869 5894 15875 5896
rect 15882 5894 15990 5910
rect 15997 5894 16003 5896
rect 16011 5894 16026 5910
rect 16092 5904 16111 5907
rect 15733 5882 15831 5884
rect 15858 5882 16026 5894
rect 16041 5884 16057 5898
rect 16092 5885 16114 5904
rect 16124 5898 16140 5899
rect 16123 5896 16140 5898
rect 16124 5891 16140 5896
rect 16114 5884 16120 5885
rect 16123 5884 16152 5891
rect 16041 5883 16152 5884
rect 16041 5882 16158 5883
rect 15717 5874 15768 5882
rect 15815 5874 15849 5882
rect 15717 5862 15742 5874
rect 15749 5862 15768 5874
rect 15822 5872 15849 5874
rect 15858 5872 16079 5882
rect 16114 5879 16120 5882
rect 15822 5868 16079 5872
rect 15717 5854 15768 5862
rect 15815 5854 16079 5868
rect 16123 5874 16158 5882
rect 15669 5806 15688 5840
rect 15733 5846 15762 5854
rect 15733 5840 15750 5846
rect 15733 5838 15767 5840
rect 15815 5838 15831 5854
rect 15832 5844 16040 5854
rect 16041 5844 16057 5854
rect 16105 5850 16120 5865
rect 16123 5862 16124 5874
rect 16131 5862 16158 5874
rect 16123 5854 16158 5862
rect 16123 5853 16152 5854
rect 15843 5840 16057 5844
rect 15858 5838 16057 5840
rect 16092 5840 16105 5850
rect 16123 5840 16140 5853
rect 16092 5838 16140 5840
rect 15734 5834 15767 5838
rect 15730 5832 15767 5834
rect 15730 5831 15797 5832
rect 15730 5826 15761 5831
rect 15767 5826 15797 5831
rect 15730 5822 15797 5826
rect 15703 5819 15797 5822
rect 15703 5812 15752 5819
rect 15703 5806 15733 5812
rect 15752 5807 15757 5812
rect 15669 5790 15749 5806
rect 15761 5798 15797 5819
rect 15858 5814 16047 5838
rect 16092 5837 16139 5838
rect 16105 5832 16139 5837
rect 15873 5811 16047 5814
rect 15866 5808 16047 5811
rect 16075 5831 16139 5832
rect 15669 5788 15688 5790
rect 15703 5788 15737 5790
rect 15669 5772 15749 5788
rect 15669 5766 15688 5772
rect 15385 5740 15488 5750
rect 15339 5738 15488 5740
rect 15509 5738 15544 5750
rect 15178 5736 15340 5738
rect 15190 5716 15209 5736
rect 15224 5734 15254 5736
rect 15073 5708 15114 5716
rect 15196 5712 15209 5716
rect 15261 5720 15340 5736
rect 15372 5736 15544 5738
rect 15372 5720 15451 5736
rect 15458 5734 15488 5736
rect 15036 5698 15065 5708
rect 15079 5698 15108 5708
rect 15123 5698 15153 5712
rect 15196 5698 15239 5712
rect 15261 5708 15451 5720
rect 15516 5716 15522 5736
rect 15246 5698 15276 5708
rect 15277 5698 15435 5708
rect 15439 5698 15469 5708
rect 15473 5698 15503 5712
rect 15531 5698 15544 5736
rect 15616 5750 15645 5766
rect 15659 5750 15688 5766
rect 15703 5756 15733 5772
rect 15761 5750 15767 5798
rect 15770 5792 15789 5798
rect 15804 5792 15834 5800
rect 15770 5784 15834 5792
rect 15770 5768 15850 5784
rect 15866 5777 15928 5808
rect 15944 5777 16006 5808
rect 16075 5806 16124 5831
rect 16139 5806 16169 5822
rect 16038 5792 16068 5800
rect 16075 5798 16185 5806
rect 16038 5784 16083 5792
rect 15770 5766 15789 5768
rect 15804 5766 15850 5768
rect 15770 5750 15850 5766
rect 15877 5764 15912 5777
rect 15953 5774 15990 5777
rect 15953 5772 15995 5774
rect 15882 5761 15912 5764
rect 15891 5757 15898 5761
rect 15898 5756 15899 5757
rect 15857 5750 15867 5756
rect 15616 5742 15651 5750
rect 15616 5716 15617 5742
rect 15624 5716 15651 5742
rect 15559 5698 15589 5712
rect 15616 5708 15651 5716
rect 15653 5742 15694 5750
rect 15653 5716 15668 5742
rect 15675 5716 15694 5742
rect 15758 5738 15789 5750
rect 15804 5738 15907 5750
rect 15919 5740 15945 5766
rect 15960 5761 15990 5772
rect 16022 5768 16084 5784
rect 16022 5766 16068 5768
rect 16022 5750 16084 5766
rect 16096 5750 16102 5798
rect 16105 5790 16185 5798
rect 16105 5788 16124 5790
rect 16139 5788 16173 5790
rect 16105 5772 16185 5788
rect 16105 5750 16124 5772
rect 16139 5756 16169 5772
rect 16197 5766 16203 5840
rect 16206 5766 16225 5910
rect 16240 5766 16246 5910
rect 16255 5840 16268 5910
rect 16320 5906 16342 5910
rect 16313 5884 16342 5898
rect 16395 5884 16411 5898
rect 16449 5894 16455 5896
rect 16462 5894 16570 5910
rect 16577 5894 16583 5896
rect 16591 5894 16606 5910
rect 16672 5904 16691 5907
rect 16313 5882 16411 5884
rect 16438 5882 16606 5894
rect 16621 5884 16637 5898
rect 16672 5885 16694 5904
rect 16704 5898 16720 5899
rect 16703 5896 16720 5898
rect 16704 5891 16720 5896
rect 16694 5884 16700 5885
rect 16703 5884 16732 5891
rect 16621 5883 16732 5884
rect 16621 5882 16738 5883
rect 16297 5874 16348 5882
rect 16395 5874 16429 5882
rect 16297 5862 16322 5874
rect 16329 5862 16348 5874
rect 16402 5872 16429 5874
rect 16438 5872 16659 5882
rect 16694 5879 16700 5882
rect 16402 5868 16659 5872
rect 16297 5854 16348 5862
rect 16395 5854 16659 5868
rect 16703 5874 16738 5882
rect 16249 5806 16268 5840
rect 16313 5846 16342 5854
rect 16313 5840 16330 5846
rect 16313 5838 16347 5840
rect 16395 5838 16411 5854
rect 16412 5844 16620 5854
rect 16621 5844 16637 5854
rect 16685 5850 16700 5865
rect 16703 5862 16704 5874
rect 16711 5862 16738 5874
rect 16703 5854 16738 5862
rect 16703 5853 16732 5854
rect 16423 5840 16637 5844
rect 16438 5838 16637 5840
rect 16672 5840 16685 5850
rect 16703 5840 16720 5853
rect 16672 5838 16720 5840
rect 16314 5834 16347 5838
rect 16310 5832 16347 5834
rect 16310 5831 16377 5832
rect 16310 5826 16341 5831
rect 16347 5826 16377 5831
rect 16310 5822 16377 5826
rect 16283 5819 16377 5822
rect 16283 5812 16332 5819
rect 16283 5806 16313 5812
rect 16332 5807 16337 5812
rect 16249 5790 16329 5806
rect 16341 5798 16377 5819
rect 16438 5814 16627 5838
rect 16672 5837 16719 5838
rect 16685 5832 16719 5837
rect 16453 5811 16627 5814
rect 16446 5808 16627 5811
rect 16655 5831 16719 5832
rect 16249 5788 16268 5790
rect 16283 5788 16317 5790
rect 16249 5772 16329 5788
rect 16249 5766 16268 5772
rect 15965 5740 16068 5750
rect 15919 5738 16068 5740
rect 16089 5738 16124 5750
rect 15758 5736 15920 5738
rect 15770 5716 15789 5736
rect 15804 5734 15834 5736
rect 15653 5708 15694 5716
rect 15776 5712 15789 5716
rect 15841 5720 15920 5736
rect 15952 5736 16124 5738
rect 15952 5720 16031 5736
rect 16038 5734 16068 5736
rect 15616 5698 15645 5708
rect 15659 5698 15688 5708
rect 15703 5698 15733 5712
rect 15776 5698 15819 5712
rect 15841 5708 16031 5720
rect 16096 5716 16102 5736
rect 15826 5698 15856 5708
rect 15857 5698 16015 5708
rect 16019 5698 16049 5708
rect 16053 5698 16083 5712
rect 16111 5698 16124 5736
rect 16196 5750 16225 5766
rect 16239 5750 16268 5766
rect 16283 5756 16313 5772
rect 16341 5750 16347 5798
rect 16350 5792 16369 5798
rect 16384 5792 16414 5800
rect 16350 5784 16414 5792
rect 16350 5768 16430 5784
rect 16446 5777 16508 5808
rect 16524 5777 16586 5808
rect 16655 5806 16704 5831
rect 16719 5806 16749 5822
rect 16618 5792 16648 5800
rect 16655 5798 16765 5806
rect 16618 5784 16663 5792
rect 16350 5766 16369 5768
rect 16384 5766 16430 5768
rect 16350 5750 16430 5766
rect 16457 5764 16492 5777
rect 16533 5774 16570 5777
rect 16533 5772 16575 5774
rect 16462 5761 16492 5764
rect 16471 5757 16478 5761
rect 16478 5756 16479 5757
rect 16437 5750 16447 5756
rect 16196 5742 16231 5750
rect 16196 5716 16197 5742
rect 16204 5716 16231 5742
rect 16139 5698 16169 5712
rect 16196 5708 16231 5716
rect 16233 5742 16274 5750
rect 16233 5716 16248 5742
rect 16255 5716 16274 5742
rect 16338 5738 16369 5750
rect 16384 5738 16487 5750
rect 16499 5740 16525 5766
rect 16540 5761 16570 5772
rect 16602 5768 16664 5784
rect 16602 5766 16648 5768
rect 16602 5750 16664 5766
rect 16676 5750 16682 5798
rect 16685 5790 16765 5798
rect 16685 5788 16704 5790
rect 16719 5788 16753 5790
rect 16685 5772 16765 5788
rect 16685 5750 16704 5772
rect 16719 5756 16749 5772
rect 16777 5766 16783 5840
rect 16786 5766 16805 5910
rect 16820 5766 16826 5910
rect 16835 5840 16848 5910
rect 16900 5906 16922 5910
rect 16893 5884 16922 5898
rect 16975 5884 16991 5898
rect 17029 5894 17035 5896
rect 17042 5894 17150 5910
rect 17157 5894 17163 5896
rect 17171 5894 17186 5910
rect 17252 5904 17271 5907
rect 16893 5882 16991 5884
rect 17018 5882 17186 5894
rect 17201 5884 17217 5898
rect 17252 5885 17274 5904
rect 17284 5898 17300 5899
rect 17283 5896 17300 5898
rect 17284 5891 17300 5896
rect 17274 5884 17280 5885
rect 17283 5884 17312 5891
rect 17201 5883 17312 5884
rect 17201 5882 17318 5883
rect 16877 5874 16928 5882
rect 16975 5874 17009 5882
rect 16877 5862 16902 5874
rect 16909 5862 16928 5874
rect 16982 5872 17009 5874
rect 17018 5872 17239 5882
rect 17274 5879 17280 5882
rect 16982 5868 17239 5872
rect 16877 5854 16928 5862
rect 16975 5854 17239 5868
rect 17283 5874 17318 5882
rect 16829 5806 16848 5840
rect 16893 5846 16922 5854
rect 16893 5840 16910 5846
rect 16893 5838 16927 5840
rect 16975 5838 16991 5854
rect 16992 5844 17200 5854
rect 17201 5844 17217 5854
rect 17265 5850 17280 5865
rect 17283 5862 17284 5874
rect 17291 5862 17318 5874
rect 17283 5854 17318 5862
rect 17283 5853 17312 5854
rect 17003 5840 17217 5844
rect 17018 5838 17217 5840
rect 17252 5840 17265 5850
rect 17283 5840 17300 5853
rect 17252 5838 17300 5840
rect 16894 5834 16927 5838
rect 16890 5832 16927 5834
rect 16890 5831 16957 5832
rect 16890 5826 16921 5831
rect 16927 5826 16957 5831
rect 16890 5822 16957 5826
rect 16863 5819 16957 5822
rect 16863 5812 16912 5819
rect 16863 5806 16893 5812
rect 16912 5807 16917 5812
rect 16829 5790 16909 5806
rect 16921 5798 16957 5819
rect 17018 5814 17207 5838
rect 17252 5837 17299 5838
rect 17265 5832 17299 5837
rect 17033 5811 17207 5814
rect 17026 5808 17207 5811
rect 17235 5831 17299 5832
rect 16829 5788 16848 5790
rect 16863 5788 16897 5790
rect 16829 5772 16909 5788
rect 16829 5766 16848 5772
rect 16545 5740 16648 5750
rect 16499 5738 16648 5740
rect 16669 5738 16704 5750
rect 16338 5736 16500 5738
rect 16350 5716 16369 5736
rect 16384 5734 16414 5736
rect 16233 5708 16274 5716
rect 16356 5712 16369 5716
rect 16421 5720 16500 5736
rect 16532 5736 16704 5738
rect 16532 5720 16611 5736
rect 16618 5734 16648 5736
rect 16196 5698 16225 5708
rect 16239 5698 16268 5708
rect 16283 5698 16313 5712
rect 16356 5698 16399 5712
rect 16421 5708 16611 5720
rect 16676 5716 16682 5736
rect 16406 5698 16436 5708
rect 16437 5698 16595 5708
rect 16599 5698 16629 5708
rect 16633 5698 16663 5712
rect 16691 5698 16704 5736
rect 16776 5750 16805 5766
rect 16819 5750 16848 5766
rect 16863 5756 16893 5772
rect 16921 5750 16927 5798
rect 16930 5792 16949 5798
rect 16964 5792 16994 5800
rect 16930 5784 16994 5792
rect 16930 5768 17010 5784
rect 17026 5777 17088 5808
rect 17104 5777 17166 5808
rect 17235 5806 17284 5831
rect 17299 5806 17329 5822
rect 17198 5792 17228 5800
rect 17235 5798 17345 5806
rect 17198 5784 17243 5792
rect 16930 5766 16949 5768
rect 16964 5766 17010 5768
rect 16930 5750 17010 5766
rect 17037 5764 17072 5777
rect 17113 5774 17150 5777
rect 17113 5772 17155 5774
rect 17042 5761 17072 5764
rect 17051 5757 17058 5761
rect 17058 5756 17059 5757
rect 17017 5750 17027 5756
rect 16776 5742 16811 5750
rect 16776 5716 16777 5742
rect 16784 5716 16811 5742
rect 16719 5698 16749 5712
rect 16776 5708 16811 5716
rect 16813 5742 16854 5750
rect 16813 5716 16828 5742
rect 16835 5716 16854 5742
rect 16918 5738 16949 5750
rect 16964 5738 17067 5750
rect 17079 5740 17105 5766
rect 17120 5761 17150 5772
rect 17182 5768 17244 5784
rect 17182 5766 17228 5768
rect 17182 5750 17244 5766
rect 17256 5750 17262 5798
rect 17265 5790 17345 5798
rect 17265 5788 17284 5790
rect 17299 5788 17333 5790
rect 17265 5772 17345 5788
rect 17265 5750 17284 5772
rect 17299 5756 17329 5772
rect 17357 5766 17363 5840
rect 17366 5766 17385 5910
rect 17400 5766 17406 5910
rect 17415 5840 17428 5910
rect 17480 5906 17502 5910
rect 17473 5884 17502 5898
rect 17555 5884 17571 5898
rect 17609 5894 17615 5896
rect 17622 5894 17730 5910
rect 17737 5894 17743 5896
rect 17751 5894 17766 5910
rect 17832 5904 17851 5907
rect 17473 5882 17571 5884
rect 17598 5882 17766 5894
rect 17781 5884 17797 5898
rect 17832 5885 17854 5904
rect 17864 5898 17880 5899
rect 17863 5896 17880 5898
rect 17864 5891 17880 5896
rect 17854 5884 17860 5885
rect 17863 5884 17892 5891
rect 17781 5883 17892 5884
rect 17781 5882 17898 5883
rect 17457 5874 17508 5882
rect 17555 5874 17589 5882
rect 17457 5862 17482 5874
rect 17489 5862 17508 5874
rect 17562 5872 17589 5874
rect 17598 5872 17819 5882
rect 17854 5879 17860 5882
rect 17562 5868 17819 5872
rect 17457 5854 17508 5862
rect 17555 5854 17819 5868
rect 17863 5874 17898 5882
rect 17409 5806 17428 5840
rect 17473 5846 17502 5854
rect 17473 5840 17490 5846
rect 17473 5838 17507 5840
rect 17555 5838 17571 5854
rect 17572 5844 17780 5854
rect 17781 5844 17797 5854
rect 17845 5850 17860 5865
rect 17863 5862 17864 5874
rect 17871 5862 17898 5874
rect 17863 5854 17898 5862
rect 17863 5853 17892 5854
rect 17583 5840 17797 5844
rect 17598 5838 17797 5840
rect 17832 5840 17845 5850
rect 17863 5840 17880 5853
rect 17832 5838 17880 5840
rect 17474 5834 17507 5838
rect 17470 5832 17507 5834
rect 17470 5831 17537 5832
rect 17470 5826 17501 5831
rect 17507 5826 17537 5831
rect 17470 5822 17537 5826
rect 17443 5819 17537 5822
rect 17443 5812 17492 5819
rect 17443 5806 17473 5812
rect 17492 5807 17497 5812
rect 17409 5790 17489 5806
rect 17501 5798 17537 5819
rect 17598 5814 17787 5838
rect 17832 5837 17879 5838
rect 17845 5832 17879 5837
rect 17613 5811 17787 5814
rect 17606 5808 17787 5811
rect 17815 5831 17879 5832
rect 17409 5788 17428 5790
rect 17443 5788 17477 5790
rect 17409 5772 17489 5788
rect 17409 5766 17428 5772
rect 17125 5740 17228 5750
rect 17079 5738 17228 5740
rect 17249 5738 17284 5750
rect 16918 5736 17080 5738
rect 16930 5716 16949 5736
rect 16964 5734 16994 5736
rect 16813 5708 16854 5716
rect 16936 5712 16949 5716
rect 17001 5720 17080 5736
rect 17112 5736 17284 5738
rect 17112 5720 17191 5736
rect 17198 5734 17228 5736
rect 16776 5698 16805 5708
rect 16819 5698 16848 5708
rect 16863 5698 16893 5712
rect 16936 5698 16979 5712
rect 17001 5708 17191 5720
rect 17256 5716 17262 5736
rect 16986 5698 17016 5708
rect 17017 5698 17175 5708
rect 17179 5698 17209 5708
rect 17213 5698 17243 5712
rect 17271 5698 17284 5736
rect 17356 5750 17385 5766
rect 17399 5750 17428 5766
rect 17443 5756 17473 5772
rect 17501 5750 17507 5798
rect 17510 5792 17529 5798
rect 17544 5792 17574 5800
rect 17510 5784 17574 5792
rect 17510 5768 17590 5784
rect 17606 5777 17668 5808
rect 17684 5777 17746 5808
rect 17815 5806 17864 5831
rect 17879 5806 17909 5822
rect 17778 5792 17808 5800
rect 17815 5798 17925 5806
rect 17778 5784 17823 5792
rect 17510 5766 17529 5768
rect 17544 5766 17590 5768
rect 17510 5750 17590 5766
rect 17617 5764 17652 5777
rect 17693 5774 17730 5777
rect 17693 5772 17735 5774
rect 17622 5761 17652 5764
rect 17631 5757 17638 5761
rect 17638 5756 17639 5757
rect 17597 5750 17607 5756
rect 17356 5742 17391 5750
rect 17356 5716 17357 5742
rect 17364 5716 17391 5742
rect 17299 5698 17329 5712
rect 17356 5708 17391 5716
rect 17393 5742 17434 5750
rect 17393 5716 17408 5742
rect 17415 5716 17434 5742
rect 17498 5738 17529 5750
rect 17544 5738 17647 5750
rect 17659 5740 17685 5766
rect 17700 5761 17730 5772
rect 17762 5768 17824 5784
rect 17762 5766 17808 5768
rect 17762 5750 17824 5766
rect 17836 5750 17842 5798
rect 17845 5790 17925 5798
rect 17845 5788 17864 5790
rect 17879 5788 17913 5790
rect 17845 5772 17925 5788
rect 17845 5750 17864 5772
rect 17879 5756 17909 5772
rect 17937 5766 17943 5840
rect 17946 5766 17965 5910
rect 17980 5766 17986 5910
rect 17995 5840 18008 5910
rect 18060 5906 18082 5910
rect 18053 5884 18082 5898
rect 18135 5884 18151 5898
rect 18189 5894 18195 5896
rect 18202 5894 18310 5910
rect 18317 5894 18323 5896
rect 18331 5894 18346 5910
rect 18412 5904 18431 5907
rect 18053 5882 18151 5884
rect 18178 5882 18346 5894
rect 18361 5884 18377 5898
rect 18412 5885 18434 5904
rect 18444 5898 18460 5899
rect 18443 5896 18460 5898
rect 18444 5891 18460 5896
rect 18434 5884 18440 5885
rect 18443 5884 18472 5891
rect 18361 5883 18472 5884
rect 18361 5882 18478 5883
rect 18037 5874 18088 5882
rect 18135 5874 18169 5882
rect 18037 5862 18062 5874
rect 18069 5862 18088 5874
rect 18142 5872 18169 5874
rect 18178 5872 18399 5882
rect 18434 5879 18440 5882
rect 18142 5868 18399 5872
rect 18037 5854 18088 5862
rect 18135 5854 18399 5868
rect 18443 5874 18478 5882
rect 17989 5806 18008 5840
rect 18053 5846 18082 5854
rect 18053 5840 18070 5846
rect 18053 5838 18087 5840
rect 18135 5838 18151 5854
rect 18152 5844 18360 5854
rect 18361 5844 18377 5854
rect 18425 5850 18440 5865
rect 18443 5862 18444 5874
rect 18451 5862 18478 5874
rect 18443 5854 18478 5862
rect 18443 5853 18472 5854
rect 18163 5840 18377 5844
rect 18178 5838 18377 5840
rect 18412 5840 18425 5850
rect 18443 5840 18460 5853
rect 18412 5838 18460 5840
rect 18054 5834 18087 5838
rect 18050 5832 18087 5834
rect 18050 5831 18117 5832
rect 18050 5826 18081 5831
rect 18087 5826 18117 5831
rect 18050 5822 18117 5826
rect 18023 5819 18117 5822
rect 18023 5812 18072 5819
rect 18023 5806 18053 5812
rect 18072 5807 18077 5812
rect 17989 5790 18069 5806
rect 18081 5798 18117 5819
rect 18178 5814 18367 5838
rect 18412 5837 18459 5838
rect 18425 5832 18459 5837
rect 18193 5811 18367 5814
rect 18186 5808 18367 5811
rect 18395 5831 18459 5832
rect 17989 5788 18008 5790
rect 18023 5788 18057 5790
rect 17989 5772 18069 5788
rect 17989 5766 18008 5772
rect 17705 5740 17808 5750
rect 17659 5738 17808 5740
rect 17829 5738 17864 5750
rect 17498 5736 17660 5738
rect 17510 5716 17529 5736
rect 17544 5734 17574 5736
rect 17393 5708 17434 5716
rect 17516 5712 17529 5716
rect 17581 5720 17660 5736
rect 17692 5736 17864 5738
rect 17692 5720 17771 5736
rect 17778 5734 17808 5736
rect 17356 5698 17385 5708
rect 17399 5698 17428 5708
rect 17443 5698 17473 5712
rect 17516 5698 17559 5712
rect 17581 5708 17771 5720
rect 17836 5716 17842 5736
rect 17566 5698 17596 5708
rect 17597 5698 17755 5708
rect 17759 5698 17789 5708
rect 17793 5698 17823 5712
rect 17851 5698 17864 5736
rect 17936 5750 17965 5766
rect 17979 5750 18008 5766
rect 18023 5756 18053 5772
rect 18081 5750 18087 5798
rect 18090 5792 18109 5798
rect 18124 5792 18154 5800
rect 18090 5784 18154 5792
rect 18090 5768 18170 5784
rect 18186 5777 18248 5808
rect 18264 5777 18326 5808
rect 18395 5806 18444 5831
rect 18459 5806 18489 5822
rect 18358 5792 18388 5800
rect 18395 5798 18505 5806
rect 18358 5784 18403 5792
rect 18090 5766 18109 5768
rect 18124 5766 18170 5768
rect 18090 5750 18170 5766
rect 18197 5764 18232 5777
rect 18273 5774 18310 5777
rect 18273 5772 18315 5774
rect 18202 5761 18232 5764
rect 18211 5757 18218 5761
rect 18218 5756 18219 5757
rect 18177 5750 18187 5756
rect 17936 5742 17971 5750
rect 17936 5716 17937 5742
rect 17944 5716 17971 5742
rect 17879 5698 17909 5712
rect 17936 5708 17971 5716
rect 17973 5742 18014 5750
rect 17973 5716 17988 5742
rect 17995 5716 18014 5742
rect 18078 5738 18109 5750
rect 18124 5738 18227 5750
rect 18239 5740 18265 5766
rect 18280 5761 18310 5772
rect 18342 5768 18404 5784
rect 18342 5766 18388 5768
rect 18342 5750 18404 5766
rect 18416 5750 18422 5798
rect 18425 5790 18505 5798
rect 18425 5788 18444 5790
rect 18459 5788 18493 5790
rect 18425 5772 18505 5788
rect 18425 5750 18444 5772
rect 18459 5756 18489 5772
rect 18517 5766 18523 5840
rect 18532 5766 18545 5910
rect 18285 5740 18388 5750
rect 18239 5738 18388 5740
rect 18409 5738 18444 5750
rect 18078 5736 18240 5738
rect 18090 5716 18109 5736
rect 18124 5734 18154 5736
rect 17973 5708 18014 5716
rect 18096 5712 18109 5716
rect 18161 5720 18240 5736
rect 18272 5736 18444 5738
rect 18272 5720 18351 5736
rect 18358 5734 18388 5736
rect 17936 5698 17965 5708
rect 17979 5698 18008 5708
rect 18023 5698 18053 5712
rect 18096 5698 18139 5712
rect 18161 5708 18351 5720
rect 18416 5716 18422 5736
rect 18146 5698 18176 5708
rect 18177 5698 18335 5708
rect 18339 5698 18369 5708
rect 18373 5698 18403 5712
rect 18431 5698 18444 5736
rect 18516 5750 18545 5766
rect 18516 5742 18551 5750
rect 18516 5716 18517 5742
rect 18524 5716 18551 5742
rect 18459 5698 18489 5712
rect 18516 5708 18551 5716
rect 18516 5698 18545 5708
rect -1 5692 18545 5698
rect 0 5684 18545 5692
rect 15 5654 28 5684
rect 43 5670 73 5684
rect 116 5670 159 5684
rect 166 5670 386 5684
rect 393 5670 423 5684
rect 83 5656 98 5668
rect 117 5656 130 5670
rect 198 5666 351 5670
rect 80 5654 102 5656
rect 180 5654 372 5666
rect 451 5654 464 5684
rect 479 5670 509 5684
rect 546 5654 565 5684
rect 580 5654 586 5684
rect 595 5654 608 5684
rect 623 5670 653 5684
rect 696 5670 739 5684
rect 746 5670 966 5684
rect 973 5670 1003 5684
rect 663 5656 678 5668
rect 697 5656 710 5670
rect 778 5666 931 5670
rect 660 5654 682 5656
rect 760 5654 952 5666
rect 1031 5654 1044 5684
rect 1059 5670 1089 5684
rect 1126 5654 1145 5684
rect 1160 5654 1166 5684
rect 1175 5654 1188 5684
rect 1203 5670 1233 5684
rect 1276 5670 1319 5684
rect 1326 5670 1546 5684
rect 1553 5670 1583 5684
rect 1243 5656 1258 5668
rect 1277 5656 1290 5670
rect 1358 5666 1511 5670
rect 1240 5654 1262 5656
rect 1340 5654 1532 5666
rect 1611 5654 1624 5684
rect 1639 5670 1669 5684
rect 1706 5654 1725 5684
rect 1740 5654 1746 5684
rect 1755 5654 1768 5684
rect 1783 5670 1813 5684
rect 1856 5670 1899 5684
rect 1906 5670 2126 5684
rect 2133 5670 2163 5684
rect 1823 5656 1838 5668
rect 1857 5656 1870 5670
rect 1938 5666 2091 5670
rect 1820 5654 1842 5656
rect 1920 5654 2112 5666
rect 2191 5654 2204 5684
rect 2219 5670 2249 5684
rect 2286 5654 2305 5684
rect 2320 5654 2326 5684
rect 2335 5654 2348 5684
rect 2363 5670 2393 5684
rect 2436 5670 2479 5684
rect 2486 5670 2706 5684
rect 2713 5670 2743 5684
rect 2403 5656 2418 5668
rect 2437 5656 2450 5670
rect 2518 5666 2671 5670
rect 2400 5654 2422 5656
rect 2500 5654 2692 5666
rect 2771 5654 2784 5684
rect 2799 5670 2829 5684
rect 2866 5654 2885 5684
rect 2900 5654 2906 5684
rect 2915 5654 2928 5684
rect 2943 5670 2973 5684
rect 3016 5670 3059 5684
rect 3066 5670 3286 5684
rect 3293 5670 3323 5684
rect 2983 5656 2998 5668
rect 3017 5656 3030 5670
rect 3098 5666 3251 5670
rect 2980 5654 3002 5656
rect 3080 5654 3272 5666
rect 3351 5654 3364 5684
rect 3379 5670 3409 5684
rect 3446 5654 3465 5684
rect 3480 5654 3486 5684
rect 3495 5654 3508 5684
rect 3523 5670 3553 5684
rect 3596 5670 3639 5684
rect 3646 5670 3866 5684
rect 3873 5670 3903 5684
rect 3563 5656 3578 5668
rect 3597 5656 3610 5670
rect 3678 5666 3831 5670
rect 3560 5654 3582 5656
rect 3660 5654 3852 5666
rect 3931 5654 3944 5684
rect 3959 5670 3989 5684
rect 4026 5654 4045 5684
rect 4060 5654 4066 5684
rect 4075 5654 4088 5684
rect 4103 5670 4133 5684
rect 4176 5670 4219 5684
rect 4226 5670 4446 5684
rect 4453 5670 4483 5684
rect 4143 5656 4158 5668
rect 4177 5656 4190 5670
rect 4258 5666 4411 5670
rect 4140 5654 4162 5656
rect 4240 5654 4432 5666
rect 4511 5654 4524 5684
rect 4539 5670 4569 5684
rect 4606 5654 4625 5684
rect 4640 5654 4646 5684
rect 4655 5654 4668 5684
rect 4683 5670 4713 5684
rect 4756 5670 4799 5684
rect 4806 5670 5026 5684
rect 5033 5670 5063 5684
rect 4723 5656 4738 5668
rect 4757 5656 4770 5670
rect 4838 5666 4991 5670
rect 4720 5654 4742 5656
rect 4820 5654 5012 5666
rect 5091 5654 5104 5684
rect 5119 5670 5149 5684
rect 5186 5654 5205 5684
rect 5220 5654 5226 5684
rect 5235 5654 5248 5684
rect 5263 5670 5293 5684
rect 5336 5670 5379 5684
rect 5386 5670 5606 5684
rect 5613 5670 5643 5684
rect 5303 5656 5318 5668
rect 5337 5656 5350 5670
rect 5418 5666 5571 5670
rect 5300 5654 5322 5656
rect 5400 5654 5592 5666
rect 5671 5654 5684 5684
rect 5699 5670 5729 5684
rect 5766 5654 5785 5684
rect 5800 5654 5806 5684
rect 5815 5654 5828 5684
rect 5843 5670 5873 5684
rect 5916 5670 5959 5684
rect 5966 5670 6186 5684
rect 6193 5670 6223 5684
rect 5883 5656 5898 5668
rect 5917 5656 5930 5670
rect 5998 5666 6151 5670
rect 5880 5654 5902 5656
rect 5980 5654 6172 5666
rect 6251 5654 6264 5684
rect 6279 5670 6309 5684
rect 6346 5654 6365 5684
rect 6380 5654 6386 5684
rect 6395 5654 6408 5684
rect 6423 5670 6453 5684
rect 6496 5670 6539 5684
rect 6546 5670 6766 5684
rect 6773 5670 6803 5684
rect 6463 5656 6478 5668
rect 6497 5656 6510 5670
rect 6578 5666 6731 5670
rect 6460 5654 6482 5656
rect 6560 5654 6752 5666
rect 6831 5654 6844 5684
rect 6859 5670 6889 5684
rect 6926 5654 6945 5684
rect 6960 5654 6966 5684
rect 6975 5654 6988 5684
rect 7003 5670 7033 5684
rect 7076 5670 7119 5684
rect 7126 5670 7346 5684
rect 7353 5670 7383 5684
rect 7043 5656 7058 5668
rect 7077 5656 7090 5670
rect 7158 5666 7311 5670
rect 7040 5654 7062 5656
rect 7140 5654 7332 5666
rect 7411 5654 7424 5684
rect 7439 5670 7469 5684
rect 7506 5654 7525 5684
rect 7540 5654 7546 5684
rect 7555 5654 7568 5684
rect 7583 5670 7613 5684
rect 7656 5670 7699 5684
rect 7706 5670 7926 5684
rect 7933 5670 7963 5684
rect 7623 5656 7638 5668
rect 7657 5656 7670 5670
rect 7738 5666 7891 5670
rect 7620 5654 7642 5656
rect 7720 5654 7912 5666
rect 7991 5654 8004 5684
rect 8019 5670 8049 5684
rect 8086 5654 8105 5684
rect 8120 5654 8126 5684
rect 8135 5654 8148 5684
rect 8163 5670 8193 5684
rect 8236 5670 8279 5684
rect 8286 5670 8506 5684
rect 8513 5670 8543 5684
rect 8203 5656 8218 5668
rect 8237 5656 8250 5670
rect 8318 5666 8471 5670
rect 8200 5654 8222 5656
rect 8300 5654 8492 5666
rect 8571 5654 8584 5684
rect 8599 5670 8629 5684
rect 8666 5654 8685 5684
rect 8700 5654 8706 5684
rect 8715 5654 8728 5684
rect 8743 5670 8773 5684
rect 8816 5670 8859 5684
rect 8866 5670 9086 5684
rect 9093 5670 9123 5684
rect 8783 5656 8798 5668
rect 8817 5656 8830 5670
rect 8898 5666 9051 5670
rect 8780 5654 8802 5656
rect 8880 5654 9072 5666
rect 9151 5654 9164 5684
rect 9179 5670 9209 5684
rect 9246 5654 9265 5684
rect 9280 5654 9286 5684
rect 9295 5654 9308 5684
rect 9323 5670 9353 5684
rect 9396 5670 9439 5684
rect 9446 5670 9666 5684
rect 9673 5670 9703 5684
rect 9363 5656 9378 5668
rect 9397 5656 9410 5670
rect 9478 5666 9631 5670
rect 9360 5654 9382 5656
rect 9460 5654 9652 5666
rect 9731 5654 9744 5684
rect 9759 5670 9789 5684
rect 9826 5654 9845 5684
rect 9860 5654 9866 5684
rect 9875 5654 9888 5684
rect 9903 5670 9933 5684
rect 9976 5670 10019 5684
rect 10026 5670 10246 5684
rect 10253 5670 10283 5684
rect 9943 5656 9958 5668
rect 9977 5656 9990 5670
rect 10058 5666 10211 5670
rect 9940 5654 9962 5656
rect 10040 5654 10232 5666
rect 10311 5654 10324 5684
rect 10339 5670 10369 5684
rect 10406 5654 10425 5684
rect 10440 5654 10446 5684
rect 10455 5654 10468 5684
rect 10483 5670 10513 5684
rect 10556 5670 10599 5684
rect 10606 5670 10826 5684
rect 10833 5670 10863 5684
rect 10523 5656 10538 5668
rect 10557 5656 10570 5670
rect 10638 5666 10791 5670
rect 10520 5654 10542 5656
rect 10620 5654 10812 5666
rect 10891 5654 10904 5684
rect 10919 5670 10949 5684
rect 10986 5654 11005 5684
rect 11020 5654 11026 5684
rect 11035 5654 11048 5684
rect 11063 5670 11093 5684
rect 11136 5670 11179 5684
rect 11186 5670 11406 5684
rect 11413 5670 11443 5684
rect 11103 5656 11118 5668
rect 11137 5656 11150 5670
rect 11218 5666 11371 5670
rect 11100 5654 11122 5656
rect 11200 5654 11392 5666
rect 11471 5654 11484 5684
rect 11499 5670 11529 5684
rect 11566 5654 11585 5684
rect 11600 5654 11606 5684
rect 11615 5654 11628 5684
rect 11643 5670 11673 5684
rect 11716 5670 11759 5684
rect 11766 5670 11986 5684
rect 11993 5670 12023 5684
rect 11683 5656 11698 5668
rect 11717 5656 11730 5670
rect 11798 5666 11951 5670
rect 11680 5654 11702 5656
rect 11780 5654 11972 5666
rect 12051 5654 12064 5684
rect 12079 5670 12109 5684
rect 12146 5654 12165 5684
rect 12180 5654 12186 5684
rect 12195 5654 12208 5684
rect 12223 5670 12253 5684
rect 12296 5670 12339 5684
rect 12346 5670 12566 5684
rect 12573 5670 12603 5684
rect 12263 5656 12278 5668
rect 12297 5656 12310 5670
rect 12378 5666 12531 5670
rect 12260 5654 12282 5656
rect 12360 5654 12552 5666
rect 12631 5654 12644 5684
rect 12659 5670 12689 5684
rect 12726 5654 12745 5684
rect 12760 5654 12766 5684
rect 12775 5654 12788 5684
rect 12803 5670 12833 5684
rect 12876 5670 12919 5684
rect 12926 5670 13146 5684
rect 13153 5670 13183 5684
rect 12843 5656 12858 5668
rect 12877 5656 12890 5670
rect 12958 5666 13111 5670
rect 12840 5654 12862 5656
rect 12940 5654 13132 5666
rect 13211 5654 13224 5684
rect 13239 5670 13269 5684
rect 13306 5654 13325 5684
rect 13340 5654 13346 5684
rect 13355 5654 13368 5684
rect 13383 5670 13413 5684
rect 13456 5670 13499 5684
rect 13506 5670 13726 5684
rect 13733 5670 13763 5684
rect 13423 5656 13438 5668
rect 13457 5656 13470 5670
rect 13538 5666 13691 5670
rect 13420 5654 13442 5656
rect 13520 5654 13712 5666
rect 13791 5654 13804 5684
rect 13819 5670 13849 5684
rect 13886 5654 13905 5684
rect 13920 5654 13926 5684
rect 13935 5654 13948 5684
rect 13963 5670 13993 5684
rect 14036 5670 14079 5684
rect 14086 5670 14306 5684
rect 14313 5670 14343 5684
rect 14003 5656 14018 5668
rect 14037 5656 14050 5670
rect 14118 5666 14271 5670
rect 14000 5654 14022 5656
rect 14100 5654 14292 5666
rect 14371 5654 14384 5684
rect 14399 5670 14429 5684
rect 14466 5654 14485 5684
rect 14500 5654 14506 5684
rect 14515 5654 14528 5684
rect 14543 5670 14573 5684
rect 14616 5670 14659 5684
rect 14666 5670 14886 5684
rect 14893 5670 14923 5684
rect 14583 5656 14598 5668
rect 14617 5656 14630 5670
rect 14698 5666 14851 5670
rect 14580 5654 14602 5656
rect 14680 5654 14872 5666
rect 14951 5654 14964 5684
rect 14979 5670 15009 5684
rect 15046 5654 15065 5684
rect 15080 5654 15086 5684
rect 15095 5654 15108 5684
rect 15123 5670 15153 5684
rect 15196 5670 15239 5684
rect 15246 5670 15466 5684
rect 15473 5670 15503 5684
rect 15163 5656 15178 5668
rect 15197 5656 15210 5670
rect 15278 5666 15431 5670
rect 15160 5654 15182 5656
rect 15260 5654 15452 5666
rect 15531 5654 15544 5684
rect 15559 5670 15589 5684
rect 15626 5654 15645 5684
rect 15660 5654 15666 5684
rect 15675 5654 15688 5684
rect 15703 5670 15733 5684
rect 15776 5670 15819 5684
rect 15826 5670 16046 5684
rect 16053 5670 16083 5684
rect 15743 5656 15758 5668
rect 15777 5656 15790 5670
rect 15858 5666 16011 5670
rect 15740 5654 15762 5656
rect 15840 5654 16032 5666
rect 16111 5654 16124 5684
rect 16139 5670 16169 5684
rect 16206 5654 16225 5684
rect 16240 5654 16246 5684
rect 16255 5654 16268 5684
rect 16283 5670 16313 5684
rect 16356 5670 16399 5684
rect 16406 5670 16626 5684
rect 16633 5670 16663 5684
rect 16323 5656 16338 5668
rect 16357 5656 16370 5670
rect 16438 5666 16591 5670
rect 16320 5654 16342 5656
rect 16420 5654 16612 5666
rect 16691 5654 16704 5684
rect 16719 5670 16749 5684
rect 16786 5654 16805 5684
rect 16820 5654 16826 5684
rect 16835 5654 16848 5684
rect 16863 5670 16893 5684
rect 16936 5670 16979 5684
rect 16986 5670 17206 5684
rect 17213 5670 17243 5684
rect 16903 5656 16918 5668
rect 16937 5656 16950 5670
rect 17018 5666 17171 5670
rect 16900 5654 16922 5656
rect 17000 5654 17192 5666
rect 17271 5654 17284 5684
rect 17299 5670 17329 5684
rect 17366 5654 17385 5684
rect 17400 5654 17406 5684
rect 17415 5654 17428 5684
rect 17443 5670 17473 5684
rect 17516 5670 17559 5684
rect 17566 5670 17786 5684
rect 17793 5670 17823 5684
rect 17483 5656 17498 5668
rect 17517 5656 17530 5670
rect 17598 5666 17751 5670
rect 17480 5654 17502 5656
rect 17580 5654 17772 5666
rect 17851 5654 17864 5684
rect 17879 5670 17909 5684
rect 17946 5654 17965 5684
rect 17980 5654 17986 5684
rect 17995 5654 18008 5684
rect 18023 5670 18053 5684
rect 18096 5670 18139 5684
rect 18146 5670 18366 5684
rect 18373 5670 18403 5684
rect 18063 5656 18078 5668
rect 18097 5656 18110 5670
rect 18178 5666 18331 5670
rect 18060 5654 18082 5656
rect 18160 5654 18352 5666
rect 18431 5654 18444 5684
rect 18459 5670 18489 5684
rect 18532 5654 18545 5684
rect 0 5640 18545 5654
rect 15 5570 28 5640
rect 80 5636 102 5640
rect 73 5614 102 5628
rect 155 5614 171 5628
rect 209 5624 215 5626
rect 222 5624 330 5640
rect 337 5624 343 5626
rect 351 5624 366 5640
rect 432 5634 451 5637
rect 73 5612 171 5614
rect 198 5612 366 5624
rect 381 5614 397 5628
rect 432 5615 454 5634
rect 464 5628 480 5629
rect 463 5626 480 5628
rect 464 5621 480 5626
rect 454 5614 460 5615
rect 463 5614 492 5621
rect 381 5613 492 5614
rect 381 5612 498 5613
rect 57 5604 108 5612
rect 155 5604 189 5612
rect 57 5592 82 5604
rect 89 5592 108 5604
rect 162 5602 189 5604
rect 198 5602 419 5612
rect 454 5609 460 5612
rect 162 5598 419 5602
rect 57 5584 108 5592
rect 155 5584 419 5598
rect 463 5604 498 5612
rect 9 5536 28 5570
rect 73 5576 102 5584
rect 73 5570 90 5576
rect 73 5568 107 5570
rect 155 5568 171 5584
rect 172 5574 380 5584
rect 381 5574 397 5584
rect 445 5580 460 5595
rect 463 5592 464 5604
rect 471 5592 498 5604
rect 463 5584 498 5592
rect 463 5583 492 5584
rect 183 5570 397 5574
rect 198 5568 397 5570
rect 432 5570 445 5580
rect 463 5570 480 5583
rect 432 5568 480 5570
rect 74 5564 107 5568
rect 70 5562 107 5564
rect 70 5561 137 5562
rect 70 5556 101 5561
rect 107 5556 137 5561
rect 70 5552 137 5556
rect 43 5549 137 5552
rect 43 5542 92 5549
rect 43 5536 73 5542
rect 92 5537 97 5542
rect 9 5520 89 5536
rect 101 5528 137 5549
rect 198 5544 387 5568
rect 432 5567 479 5568
rect 445 5562 479 5567
rect 213 5541 387 5544
rect 206 5538 387 5541
rect 415 5561 479 5562
rect 9 5518 28 5520
rect 43 5518 77 5520
rect 9 5502 89 5518
rect 9 5496 28 5502
rect -1 5480 28 5496
rect 43 5486 73 5502
rect 101 5480 107 5528
rect 110 5522 129 5528
rect 144 5522 174 5530
rect 110 5514 174 5522
rect 110 5498 190 5514
rect 206 5507 268 5538
rect 284 5507 346 5538
rect 415 5536 464 5561
rect 479 5536 509 5552
rect 378 5522 408 5530
rect 415 5528 525 5536
rect 378 5514 423 5522
rect 110 5496 129 5498
rect 144 5496 190 5498
rect 110 5480 190 5496
rect 217 5494 252 5507
rect 293 5504 330 5507
rect 293 5502 335 5504
rect 222 5491 252 5494
rect 231 5487 238 5491
rect 238 5486 239 5487
rect 197 5480 207 5486
rect -7 5472 34 5480
rect -7 5446 8 5472
rect 15 5446 34 5472
rect 98 5468 129 5480
rect 144 5468 247 5480
rect 259 5470 285 5496
rect 300 5491 330 5502
rect 362 5498 424 5514
rect 362 5496 408 5498
rect 362 5480 424 5496
rect 436 5480 442 5528
rect 445 5520 525 5528
rect 445 5518 464 5520
rect 479 5518 513 5520
rect 445 5502 525 5518
rect 445 5480 464 5502
rect 479 5486 509 5502
rect 537 5496 543 5570
rect 546 5496 565 5640
rect 580 5496 586 5640
rect 595 5570 608 5640
rect 660 5636 682 5640
rect 653 5614 682 5628
rect 735 5614 751 5628
rect 789 5624 795 5626
rect 802 5624 910 5640
rect 917 5624 923 5626
rect 931 5624 946 5640
rect 1012 5634 1031 5637
rect 653 5612 751 5614
rect 778 5612 946 5624
rect 961 5614 977 5628
rect 1012 5615 1034 5634
rect 1044 5628 1060 5629
rect 1043 5626 1060 5628
rect 1044 5621 1060 5626
rect 1034 5614 1040 5615
rect 1043 5614 1072 5621
rect 961 5613 1072 5614
rect 961 5612 1078 5613
rect 637 5604 688 5612
rect 735 5604 769 5612
rect 637 5592 662 5604
rect 669 5592 688 5604
rect 742 5602 769 5604
rect 778 5602 999 5612
rect 1034 5609 1040 5612
rect 742 5598 999 5602
rect 637 5584 688 5592
rect 735 5584 999 5598
rect 1043 5604 1078 5612
rect 589 5536 608 5570
rect 653 5576 682 5584
rect 653 5570 670 5576
rect 653 5568 687 5570
rect 735 5568 751 5584
rect 752 5574 960 5584
rect 961 5574 977 5584
rect 1025 5580 1040 5595
rect 1043 5592 1044 5604
rect 1051 5592 1078 5604
rect 1043 5584 1078 5592
rect 1043 5583 1072 5584
rect 763 5570 977 5574
rect 778 5568 977 5570
rect 1012 5570 1025 5580
rect 1043 5570 1060 5583
rect 1012 5568 1060 5570
rect 654 5564 687 5568
rect 650 5562 687 5564
rect 650 5561 717 5562
rect 650 5556 681 5561
rect 687 5556 717 5561
rect 650 5552 717 5556
rect 623 5549 717 5552
rect 623 5542 672 5549
rect 623 5536 653 5542
rect 672 5537 677 5542
rect 589 5520 669 5536
rect 681 5528 717 5549
rect 778 5544 967 5568
rect 1012 5567 1059 5568
rect 1025 5562 1059 5567
rect 793 5541 967 5544
rect 786 5538 967 5541
rect 995 5561 1059 5562
rect 589 5518 608 5520
rect 623 5518 657 5520
rect 589 5502 669 5518
rect 589 5496 608 5502
rect 305 5470 408 5480
rect 259 5468 408 5470
rect 429 5468 464 5480
rect 98 5466 260 5468
rect 110 5446 129 5466
rect 144 5464 174 5466
rect -7 5438 34 5446
rect 116 5442 129 5446
rect 181 5450 260 5466
rect 292 5466 464 5468
rect 292 5450 371 5466
rect 378 5464 408 5466
rect -1 5428 28 5438
rect 43 5428 73 5442
rect 116 5428 159 5442
rect 181 5438 371 5450
rect 436 5446 442 5466
rect 166 5428 196 5438
rect 197 5428 355 5438
rect 359 5428 389 5438
rect 393 5428 423 5442
rect 451 5428 464 5466
rect 536 5480 565 5496
rect 579 5480 608 5496
rect 623 5486 653 5502
rect 681 5480 687 5528
rect 690 5522 709 5528
rect 724 5522 754 5530
rect 690 5514 754 5522
rect 690 5498 770 5514
rect 786 5507 848 5538
rect 864 5507 926 5538
rect 995 5536 1044 5561
rect 1059 5536 1089 5552
rect 958 5522 988 5530
rect 995 5528 1105 5536
rect 958 5514 1003 5522
rect 690 5496 709 5498
rect 724 5496 770 5498
rect 690 5480 770 5496
rect 797 5494 832 5507
rect 873 5504 910 5507
rect 873 5502 915 5504
rect 802 5491 832 5494
rect 811 5487 818 5491
rect 818 5486 819 5487
rect 777 5480 787 5486
rect 536 5472 571 5480
rect 536 5446 537 5472
rect 544 5446 571 5472
rect 479 5428 509 5442
rect 536 5438 571 5446
rect 573 5472 614 5480
rect 573 5446 588 5472
rect 595 5446 614 5472
rect 678 5468 709 5480
rect 724 5468 827 5480
rect 839 5470 865 5496
rect 880 5491 910 5502
rect 942 5498 1004 5514
rect 942 5496 988 5498
rect 942 5480 1004 5496
rect 1016 5480 1022 5528
rect 1025 5520 1105 5528
rect 1025 5518 1044 5520
rect 1059 5518 1093 5520
rect 1025 5502 1105 5518
rect 1025 5480 1044 5502
rect 1059 5486 1089 5502
rect 1117 5496 1123 5570
rect 1126 5496 1145 5640
rect 1160 5496 1166 5640
rect 1175 5570 1188 5640
rect 1240 5636 1262 5640
rect 1233 5614 1262 5628
rect 1315 5614 1331 5628
rect 1369 5624 1375 5626
rect 1382 5624 1490 5640
rect 1497 5624 1503 5626
rect 1511 5624 1526 5640
rect 1592 5634 1611 5637
rect 1233 5612 1331 5614
rect 1358 5612 1526 5624
rect 1541 5614 1557 5628
rect 1592 5615 1614 5634
rect 1624 5628 1640 5629
rect 1623 5626 1640 5628
rect 1624 5621 1640 5626
rect 1614 5614 1620 5615
rect 1623 5614 1652 5621
rect 1541 5613 1652 5614
rect 1541 5612 1658 5613
rect 1217 5604 1268 5612
rect 1315 5604 1349 5612
rect 1217 5592 1242 5604
rect 1249 5592 1268 5604
rect 1322 5602 1349 5604
rect 1358 5602 1579 5612
rect 1614 5609 1620 5612
rect 1322 5598 1579 5602
rect 1217 5584 1268 5592
rect 1315 5584 1579 5598
rect 1623 5604 1658 5612
rect 1169 5536 1188 5570
rect 1233 5576 1262 5584
rect 1233 5570 1250 5576
rect 1233 5568 1267 5570
rect 1315 5568 1331 5584
rect 1332 5574 1540 5584
rect 1541 5574 1557 5584
rect 1605 5580 1620 5595
rect 1623 5592 1624 5604
rect 1631 5592 1658 5604
rect 1623 5584 1658 5592
rect 1623 5583 1652 5584
rect 1343 5570 1557 5574
rect 1358 5568 1557 5570
rect 1592 5570 1605 5580
rect 1623 5570 1640 5583
rect 1592 5568 1640 5570
rect 1234 5564 1267 5568
rect 1230 5562 1267 5564
rect 1230 5561 1297 5562
rect 1230 5556 1261 5561
rect 1267 5556 1297 5561
rect 1230 5552 1297 5556
rect 1203 5549 1297 5552
rect 1203 5542 1252 5549
rect 1203 5536 1233 5542
rect 1252 5537 1257 5542
rect 1169 5520 1249 5536
rect 1261 5528 1297 5549
rect 1358 5544 1547 5568
rect 1592 5567 1639 5568
rect 1605 5562 1639 5567
rect 1373 5541 1547 5544
rect 1366 5538 1547 5541
rect 1575 5561 1639 5562
rect 1169 5518 1188 5520
rect 1203 5518 1237 5520
rect 1169 5502 1249 5518
rect 1169 5496 1188 5502
rect 885 5470 988 5480
rect 839 5468 988 5470
rect 1009 5468 1044 5480
rect 678 5466 840 5468
rect 690 5446 709 5466
rect 724 5464 754 5466
rect 573 5438 614 5446
rect 696 5442 709 5446
rect 761 5450 840 5466
rect 872 5466 1044 5468
rect 872 5450 951 5466
rect 958 5464 988 5466
rect 536 5428 565 5438
rect 579 5428 608 5438
rect 623 5428 653 5442
rect 696 5428 739 5442
rect 761 5438 951 5450
rect 1016 5446 1022 5466
rect 746 5428 776 5438
rect 777 5428 935 5438
rect 939 5428 969 5438
rect 973 5428 1003 5442
rect 1031 5428 1044 5466
rect 1116 5480 1145 5496
rect 1159 5480 1188 5496
rect 1203 5486 1233 5502
rect 1261 5480 1267 5528
rect 1270 5522 1289 5528
rect 1304 5522 1334 5530
rect 1270 5514 1334 5522
rect 1270 5498 1350 5514
rect 1366 5507 1428 5538
rect 1444 5507 1506 5538
rect 1575 5536 1624 5561
rect 1639 5536 1669 5552
rect 1538 5522 1568 5530
rect 1575 5528 1685 5536
rect 1538 5514 1583 5522
rect 1270 5496 1289 5498
rect 1304 5496 1350 5498
rect 1270 5480 1350 5496
rect 1377 5494 1412 5507
rect 1453 5504 1490 5507
rect 1453 5502 1495 5504
rect 1382 5491 1412 5494
rect 1391 5487 1398 5491
rect 1398 5486 1399 5487
rect 1357 5480 1367 5486
rect 1116 5472 1151 5480
rect 1116 5446 1117 5472
rect 1124 5446 1151 5472
rect 1059 5428 1089 5442
rect 1116 5438 1151 5446
rect 1153 5472 1194 5480
rect 1153 5446 1168 5472
rect 1175 5446 1194 5472
rect 1258 5468 1289 5480
rect 1304 5468 1407 5480
rect 1419 5470 1445 5496
rect 1460 5491 1490 5502
rect 1522 5498 1584 5514
rect 1522 5496 1568 5498
rect 1522 5480 1584 5496
rect 1596 5480 1602 5528
rect 1605 5520 1685 5528
rect 1605 5518 1624 5520
rect 1639 5518 1673 5520
rect 1605 5502 1685 5518
rect 1605 5480 1624 5502
rect 1639 5486 1669 5502
rect 1697 5496 1703 5570
rect 1706 5496 1725 5640
rect 1740 5496 1746 5640
rect 1755 5570 1768 5640
rect 1820 5636 1842 5640
rect 1813 5614 1842 5628
rect 1895 5614 1911 5628
rect 1949 5624 1955 5626
rect 1962 5624 2070 5640
rect 2077 5624 2083 5626
rect 2091 5624 2106 5640
rect 2172 5634 2191 5637
rect 1813 5612 1911 5614
rect 1938 5612 2106 5624
rect 2121 5614 2137 5628
rect 2172 5615 2194 5634
rect 2204 5628 2220 5629
rect 2203 5626 2220 5628
rect 2204 5621 2220 5626
rect 2194 5614 2200 5615
rect 2203 5614 2232 5621
rect 2121 5613 2232 5614
rect 2121 5612 2238 5613
rect 1797 5604 1848 5612
rect 1895 5604 1929 5612
rect 1797 5592 1822 5604
rect 1829 5592 1848 5604
rect 1902 5602 1929 5604
rect 1938 5602 2159 5612
rect 2194 5609 2200 5612
rect 1902 5598 2159 5602
rect 1797 5584 1848 5592
rect 1895 5584 2159 5598
rect 2203 5604 2238 5612
rect 1749 5536 1768 5570
rect 1813 5576 1842 5584
rect 1813 5570 1830 5576
rect 1813 5568 1847 5570
rect 1895 5568 1911 5584
rect 1912 5574 2120 5584
rect 2121 5574 2137 5584
rect 2185 5580 2200 5595
rect 2203 5592 2204 5604
rect 2211 5592 2238 5604
rect 2203 5584 2238 5592
rect 2203 5583 2232 5584
rect 1923 5570 2137 5574
rect 1938 5568 2137 5570
rect 2172 5570 2185 5580
rect 2203 5570 2220 5583
rect 2172 5568 2220 5570
rect 1814 5564 1847 5568
rect 1810 5562 1847 5564
rect 1810 5561 1877 5562
rect 1810 5556 1841 5561
rect 1847 5556 1877 5561
rect 1810 5552 1877 5556
rect 1783 5549 1877 5552
rect 1783 5542 1832 5549
rect 1783 5536 1813 5542
rect 1832 5537 1837 5542
rect 1749 5520 1829 5536
rect 1841 5528 1877 5549
rect 1938 5544 2127 5568
rect 2172 5567 2219 5568
rect 2185 5562 2219 5567
rect 1953 5541 2127 5544
rect 1946 5538 2127 5541
rect 2155 5561 2219 5562
rect 1749 5518 1768 5520
rect 1783 5518 1817 5520
rect 1749 5502 1829 5518
rect 1749 5496 1768 5502
rect 1465 5470 1568 5480
rect 1419 5468 1568 5470
rect 1589 5468 1624 5480
rect 1258 5466 1420 5468
rect 1270 5446 1289 5466
rect 1304 5464 1334 5466
rect 1153 5438 1194 5446
rect 1276 5442 1289 5446
rect 1341 5450 1420 5466
rect 1452 5466 1624 5468
rect 1452 5450 1531 5466
rect 1538 5464 1568 5466
rect 1116 5428 1145 5438
rect 1159 5428 1188 5438
rect 1203 5428 1233 5442
rect 1276 5428 1319 5442
rect 1341 5438 1531 5450
rect 1596 5446 1602 5466
rect 1326 5428 1356 5438
rect 1357 5428 1515 5438
rect 1519 5428 1549 5438
rect 1553 5428 1583 5442
rect 1611 5428 1624 5466
rect 1696 5480 1725 5496
rect 1739 5480 1768 5496
rect 1783 5486 1813 5502
rect 1841 5480 1847 5528
rect 1850 5522 1869 5528
rect 1884 5522 1914 5530
rect 1850 5514 1914 5522
rect 1850 5498 1930 5514
rect 1946 5507 2008 5538
rect 2024 5507 2086 5538
rect 2155 5536 2204 5561
rect 2219 5536 2249 5552
rect 2118 5522 2148 5530
rect 2155 5528 2265 5536
rect 2118 5514 2163 5522
rect 1850 5496 1869 5498
rect 1884 5496 1930 5498
rect 1850 5480 1930 5496
rect 1957 5494 1992 5507
rect 2033 5504 2070 5507
rect 2033 5502 2075 5504
rect 1962 5491 1992 5494
rect 1971 5487 1978 5491
rect 1978 5486 1979 5487
rect 1937 5480 1947 5486
rect 1696 5472 1731 5480
rect 1696 5446 1697 5472
rect 1704 5446 1731 5472
rect 1639 5428 1669 5442
rect 1696 5438 1731 5446
rect 1733 5472 1774 5480
rect 1733 5446 1748 5472
rect 1755 5446 1774 5472
rect 1838 5468 1869 5480
rect 1884 5468 1987 5480
rect 1999 5470 2025 5496
rect 2040 5491 2070 5502
rect 2102 5498 2164 5514
rect 2102 5496 2148 5498
rect 2102 5480 2164 5496
rect 2176 5480 2182 5528
rect 2185 5520 2265 5528
rect 2185 5518 2204 5520
rect 2219 5518 2253 5520
rect 2185 5502 2265 5518
rect 2185 5480 2204 5502
rect 2219 5486 2249 5502
rect 2277 5496 2283 5570
rect 2286 5496 2305 5640
rect 2320 5496 2326 5640
rect 2335 5570 2348 5640
rect 2400 5636 2422 5640
rect 2393 5614 2422 5628
rect 2475 5614 2491 5628
rect 2529 5624 2535 5626
rect 2542 5624 2650 5640
rect 2657 5624 2663 5626
rect 2671 5624 2686 5640
rect 2752 5634 2771 5637
rect 2393 5612 2491 5614
rect 2518 5612 2686 5624
rect 2701 5614 2717 5628
rect 2752 5615 2774 5634
rect 2784 5628 2800 5629
rect 2783 5626 2800 5628
rect 2784 5621 2800 5626
rect 2774 5614 2780 5615
rect 2783 5614 2812 5621
rect 2701 5613 2812 5614
rect 2701 5612 2818 5613
rect 2377 5604 2428 5612
rect 2475 5604 2509 5612
rect 2377 5592 2402 5604
rect 2409 5592 2428 5604
rect 2482 5602 2509 5604
rect 2518 5602 2739 5612
rect 2774 5609 2780 5612
rect 2482 5598 2739 5602
rect 2377 5584 2428 5592
rect 2475 5584 2739 5598
rect 2783 5604 2818 5612
rect 2329 5536 2348 5570
rect 2393 5576 2422 5584
rect 2393 5570 2410 5576
rect 2393 5568 2427 5570
rect 2475 5568 2491 5584
rect 2492 5574 2700 5584
rect 2701 5574 2717 5584
rect 2765 5580 2780 5595
rect 2783 5592 2784 5604
rect 2791 5592 2818 5604
rect 2783 5584 2818 5592
rect 2783 5583 2812 5584
rect 2503 5570 2717 5574
rect 2518 5568 2717 5570
rect 2752 5570 2765 5580
rect 2783 5570 2800 5583
rect 2752 5568 2800 5570
rect 2394 5564 2427 5568
rect 2390 5562 2427 5564
rect 2390 5561 2457 5562
rect 2390 5556 2421 5561
rect 2427 5556 2457 5561
rect 2390 5552 2457 5556
rect 2363 5549 2457 5552
rect 2363 5542 2412 5549
rect 2363 5536 2393 5542
rect 2412 5537 2417 5542
rect 2329 5520 2409 5536
rect 2421 5528 2457 5549
rect 2518 5544 2707 5568
rect 2752 5567 2799 5568
rect 2765 5562 2799 5567
rect 2533 5541 2707 5544
rect 2526 5538 2707 5541
rect 2735 5561 2799 5562
rect 2329 5518 2348 5520
rect 2363 5518 2397 5520
rect 2329 5502 2409 5518
rect 2329 5496 2348 5502
rect 2045 5470 2148 5480
rect 1999 5468 2148 5470
rect 2169 5468 2204 5480
rect 1838 5466 2000 5468
rect 1850 5446 1869 5466
rect 1884 5464 1914 5466
rect 1733 5438 1774 5446
rect 1856 5442 1869 5446
rect 1921 5450 2000 5466
rect 2032 5466 2204 5468
rect 2032 5450 2111 5466
rect 2118 5464 2148 5466
rect 1696 5428 1725 5438
rect 1739 5428 1768 5438
rect 1783 5428 1813 5442
rect 1856 5428 1899 5442
rect 1921 5438 2111 5450
rect 2176 5446 2182 5466
rect 1906 5428 1936 5438
rect 1937 5428 2095 5438
rect 2099 5428 2129 5438
rect 2133 5428 2163 5442
rect 2191 5428 2204 5466
rect 2276 5480 2305 5496
rect 2319 5480 2348 5496
rect 2363 5486 2393 5502
rect 2421 5480 2427 5528
rect 2430 5522 2449 5528
rect 2464 5522 2494 5530
rect 2430 5514 2494 5522
rect 2430 5498 2510 5514
rect 2526 5507 2588 5538
rect 2604 5507 2666 5538
rect 2735 5536 2784 5561
rect 2799 5536 2829 5552
rect 2698 5522 2728 5530
rect 2735 5528 2845 5536
rect 2698 5514 2743 5522
rect 2430 5496 2449 5498
rect 2464 5496 2510 5498
rect 2430 5480 2510 5496
rect 2537 5494 2572 5507
rect 2613 5504 2650 5507
rect 2613 5502 2655 5504
rect 2542 5491 2572 5494
rect 2551 5487 2558 5491
rect 2558 5486 2559 5487
rect 2517 5480 2527 5486
rect 2276 5472 2311 5480
rect 2276 5446 2277 5472
rect 2284 5446 2311 5472
rect 2219 5428 2249 5442
rect 2276 5438 2311 5446
rect 2313 5472 2354 5480
rect 2313 5446 2328 5472
rect 2335 5446 2354 5472
rect 2418 5468 2449 5480
rect 2464 5468 2567 5480
rect 2579 5470 2605 5496
rect 2620 5491 2650 5502
rect 2682 5498 2744 5514
rect 2682 5496 2728 5498
rect 2682 5480 2744 5496
rect 2756 5480 2762 5528
rect 2765 5520 2845 5528
rect 2765 5518 2784 5520
rect 2799 5518 2833 5520
rect 2765 5502 2845 5518
rect 2765 5480 2784 5502
rect 2799 5486 2829 5502
rect 2857 5496 2863 5570
rect 2866 5496 2885 5640
rect 2900 5496 2906 5640
rect 2915 5570 2928 5640
rect 2980 5636 3002 5640
rect 2973 5614 3002 5628
rect 3055 5614 3071 5628
rect 3109 5624 3115 5626
rect 3122 5624 3230 5640
rect 3237 5624 3243 5626
rect 3251 5624 3266 5640
rect 3332 5634 3351 5637
rect 2973 5612 3071 5614
rect 3098 5612 3266 5624
rect 3281 5614 3297 5628
rect 3332 5615 3354 5634
rect 3364 5628 3380 5629
rect 3363 5626 3380 5628
rect 3364 5621 3380 5626
rect 3354 5614 3360 5615
rect 3363 5614 3392 5621
rect 3281 5613 3392 5614
rect 3281 5612 3398 5613
rect 2957 5604 3008 5612
rect 3055 5604 3089 5612
rect 2957 5592 2982 5604
rect 2989 5592 3008 5604
rect 3062 5602 3089 5604
rect 3098 5602 3319 5612
rect 3354 5609 3360 5612
rect 3062 5598 3319 5602
rect 2957 5584 3008 5592
rect 3055 5584 3319 5598
rect 3363 5604 3398 5612
rect 2909 5536 2928 5570
rect 2973 5576 3002 5584
rect 2973 5570 2990 5576
rect 2973 5568 3007 5570
rect 3055 5568 3071 5584
rect 3072 5574 3280 5584
rect 3281 5574 3297 5584
rect 3345 5580 3360 5595
rect 3363 5592 3364 5604
rect 3371 5592 3398 5604
rect 3363 5584 3398 5592
rect 3363 5583 3392 5584
rect 3083 5570 3297 5574
rect 3098 5568 3297 5570
rect 3332 5570 3345 5580
rect 3363 5570 3380 5583
rect 3332 5568 3380 5570
rect 2974 5564 3007 5568
rect 2970 5562 3007 5564
rect 2970 5561 3037 5562
rect 2970 5556 3001 5561
rect 3007 5556 3037 5561
rect 2970 5552 3037 5556
rect 2943 5549 3037 5552
rect 2943 5542 2992 5549
rect 2943 5536 2973 5542
rect 2992 5537 2997 5542
rect 2909 5520 2989 5536
rect 3001 5528 3037 5549
rect 3098 5544 3287 5568
rect 3332 5567 3379 5568
rect 3345 5562 3379 5567
rect 3113 5541 3287 5544
rect 3106 5538 3287 5541
rect 3315 5561 3379 5562
rect 2909 5518 2928 5520
rect 2943 5518 2977 5520
rect 2909 5502 2989 5518
rect 2909 5496 2928 5502
rect 2625 5470 2728 5480
rect 2579 5468 2728 5470
rect 2749 5468 2784 5480
rect 2418 5466 2580 5468
rect 2430 5446 2449 5466
rect 2464 5464 2494 5466
rect 2313 5438 2354 5446
rect 2436 5442 2449 5446
rect 2501 5450 2580 5466
rect 2612 5466 2784 5468
rect 2612 5450 2691 5466
rect 2698 5464 2728 5466
rect 2276 5428 2305 5438
rect 2319 5428 2348 5438
rect 2363 5428 2393 5442
rect 2436 5428 2479 5442
rect 2501 5438 2691 5450
rect 2756 5446 2762 5466
rect 2486 5428 2516 5438
rect 2517 5428 2675 5438
rect 2679 5428 2709 5438
rect 2713 5428 2743 5442
rect 2771 5428 2784 5466
rect 2856 5480 2885 5496
rect 2899 5480 2928 5496
rect 2943 5486 2973 5502
rect 3001 5480 3007 5528
rect 3010 5522 3029 5528
rect 3044 5522 3074 5530
rect 3010 5514 3074 5522
rect 3010 5498 3090 5514
rect 3106 5507 3168 5538
rect 3184 5507 3246 5538
rect 3315 5536 3364 5561
rect 3379 5536 3409 5552
rect 3278 5522 3308 5530
rect 3315 5528 3425 5536
rect 3278 5514 3323 5522
rect 3010 5496 3029 5498
rect 3044 5496 3090 5498
rect 3010 5480 3090 5496
rect 3117 5494 3152 5507
rect 3193 5504 3230 5507
rect 3193 5502 3235 5504
rect 3122 5491 3152 5494
rect 3131 5487 3138 5491
rect 3138 5486 3139 5487
rect 3097 5480 3107 5486
rect 2856 5472 2891 5480
rect 2856 5446 2857 5472
rect 2864 5446 2891 5472
rect 2799 5428 2829 5442
rect 2856 5438 2891 5446
rect 2893 5472 2934 5480
rect 2893 5446 2908 5472
rect 2915 5446 2934 5472
rect 2998 5468 3029 5480
rect 3044 5468 3147 5480
rect 3159 5470 3185 5496
rect 3200 5491 3230 5502
rect 3262 5498 3324 5514
rect 3262 5496 3308 5498
rect 3262 5480 3324 5496
rect 3336 5480 3342 5528
rect 3345 5520 3425 5528
rect 3345 5518 3364 5520
rect 3379 5518 3413 5520
rect 3345 5502 3425 5518
rect 3345 5480 3364 5502
rect 3379 5486 3409 5502
rect 3437 5496 3443 5570
rect 3446 5496 3465 5640
rect 3480 5496 3486 5640
rect 3495 5570 3508 5640
rect 3560 5636 3582 5640
rect 3553 5614 3582 5628
rect 3635 5614 3651 5628
rect 3689 5624 3695 5626
rect 3702 5624 3810 5640
rect 3817 5624 3823 5626
rect 3831 5624 3846 5640
rect 3912 5634 3931 5637
rect 3553 5612 3651 5614
rect 3678 5612 3846 5624
rect 3861 5614 3877 5628
rect 3912 5615 3934 5634
rect 3944 5628 3960 5629
rect 3943 5626 3960 5628
rect 3944 5621 3960 5626
rect 3934 5614 3940 5615
rect 3943 5614 3972 5621
rect 3861 5613 3972 5614
rect 3861 5612 3978 5613
rect 3537 5604 3588 5612
rect 3635 5604 3669 5612
rect 3537 5592 3562 5604
rect 3569 5592 3588 5604
rect 3642 5602 3669 5604
rect 3678 5602 3899 5612
rect 3934 5609 3940 5612
rect 3642 5598 3899 5602
rect 3537 5584 3588 5592
rect 3635 5584 3899 5598
rect 3943 5604 3978 5612
rect 3489 5536 3508 5570
rect 3553 5576 3582 5584
rect 3553 5570 3570 5576
rect 3553 5568 3587 5570
rect 3635 5568 3651 5584
rect 3652 5574 3860 5584
rect 3861 5574 3877 5584
rect 3925 5580 3940 5595
rect 3943 5592 3944 5604
rect 3951 5592 3978 5604
rect 3943 5584 3978 5592
rect 3943 5583 3972 5584
rect 3663 5570 3877 5574
rect 3678 5568 3877 5570
rect 3912 5570 3925 5580
rect 3943 5570 3960 5583
rect 3912 5568 3960 5570
rect 3554 5564 3587 5568
rect 3550 5562 3587 5564
rect 3550 5561 3617 5562
rect 3550 5556 3581 5561
rect 3587 5556 3617 5561
rect 3550 5552 3617 5556
rect 3523 5549 3617 5552
rect 3523 5542 3572 5549
rect 3523 5536 3553 5542
rect 3572 5537 3577 5542
rect 3489 5520 3569 5536
rect 3581 5528 3617 5549
rect 3678 5544 3867 5568
rect 3912 5567 3959 5568
rect 3925 5562 3959 5567
rect 3693 5541 3867 5544
rect 3686 5538 3867 5541
rect 3895 5561 3959 5562
rect 3489 5518 3508 5520
rect 3523 5518 3557 5520
rect 3489 5502 3569 5518
rect 3489 5496 3508 5502
rect 3205 5470 3308 5480
rect 3159 5468 3308 5470
rect 3329 5468 3364 5480
rect 2998 5466 3160 5468
rect 3010 5446 3029 5466
rect 3044 5464 3074 5466
rect 2893 5438 2934 5446
rect 3016 5442 3029 5446
rect 3081 5450 3160 5466
rect 3192 5466 3364 5468
rect 3192 5450 3271 5466
rect 3278 5464 3308 5466
rect 2856 5428 2885 5438
rect 2899 5428 2928 5438
rect 2943 5428 2973 5442
rect 3016 5428 3059 5442
rect 3081 5438 3271 5450
rect 3336 5446 3342 5466
rect 3066 5428 3096 5438
rect 3097 5428 3255 5438
rect 3259 5428 3289 5438
rect 3293 5428 3323 5442
rect 3351 5428 3364 5466
rect 3436 5480 3465 5496
rect 3479 5480 3508 5496
rect 3523 5486 3553 5502
rect 3581 5480 3587 5528
rect 3590 5522 3609 5528
rect 3624 5522 3654 5530
rect 3590 5514 3654 5522
rect 3590 5498 3670 5514
rect 3686 5507 3748 5538
rect 3764 5507 3826 5538
rect 3895 5536 3944 5561
rect 3959 5536 3989 5552
rect 3858 5522 3888 5530
rect 3895 5528 4005 5536
rect 3858 5514 3903 5522
rect 3590 5496 3609 5498
rect 3624 5496 3670 5498
rect 3590 5480 3670 5496
rect 3697 5494 3732 5507
rect 3773 5504 3810 5507
rect 3773 5502 3815 5504
rect 3702 5491 3732 5494
rect 3711 5487 3718 5491
rect 3718 5486 3719 5487
rect 3677 5480 3687 5486
rect 3436 5472 3471 5480
rect 3436 5446 3437 5472
rect 3444 5446 3471 5472
rect 3379 5428 3409 5442
rect 3436 5438 3471 5446
rect 3473 5472 3514 5480
rect 3473 5446 3488 5472
rect 3495 5446 3514 5472
rect 3578 5468 3609 5480
rect 3624 5468 3727 5480
rect 3739 5470 3765 5496
rect 3780 5491 3810 5502
rect 3842 5498 3904 5514
rect 3842 5496 3888 5498
rect 3842 5480 3904 5496
rect 3916 5480 3922 5528
rect 3925 5520 4005 5528
rect 3925 5518 3944 5520
rect 3959 5518 3993 5520
rect 3925 5502 4005 5518
rect 3925 5480 3944 5502
rect 3959 5486 3989 5502
rect 4017 5496 4023 5570
rect 4026 5496 4045 5640
rect 4060 5496 4066 5640
rect 4075 5570 4088 5640
rect 4140 5636 4162 5640
rect 4133 5614 4162 5628
rect 4215 5614 4231 5628
rect 4269 5624 4275 5626
rect 4282 5624 4390 5640
rect 4397 5624 4403 5626
rect 4411 5624 4426 5640
rect 4492 5634 4511 5637
rect 4133 5612 4231 5614
rect 4258 5612 4426 5624
rect 4441 5614 4457 5628
rect 4492 5615 4514 5634
rect 4524 5628 4540 5629
rect 4523 5626 4540 5628
rect 4524 5621 4540 5626
rect 4514 5614 4520 5615
rect 4523 5614 4552 5621
rect 4441 5613 4552 5614
rect 4441 5612 4558 5613
rect 4117 5604 4168 5612
rect 4215 5604 4249 5612
rect 4117 5592 4142 5604
rect 4149 5592 4168 5604
rect 4222 5602 4249 5604
rect 4258 5602 4479 5612
rect 4514 5609 4520 5612
rect 4222 5598 4479 5602
rect 4117 5584 4168 5592
rect 4215 5584 4479 5598
rect 4523 5604 4558 5612
rect 4069 5536 4088 5570
rect 4133 5576 4162 5584
rect 4133 5570 4150 5576
rect 4133 5568 4167 5570
rect 4215 5568 4231 5584
rect 4232 5574 4440 5584
rect 4441 5574 4457 5584
rect 4505 5580 4520 5595
rect 4523 5592 4524 5604
rect 4531 5592 4558 5604
rect 4523 5584 4558 5592
rect 4523 5583 4552 5584
rect 4243 5570 4457 5574
rect 4258 5568 4457 5570
rect 4492 5570 4505 5580
rect 4523 5570 4540 5583
rect 4492 5568 4540 5570
rect 4134 5564 4167 5568
rect 4130 5562 4167 5564
rect 4130 5561 4197 5562
rect 4130 5556 4161 5561
rect 4167 5556 4197 5561
rect 4130 5552 4197 5556
rect 4103 5549 4197 5552
rect 4103 5542 4152 5549
rect 4103 5536 4133 5542
rect 4152 5537 4157 5542
rect 4069 5520 4149 5536
rect 4161 5528 4197 5549
rect 4258 5544 4447 5568
rect 4492 5567 4539 5568
rect 4505 5562 4539 5567
rect 4273 5541 4447 5544
rect 4266 5538 4447 5541
rect 4475 5561 4539 5562
rect 4069 5518 4088 5520
rect 4103 5518 4137 5520
rect 4069 5502 4149 5518
rect 4069 5496 4088 5502
rect 3785 5470 3888 5480
rect 3739 5468 3888 5470
rect 3909 5468 3944 5480
rect 3578 5466 3740 5468
rect 3590 5446 3609 5466
rect 3624 5464 3654 5466
rect 3473 5438 3514 5446
rect 3596 5442 3609 5446
rect 3661 5450 3740 5466
rect 3772 5466 3944 5468
rect 3772 5450 3851 5466
rect 3858 5464 3888 5466
rect 3436 5428 3465 5438
rect 3479 5428 3508 5438
rect 3523 5428 3553 5442
rect 3596 5428 3639 5442
rect 3661 5438 3851 5450
rect 3916 5446 3922 5466
rect 3646 5428 3676 5438
rect 3677 5428 3835 5438
rect 3839 5428 3869 5438
rect 3873 5428 3903 5442
rect 3931 5428 3944 5466
rect 4016 5480 4045 5496
rect 4059 5480 4088 5496
rect 4103 5486 4133 5502
rect 4161 5480 4167 5528
rect 4170 5522 4189 5528
rect 4204 5522 4234 5530
rect 4170 5514 4234 5522
rect 4170 5498 4250 5514
rect 4266 5507 4328 5538
rect 4344 5507 4406 5538
rect 4475 5536 4524 5561
rect 4539 5536 4569 5552
rect 4438 5522 4468 5530
rect 4475 5528 4585 5536
rect 4438 5514 4483 5522
rect 4170 5496 4189 5498
rect 4204 5496 4250 5498
rect 4170 5480 4250 5496
rect 4277 5494 4312 5507
rect 4353 5504 4390 5507
rect 4353 5502 4395 5504
rect 4282 5491 4312 5494
rect 4291 5487 4298 5491
rect 4298 5486 4299 5487
rect 4257 5480 4267 5486
rect 4016 5472 4051 5480
rect 4016 5446 4017 5472
rect 4024 5446 4051 5472
rect 3959 5428 3989 5442
rect 4016 5438 4051 5446
rect 4053 5472 4094 5480
rect 4053 5446 4068 5472
rect 4075 5446 4094 5472
rect 4158 5468 4189 5480
rect 4204 5468 4307 5480
rect 4319 5470 4345 5496
rect 4360 5491 4390 5502
rect 4422 5498 4484 5514
rect 4422 5496 4468 5498
rect 4422 5480 4484 5496
rect 4496 5480 4502 5528
rect 4505 5520 4585 5528
rect 4505 5518 4524 5520
rect 4539 5518 4573 5520
rect 4505 5502 4585 5518
rect 4505 5480 4524 5502
rect 4539 5486 4569 5502
rect 4597 5496 4603 5570
rect 4606 5496 4625 5640
rect 4640 5496 4646 5640
rect 4655 5570 4668 5640
rect 4720 5636 4742 5640
rect 4713 5614 4742 5628
rect 4795 5614 4811 5628
rect 4849 5624 4855 5626
rect 4862 5624 4970 5640
rect 4977 5624 4983 5626
rect 4991 5624 5006 5640
rect 5072 5634 5091 5637
rect 4713 5612 4811 5614
rect 4838 5612 5006 5624
rect 5021 5614 5037 5628
rect 5072 5615 5094 5634
rect 5104 5628 5120 5629
rect 5103 5626 5120 5628
rect 5104 5621 5120 5626
rect 5094 5614 5100 5615
rect 5103 5614 5132 5621
rect 5021 5613 5132 5614
rect 5021 5612 5138 5613
rect 4697 5604 4748 5612
rect 4795 5604 4829 5612
rect 4697 5592 4722 5604
rect 4729 5592 4748 5604
rect 4802 5602 4829 5604
rect 4838 5602 5059 5612
rect 5094 5609 5100 5612
rect 4802 5598 5059 5602
rect 4697 5584 4748 5592
rect 4795 5584 5059 5598
rect 5103 5604 5138 5612
rect 4649 5536 4668 5570
rect 4713 5576 4742 5584
rect 4713 5570 4730 5576
rect 4713 5568 4747 5570
rect 4795 5568 4811 5584
rect 4812 5574 5020 5584
rect 5021 5574 5037 5584
rect 5085 5580 5100 5595
rect 5103 5592 5104 5604
rect 5111 5592 5138 5604
rect 5103 5584 5138 5592
rect 5103 5583 5132 5584
rect 4823 5570 5037 5574
rect 4838 5568 5037 5570
rect 5072 5570 5085 5580
rect 5103 5570 5120 5583
rect 5072 5568 5120 5570
rect 4714 5564 4747 5568
rect 4710 5562 4747 5564
rect 4710 5561 4777 5562
rect 4710 5556 4741 5561
rect 4747 5556 4777 5561
rect 4710 5552 4777 5556
rect 4683 5549 4777 5552
rect 4683 5542 4732 5549
rect 4683 5536 4713 5542
rect 4732 5537 4737 5542
rect 4649 5520 4729 5536
rect 4741 5528 4777 5549
rect 4838 5544 5027 5568
rect 5072 5567 5119 5568
rect 5085 5562 5119 5567
rect 4853 5541 5027 5544
rect 4846 5538 5027 5541
rect 5055 5561 5119 5562
rect 4649 5518 4668 5520
rect 4683 5518 4717 5520
rect 4649 5502 4729 5518
rect 4649 5496 4668 5502
rect 4365 5470 4468 5480
rect 4319 5468 4468 5470
rect 4489 5468 4524 5480
rect 4158 5466 4320 5468
rect 4170 5446 4189 5466
rect 4204 5464 4234 5466
rect 4053 5438 4094 5446
rect 4176 5442 4189 5446
rect 4241 5450 4320 5466
rect 4352 5466 4524 5468
rect 4352 5450 4431 5466
rect 4438 5464 4468 5466
rect 4016 5428 4045 5438
rect 4059 5428 4088 5438
rect 4103 5428 4133 5442
rect 4176 5428 4219 5442
rect 4241 5438 4431 5450
rect 4496 5446 4502 5466
rect 4226 5428 4256 5438
rect 4257 5428 4415 5438
rect 4419 5428 4449 5438
rect 4453 5428 4483 5442
rect 4511 5428 4524 5466
rect 4596 5480 4625 5496
rect 4639 5480 4668 5496
rect 4683 5486 4713 5502
rect 4741 5480 4747 5528
rect 4750 5522 4769 5528
rect 4784 5522 4814 5530
rect 4750 5514 4814 5522
rect 4750 5498 4830 5514
rect 4846 5507 4908 5538
rect 4924 5507 4986 5538
rect 5055 5536 5104 5561
rect 5119 5536 5149 5552
rect 5018 5522 5048 5530
rect 5055 5528 5165 5536
rect 5018 5514 5063 5522
rect 4750 5496 4769 5498
rect 4784 5496 4830 5498
rect 4750 5480 4830 5496
rect 4857 5494 4892 5507
rect 4933 5504 4970 5507
rect 4933 5502 4975 5504
rect 4862 5491 4892 5494
rect 4871 5487 4878 5491
rect 4878 5486 4879 5487
rect 4837 5480 4847 5486
rect 4596 5472 4631 5480
rect 4596 5446 4597 5472
rect 4604 5446 4631 5472
rect 4539 5428 4569 5442
rect 4596 5438 4631 5446
rect 4633 5472 4674 5480
rect 4633 5446 4648 5472
rect 4655 5446 4674 5472
rect 4738 5468 4769 5480
rect 4784 5468 4887 5480
rect 4899 5470 4925 5496
rect 4940 5491 4970 5502
rect 5002 5498 5064 5514
rect 5002 5496 5048 5498
rect 5002 5480 5064 5496
rect 5076 5480 5082 5528
rect 5085 5520 5165 5528
rect 5085 5518 5104 5520
rect 5119 5518 5153 5520
rect 5085 5502 5165 5518
rect 5085 5480 5104 5502
rect 5119 5486 5149 5502
rect 5177 5496 5183 5570
rect 5186 5496 5205 5640
rect 5220 5496 5226 5640
rect 5235 5570 5248 5640
rect 5300 5636 5322 5640
rect 5293 5614 5322 5628
rect 5375 5614 5391 5628
rect 5429 5624 5435 5626
rect 5442 5624 5550 5640
rect 5557 5624 5563 5626
rect 5571 5624 5586 5640
rect 5652 5634 5671 5637
rect 5293 5612 5391 5614
rect 5418 5612 5586 5624
rect 5601 5614 5617 5628
rect 5652 5615 5674 5634
rect 5684 5628 5700 5629
rect 5683 5626 5700 5628
rect 5684 5621 5700 5626
rect 5674 5614 5680 5615
rect 5683 5614 5712 5621
rect 5601 5613 5712 5614
rect 5601 5612 5718 5613
rect 5277 5604 5328 5612
rect 5375 5604 5409 5612
rect 5277 5592 5302 5604
rect 5309 5592 5328 5604
rect 5382 5602 5409 5604
rect 5418 5602 5639 5612
rect 5674 5609 5680 5612
rect 5382 5598 5639 5602
rect 5277 5584 5328 5592
rect 5375 5584 5639 5598
rect 5683 5604 5718 5612
rect 5229 5536 5248 5570
rect 5293 5576 5322 5584
rect 5293 5570 5310 5576
rect 5293 5568 5327 5570
rect 5375 5568 5391 5584
rect 5392 5574 5600 5584
rect 5601 5574 5617 5584
rect 5665 5580 5680 5595
rect 5683 5592 5684 5604
rect 5691 5592 5718 5604
rect 5683 5584 5718 5592
rect 5683 5583 5712 5584
rect 5403 5570 5617 5574
rect 5418 5568 5617 5570
rect 5652 5570 5665 5580
rect 5683 5570 5700 5583
rect 5652 5568 5700 5570
rect 5294 5564 5327 5568
rect 5290 5562 5327 5564
rect 5290 5561 5357 5562
rect 5290 5556 5321 5561
rect 5327 5556 5357 5561
rect 5290 5552 5357 5556
rect 5263 5549 5357 5552
rect 5263 5542 5312 5549
rect 5263 5536 5293 5542
rect 5312 5537 5317 5542
rect 5229 5520 5309 5536
rect 5321 5528 5357 5549
rect 5418 5544 5607 5568
rect 5652 5567 5699 5568
rect 5665 5562 5699 5567
rect 5433 5541 5607 5544
rect 5426 5538 5607 5541
rect 5635 5561 5699 5562
rect 5229 5518 5248 5520
rect 5263 5518 5297 5520
rect 5229 5502 5309 5518
rect 5229 5496 5248 5502
rect 4945 5470 5048 5480
rect 4899 5468 5048 5470
rect 5069 5468 5104 5480
rect 4738 5466 4900 5468
rect 4750 5446 4769 5466
rect 4784 5464 4814 5466
rect 4633 5438 4674 5446
rect 4756 5442 4769 5446
rect 4821 5450 4900 5466
rect 4932 5466 5104 5468
rect 4932 5450 5011 5466
rect 5018 5464 5048 5466
rect 4596 5428 4625 5438
rect 4639 5428 4668 5438
rect 4683 5428 4713 5442
rect 4756 5428 4799 5442
rect 4821 5438 5011 5450
rect 5076 5446 5082 5466
rect 4806 5428 4836 5438
rect 4837 5428 4995 5438
rect 4999 5428 5029 5438
rect 5033 5428 5063 5442
rect 5091 5428 5104 5466
rect 5176 5480 5205 5496
rect 5219 5480 5248 5496
rect 5263 5486 5293 5502
rect 5321 5480 5327 5528
rect 5330 5522 5349 5528
rect 5364 5522 5394 5530
rect 5330 5514 5394 5522
rect 5330 5498 5410 5514
rect 5426 5507 5488 5538
rect 5504 5507 5566 5538
rect 5635 5536 5684 5561
rect 5699 5536 5729 5552
rect 5598 5522 5628 5530
rect 5635 5528 5745 5536
rect 5598 5514 5643 5522
rect 5330 5496 5349 5498
rect 5364 5496 5410 5498
rect 5330 5480 5410 5496
rect 5437 5494 5472 5507
rect 5513 5504 5550 5507
rect 5513 5502 5555 5504
rect 5442 5491 5472 5494
rect 5451 5487 5458 5491
rect 5458 5486 5459 5487
rect 5417 5480 5427 5486
rect 5176 5472 5211 5480
rect 5176 5446 5177 5472
rect 5184 5446 5211 5472
rect 5119 5428 5149 5442
rect 5176 5438 5211 5446
rect 5213 5472 5254 5480
rect 5213 5446 5228 5472
rect 5235 5446 5254 5472
rect 5318 5468 5349 5480
rect 5364 5468 5467 5480
rect 5479 5470 5505 5496
rect 5520 5491 5550 5502
rect 5582 5498 5644 5514
rect 5582 5496 5628 5498
rect 5582 5480 5644 5496
rect 5656 5480 5662 5528
rect 5665 5520 5745 5528
rect 5665 5518 5684 5520
rect 5699 5518 5733 5520
rect 5665 5502 5745 5518
rect 5665 5480 5684 5502
rect 5699 5486 5729 5502
rect 5757 5496 5763 5570
rect 5766 5496 5785 5640
rect 5800 5496 5806 5640
rect 5815 5570 5828 5640
rect 5880 5636 5902 5640
rect 5873 5614 5902 5628
rect 5955 5614 5971 5628
rect 6009 5624 6015 5626
rect 6022 5624 6130 5640
rect 6137 5624 6143 5626
rect 6151 5624 6166 5640
rect 6232 5634 6251 5637
rect 5873 5612 5971 5614
rect 5998 5612 6166 5624
rect 6181 5614 6197 5628
rect 6232 5615 6254 5634
rect 6264 5628 6280 5629
rect 6263 5626 6280 5628
rect 6264 5621 6280 5626
rect 6254 5614 6260 5615
rect 6263 5614 6292 5621
rect 6181 5613 6292 5614
rect 6181 5612 6298 5613
rect 5857 5604 5908 5612
rect 5955 5604 5989 5612
rect 5857 5592 5882 5604
rect 5889 5592 5908 5604
rect 5962 5602 5989 5604
rect 5998 5602 6219 5612
rect 6254 5609 6260 5612
rect 5962 5598 6219 5602
rect 5857 5584 5908 5592
rect 5955 5584 6219 5598
rect 6263 5604 6298 5612
rect 5809 5536 5828 5570
rect 5873 5576 5902 5584
rect 5873 5570 5890 5576
rect 5873 5568 5907 5570
rect 5955 5568 5971 5584
rect 5972 5574 6180 5584
rect 6181 5574 6197 5584
rect 6245 5580 6260 5595
rect 6263 5592 6264 5604
rect 6271 5592 6298 5604
rect 6263 5584 6298 5592
rect 6263 5583 6292 5584
rect 5983 5570 6197 5574
rect 5998 5568 6197 5570
rect 6232 5570 6245 5580
rect 6263 5570 6280 5583
rect 6232 5568 6280 5570
rect 5874 5564 5907 5568
rect 5870 5562 5907 5564
rect 5870 5561 5937 5562
rect 5870 5556 5901 5561
rect 5907 5556 5937 5561
rect 5870 5552 5937 5556
rect 5843 5549 5937 5552
rect 5843 5542 5892 5549
rect 5843 5536 5873 5542
rect 5892 5537 5897 5542
rect 5809 5520 5889 5536
rect 5901 5528 5937 5549
rect 5998 5544 6187 5568
rect 6232 5567 6279 5568
rect 6245 5562 6279 5567
rect 6013 5541 6187 5544
rect 6006 5538 6187 5541
rect 6215 5561 6279 5562
rect 5809 5518 5828 5520
rect 5843 5518 5877 5520
rect 5809 5502 5889 5518
rect 5809 5496 5828 5502
rect 5525 5470 5628 5480
rect 5479 5468 5628 5470
rect 5649 5468 5684 5480
rect 5318 5466 5480 5468
rect 5330 5446 5349 5466
rect 5364 5464 5394 5466
rect 5213 5438 5254 5446
rect 5336 5442 5349 5446
rect 5401 5450 5480 5466
rect 5512 5466 5684 5468
rect 5512 5450 5591 5466
rect 5598 5464 5628 5466
rect 5176 5428 5205 5438
rect 5219 5428 5248 5438
rect 5263 5428 5293 5442
rect 5336 5428 5379 5442
rect 5401 5438 5591 5450
rect 5656 5446 5662 5466
rect 5386 5428 5416 5438
rect 5417 5428 5575 5438
rect 5579 5428 5609 5438
rect 5613 5428 5643 5442
rect 5671 5428 5684 5466
rect 5756 5480 5785 5496
rect 5799 5480 5828 5496
rect 5843 5486 5873 5502
rect 5901 5480 5907 5528
rect 5910 5522 5929 5528
rect 5944 5522 5974 5530
rect 5910 5514 5974 5522
rect 5910 5498 5990 5514
rect 6006 5507 6068 5538
rect 6084 5507 6146 5538
rect 6215 5536 6264 5561
rect 6279 5536 6309 5552
rect 6178 5522 6208 5530
rect 6215 5528 6325 5536
rect 6178 5514 6223 5522
rect 5910 5496 5929 5498
rect 5944 5496 5990 5498
rect 5910 5480 5990 5496
rect 6017 5494 6052 5507
rect 6093 5504 6130 5507
rect 6093 5502 6135 5504
rect 6022 5491 6052 5494
rect 6031 5487 6038 5491
rect 6038 5486 6039 5487
rect 5997 5480 6007 5486
rect 5756 5472 5791 5480
rect 5756 5446 5757 5472
rect 5764 5446 5791 5472
rect 5699 5428 5729 5442
rect 5756 5438 5791 5446
rect 5793 5472 5834 5480
rect 5793 5446 5808 5472
rect 5815 5446 5834 5472
rect 5898 5468 5929 5480
rect 5944 5468 6047 5480
rect 6059 5470 6085 5496
rect 6100 5491 6130 5502
rect 6162 5498 6224 5514
rect 6162 5496 6208 5498
rect 6162 5480 6224 5496
rect 6236 5480 6242 5528
rect 6245 5520 6325 5528
rect 6245 5518 6264 5520
rect 6279 5518 6313 5520
rect 6245 5502 6325 5518
rect 6245 5480 6264 5502
rect 6279 5486 6309 5502
rect 6337 5496 6343 5570
rect 6346 5496 6365 5640
rect 6380 5496 6386 5640
rect 6395 5570 6408 5640
rect 6460 5636 6482 5640
rect 6453 5614 6482 5628
rect 6535 5614 6551 5628
rect 6589 5624 6595 5626
rect 6602 5624 6710 5640
rect 6717 5624 6723 5626
rect 6731 5624 6746 5640
rect 6812 5634 6831 5637
rect 6453 5612 6551 5614
rect 6578 5612 6746 5624
rect 6761 5614 6777 5628
rect 6812 5615 6834 5634
rect 6844 5628 6860 5629
rect 6843 5626 6860 5628
rect 6844 5621 6860 5626
rect 6834 5614 6840 5615
rect 6843 5614 6872 5621
rect 6761 5613 6872 5614
rect 6761 5612 6878 5613
rect 6437 5604 6488 5612
rect 6535 5604 6569 5612
rect 6437 5592 6462 5604
rect 6469 5592 6488 5604
rect 6542 5602 6569 5604
rect 6578 5602 6799 5612
rect 6834 5609 6840 5612
rect 6542 5598 6799 5602
rect 6437 5584 6488 5592
rect 6535 5584 6799 5598
rect 6843 5604 6878 5612
rect 6389 5536 6408 5570
rect 6453 5576 6482 5584
rect 6453 5570 6470 5576
rect 6453 5568 6487 5570
rect 6535 5568 6551 5584
rect 6552 5574 6760 5584
rect 6761 5574 6777 5584
rect 6825 5580 6840 5595
rect 6843 5592 6844 5604
rect 6851 5592 6878 5604
rect 6843 5584 6878 5592
rect 6843 5583 6872 5584
rect 6563 5570 6777 5574
rect 6578 5568 6777 5570
rect 6812 5570 6825 5580
rect 6843 5570 6860 5583
rect 6812 5568 6860 5570
rect 6454 5564 6487 5568
rect 6450 5562 6487 5564
rect 6450 5561 6517 5562
rect 6450 5556 6481 5561
rect 6487 5556 6517 5561
rect 6450 5552 6517 5556
rect 6423 5549 6517 5552
rect 6423 5542 6472 5549
rect 6423 5536 6453 5542
rect 6472 5537 6477 5542
rect 6389 5520 6469 5536
rect 6481 5528 6517 5549
rect 6578 5544 6767 5568
rect 6812 5567 6859 5568
rect 6825 5562 6859 5567
rect 6593 5541 6767 5544
rect 6586 5538 6767 5541
rect 6795 5561 6859 5562
rect 6389 5518 6408 5520
rect 6423 5518 6457 5520
rect 6389 5502 6469 5518
rect 6389 5496 6408 5502
rect 6105 5470 6208 5480
rect 6059 5468 6208 5470
rect 6229 5468 6264 5480
rect 5898 5466 6060 5468
rect 5910 5446 5929 5466
rect 5944 5464 5974 5466
rect 5793 5438 5834 5446
rect 5916 5442 5929 5446
rect 5981 5450 6060 5466
rect 6092 5466 6264 5468
rect 6092 5450 6171 5466
rect 6178 5464 6208 5466
rect 5756 5428 5785 5438
rect 5799 5428 5828 5438
rect 5843 5428 5873 5442
rect 5916 5428 5959 5442
rect 5981 5438 6171 5450
rect 6236 5446 6242 5466
rect 5966 5428 5996 5438
rect 5997 5428 6155 5438
rect 6159 5428 6189 5438
rect 6193 5428 6223 5442
rect 6251 5428 6264 5466
rect 6336 5480 6365 5496
rect 6379 5480 6408 5496
rect 6423 5486 6453 5502
rect 6481 5480 6487 5528
rect 6490 5522 6509 5528
rect 6524 5522 6554 5530
rect 6490 5514 6554 5522
rect 6490 5498 6570 5514
rect 6586 5507 6648 5538
rect 6664 5507 6726 5538
rect 6795 5536 6844 5561
rect 6859 5536 6889 5552
rect 6758 5522 6788 5530
rect 6795 5528 6905 5536
rect 6758 5514 6803 5522
rect 6490 5496 6509 5498
rect 6524 5496 6570 5498
rect 6490 5480 6570 5496
rect 6597 5494 6632 5507
rect 6673 5504 6710 5507
rect 6673 5502 6715 5504
rect 6602 5491 6632 5494
rect 6611 5487 6618 5491
rect 6618 5486 6619 5487
rect 6577 5480 6587 5486
rect 6336 5472 6371 5480
rect 6336 5446 6337 5472
rect 6344 5446 6371 5472
rect 6279 5428 6309 5442
rect 6336 5438 6371 5446
rect 6373 5472 6414 5480
rect 6373 5446 6388 5472
rect 6395 5446 6414 5472
rect 6478 5468 6509 5480
rect 6524 5468 6627 5480
rect 6639 5470 6665 5496
rect 6680 5491 6710 5502
rect 6742 5498 6804 5514
rect 6742 5496 6788 5498
rect 6742 5480 6804 5496
rect 6816 5480 6822 5528
rect 6825 5520 6905 5528
rect 6825 5518 6844 5520
rect 6859 5518 6893 5520
rect 6825 5502 6905 5518
rect 6825 5480 6844 5502
rect 6859 5486 6889 5502
rect 6917 5496 6923 5570
rect 6926 5496 6945 5640
rect 6960 5496 6966 5640
rect 6975 5570 6988 5640
rect 7040 5636 7062 5640
rect 7033 5614 7062 5628
rect 7115 5614 7131 5628
rect 7169 5624 7175 5626
rect 7182 5624 7290 5640
rect 7297 5624 7303 5626
rect 7311 5624 7326 5640
rect 7392 5634 7411 5637
rect 7033 5612 7131 5614
rect 7158 5612 7326 5624
rect 7341 5614 7357 5628
rect 7392 5615 7414 5634
rect 7424 5628 7440 5629
rect 7423 5626 7440 5628
rect 7424 5621 7440 5626
rect 7414 5614 7420 5615
rect 7423 5614 7452 5621
rect 7341 5613 7452 5614
rect 7341 5612 7458 5613
rect 7017 5604 7068 5612
rect 7115 5604 7149 5612
rect 7017 5592 7042 5604
rect 7049 5592 7068 5604
rect 7122 5602 7149 5604
rect 7158 5602 7379 5612
rect 7414 5609 7420 5612
rect 7122 5598 7379 5602
rect 7017 5584 7068 5592
rect 7115 5584 7379 5598
rect 7423 5604 7458 5612
rect 6969 5536 6988 5570
rect 7033 5576 7062 5584
rect 7033 5570 7050 5576
rect 7033 5568 7067 5570
rect 7115 5568 7131 5584
rect 7132 5574 7340 5584
rect 7341 5574 7357 5584
rect 7405 5580 7420 5595
rect 7423 5592 7424 5604
rect 7431 5592 7458 5604
rect 7423 5584 7458 5592
rect 7423 5583 7452 5584
rect 7143 5570 7357 5574
rect 7158 5568 7357 5570
rect 7392 5570 7405 5580
rect 7423 5570 7440 5583
rect 7392 5568 7440 5570
rect 7034 5564 7067 5568
rect 7030 5562 7067 5564
rect 7030 5561 7097 5562
rect 7030 5556 7061 5561
rect 7067 5556 7097 5561
rect 7030 5552 7097 5556
rect 7003 5549 7097 5552
rect 7003 5542 7052 5549
rect 7003 5536 7033 5542
rect 7052 5537 7057 5542
rect 6969 5520 7049 5536
rect 7061 5528 7097 5549
rect 7158 5544 7347 5568
rect 7392 5567 7439 5568
rect 7405 5562 7439 5567
rect 7173 5541 7347 5544
rect 7166 5538 7347 5541
rect 7375 5561 7439 5562
rect 6969 5518 6988 5520
rect 7003 5518 7037 5520
rect 6969 5502 7049 5518
rect 6969 5496 6988 5502
rect 6685 5470 6788 5480
rect 6639 5468 6788 5470
rect 6809 5468 6844 5480
rect 6478 5466 6640 5468
rect 6490 5446 6509 5466
rect 6524 5464 6554 5466
rect 6373 5438 6414 5446
rect 6496 5442 6509 5446
rect 6561 5450 6640 5466
rect 6672 5466 6844 5468
rect 6672 5450 6751 5466
rect 6758 5464 6788 5466
rect 6336 5428 6365 5438
rect 6379 5428 6408 5438
rect 6423 5428 6453 5442
rect 6496 5428 6539 5442
rect 6561 5438 6751 5450
rect 6816 5446 6822 5466
rect 6546 5428 6576 5438
rect 6577 5428 6735 5438
rect 6739 5428 6769 5438
rect 6773 5428 6803 5442
rect 6831 5428 6844 5466
rect 6916 5480 6945 5496
rect 6959 5480 6988 5496
rect 7003 5486 7033 5502
rect 7061 5480 7067 5528
rect 7070 5522 7089 5528
rect 7104 5522 7134 5530
rect 7070 5514 7134 5522
rect 7070 5498 7150 5514
rect 7166 5507 7228 5538
rect 7244 5507 7306 5538
rect 7375 5536 7424 5561
rect 7439 5536 7469 5552
rect 7338 5522 7368 5530
rect 7375 5528 7485 5536
rect 7338 5514 7383 5522
rect 7070 5496 7089 5498
rect 7104 5496 7150 5498
rect 7070 5480 7150 5496
rect 7177 5494 7212 5507
rect 7253 5504 7290 5507
rect 7253 5502 7295 5504
rect 7182 5491 7212 5494
rect 7191 5487 7198 5491
rect 7198 5486 7199 5487
rect 7157 5480 7167 5486
rect 6916 5472 6951 5480
rect 6916 5446 6917 5472
rect 6924 5446 6951 5472
rect 6859 5428 6889 5442
rect 6916 5438 6951 5446
rect 6953 5472 6994 5480
rect 6953 5446 6968 5472
rect 6975 5446 6994 5472
rect 7058 5468 7089 5480
rect 7104 5468 7207 5480
rect 7219 5470 7245 5496
rect 7260 5491 7290 5502
rect 7322 5498 7384 5514
rect 7322 5496 7368 5498
rect 7322 5480 7384 5496
rect 7396 5480 7402 5528
rect 7405 5520 7485 5528
rect 7405 5518 7424 5520
rect 7439 5518 7473 5520
rect 7405 5502 7485 5518
rect 7405 5480 7424 5502
rect 7439 5486 7469 5502
rect 7497 5496 7503 5570
rect 7506 5496 7525 5640
rect 7540 5496 7546 5640
rect 7555 5570 7568 5640
rect 7620 5636 7642 5640
rect 7613 5614 7642 5628
rect 7695 5614 7711 5628
rect 7749 5624 7755 5626
rect 7762 5624 7870 5640
rect 7877 5624 7883 5626
rect 7891 5624 7906 5640
rect 7972 5634 7991 5637
rect 7613 5612 7711 5614
rect 7738 5612 7906 5624
rect 7921 5614 7937 5628
rect 7972 5615 7994 5634
rect 8004 5628 8020 5629
rect 8003 5626 8020 5628
rect 8004 5621 8020 5626
rect 7994 5614 8000 5615
rect 8003 5614 8032 5621
rect 7921 5613 8032 5614
rect 7921 5612 8038 5613
rect 7597 5604 7648 5612
rect 7695 5604 7729 5612
rect 7597 5592 7622 5604
rect 7629 5592 7648 5604
rect 7702 5602 7729 5604
rect 7738 5602 7959 5612
rect 7994 5609 8000 5612
rect 7702 5598 7959 5602
rect 7597 5584 7648 5592
rect 7695 5584 7959 5598
rect 8003 5604 8038 5612
rect 7549 5536 7568 5570
rect 7613 5576 7642 5584
rect 7613 5570 7630 5576
rect 7613 5568 7647 5570
rect 7695 5568 7711 5584
rect 7712 5574 7920 5584
rect 7921 5574 7937 5584
rect 7985 5580 8000 5595
rect 8003 5592 8004 5604
rect 8011 5592 8038 5604
rect 8003 5584 8038 5592
rect 8003 5583 8032 5584
rect 7723 5570 7937 5574
rect 7738 5568 7937 5570
rect 7972 5570 7985 5580
rect 8003 5570 8020 5583
rect 7972 5568 8020 5570
rect 7614 5564 7647 5568
rect 7610 5562 7647 5564
rect 7610 5561 7677 5562
rect 7610 5556 7641 5561
rect 7647 5556 7677 5561
rect 7610 5552 7677 5556
rect 7583 5549 7677 5552
rect 7583 5542 7632 5549
rect 7583 5536 7613 5542
rect 7632 5537 7637 5542
rect 7549 5520 7629 5536
rect 7641 5528 7677 5549
rect 7738 5544 7927 5568
rect 7972 5567 8019 5568
rect 7985 5562 8019 5567
rect 7753 5541 7927 5544
rect 7746 5538 7927 5541
rect 7955 5561 8019 5562
rect 7549 5518 7568 5520
rect 7583 5518 7617 5520
rect 7549 5502 7629 5518
rect 7549 5496 7568 5502
rect 7265 5470 7368 5480
rect 7219 5468 7368 5470
rect 7389 5468 7424 5480
rect 7058 5466 7220 5468
rect 7070 5446 7089 5466
rect 7104 5464 7134 5466
rect 6953 5438 6994 5446
rect 7076 5442 7089 5446
rect 7141 5450 7220 5466
rect 7252 5466 7424 5468
rect 7252 5450 7331 5466
rect 7338 5464 7368 5466
rect 6916 5428 6945 5438
rect 6959 5428 6988 5438
rect 7003 5428 7033 5442
rect 7076 5428 7119 5442
rect 7141 5438 7331 5450
rect 7396 5446 7402 5466
rect 7126 5428 7156 5438
rect 7157 5428 7315 5438
rect 7319 5428 7349 5438
rect 7353 5428 7383 5442
rect 7411 5428 7424 5466
rect 7496 5480 7525 5496
rect 7539 5480 7568 5496
rect 7583 5486 7613 5502
rect 7641 5480 7647 5528
rect 7650 5522 7669 5528
rect 7684 5522 7714 5530
rect 7650 5514 7714 5522
rect 7650 5498 7730 5514
rect 7746 5507 7808 5538
rect 7824 5507 7886 5538
rect 7955 5536 8004 5561
rect 8019 5536 8049 5552
rect 7918 5522 7948 5530
rect 7955 5528 8065 5536
rect 7918 5514 7963 5522
rect 7650 5496 7669 5498
rect 7684 5496 7730 5498
rect 7650 5480 7730 5496
rect 7757 5494 7792 5507
rect 7833 5504 7870 5507
rect 7833 5502 7875 5504
rect 7762 5491 7792 5494
rect 7771 5487 7778 5491
rect 7778 5486 7779 5487
rect 7737 5480 7747 5486
rect 7496 5472 7531 5480
rect 7496 5446 7497 5472
rect 7504 5446 7531 5472
rect 7439 5428 7469 5442
rect 7496 5438 7531 5446
rect 7533 5472 7574 5480
rect 7533 5446 7548 5472
rect 7555 5446 7574 5472
rect 7638 5468 7669 5480
rect 7684 5468 7787 5480
rect 7799 5470 7825 5496
rect 7840 5491 7870 5502
rect 7902 5498 7964 5514
rect 7902 5496 7948 5498
rect 7902 5480 7964 5496
rect 7976 5480 7982 5528
rect 7985 5520 8065 5528
rect 7985 5518 8004 5520
rect 8019 5518 8053 5520
rect 7985 5502 8065 5518
rect 7985 5480 8004 5502
rect 8019 5486 8049 5502
rect 8077 5496 8083 5570
rect 8086 5496 8105 5640
rect 8120 5496 8126 5640
rect 8135 5570 8148 5640
rect 8200 5636 8222 5640
rect 8193 5614 8222 5628
rect 8275 5614 8291 5628
rect 8329 5624 8335 5626
rect 8342 5624 8450 5640
rect 8457 5624 8463 5626
rect 8471 5624 8486 5640
rect 8552 5634 8571 5637
rect 8193 5612 8291 5614
rect 8318 5612 8486 5624
rect 8501 5614 8517 5628
rect 8552 5615 8574 5634
rect 8584 5628 8600 5629
rect 8583 5626 8600 5628
rect 8584 5621 8600 5626
rect 8574 5614 8580 5615
rect 8583 5614 8612 5621
rect 8501 5613 8612 5614
rect 8501 5612 8618 5613
rect 8177 5604 8228 5612
rect 8275 5604 8309 5612
rect 8177 5592 8202 5604
rect 8209 5592 8228 5604
rect 8282 5602 8309 5604
rect 8318 5602 8539 5612
rect 8574 5609 8580 5612
rect 8282 5598 8539 5602
rect 8177 5584 8228 5592
rect 8275 5584 8539 5598
rect 8583 5604 8618 5612
rect 8129 5536 8148 5570
rect 8193 5576 8222 5584
rect 8193 5570 8210 5576
rect 8193 5568 8227 5570
rect 8275 5568 8291 5584
rect 8292 5574 8500 5584
rect 8501 5574 8517 5584
rect 8565 5580 8580 5595
rect 8583 5592 8584 5604
rect 8591 5592 8618 5604
rect 8583 5584 8618 5592
rect 8583 5583 8612 5584
rect 8303 5570 8517 5574
rect 8318 5568 8517 5570
rect 8552 5570 8565 5580
rect 8583 5570 8600 5583
rect 8552 5568 8600 5570
rect 8194 5564 8227 5568
rect 8190 5562 8227 5564
rect 8190 5561 8257 5562
rect 8190 5556 8221 5561
rect 8227 5556 8257 5561
rect 8190 5552 8257 5556
rect 8163 5549 8257 5552
rect 8163 5542 8212 5549
rect 8163 5536 8193 5542
rect 8212 5537 8217 5542
rect 8129 5520 8209 5536
rect 8221 5528 8257 5549
rect 8318 5544 8507 5568
rect 8552 5567 8599 5568
rect 8565 5562 8599 5567
rect 8333 5541 8507 5544
rect 8326 5538 8507 5541
rect 8535 5561 8599 5562
rect 8129 5518 8148 5520
rect 8163 5518 8197 5520
rect 8129 5502 8209 5518
rect 8129 5496 8148 5502
rect 7845 5470 7948 5480
rect 7799 5468 7948 5470
rect 7969 5468 8004 5480
rect 7638 5466 7800 5468
rect 7650 5446 7669 5466
rect 7684 5464 7714 5466
rect 7533 5438 7574 5446
rect 7656 5442 7669 5446
rect 7721 5450 7800 5466
rect 7832 5466 8004 5468
rect 7832 5450 7911 5466
rect 7918 5464 7948 5466
rect 7496 5428 7525 5438
rect 7539 5428 7568 5438
rect 7583 5428 7613 5442
rect 7656 5428 7699 5442
rect 7721 5438 7911 5450
rect 7976 5446 7982 5466
rect 7706 5428 7736 5438
rect 7737 5428 7895 5438
rect 7899 5428 7929 5438
rect 7933 5428 7963 5442
rect 7991 5428 8004 5466
rect 8076 5480 8105 5496
rect 8119 5480 8148 5496
rect 8163 5486 8193 5502
rect 8221 5480 8227 5528
rect 8230 5522 8249 5528
rect 8264 5522 8294 5530
rect 8230 5514 8294 5522
rect 8230 5498 8310 5514
rect 8326 5507 8388 5538
rect 8404 5507 8466 5538
rect 8535 5536 8584 5561
rect 8599 5536 8629 5552
rect 8498 5522 8528 5530
rect 8535 5528 8645 5536
rect 8498 5514 8543 5522
rect 8230 5496 8249 5498
rect 8264 5496 8310 5498
rect 8230 5480 8310 5496
rect 8337 5494 8372 5507
rect 8413 5504 8450 5507
rect 8413 5502 8455 5504
rect 8342 5491 8372 5494
rect 8351 5487 8358 5491
rect 8358 5486 8359 5487
rect 8317 5480 8327 5486
rect 8076 5472 8111 5480
rect 8076 5446 8077 5472
rect 8084 5446 8111 5472
rect 8019 5428 8049 5442
rect 8076 5438 8111 5446
rect 8113 5472 8154 5480
rect 8113 5446 8128 5472
rect 8135 5446 8154 5472
rect 8218 5468 8249 5480
rect 8264 5468 8367 5480
rect 8379 5470 8405 5496
rect 8420 5491 8450 5502
rect 8482 5498 8544 5514
rect 8482 5496 8528 5498
rect 8482 5480 8544 5496
rect 8556 5480 8562 5528
rect 8565 5520 8645 5528
rect 8565 5518 8584 5520
rect 8599 5518 8633 5520
rect 8565 5502 8645 5518
rect 8565 5480 8584 5502
rect 8599 5486 8629 5502
rect 8657 5496 8663 5570
rect 8666 5496 8685 5640
rect 8700 5496 8706 5640
rect 8715 5570 8728 5640
rect 8780 5636 8802 5640
rect 8773 5614 8802 5628
rect 8855 5614 8871 5628
rect 8909 5624 8915 5626
rect 8922 5624 9030 5640
rect 9037 5624 9043 5626
rect 9051 5624 9066 5640
rect 9132 5634 9151 5637
rect 8773 5612 8871 5614
rect 8898 5612 9066 5624
rect 9081 5614 9097 5628
rect 9132 5615 9154 5634
rect 9164 5628 9180 5629
rect 9163 5626 9180 5628
rect 9164 5621 9180 5626
rect 9154 5614 9160 5615
rect 9163 5614 9192 5621
rect 9081 5613 9192 5614
rect 9081 5612 9198 5613
rect 8757 5604 8808 5612
rect 8855 5604 8889 5612
rect 8757 5592 8782 5604
rect 8789 5592 8808 5604
rect 8862 5602 8889 5604
rect 8898 5602 9119 5612
rect 9154 5609 9160 5612
rect 8862 5598 9119 5602
rect 8757 5584 8808 5592
rect 8855 5584 9119 5598
rect 9163 5604 9198 5612
rect 8709 5536 8728 5570
rect 8773 5576 8802 5584
rect 8773 5570 8790 5576
rect 8773 5568 8807 5570
rect 8855 5568 8871 5584
rect 8872 5574 9080 5584
rect 9081 5574 9097 5584
rect 9145 5580 9160 5595
rect 9163 5592 9164 5604
rect 9171 5592 9198 5604
rect 9163 5584 9198 5592
rect 9163 5583 9192 5584
rect 8883 5570 9097 5574
rect 8898 5568 9097 5570
rect 9132 5570 9145 5580
rect 9163 5570 9180 5583
rect 9132 5568 9180 5570
rect 8774 5564 8807 5568
rect 8770 5562 8807 5564
rect 8770 5561 8837 5562
rect 8770 5556 8801 5561
rect 8807 5556 8837 5561
rect 8770 5552 8837 5556
rect 8743 5549 8837 5552
rect 8743 5542 8792 5549
rect 8743 5536 8773 5542
rect 8792 5537 8797 5542
rect 8709 5520 8789 5536
rect 8801 5528 8837 5549
rect 8898 5544 9087 5568
rect 9132 5567 9179 5568
rect 9145 5562 9179 5567
rect 8913 5541 9087 5544
rect 8906 5538 9087 5541
rect 9115 5561 9179 5562
rect 8709 5518 8728 5520
rect 8743 5518 8777 5520
rect 8709 5502 8789 5518
rect 8709 5496 8728 5502
rect 8425 5470 8528 5480
rect 8379 5468 8528 5470
rect 8549 5468 8584 5480
rect 8218 5466 8380 5468
rect 8230 5446 8249 5466
rect 8264 5464 8294 5466
rect 8113 5438 8154 5446
rect 8236 5442 8249 5446
rect 8301 5450 8380 5466
rect 8412 5466 8584 5468
rect 8412 5450 8491 5466
rect 8498 5464 8528 5466
rect 8076 5428 8105 5438
rect 8119 5428 8148 5438
rect 8163 5428 8193 5442
rect 8236 5428 8279 5442
rect 8301 5438 8491 5450
rect 8556 5446 8562 5466
rect 8286 5428 8316 5438
rect 8317 5428 8475 5438
rect 8479 5428 8509 5438
rect 8513 5428 8543 5442
rect 8571 5428 8584 5466
rect 8656 5480 8685 5496
rect 8699 5480 8728 5496
rect 8743 5486 8773 5502
rect 8801 5480 8807 5528
rect 8810 5522 8829 5528
rect 8844 5522 8874 5530
rect 8810 5514 8874 5522
rect 8810 5498 8890 5514
rect 8906 5507 8968 5538
rect 8984 5507 9046 5538
rect 9115 5536 9164 5561
rect 9179 5536 9209 5552
rect 9078 5522 9108 5530
rect 9115 5528 9225 5536
rect 9078 5514 9123 5522
rect 8810 5496 8829 5498
rect 8844 5496 8890 5498
rect 8810 5480 8890 5496
rect 8917 5494 8952 5507
rect 8993 5504 9030 5507
rect 8993 5502 9035 5504
rect 8922 5491 8952 5494
rect 8931 5487 8938 5491
rect 8938 5486 8939 5487
rect 8897 5480 8907 5486
rect 8656 5472 8691 5480
rect 8656 5446 8657 5472
rect 8664 5446 8691 5472
rect 8599 5428 8629 5442
rect 8656 5438 8691 5446
rect 8693 5472 8734 5480
rect 8693 5446 8708 5472
rect 8715 5446 8734 5472
rect 8798 5468 8829 5480
rect 8844 5468 8947 5480
rect 8959 5470 8985 5496
rect 9000 5491 9030 5502
rect 9062 5498 9124 5514
rect 9062 5496 9108 5498
rect 9062 5480 9124 5496
rect 9136 5480 9142 5528
rect 9145 5520 9225 5528
rect 9145 5518 9164 5520
rect 9179 5518 9213 5520
rect 9145 5502 9225 5518
rect 9145 5480 9164 5502
rect 9179 5486 9209 5502
rect 9237 5496 9243 5570
rect 9246 5496 9265 5640
rect 9280 5496 9286 5640
rect 9295 5570 9308 5640
rect 9360 5636 9382 5640
rect 9353 5614 9382 5628
rect 9435 5614 9451 5628
rect 9489 5624 9495 5626
rect 9502 5624 9610 5640
rect 9617 5624 9623 5626
rect 9631 5624 9646 5640
rect 9712 5634 9731 5637
rect 9353 5612 9451 5614
rect 9478 5612 9646 5624
rect 9661 5614 9677 5628
rect 9712 5615 9734 5634
rect 9744 5628 9760 5629
rect 9743 5626 9760 5628
rect 9744 5621 9760 5626
rect 9734 5614 9740 5615
rect 9743 5614 9772 5621
rect 9661 5613 9772 5614
rect 9661 5612 9778 5613
rect 9337 5604 9388 5612
rect 9435 5604 9469 5612
rect 9337 5592 9362 5604
rect 9369 5592 9388 5604
rect 9442 5602 9469 5604
rect 9478 5602 9699 5612
rect 9734 5609 9740 5612
rect 9442 5598 9699 5602
rect 9337 5584 9388 5592
rect 9435 5584 9699 5598
rect 9743 5604 9778 5612
rect 9289 5536 9308 5570
rect 9353 5576 9382 5584
rect 9353 5570 9370 5576
rect 9353 5568 9387 5570
rect 9435 5568 9451 5584
rect 9452 5574 9660 5584
rect 9661 5574 9677 5584
rect 9725 5580 9740 5595
rect 9743 5592 9744 5604
rect 9751 5592 9778 5604
rect 9743 5584 9778 5592
rect 9743 5583 9772 5584
rect 9463 5570 9677 5574
rect 9478 5568 9677 5570
rect 9712 5570 9725 5580
rect 9743 5570 9760 5583
rect 9712 5568 9760 5570
rect 9354 5564 9387 5568
rect 9350 5562 9387 5564
rect 9350 5561 9417 5562
rect 9350 5556 9381 5561
rect 9387 5556 9417 5561
rect 9350 5552 9417 5556
rect 9323 5549 9417 5552
rect 9323 5542 9372 5549
rect 9323 5536 9353 5542
rect 9372 5537 9377 5542
rect 9289 5520 9369 5536
rect 9381 5528 9417 5549
rect 9478 5544 9667 5568
rect 9712 5567 9759 5568
rect 9725 5562 9759 5567
rect 9493 5541 9667 5544
rect 9486 5538 9667 5541
rect 9695 5561 9759 5562
rect 9289 5518 9308 5520
rect 9323 5518 9357 5520
rect 9289 5502 9369 5518
rect 9289 5496 9308 5502
rect 9005 5470 9108 5480
rect 8959 5468 9108 5470
rect 9129 5468 9164 5480
rect 8798 5466 8960 5468
rect 8810 5446 8829 5466
rect 8844 5464 8874 5466
rect 8693 5438 8734 5446
rect 8816 5442 8829 5446
rect 8881 5450 8960 5466
rect 8992 5466 9164 5468
rect 8992 5450 9071 5466
rect 9078 5464 9108 5466
rect 8656 5428 8685 5438
rect 8699 5428 8728 5438
rect 8743 5428 8773 5442
rect 8816 5428 8859 5442
rect 8881 5438 9071 5450
rect 9136 5446 9142 5466
rect 8866 5428 8896 5438
rect 8897 5428 9055 5438
rect 9059 5428 9089 5438
rect 9093 5428 9123 5442
rect 9151 5428 9164 5466
rect 9236 5480 9265 5496
rect 9279 5480 9308 5496
rect 9323 5486 9353 5502
rect 9381 5480 9387 5528
rect 9390 5522 9409 5528
rect 9424 5522 9454 5530
rect 9390 5514 9454 5522
rect 9390 5498 9470 5514
rect 9486 5507 9548 5538
rect 9564 5507 9626 5538
rect 9695 5536 9744 5561
rect 9759 5536 9789 5552
rect 9658 5522 9688 5530
rect 9695 5528 9805 5536
rect 9658 5514 9703 5522
rect 9390 5496 9409 5498
rect 9424 5496 9470 5498
rect 9390 5480 9470 5496
rect 9497 5494 9532 5507
rect 9573 5504 9610 5507
rect 9573 5502 9615 5504
rect 9502 5491 9532 5494
rect 9511 5487 9518 5491
rect 9518 5486 9519 5487
rect 9477 5480 9487 5486
rect 9236 5472 9271 5480
rect 9236 5446 9237 5472
rect 9244 5446 9271 5472
rect 9179 5428 9209 5442
rect 9236 5438 9271 5446
rect 9273 5472 9314 5480
rect 9273 5446 9288 5472
rect 9295 5446 9314 5472
rect 9378 5468 9409 5480
rect 9424 5468 9527 5480
rect 9539 5470 9565 5496
rect 9580 5491 9610 5502
rect 9642 5498 9704 5514
rect 9642 5496 9688 5498
rect 9642 5480 9704 5496
rect 9716 5480 9722 5528
rect 9725 5520 9805 5528
rect 9725 5518 9744 5520
rect 9759 5518 9793 5520
rect 9725 5502 9805 5518
rect 9725 5480 9744 5502
rect 9759 5486 9789 5502
rect 9817 5496 9823 5570
rect 9826 5496 9845 5640
rect 9860 5496 9866 5640
rect 9875 5570 9888 5640
rect 9940 5636 9962 5640
rect 9933 5614 9962 5628
rect 10015 5614 10031 5628
rect 10069 5624 10075 5626
rect 10082 5624 10190 5640
rect 10197 5624 10203 5626
rect 10211 5624 10226 5640
rect 10292 5634 10311 5637
rect 9933 5612 10031 5614
rect 10058 5612 10226 5624
rect 10241 5614 10257 5628
rect 10292 5615 10314 5634
rect 10324 5628 10340 5629
rect 10323 5626 10340 5628
rect 10324 5621 10340 5626
rect 10314 5614 10320 5615
rect 10323 5614 10352 5621
rect 10241 5613 10352 5614
rect 10241 5612 10358 5613
rect 9917 5604 9968 5612
rect 10015 5604 10049 5612
rect 9917 5592 9942 5604
rect 9949 5592 9968 5604
rect 10022 5602 10049 5604
rect 10058 5602 10279 5612
rect 10314 5609 10320 5612
rect 10022 5598 10279 5602
rect 9917 5584 9968 5592
rect 10015 5584 10279 5598
rect 10323 5604 10358 5612
rect 9869 5536 9888 5570
rect 9933 5576 9962 5584
rect 9933 5570 9950 5576
rect 9933 5568 9967 5570
rect 10015 5568 10031 5584
rect 10032 5574 10240 5584
rect 10241 5574 10257 5584
rect 10305 5580 10320 5595
rect 10323 5592 10324 5604
rect 10331 5592 10358 5604
rect 10323 5584 10358 5592
rect 10323 5583 10352 5584
rect 10043 5570 10257 5574
rect 10058 5568 10257 5570
rect 10292 5570 10305 5580
rect 10323 5570 10340 5583
rect 10292 5568 10340 5570
rect 9934 5564 9967 5568
rect 9930 5562 9967 5564
rect 9930 5561 9997 5562
rect 9930 5556 9961 5561
rect 9967 5556 9997 5561
rect 9930 5552 9997 5556
rect 9903 5549 9997 5552
rect 9903 5542 9952 5549
rect 9903 5536 9933 5542
rect 9952 5537 9957 5542
rect 9869 5520 9949 5536
rect 9961 5528 9997 5549
rect 10058 5544 10247 5568
rect 10292 5567 10339 5568
rect 10305 5562 10339 5567
rect 10073 5541 10247 5544
rect 10066 5538 10247 5541
rect 10275 5561 10339 5562
rect 9869 5518 9888 5520
rect 9903 5518 9937 5520
rect 9869 5502 9949 5518
rect 9869 5496 9888 5502
rect 9585 5470 9688 5480
rect 9539 5468 9688 5470
rect 9709 5468 9744 5480
rect 9378 5466 9540 5468
rect 9390 5446 9409 5466
rect 9424 5464 9454 5466
rect 9273 5438 9314 5446
rect 9396 5442 9409 5446
rect 9461 5450 9540 5466
rect 9572 5466 9744 5468
rect 9572 5450 9651 5466
rect 9658 5464 9688 5466
rect 9236 5428 9265 5438
rect 9279 5428 9308 5438
rect 9323 5428 9353 5442
rect 9396 5428 9439 5442
rect 9461 5438 9651 5450
rect 9716 5446 9722 5466
rect 9446 5428 9476 5438
rect 9477 5428 9635 5438
rect 9639 5428 9669 5438
rect 9673 5428 9703 5442
rect 9731 5428 9744 5466
rect 9816 5480 9845 5496
rect 9859 5480 9888 5496
rect 9903 5486 9933 5502
rect 9961 5480 9967 5528
rect 9970 5522 9989 5528
rect 10004 5522 10034 5530
rect 9970 5514 10034 5522
rect 9970 5498 10050 5514
rect 10066 5507 10128 5538
rect 10144 5507 10206 5538
rect 10275 5536 10324 5561
rect 10339 5536 10369 5552
rect 10238 5522 10268 5530
rect 10275 5528 10385 5536
rect 10238 5514 10283 5522
rect 9970 5496 9989 5498
rect 10004 5496 10050 5498
rect 9970 5480 10050 5496
rect 10077 5494 10112 5507
rect 10153 5504 10190 5507
rect 10153 5502 10195 5504
rect 10082 5491 10112 5494
rect 10091 5487 10098 5491
rect 10098 5486 10099 5487
rect 10057 5480 10067 5486
rect 9816 5472 9851 5480
rect 9816 5446 9817 5472
rect 9824 5446 9851 5472
rect 9759 5428 9789 5442
rect 9816 5438 9851 5446
rect 9853 5472 9894 5480
rect 9853 5446 9868 5472
rect 9875 5446 9894 5472
rect 9958 5468 9989 5480
rect 10004 5468 10107 5480
rect 10119 5470 10145 5496
rect 10160 5491 10190 5502
rect 10222 5498 10284 5514
rect 10222 5496 10268 5498
rect 10222 5480 10284 5496
rect 10296 5480 10302 5528
rect 10305 5520 10385 5528
rect 10305 5518 10324 5520
rect 10339 5518 10373 5520
rect 10305 5502 10385 5518
rect 10305 5480 10324 5502
rect 10339 5486 10369 5502
rect 10397 5496 10403 5570
rect 10406 5496 10425 5640
rect 10440 5496 10446 5640
rect 10455 5570 10468 5640
rect 10520 5636 10542 5640
rect 10513 5614 10542 5628
rect 10595 5614 10611 5628
rect 10649 5624 10655 5626
rect 10662 5624 10770 5640
rect 10777 5624 10783 5626
rect 10791 5624 10806 5640
rect 10872 5634 10891 5637
rect 10513 5612 10611 5614
rect 10638 5612 10806 5624
rect 10821 5614 10837 5628
rect 10872 5615 10894 5634
rect 10904 5628 10920 5629
rect 10903 5626 10920 5628
rect 10904 5621 10920 5626
rect 10894 5614 10900 5615
rect 10903 5614 10932 5621
rect 10821 5613 10932 5614
rect 10821 5612 10938 5613
rect 10497 5604 10548 5612
rect 10595 5604 10629 5612
rect 10497 5592 10522 5604
rect 10529 5592 10548 5604
rect 10602 5602 10629 5604
rect 10638 5602 10859 5612
rect 10894 5609 10900 5612
rect 10602 5598 10859 5602
rect 10497 5584 10548 5592
rect 10595 5584 10859 5598
rect 10903 5604 10938 5612
rect 10449 5536 10468 5570
rect 10513 5576 10542 5584
rect 10513 5570 10530 5576
rect 10513 5568 10547 5570
rect 10595 5568 10611 5584
rect 10612 5574 10820 5584
rect 10821 5574 10837 5584
rect 10885 5580 10900 5595
rect 10903 5592 10904 5604
rect 10911 5592 10938 5604
rect 10903 5584 10938 5592
rect 10903 5583 10932 5584
rect 10623 5570 10837 5574
rect 10638 5568 10837 5570
rect 10872 5570 10885 5580
rect 10903 5570 10920 5583
rect 10872 5568 10920 5570
rect 10514 5564 10547 5568
rect 10510 5562 10547 5564
rect 10510 5561 10577 5562
rect 10510 5556 10541 5561
rect 10547 5556 10577 5561
rect 10510 5552 10577 5556
rect 10483 5549 10577 5552
rect 10483 5542 10532 5549
rect 10483 5536 10513 5542
rect 10532 5537 10537 5542
rect 10449 5520 10529 5536
rect 10541 5528 10577 5549
rect 10638 5544 10827 5568
rect 10872 5567 10919 5568
rect 10885 5562 10919 5567
rect 10653 5541 10827 5544
rect 10646 5538 10827 5541
rect 10855 5561 10919 5562
rect 10449 5518 10468 5520
rect 10483 5518 10517 5520
rect 10449 5502 10529 5518
rect 10449 5496 10468 5502
rect 10165 5470 10268 5480
rect 10119 5468 10268 5470
rect 10289 5468 10324 5480
rect 9958 5466 10120 5468
rect 9970 5446 9989 5466
rect 10004 5464 10034 5466
rect 9853 5438 9894 5446
rect 9976 5442 9989 5446
rect 10041 5450 10120 5466
rect 10152 5466 10324 5468
rect 10152 5450 10231 5466
rect 10238 5464 10268 5466
rect 9816 5428 9845 5438
rect 9859 5428 9888 5438
rect 9903 5428 9933 5442
rect 9976 5428 10019 5442
rect 10041 5438 10231 5450
rect 10296 5446 10302 5466
rect 10026 5428 10056 5438
rect 10057 5428 10215 5438
rect 10219 5428 10249 5438
rect 10253 5428 10283 5442
rect 10311 5428 10324 5466
rect 10396 5480 10425 5496
rect 10439 5480 10468 5496
rect 10483 5486 10513 5502
rect 10541 5480 10547 5528
rect 10550 5522 10569 5528
rect 10584 5522 10614 5530
rect 10550 5514 10614 5522
rect 10550 5498 10630 5514
rect 10646 5507 10708 5538
rect 10724 5507 10786 5538
rect 10855 5536 10904 5561
rect 10919 5536 10949 5552
rect 10818 5522 10848 5530
rect 10855 5528 10965 5536
rect 10818 5514 10863 5522
rect 10550 5496 10569 5498
rect 10584 5496 10630 5498
rect 10550 5480 10630 5496
rect 10657 5494 10692 5507
rect 10733 5504 10770 5507
rect 10733 5502 10775 5504
rect 10662 5491 10692 5494
rect 10671 5487 10678 5491
rect 10678 5486 10679 5487
rect 10637 5480 10647 5486
rect 10396 5472 10431 5480
rect 10396 5446 10397 5472
rect 10404 5446 10431 5472
rect 10339 5428 10369 5442
rect 10396 5438 10431 5446
rect 10433 5472 10474 5480
rect 10433 5446 10448 5472
rect 10455 5446 10474 5472
rect 10538 5468 10569 5480
rect 10584 5468 10687 5480
rect 10699 5470 10725 5496
rect 10740 5491 10770 5502
rect 10802 5498 10864 5514
rect 10802 5496 10848 5498
rect 10802 5480 10864 5496
rect 10876 5480 10882 5528
rect 10885 5520 10965 5528
rect 10885 5518 10904 5520
rect 10919 5518 10953 5520
rect 10885 5502 10965 5518
rect 10885 5480 10904 5502
rect 10919 5486 10949 5502
rect 10977 5496 10983 5570
rect 10986 5496 11005 5640
rect 11020 5496 11026 5640
rect 11035 5570 11048 5640
rect 11100 5636 11122 5640
rect 11093 5614 11122 5628
rect 11175 5614 11191 5628
rect 11229 5624 11235 5626
rect 11242 5624 11350 5640
rect 11357 5624 11363 5626
rect 11371 5624 11386 5640
rect 11452 5634 11471 5637
rect 11093 5612 11191 5614
rect 11218 5612 11386 5624
rect 11401 5614 11417 5628
rect 11452 5615 11474 5634
rect 11484 5628 11500 5629
rect 11483 5626 11500 5628
rect 11484 5621 11500 5626
rect 11474 5614 11480 5615
rect 11483 5614 11512 5621
rect 11401 5613 11512 5614
rect 11401 5612 11518 5613
rect 11077 5604 11128 5612
rect 11175 5604 11209 5612
rect 11077 5592 11102 5604
rect 11109 5592 11128 5604
rect 11182 5602 11209 5604
rect 11218 5602 11439 5612
rect 11474 5609 11480 5612
rect 11182 5598 11439 5602
rect 11077 5584 11128 5592
rect 11175 5584 11439 5598
rect 11483 5604 11518 5612
rect 11029 5536 11048 5570
rect 11093 5576 11122 5584
rect 11093 5570 11110 5576
rect 11093 5568 11127 5570
rect 11175 5568 11191 5584
rect 11192 5574 11400 5584
rect 11401 5574 11417 5584
rect 11465 5580 11480 5595
rect 11483 5592 11484 5604
rect 11491 5592 11518 5604
rect 11483 5584 11518 5592
rect 11483 5583 11512 5584
rect 11203 5570 11417 5574
rect 11218 5568 11417 5570
rect 11452 5570 11465 5580
rect 11483 5570 11500 5583
rect 11452 5568 11500 5570
rect 11094 5564 11127 5568
rect 11090 5562 11127 5564
rect 11090 5561 11157 5562
rect 11090 5556 11121 5561
rect 11127 5556 11157 5561
rect 11090 5552 11157 5556
rect 11063 5549 11157 5552
rect 11063 5542 11112 5549
rect 11063 5536 11093 5542
rect 11112 5537 11117 5542
rect 11029 5520 11109 5536
rect 11121 5528 11157 5549
rect 11218 5544 11407 5568
rect 11452 5567 11499 5568
rect 11465 5562 11499 5567
rect 11233 5541 11407 5544
rect 11226 5538 11407 5541
rect 11435 5561 11499 5562
rect 11029 5518 11048 5520
rect 11063 5518 11097 5520
rect 11029 5502 11109 5518
rect 11029 5496 11048 5502
rect 10745 5470 10848 5480
rect 10699 5468 10848 5470
rect 10869 5468 10904 5480
rect 10538 5466 10700 5468
rect 10550 5446 10569 5466
rect 10584 5464 10614 5466
rect 10433 5438 10474 5446
rect 10556 5442 10569 5446
rect 10621 5450 10700 5466
rect 10732 5466 10904 5468
rect 10732 5450 10811 5466
rect 10818 5464 10848 5466
rect 10396 5428 10425 5438
rect 10439 5428 10468 5438
rect 10483 5428 10513 5442
rect 10556 5428 10599 5442
rect 10621 5438 10811 5450
rect 10876 5446 10882 5466
rect 10606 5428 10636 5438
rect 10637 5428 10795 5438
rect 10799 5428 10829 5438
rect 10833 5428 10863 5442
rect 10891 5428 10904 5466
rect 10976 5480 11005 5496
rect 11019 5480 11048 5496
rect 11063 5486 11093 5502
rect 11121 5480 11127 5528
rect 11130 5522 11149 5528
rect 11164 5522 11194 5530
rect 11130 5514 11194 5522
rect 11130 5498 11210 5514
rect 11226 5507 11288 5538
rect 11304 5507 11366 5538
rect 11435 5536 11484 5561
rect 11499 5536 11529 5552
rect 11398 5522 11428 5530
rect 11435 5528 11545 5536
rect 11398 5514 11443 5522
rect 11130 5496 11149 5498
rect 11164 5496 11210 5498
rect 11130 5480 11210 5496
rect 11237 5494 11272 5507
rect 11313 5504 11350 5507
rect 11313 5502 11355 5504
rect 11242 5491 11272 5494
rect 11251 5487 11258 5491
rect 11258 5486 11259 5487
rect 11217 5480 11227 5486
rect 10976 5472 11011 5480
rect 10976 5446 10977 5472
rect 10984 5446 11011 5472
rect 10919 5428 10949 5442
rect 10976 5438 11011 5446
rect 11013 5472 11054 5480
rect 11013 5446 11028 5472
rect 11035 5446 11054 5472
rect 11118 5468 11149 5480
rect 11164 5468 11267 5480
rect 11279 5470 11305 5496
rect 11320 5491 11350 5502
rect 11382 5498 11444 5514
rect 11382 5496 11428 5498
rect 11382 5480 11444 5496
rect 11456 5480 11462 5528
rect 11465 5520 11545 5528
rect 11465 5518 11484 5520
rect 11499 5518 11533 5520
rect 11465 5502 11545 5518
rect 11465 5480 11484 5502
rect 11499 5486 11529 5502
rect 11557 5496 11563 5570
rect 11566 5496 11585 5640
rect 11600 5496 11606 5640
rect 11615 5570 11628 5640
rect 11680 5636 11702 5640
rect 11673 5614 11702 5628
rect 11755 5614 11771 5628
rect 11809 5624 11815 5626
rect 11822 5624 11930 5640
rect 11937 5624 11943 5626
rect 11951 5624 11966 5640
rect 12032 5634 12051 5637
rect 11673 5612 11771 5614
rect 11798 5612 11966 5624
rect 11981 5614 11997 5628
rect 12032 5615 12054 5634
rect 12064 5628 12080 5629
rect 12063 5626 12080 5628
rect 12064 5621 12080 5626
rect 12054 5614 12060 5615
rect 12063 5614 12092 5621
rect 11981 5613 12092 5614
rect 11981 5612 12098 5613
rect 11657 5604 11708 5612
rect 11755 5604 11789 5612
rect 11657 5592 11682 5604
rect 11689 5592 11708 5604
rect 11762 5602 11789 5604
rect 11798 5602 12019 5612
rect 12054 5609 12060 5612
rect 11762 5598 12019 5602
rect 11657 5584 11708 5592
rect 11755 5584 12019 5598
rect 12063 5604 12098 5612
rect 11609 5536 11628 5570
rect 11673 5576 11702 5584
rect 11673 5570 11690 5576
rect 11673 5568 11707 5570
rect 11755 5568 11771 5584
rect 11772 5574 11980 5584
rect 11981 5574 11997 5584
rect 12045 5580 12060 5595
rect 12063 5592 12064 5604
rect 12071 5592 12098 5604
rect 12063 5584 12098 5592
rect 12063 5583 12092 5584
rect 11783 5570 11997 5574
rect 11798 5568 11997 5570
rect 12032 5570 12045 5580
rect 12063 5570 12080 5583
rect 12032 5568 12080 5570
rect 11674 5564 11707 5568
rect 11670 5562 11707 5564
rect 11670 5561 11737 5562
rect 11670 5556 11701 5561
rect 11707 5556 11737 5561
rect 11670 5552 11737 5556
rect 11643 5549 11737 5552
rect 11643 5542 11692 5549
rect 11643 5536 11673 5542
rect 11692 5537 11697 5542
rect 11609 5520 11689 5536
rect 11701 5528 11737 5549
rect 11798 5544 11987 5568
rect 12032 5567 12079 5568
rect 12045 5562 12079 5567
rect 11813 5541 11987 5544
rect 11806 5538 11987 5541
rect 12015 5561 12079 5562
rect 11609 5518 11628 5520
rect 11643 5518 11677 5520
rect 11609 5502 11689 5518
rect 11609 5496 11628 5502
rect 11325 5470 11428 5480
rect 11279 5468 11428 5470
rect 11449 5468 11484 5480
rect 11118 5466 11280 5468
rect 11130 5446 11149 5466
rect 11164 5464 11194 5466
rect 11013 5438 11054 5446
rect 11136 5442 11149 5446
rect 11201 5450 11280 5466
rect 11312 5466 11484 5468
rect 11312 5450 11391 5466
rect 11398 5464 11428 5466
rect 10976 5428 11005 5438
rect 11019 5428 11048 5438
rect 11063 5428 11093 5442
rect 11136 5428 11179 5442
rect 11201 5438 11391 5450
rect 11456 5446 11462 5466
rect 11186 5428 11216 5438
rect 11217 5428 11375 5438
rect 11379 5428 11409 5438
rect 11413 5428 11443 5442
rect 11471 5428 11484 5466
rect 11556 5480 11585 5496
rect 11599 5480 11628 5496
rect 11643 5486 11673 5502
rect 11701 5480 11707 5528
rect 11710 5522 11729 5528
rect 11744 5522 11774 5530
rect 11710 5514 11774 5522
rect 11710 5498 11790 5514
rect 11806 5507 11868 5538
rect 11884 5507 11946 5538
rect 12015 5536 12064 5561
rect 12079 5536 12109 5552
rect 11978 5522 12008 5530
rect 12015 5528 12125 5536
rect 11978 5514 12023 5522
rect 11710 5496 11729 5498
rect 11744 5496 11790 5498
rect 11710 5480 11790 5496
rect 11817 5494 11852 5507
rect 11893 5504 11930 5507
rect 11893 5502 11935 5504
rect 11822 5491 11852 5494
rect 11831 5487 11838 5491
rect 11838 5486 11839 5487
rect 11797 5480 11807 5486
rect 11556 5472 11591 5480
rect 11556 5446 11557 5472
rect 11564 5446 11591 5472
rect 11499 5428 11529 5442
rect 11556 5438 11591 5446
rect 11593 5472 11634 5480
rect 11593 5446 11608 5472
rect 11615 5446 11634 5472
rect 11698 5468 11729 5480
rect 11744 5468 11847 5480
rect 11859 5470 11885 5496
rect 11900 5491 11930 5502
rect 11962 5498 12024 5514
rect 11962 5496 12008 5498
rect 11962 5480 12024 5496
rect 12036 5480 12042 5528
rect 12045 5520 12125 5528
rect 12045 5518 12064 5520
rect 12079 5518 12113 5520
rect 12045 5502 12125 5518
rect 12045 5480 12064 5502
rect 12079 5486 12109 5502
rect 12137 5496 12143 5570
rect 12146 5496 12165 5640
rect 12180 5496 12186 5640
rect 12195 5570 12208 5640
rect 12260 5636 12282 5640
rect 12253 5614 12282 5628
rect 12335 5614 12351 5628
rect 12389 5624 12395 5626
rect 12402 5624 12510 5640
rect 12517 5624 12523 5626
rect 12531 5624 12546 5640
rect 12612 5634 12631 5637
rect 12253 5612 12351 5614
rect 12378 5612 12546 5624
rect 12561 5614 12577 5628
rect 12612 5615 12634 5634
rect 12644 5628 12660 5629
rect 12643 5626 12660 5628
rect 12644 5621 12660 5626
rect 12634 5614 12640 5615
rect 12643 5614 12672 5621
rect 12561 5613 12672 5614
rect 12561 5612 12678 5613
rect 12237 5604 12288 5612
rect 12335 5604 12369 5612
rect 12237 5592 12262 5604
rect 12269 5592 12288 5604
rect 12342 5602 12369 5604
rect 12378 5602 12599 5612
rect 12634 5609 12640 5612
rect 12342 5598 12599 5602
rect 12237 5584 12288 5592
rect 12335 5584 12599 5598
rect 12643 5604 12678 5612
rect 12189 5536 12208 5570
rect 12253 5576 12282 5584
rect 12253 5570 12270 5576
rect 12253 5568 12287 5570
rect 12335 5568 12351 5584
rect 12352 5574 12560 5584
rect 12561 5574 12577 5584
rect 12625 5580 12640 5595
rect 12643 5592 12644 5604
rect 12651 5592 12678 5604
rect 12643 5584 12678 5592
rect 12643 5583 12672 5584
rect 12363 5570 12577 5574
rect 12378 5568 12577 5570
rect 12612 5570 12625 5580
rect 12643 5570 12660 5583
rect 12612 5568 12660 5570
rect 12254 5564 12287 5568
rect 12250 5562 12287 5564
rect 12250 5561 12317 5562
rect 12250 5556 12281 5561
rect 12287 5556 12317 5561
rect 12250 5552 12317 5556
rect 12223 5549 12317 5552
rect 12223 5542 12272 5549
rect 12223 5536 12253 5542
rect 12272 5537 12277 5542
rect 12189 5520 12269 5536
rect 12281 5528 12317 5549
rect 12378 5544 12567 5568
rect 12612 5567 12659 5568
rect 12625 5562 12659 5567
rect 12393 5541 12567 5544
rect 12386 5538 12567 5541
rect 12595 5561 12659 5562
rect 12189 5518 12208 5520
rect 12223 5518 12257 5520
rect 12189 5502 12269 5518
rect 12189 5496 12208 5502
rect 11905 5470 12008 5480
rect 11859 5468 12008 5470
rect 12029 5468 12064 5480
rect 11698 5466 11860 5468
rect 11710 5446 11729 5466
rect 11744 5464 11774 5466
rect 11593 5438 11634 5446
rect 11716 5442 11729 5446
rect 11781 5450 11860 5466
rect 11892 5466 12064 5468
rect 11892 5450 11971 5466
rect 11978 5464 12008 5466
rect 11556 5428 11585 5438
rect 11599 5428 11628 5438
rect 11643 5428 11673 5442
rect 11716 5428 11759 5442
rect 11781 5438 11971 5450
rect 12036 5446 12042 5466
rect 11766 5428 11796 5438
rect 11797 5428 11955 5438
rect 11959 5428 11989 5438
rect 11993 5428 12023 5442
rect 12051 5428 12064 5466
rect 12136 5480 12165 5496
rect 12179 5480 12208 5496
rect 12223 5486 12253 5502
rect 12281 5480 12287 5528
rect 12290 5522 12309 5528
rect 12324 5522 12354 5530
rect 12290 5514 12354 5522
rect 12290 5498 12370 5514
rect 12386 5507 12448 5538
rect 12464 5507 12526 5538
rect 12595 5536 12644 5561
rect 12659 5536 12689 5552
rect 12558 5522 12588 5530
rect 12595 5528 12705 5536
rect 12558 5514 12603 5522
rect 12290 5496 12309 5498
rect 12324 5496 12370 5498
rect 12290 5480 12370 5496
rect 12397 5494 12432 5507
rect 12473 5504 12510 5507
rect 12473 5502 12515 5504
rect 12402 5491 12432 5494
rect 12411 5487 12418 5491
rect 12418 5486 12419 5487
rect 12377 5480 12387 5486
rect 12136 5472 12171 5480
rect 12136 5446 12137 5472
rect 12144 5446 12171 5472
rect 12079 5428 12109 5442
rect 12136 5438 12171 5446
rect 12173 5472 12214 5480
rect 12173 5446 12188 5472
rect 12195 5446 12214 5472
rect 12278 5468 12309 5480
rect 12324 5468 12427 5480
rect 12439 5470 12465 5496
rect 12480 5491 12510 5502
rect 12542 5498 12604 5514
rect 12542 5496 12588 5498
rect 12542 5480 12604 5496
rect 12616 5480 12622 5528
rect 12625 5520 12705 5528
rect 12625 5518 12644 5520
rect 12659 5518 12693 5520
rect 12625 5502 12705 5518
rect 12625 5480 12644 5502
rect 12659 5486 12689 5502
rect 12717 5496 12723 5570
rect 12726 5496 12745 5640
rect 12760 5496 12766 5640
rect 12775 5570 12788 5640
rect 12840 5636 12862 5640
rect 12833 5614 12862 5628
rect 12915 5614 12931 5628
rect 12969 5624 12975 5626
rect 12982 5624 13090 5640
rect 13097 5624 13103 5626
rect 13111 5624 13126 5640
rect 13192 5634 13211 5637
rect 12833 5612 12931 5614
rect 12958 5612 13126 5624
rect 13141 5614 13157 5628
rect 13192 5615 13214 5634
rect 13224 5628 13240 5629
rect 13223 5626 13240 5628
rect 13224 5621 13240 5626
rect 13214 5614 13220 5615
rect 13223 5614 13252 5621
rect 13141 5613 13252 5614
rect 13141 5612 13258 5613
rect 12817 5604 12868 5612
rect 12915 5604 12949 5612
rect 12817 5592 12842 5604
rect 12849 5592 12868 5604
rect 12922 5602 12949 5604
rect 12958 5602 13179 5612
rect 13214 5609 13220 5612
rect 12922 5598 13179 5602
rect 12817 5584 12868 5592
rect 12915 5584 13179 5598
rect 13223 5604 13258 5612
rect 12769 5536 12788 5570
rect 12833 5576 12862 5584
rect 12833 5570 12850 5576
rect 12833 5568 12867 5570
rect 12915 5568 12931 5584
rect 12932 5574 13140 5584
rect 13141 5574 13157 5584
rect 13205 5580 13220 5595
rect 13223 5592 13224 5604
rect 13231 5592 13258 5604
rect 13223 5584 13258 5592
rect 13223 5583 13252 5584
rect 12943 5570 13157 5574
rect 12958 5568 13157 5570
rect 13192 5570 13205 5580
rect 13223 5570 13240 5583
rect 13192 5568 13240 5570
rect 12834 5564 12867 5568
rect 12830 5562 12867 5564
rect 12830 5561 12897 5562
rect 12830 5556 12861 5561
rect 12867 5556 12897 5561
rect 12830 5552 12897 5556
rect 12803 5549 12897 5552
rect 12803 5542 12852 5549
rect 12803 5536 12833 5542
rect 12852 5537 12857 5542
rect 12769 5520 12849 5536
rect 12861 5528 12897 5549
rect 12958 5544 13147 5568
rect 13192 5567 13239 5568
rect 13205 5562 13239 5567
rect 12973 5541 13147 5544
rect 12966 5538 13147 5541
rect 13175 5561 13239 5562
rect 12769 5518 12788 5520
rect 12803 5518 12837 5520
rect 12769 5502 12849 5518
rect 12769 5496 12788 5502
rect 12485 5470 12588 5480
rect 12439 5468 12588 5470
rect 12609 5468 12644 5480
rect 12278 5466 12440 5468
rect 12290 5446 12309 5466
rect 12324 5464 12354 5466
rect 12173 5438 12214 5446
rect 12296 5442 12309 5446
rect 12361 5450 12440 5466
rect 12472 5466 12644 5468
rect 12472 5450 12551 5466
rect 12558 5464 12588 5466
rect 12136 5428 12165 5438
rect 12179 5428 12208 5438
rect 12223 5428 12253 5442
rect 12296 5428 12339 5442
rect 12361 5438 12551 5450
rect 12616 5446 12622 5466
rect 12346 5428 12376 5438
rect 12377 5428 12535 5438
rect 12539 5428 12569 5438
rect 12573 5428 12603 5442
rect 12631 5428 12644 5466
rect 12716 5480 12745 5496
rect 12759 5480 12788 5496
rect 12803 5486 12833 5502
rect 12861 5480 12867 5528
rect 12870 5522 12889 5528
rect 12904 5522 12934 5530
rect 12870 5514 12934 5522
rect 12870 5498 12950 5514
rect 12966 5507 13028 5538
rect 13044 5507 13106 5538
rect 13175 5536 13224 5561
rect 13239 5536 13269 5552
rect 13138 5522 13168 5530
rect 13175 5528 13285 5536
rect 13138 5514 13183 5522
rect 12870 5496 12889 5498
rect 12904 5496 12950 5498
rect 12870 5480 12950 5496
rect 12977 5494 13012 5507
rect 13053 5504 13090 5507
rect 13053 5502 13095 5504
rect 12982 5491 13012 5494
rect 12991 5487 12998 5491
rect 12998 5486 12999 5487
rect 12957 5480 12967 5486
rect 12716 5472 12751 5480
rect 12716 5446 12717 5472
rect 12724 5446 12751 5472
rect 12659 5428 12689 5442
rect 12716 5438 12751 5446
rect 12753 5472 12794 5480
rect 12753 5446 12768 5472
rect 12775 5446 12794 5472
rect 12858 5468 12889 5480
rect 12904 5468 13007 5480
rect 13019 5470 13045 5496
rect 13060 5491 13090 5502
rect 13122 5498 13184 5514
rect 13122 5496 13168 5498
rect 13122 5480 13184 5496
rect 13196 5480 13202 5528
rect 13205 5520 13285 5528
rect 13205 5518 13224 5520
rect 13239 5518 13273 5520
rect 13205 5502 13285 5518
rect 13205 5480 13224 5502
rect 13239 5486 13269 5502
rect 13297 5496 13303 5570
rect 13306 5496 13325 5640
rect 13340 5496 13346 5640
rect 13355 5570 13368 5640
rect 13420 5636 13442 5640
rect 13413 5614 13442 5628
rect 13495 5614 13511 5628
rect 13549 5624 13555 5626
rect 13562 5624 13670 5640
rect 13677 5624 13683 5626
rect 13691 5624 13706 5640
rect 13772 5634 13791 5637
rect 13413 5612 13511 5614
rect 13538 5612 13706 5624
rect 13721 5614 13737 5628
rect 13772 5615 13794 5634
rect 13804 5628 13820 5629
rect 13803 5626 13820 5628
rect 13804 5621 13820 5626
rect 13794 5614 13800 5615
rect 13803 5614 13832 5621
rect 13721 5613 13832 5614
rect 13721 5612 13838 5613
rect 13397 5604 13448 5612
rect 13495 5604 13529 5612
rect 13397 5592 13422 5604
rect 13429 5592 13448 5604
rect 13502 5602 13529 5604
rect 13538 5602 13759 5612
rect 13794 5609 13800 5612
rect 13502 5598 13759 5602
rect 13397 5584 13448 5592
rect 13495 5584 13759 5598
rect 13803 5604 13838 5612
rect 13349 5536 13368 5570
rect 13413 5576 13442 5584
rect 13413 5570 13430 5576
rect 13413 5568 13447 5570
rect 13495 5568 13511 5584
rect 13512 5574 13720 5584
rect 13721 5574 13737 5584
rect 13785 5580 13800 5595
rect 13803 5592 13804 5604
rect 13811 5592 13838 5604
rect 13803 5584 13838 5592
rect 13803 5583 13832 5584
rect 13523 5570 13737 5574
rect 13538 5568 13737 5570
rect 13772 5570 13785 5580
rect 13803 5570 13820 5583
rect 13772 5568 13820 5570
rect 13414 5564 13447 5568
rect 13410 5562 13447 5564
rect 13410 5561 13477 5562
rect 13410 5556 13441 5561
rect 13447 5556 13477 5561
rect 13410 5552 13477 5556
rect 13383 5549 13477 5552
rect 13383 5542 13432 5549
rect 13383 5536 13413 5542
rect 13432 5537 13437 5542
rect 13349 5520 13429 5536
rect 13441 5528 13477 5549
rect 13538 5544 13727 5568
rect 13772 5567 13819 5568
rect 13785 5562 13819 5567
rect 13553 5541 13727 5544
rect 13546 5538 13727 5541
rect 13755 5561 13819 5562
rect 13349 5518 13368 5520
rect 13383 5518 13417 5520
rect 13349 5502 13429 5518
rect 13349 5496 13368 5502
rect 13065 5470 13168 5480
rect 13019 5468 13168 5470
rect 13189 5468 13224 5480
rect 12858 5466 13020 5468
rect 12870 5446 12889 5466
rect 12904 5464 12934 5466
rect 12753 5438 12794 5446
rect 12876 5442 12889 5446
rect 12941 5450 13020 5466
rect 13052 5466 13224 5468
rect 13052 5450 13131 5466
rect 13138 5464 13168 5466
rect 12716 5428 12745 5438
rect 12759 5428 12788 5438
rect 12803 5428 12833 5442
rect 12876 5428 12919 5442
rect 12941 5438 13131 5450
rect 13196 5446 13202 5466
rect 12926 5428 12956 5438
rect 12957 5428 13115 5438
rect 13119 5428 13149 5438
rect 13153 5428 13183 5442
rect 13211 5428 13224 5466
rect 13296 5480 13325 5496
rect 13339 5480 13368 5496
rect 13383 5486 13413 5502
rect 13441 5480 13447 5528
rect 13450 5522 13469 5528
rect 13484 5522 13514 5530
rect 13450 5514 13514 5522
rect 13450 5498 13530 5514
rect 13546 5507 13608 5538
rect 13624 5507 13686 5538
rect 13755 5536 13804 5561
rect 13819 5536 13849 5552
rect 13718 5522 13748 5530
rect 13755 5528 13865 5536
rect 13718 5514 13763 5522
rect 13450 5496 13469 5498
rect 13484 5496 13530 5498
rect 13450 5480 13530 5496
rect 13557 5494 13592 5507
rect 13633 5504 13670 5507
rect 13633 5502 13675 5504
rect 13562 5491 13592 5494
rect 13571 5487 13578 5491
rect 13578 5486 13579 5487
rect 13537 5480 13547 5486
rect 13296 5472 13331 5480
rect 13296 5446 13297 5472
rect 13304 5446 13331 5472
rect 13239 5428 13269 5442
rect 13296 5438 13331 5446
rect 13333 5472 13374 5480
rect 13333 5446 13348 5472
rect 13355 5446 13374 5472
rect 13438 5468 13469 5480
rect 13484 5468 13587 5480
rect 13599 5470 13625 5496
rect 13640 5491 13670 5502
rect 13702 5498 13764 5514
rect 13702 5496 13748 5498
rect 13702 5480 13764 5496
rect 13776 5480 13782 5528
rect 13785 5520 13865 5528
rect 13785 5518 13804 5520
rect 13819 5518 13853 5520
rect 13785 5502 13865 5518
rect 13785 5480 13804 5502
rect 13819 5486 13849 5502
rect 13877 5496 13883 5570
rect 13886 5496 13905 5640
rect 13920 5496 13926 5640
rect 13935 5570 13948 5640
rect 14000 5636 14022 5640
rect 13993 5614 14022 5628
rect 14075 5614 14091 5628
rect 14129 5624 14135 5626
rect 14142 5624 14250 5640
rect 14257 5624 14263 5626
rect 14271 5624 14286 5640
rect 14352 5634 14371 5637
rect 13993 5612 14091 5614
rect 14118 5612 14286 5624
rect 14301 5614 14317 5628
rect 14352 5615 14374 5634
rect 14384 5628 14400 5629
rect 14383 5626 14400 5628
rect 14384 5621 14400 5626
rect 14374 5614 14380 5615
rect 14383 5614 14412 5621
rect 14301 5613 14412 5614
rect 14301 5612 14418 5613
rect 13977 5604 14028 5612
rect 14075 5604 14109 5612
rect 13977 5592 14002 5604
rect 14009 5592 14028 5604
rect 14082 5602 14109 5604
rect 14118 5602 14339 5612
rect 14374 5609 14380 5612
rect 14082 5598 14339 5602
rect 13977 5584 14028 5592
rect 14075 5584 14339 5598
rect 14383 5604 14418 5612
rect 13929 5536 13948 5570
rect 13993 5576 14022 5584
rect 13993 5570 14010 5576
rect 13993 5568 14027 5570
rect 14075 5568 14091 5584
rect 14092 5574 14300 5584
rect 14301 5574 14317 5584
rect 14365 5580 14380 5595
rect 14383 5592 14384 5604
rect 14391 5592 14418 5604
rect 14383 5584 14418 5592
rect 14383 5583 14412 5584
rect 14103 5570 14317 5574
rect 14118 5568 14317 5570
rect 14352 5570 14365 5580
rect 14383 5570 14400 5583
rect 14352 5568 14400 5570
rect 13994 5564 14027 5568
rect 13990 5562 14027 5564
rect 13990 5561 14057 5562
rect 13990 5556 14021 5561
rect 14027 5556 14057 5561
rect 13990 5552 14057 5556
rect 13963 5549 14057 5552
rect 13963 5542 14012 5549
rect 13963 5536 13993 5542
rect 14012 5537 14017 5542
rect 13929 5520 14009 5536
rect 14021 5528 14057 5549
rect 14118 5544 14307 5568
rect 14352 5567 14399 5568
rect 14365 5562 14399 5567
rect 14133 5541 14307 5544
rect 14126 5538 14307 5541
rect 14335 5561 14399 5562
rect 13929 5518 13948 5520
rect 13963 5518 13997 5520
rect 13929 5502 14009 5518
rect 13929 5496 13948 5502
rect 13645 5470 13748 5480
rect 13599 5468 13748 5470
rect 13769 5468 13804 5480
rect 13438 5466 13600 5468
rect 13450 5446 13469 5466
rect 13484 5464 13514 5466
rect 13333 5438 13374 5446
rect 13456 5442 13469 5446
rect 13521 5450 13600 5466
rect 13632 5466 13804 5468
rect 13632 5450 13711 5466
rect 13718 5464 13748 5466
rect 13296 5428 13325 5438
rect 13339 5428 13368 5438
rect 13383 5428 13413 5442
rect 13456 5428 13499 5442
rect 13521 5438 13711 5450
rect 13776 5446 13782 5466
rect 13506 5428 13536 5438
rect 13537 5428 13695 5438
rect 13699 5428 13729 5438
rect 13733 5428 13763 5442
rect 13791 5428 13804 5466
rect 13876 5480 13905 5496
rect 13919 5480 13948 5496
rect 13963 5486 13993 5502
rect 14021 5480 14027 5528
rect 14030 5522 14049 5528
rect 14064 5522 14094 5530
rect 14030 5514 14094 5522
rect 14030 5498 14110 5514
rect 14126 5507 14188 5538
rect 14204 5507 14266 5538
rect 14335 5536 14384 5561
rect 14399 5536 14429 5552
rect 14298 5522 14328 5530
rect 14335 5528 14445 5536
rect 14298 5514 14343 5522
rect 14030 5496 14049 5498
rect 14064 5496 14110 5498
rect 14030 5480 14110 5496
rect 14137 5494 14172 5507
rect 14213 5504 14250 5507
rect 14213 5502 14255 5504
rect 14142 5491 14172 5494
rect 14151 5487 14158 5491
rect 14158 5486 14159 5487
rect 14117 5480 14127 5486
rect 13876 5472 13911 5480
rect 13876 5446 13877 5472
rect 13884 5446 13911 5472
rect 13819 5428 13849 5442
rect 13876 5438 13911 5446
rect 13913 5472 13954 5480
rect 13913 5446 13928 5472
rect 13935 5446 13954 5472
rect 14018 5468 14049 5480
rect 14064 5468 14167 5480
rect 14179 5470 14205 5496
rect 14220 5491 14250 5502
rect 14282 5498 14344 5514
rect 14282 5496 14328 5498
rect 14282 5480 14344 5496
rect 14356 5480 14362 5528
rect 14365 5520 14445 5528
rect 14365 5518 14384 5520
rect 14399 5518 14433 5520
rect 14365 5502 14445 5518
rect 14365 5480 14384 5502
rect 14399 5486 14429 5502
rect 14457 5496 14463 5570
rect 14466 5496 14485 5640
rect 14500 5496 14506 5640
rect 14515 5570 14528 5640
rect 14580 5636 14602 5640
rect 14573 5614 14602 5628
rect 14655 5614 14671 5628
rect 14709 5624 14715 5626
rect 14722 5624 14830 5640
rect 14837 5624 14843 5626
rect 14851 5624 14866 5640
rect 14932 5634 14951 5637
rect 14573 5612 14671 5614
rect 14698 5612 14866 5624
rect 14881 5614 14897 5628
rect 14932 5615 14954 5634
rect 14964 5628 14980 5629
rect 14963 5626 14980 5628
rect 14964 5621 14980 5626
rect 14954 5614 14960 5615
rect 14963 5614 14992 5621
rect 14881 5613 14992 5614
rect 14881 5612 14998 5613
rect 14557 5604 14608 5612
rect 14655 5604 14689 5612
rect 14557 5592 14582 5604
rect 14589 5592 14608 5604
rect 14662 5602 14689 5604
rect 14698 5602 14919 5612
rect 14954 5609 14960 5612
rect 14662 5598 14919 5602
rect 14557 5584 14608 5592
rect 14655 5584 14919 5598
rect 14963 5604 14998 5612
rect 14509 5536 14528 5570
rect 14573 5576 14602 5584
rect 14573 5570 14590 5576
rect 14573 5568 14607 5570
rect 14655 5568 14671 5584
rect 14672 5574 14880 5584
rect 14881 5574 14897 5584
rect 14945 5580 14960 5595
rect 14963 5592 14964 5604
rect 14971 5592 14998 5604
rect 14963 5584 14998 5592
rect 14963 5583 14992 5584
rect 14683 5570 14897 5574
rect 14698 5568 14897 5570
rect 14932 5570 14945 5580
rect 14963 5570 14980 5583
rect 14932 5568 14980 5570
rect 14574 5564 14607 5568
rect 14570 5562 14607 5564
rect 14570 5561 14637 5562
rect 14570 5556 14601 5561
rect 14607 5556 14637 5561
rect 14570 5552 14637 5556
rect 14543 5549 14637 5552
rect 14543 5542 14592 5549
rect 14543 5536 14573 5542
rect 14592 5537 14597 5542
rect 14509 5520 14589 5536
rect 14601 5528 14637 5549
rect 14698 5544 14887 5568
rect 14932 5567 14979 5568
rect 14945 5562 14979 5567
rect 14713 5541 14887 5544
rect 14706 5538 14887 5541
rect 14915 5561 14979 5562
rect 14509 5518 14528 5520
rect 14543 5518 14577 5520
rect 14509 5502 14589 5518
rect 14509 5496 14528 5502
rect 14225 5470 14328 5480
rect 14179 5468 14328 5470
rect 14349 5468 14384 5480
rect 14018 5466 14180 5468
rect 14030 5446 14049 5466
rect 14064 5464 14094 5466
rect 13913 5438 13954 5446
rect 14036 5442 14049 5446
rect 14101 5450 14180 5466
rect 14212 5466 14384 5468
rect 14212 5450 14291 5466
rect 14298 5464 14328 5466
rect 13876 5428 13905 5438
rect 13919 5428 13948 5438
rect 13963 5428 13993 5442
rect 14036 5428 14079 5442
rect 14101 5438 14291 5450
rect 14356 5446 14362 5466
rect 14086 5428 14116 5438
rect 14117 5428 14275 5438
rect 14279 5428 14309 5438
rect 14313 5428 14343 5442
rect 14371 5428 14384 5466
rect 14456 5480 14485 5496
rect 14499 5480 14528 5496
rect 14543 5486 14573 5502
rect 14601 5480 14607 5528
rect 14610 5522 14629 5528
rect 14644 5522 14674 5530
rect 14610 5514 14674 5522
rect 14610 5498 14690 5514
rect 14706 5507 14768 5538
rect 14784 5507 14846 5538
rect 14915 5536 14964 5561
rect 14979 5536 15009 5552
rect 14878 5522 14908 5530
rect 14915 5528 15025 5536
rect 14878 5514 14923 5522
rect 14610 5496 14629 5498
rect 14644 5496 14690 5498
rect 14610 5480 14690 5496
rect 14717 5494 14752 5507
rect 14793 5504 14830 5507
rect 14793 5502 14835 5504
rect 14722 5491 14752 5494
rect 14731 5487 14738 5491
rect 14738 5486 14739 5487
rect 14697 5480 14707 5486
rect 14456 5472 14491 5480
rect 14456 5446 14457 5472
rect 14464 5446 14491 5472
rect 14399 5428 14429 5442
rect 14456 5438 14491 5446
rect 14493 5472 14534 5480
rect 14493 5446 14508 5472
rect 14515 5446 14534 5472
rect 14598 5468 14629 5480
rect 14644 5468 14747 5480
rect 14759 5470 14785 5496
rect 14800 5491 14830 5502
rect 14862 5498 14924 5514
rect 14862 5496 14908 5498
rect 14862 5480 14924 5496
rect 14936 5480 14942 5528
rect 14945 5520 15025 5528
rect 14945 5518 14964 5520
rect 14979 5518 15013 5520
rect 14945 5502 15025 5518
rect 14945 5480 14964 5502
rect 14979 5486 15009 5502
rect 15037 5496 15043 5570
rect 15046 5496 15065 5640
rect 15080 5496 15086 5640
rect 15095 5570 15108 5640
rect 15160 5636 15182 5640
rect 15153 5614 15182 5628
rect 15235 5614 15251 5628
rect 15289 5624 15295 5626
rect 15302 5624 15410 5640
rect 15417 5624 15423 5626
rect 15431 5624 15446 5640
rect 15512 5634 15531 5637
rect 15153 5612 15251 5614
rect 15278 5612 15446 5624
rect 15461 5614 15477 5628
rect 15512 5615 15534 5634
rect 15544 5628 15560 5629
rect 15543 5626 15560 5628
rect 15544 5621 15560 5626
rect 15534 5614 15540 5615
rect 15543 5614 15572 5621
rect 15461 5613 15572 5614
rect 15461 5612 15578 5613
rect 15137 5604 15188 5612
rect 15235 5604 15269 5612
rect 15137 5592 15162 5604
rect 15169 5592 15188 5604
rect 15242 5602 15269 5604
rect 15278 5602 15499 5612
rect 15534 5609 15540 5612
rect 15242 5598 15499 5602
rect 15137 5584 15188 5592
rect 15235 5584 15499 5598
rect 15543 5604 15578 5612
rect 15089 5536 15108 5570
rect 15153 5576 15182 5584
rect 15153 5570 15170 5576
rect 15153 5568 15187 5570
rect 15235 5568 15251 5584
rect 15252 5574 15460 5584
rect 15461 5574 15477 5584
rect 15525 5580 15540 5595
rect 15543 5592 15544 5604
rect 15551 5592 15578 5604
rect 15543 5584 15578 5592
rect 15543 5583 15572 5584
rect 15263 5570 15477 5574
rect 15278 5568 15477 5570
rect 15512 5570 15525 5580
rect 15543 5570 15560 5583
rect 15512 5568 15560 5570
rect 15154 5564 15187 5568
rect 15150 5562 15187 5564
rect 15150 5561 15217 5562
rect 15150 5556 15181 5561
rect 15187 5556 15217 5561
rect 15150 5552 15217 5556
rect 15123 5549 15217 5552
rect 15123 5542 15172 5549
rect 15123 5536 15153 5542
rect 15172 5537 15177 5542
rect 15089 5520 15169 5536
rect 15181 5528 15217 5549
rect 15278 5544 15467 5568
rect 15512 5567 15559 5568
rect 15525 5562 15559 5567
rect 15293 5541 15467 5544
rect 15286 5538 15467 5541
rect 15495 5561 15559 5562
rect 15089 5518 15108 5520
rect 15123 5518 15157 5520
rect 15089 5502 15169 5518
rect 15089 5496 15108 5502
rect 14805 5470 14908 5480
rect 14759 5468 14908 5470
rect 14929 5468 14964 5480
rect 14598 5466 14760 5468
rect 14610 5446 14629 5466
rect 14644 5464 14674 5466
rect 14493 5438 14534 5446
rect 14616 5442 14629 5446
rect 14681 5450 14760 5466
rect 14792 5466 14964 5468
rect 14792 5450 14871 5466
rect 14878 5464 14908 5466
rect 14456 5428 14485 5438
rect 14499 5428 14528 5438
rect 14543 5428 14573 5442
rect 14616 5428 14659 5442
rect 14681 5438 14871 5450
rect 14936 5446 14942 5466
rect 14666 5428 14696 5438
rect 14697 5428 14855 5438
rect 14859 5428 14889 5438
rect 14893 5428 14923 5442
rect 14951 5428 14964 5466
rect 15036 5480 15065 5496
rect 15079 5480 15108 5496
rect 15123 5486 15153 5502
rect 15181 5480 15187 5528
rect 15190 5522 15209 5528
rect 15224 5522 15254 5530
rect 15190 5514 15254 5522
rect 15190 5498 15270 5514
rect 15286 5507 15348 5538
rect 15364 5507 15426 5538
rect 15495 5536 15544 5561
rect 15559 5536 15589 5552
rect 15458 5522 15488 5530
rect 15495 5528 15605 5536
rect 15458 5514 15503 5522
rect 15190 5496 15209 5498
rect 15224 5496 15270 5498
rect 15190 5480 15270 5496
rect 15297 5494 15332 5507
rect 15373 5504 15410 5507
rect 15373 5502 15415 5504
rect 15302 5491 15332 5494
rect 15311 5487 15318 5491
rect 15318 5486 15319 5487
rect 15277 5480 15287 5486
rect 15036 5472 15071 5480
rect 15036 5446 15037 5472
rect 15044 5446 15071 5472
rect 14979 5428 15009 5442
rect 15036 5438 15071 5446
rect 15073 5472 15114 5480
rect 15073 5446 15088 5472
rect 15095 5446 15114 5472
rect 15178 5468 15209 5480
rect 15224 5468 15327 5480
rect 15339 5470 15365 5496
rect 15380 5491 15410 5502
rect 15442 5498 15504 5514
rect 15442 5496 15488 5498
rect 15442 5480 15504 5496
rect 15516 5480 15522 5528
rect 15525 5520 15605 5528
rect 15525 5518 15544 5520
rect 15559 5518 15593 5520
rect 15525 5502 15605 5518
rect 15525 5480 15544 5502
rect 15559 5486 15589 5502
rect 15617 5496 15623 5570
rect 15626 5496 15645 5640
rect 15660 5496 15666 5640
rect 15675 5570 15688 5640
rect 15740 5636 15762 5640
rect 15733 5614 15762 5628
rect 15815 5614 15831 5628
rect 15869 5624 15875 5626
rect 15882 5624 15990 5640
rect 15997 5624 16003 5626
rect 16011 5624 16026 5640
rect 16092 5634 16111 5637
rect 15733 5612 15831 5614
rect 15858 5612 16026 5624
rect 16041 5614 16057 5628
rect 16092 5615 16114 5634
rect 16124 5628 16140 5629
rect 16123 5626 16140 5628
rect 16124 5621 16140 5626
rect 16114 5614 16120 5615
rect 16123 5614 16152 5621
rect 16041 5613 16152 5614
rect 16041 5612 16158 5613
rect 15717 5604 15768 5612
rect 15815 5604 15849 5612
rect 15717 5592 15742 5604
rect 15749 5592 15768 5604
rect 15822 5602 15849 5604
rect 15858 5602 16079 5612
rect 16114 5609 16120 5612
rect 15822 5598 16079 5602
rect 15717 5584 15768 5592
rect 15815 5584 16079 5598
rect 16123 5604 16158 5612
rect 15669 5536 15688 5570
rect 15733 5576 15762 5584
rect 15733 5570 15750 5576
rect 15733 5568 15767 5570
rect 15815 5568 15831 5584
rect 15832 5574 16040 5584
rect 16041 5574 16057 5584
rect 16105 5580 16120 5595
rect 16123 5592 16124 5604
rect 16131 5592 16158 5604
rect 16123 5584 16158 5592
rect 16123 5583 16152 5584
rect 15843 5570 16057 5574
rect 15858 5568 16057 5570
rect 16092 5570 16105 5580
rect 16123 5570 16140 5583
rect 16092 5568 16140 5570
rect 15734 5564 15767 5568
rect 15730 5562 15767 5564
rect 15730 5561 15797 5562
rect 15730 5556 15761 5561
rect 15767 5556 15797 5561
rect 15730 5552 15797 5556
rect 15703 5549 15797 5552
rect 15703 5542 15752 5549
rect 15703 5536 15733 5542
rect 15752 5537 15757 5542
rect 15669 5520 15749 5536
rect 15761 5528 15797 5549
rect 15858 5544 16047 5568
rect 16092 5567 16139 5568
rect 16105 5562 16139 5567
rect 15873 5541 16047 5544
rect 15866 5538 16047 5541
rect 16075 5561 16139 5562
rect 15669 5518 15688 5520
rect 15703 5518 15737 5520
rect 15669 5502 15749 5518
rect 15669 5496 15688 5502
rect 15385 5470 15488 5480
rect 15339 5468 15488 5470
rect 15509 5468 15544 5480
rect 15178 5466 15340 5468
rect 15190 5446 15209 5466
rect 15224 5464 15254 5466
rect 15073 5438 15114 5446
rect 15196 5442 15209 5446
rect 15261 5450 15340 5466
rect 15372 5466 15544 5468
rect 15372 5450 15451 5466
rect 15458 5464 15488 5466
rect 15036 5428 15065 5438
rect 15079 5428 15108 5438
rect 15123 5428 15153 5442
rect 15196 5428 15239 5442
rect 15261 5438 15451 5450
rect 15516 5446 15522 5466
rect 15246 5428 15276 5438
rect 15277 5428 15435 5438
rect 15439 5428 15469 5438
rect 15473 5428 15503 5442
rect 15531 5428 15544 5466
rect 15616 5480 15645 5496
rect 15659 5480 15688 5496
rect 15703 5486 15733 5502
rect 15761 5480 15767 5528
rect 15770 5522 15789 5528
rect 15804 5522 15834 5530
rect 15770 5514 15834 5522
rect 15770 5498 15850 5514
rect 15866 5507 15928 5538
rect 15944 5507 16006 5538
rect 16075 5536 16124 5561
rect 16139 5536 16169 5552
rect 16038 5522 16068 5530
rect 16075 5528 16185 5536
rect 16038 5514 16083 5522
rect 15770 5496 15789 5498
rect 15804 5496 15850 5498
rect 15770 5480 15850 5496
rect 15877 5494 15912 5507
rect 15953 5504 15990 5507
rect 15953 5502 15995 5504
rect 15882 5491 15912 5494
rect 15891 5487 15898 5491
rect 15898 5486 15899 5487
rect 15857 5480 15867 5486
rect 15616 5472 15651 5480
rect 15616 5446 15617 5472
rect 15624 5446 15651 5472
rect 15559 5428 15589 5442
rect 15616 5438 15651 5446
rect 15653 5472 15694 5480
rect 15653 5446 15668 5472
rect 15675 5446 15694 5472
rect 15758 5468 15789 5480
rect 15804 5468 15907 5480
rect 15919 5470 15945 5496
rect 15960 5491 15990 5502
rect 16022 5498 16084 5514
rect 16022 5496 16068 5498
rect 16022 5480 16084 5496
rect 16096 5480 16102 5528
rect 16105 5520 16185 5528
rect 16105 5518 16124 5520
rect 16139 5518 16173 5520
rect 16105 5502 16185 5518
rect 16105 5480 16124 5502
rect 16139 5486 16169 5502
rect 16197 5496 16203 5570
rect 16206 5496 16225 5640
rect 16240 5496 16246 5640
rect 16255 5570 16268 5640
rect 16320 5636 16342 5640
rect 16313 5614 16342 5628
rect 16395 5614 16411 5628
rect 16449 5624 16455 5626
rect 16462 5624 16570 5640
rect 16577 5624 16583 5626
rect 16591 5624 16606 5640
rect 16672 5634 16691 5637
rect 16313 5612 16411 5614
rect 16438 5612 16606 5624
rect 16621 5614 16637 5628
rect 16672 5615 16694 5634
rect 16704 5628 16720 5629
rect 16703 5626 16720 5628
rect 16704 5621 16720 5626
rect 16694 5614 16700 5615
rect 16703 5614 16732 5621
rect 16621 5613 16732 5614
rect 16621 5612 16738 5613
rect 16297 5604 16348 5612
rect 16395 5604 16429 5612
rect 16297 5592 16322 5604
rect 16329 5592 16348 5604
rect 16402 5602 16429 5604
rect 16438 5602 16659 5612
rect 16694 5609 16700 5612
rect 16402 5598 16659 5602
rect 16297 5584 16348 5592
rect 16395 5584 16659 5598
rect 16703 5604 16738 5612
rect 16249 5536 16268 5570
rect 16313 5576 16342 5584
rect 16313 5570 16330 5576
rect 16313 5568 16347 5570
rect 16395 5568 16411 5584
rect 16412 5574 16620 5584
rect 16621 5574 16637 5584
rect 16685 5580 16700 5595
rect 16703 5592 16704 5604
rect 16711 5592 16738 5604
rect 16703 5584 16738 5592
rect 16703 5583 16732 5584
rect 16423 5570 16637 5574
rect 16438 5568 16637 5570
rect 16672 5570 16685 5580
rect 16703 5570 16720 5583
rect 16672 5568 16720 5570
rect 16314 5564 16347 5568
rect 16310 5562 16347 5564
rect 16310 5561 16377 5562
rect 16310 5556 16341 5561
rect 16347 5556 16377 5561
rect 16310 5552 16377 5556
rect 16283 5549 16377 5552
rect 16283 5542 16332 5549
rect 16283 5536 16313 5542
rect 16332 5537 16337 5542
rect 16249 5520 16329 5536
rect 16341 5528 16377 5549
rect 16438 5544 16627 5568
rect 16672 5567 16719 5568
rect 16685 5562 16719 5567
rect 16453 5541 16627 5544
rect 16446 5538 16627 5541
rect 16655 5561 16719 5562
rect 16249 5518 16268 5520
rect 16283 5518 16317 5520
rect 16249 5502 16329 5518
rect 16249 5496 16268 5502
rect 15965 5470 16068 5480
rect 15919 5468 16068 5470
rect 16089 5468 16124 5480
rect 15758 5466 15920 5468
rect 15770 5446 15789 5466
rect 15804 5464 15834 5466
rect 15653 5438 15694 5446
rect 15776 5442 15789 5446
rect 15841 5450 15920 5466
rect 15952 5466 16124 5468
rect 15952 5450 16031 5466
rect 16038 5464 16068 5466
rect 15616 5428 15645 5438
rect 15659 5428 15688 5438
rect 15703 5428 15733 5442
rect 15776 5428 15819 5442
rect 15841 5438 16031 5450
rect 16096 5446 16102 5466
rect 15826 5428 15856 5438
rect 15857 5428 16015 5438
rect 16019 5428 16049 5438
rect 16053 5428 16083 5442
rect 16111 5428 16124 5466
rect 16196 5480 16225 5496
rect 16239 5480 16268 5496
rect 16283 5486 16313 5502
rect 16341 5480 16347 5528
rect 16350 5522 16369 5528
rect 16384 5522 16414 5530
rect 16350 5514 16414 5522
rect 16350 5498 16430 5514
rect 16446 5507 16508 5538
rect 16524 5507 16586 5538
rect 16655 5536 16704 5561
rect 16719 5536 16749 5552
rect 16618 5522 16648 5530
rect 16655 5528 16765 5536
rect 16618 5514 16663 5522
rect 16350 5496 16369 5498
rect 16384 5496 16430 5498
rect 16350 5480 16430 5496
rect 16457 5494 16492 5507
rect 16533 5504 16570 5507
rect 16533 5502 16575 5504
rect 16462 5491 16492 5494
rect 16471 5487 16478 5491
rect 16478 5486 16479 5487
rect 16437 5480 16447 5486
rect 16196 5472 16231 5480
rect 16196 5446 16197 5472
rect 16204 5446 16231 5472
rect 16139 5428 16169 5442
rect 16196 5438 16231 5446
rect 16233 5472 16274 5480
rect 16233 5446 16248 5472
rect 16255 5446 16274 5472
rect 16338 5468 16369 5480
rect 16384 5468 16487 5480
rect 16499 5470 16525 5496
rect 16540 5491 16570 5502
rect 16602 5498 16664 5514
rect 16602 5496 16648 5498
rect 16602 5480 16664 5496
rect 16676 5480 16682 5528
rect 16685 5520 16765 5528
rect 16685 5518 16704 5520
rect 16719 5518 16753 5520
rect 16685 5502 16765 5518
rect 16685 5480 16704 5502
rect 16719 5486 16749 5502
rect 16777 5496 16783 5570
rect 16786 5496 16805 5640
rect 16820 5496 16826 5640
rect 16835 5570 16848 5640
rect 16900 5636 16922 5640
rect 16893 5614 16922 5628
rect 16975 5614 16991 5628
rect 17029 5624 17035 5626
rect 17042 5624 17150 5640
rect 17157 5624 17163 5626
rect 17171 5624 17186 5640
rect 17252 5634 17271 5637
rect 16893 5612 16991 5614
rect 17018 5612 17186 5624
rect 17201 5614 17217 5628
rect 17252 5615 17274 5634
rect 17284 5628 17300 5629
rect 17283 5626 17300 5628
rect 17284 5621 17300 5626
rect 17274 5614 17280 5615
rect 17283 5614 17312 5621
rect 17201 5613 17312 5614
rect 17201 5612 17318 5613
rect 16877 5604 16928 5612
rect 16975 5604 17009 5612
rect 16877 5592 16902 5604
rect 16909 5592 16928 5604
rect 16982 5602 17009 5604
rect 17018 5602 17239 5612
rect 17274 5609 17280 5612
rect 16982 5598 17239 5602
rect 16877 5584 16928 5592
rect 16975 5584 17239 5598
rect 17283 5604 17318 5612
rect 16829 5536 16848 5570
rect 16893 5576 16922 5584
rect 16893 5570 16910 5576
rect 16893 5568 16927 5570
rect 16975 5568 16991 5584
rect 16992 5574 17200 5584
rect 17201 5574 17217 5584
rect 17265 5580 17280 5595
rect 17283 5592 17284 5604
rect 17291 5592 17318 5604
rect 17283 5584 17318 5592
rect 17283 5583 17312 5584
rect 17003 5570 17217 5574
rect 17018 5568 17217 5570
rect 17252 5570 17265 5580
rect 17283 5570 17300 5583
rect 17252 5568 17300 5570
rect 16894 5564 16927 5568
rect 16890 5562 16927 5564
rect 16890 5561 16957 5562
rect 16890 5556 16921 5561
rect 16927 5556 16957 5561
rect 16890 5552 16957 5556
rect 16863 5549 16957 5552
rect 16863 5542 16912 5549
rect 16863 5536 16893 5542
rect 16912 5537 16917 5542
rect 16829 5520 16909 5536
rect 16921 5528 16957 5549
rect 17018 5544 17207 5568
rect 17252 5567 17299 5568
rect 17265 5562 17299 5567
rect 17033 5541 17207 5544
rect 17026 5538 17207 5541
rect 17235 5561 17299 5562
rect 16829 5518 16848 5520
rect 16863 5518 16897 5520
rect 16829 5502 16909 5518
rect 16829 5496 16848 5502
rect 16545 5470 16648 5480
rect 16499 5468 16648 5470
rect 16669 5468 16704 5480
rect 16338 5466 16500 5468
rect 16350 5446 16369 5466
rect 16384 5464 16414 5466
rect 16233 5438 16274 5446
rect 16356 5442 16369 5446
rect 16421 5450 16500 5466
rect 16532 5466 16704 5468
rect 16532 5450 16611 5466
rect 16618 5464 16648 5466
rect 16196 5428 16225 5438
rect 16239 5428 16268 5438
rect 16283 5428 16313 5442
rect 16356 5428 16399 5442
rect 16421 5438 16611 5450
rect 16676 5446 16682 5466
rect 16406 5428 16436 5438
rect 16437 5428 16595 5438
rect 16599 5428 16629 5438
rect 16633 5428 16663 5442
rect 16691 5428 16704 5466
rect 16776 5480 16805 5496
rect 16819 5480 16848 5496
rect 16863 5486 16893 5502
rect 16921 5480 16927 5528
rect 16930 5522 16949 5528
rect 16964 5522 16994 5530
rect 16930 5514 16994 5522
rect 16930 5498 17010 5514
rect 17026 5507 17088 5538
rect 17104 5507 17166 5538
rect 17235 5536 17284 5561
rect 17299 5536 17329 5552
rect 17198 5522 17228 5530
rect 17235 5528 17345 5536
rect 17198 5514 17243 5522
rect 16930 5496 16949 5498
rect 16964 5496 17010 5498
rect 16930 5480 17010 5496
rect 17037 5494 17072 5507
rect 17113 5504 17150 5507
rect 17113 5502 17155 5504
rect 17042 5491 17072 5494
rect 17051 5487 17058 5491
rect 17058 5486 17059 5487
rect 17017 5480 17027 5486
rect 16776 5472 16811 5480
rect 16776 5446 16777 5472
rect 16784 5446 16811 5472
rect 16719 5428 16749 5442
rect 16776 5438 16811 5446
rect 16813 5472 16854 5480
rect 16813 5446 16828 5472
rect 16835 5446 16854 5472
rect 16918 5468 16949 5480
rect 16964 5468 17067 5480
rect 17079 5470 17105 5496
rect 17120 5491 17150 5502
rect 17182 5498 17244 5514
rect 17182 5496 17228 5498
rect 17182 5480 17244 5496
rect 17256 5480 17262 5528
rect 17265 5520 17345 5528
rect 17265 5518 17284 5520
rect 17299 5518 17333 5520
rect 17265 5502 17345 5518
rect 17265 5480 17284 5502
rect 17299 5486 17329 5502
rect 17357 5496 17363 5570
rect 17366 5496 17385 5640
rect 17400 5496 17406 5640
rect 17415 5570 17428 5640
rect 17480 5636 17502 5640
rect 17473 5614 17502 5628
rect 17555 5614 17571 5628
rect 17609 5624 17615 5626
rect 17622 5624 17730 5640
rect 17737 5624 17743 5626
rect 17751 5624 17766 5640
rect 17832 5634 17851 5637
rect 17473 5612 17571 5614
rect 17598 5612 17766 5624
rect 17781 5614 17797 5628
rect 17832 5615 17854 5634
rect 17864 5628 17880 5629
rect 17863 5626 17880 5628
rect 17864 5621 17880 5626
rect 17854 5614 17860 5615
rect 17863 5614 17892 5621
rect 17781 5613 17892 5614
rect 17781 5612 17898 5613
rect 17457 5604 17508 5612
rect 17555 5604 17589 5612
rect 17457 5592 17482 5604
rect 17489 5592 17508 5604
rect 17562 5602 17589 5604
rect 17598 5602 17819 5612
rect 17854 5609 17860 5612
rect 17562 5598 17819 5602
rect 17457 5584 17508 5592
rect 17555 5584 17819 5598
rect 17863 5604 17898 5612
rect 17409 5536 17428 5570
rect 17473 5576 17502 5584
rect 17473 5570 17490 5576
rect 17473 5568 17507 5570
rect 17555 5568 17571 5584
rect 17572 5574 17780 5584
rect 17781 5574 17797 5584
rect 17845 5580 17860 5595
rect 17863 5592 17864 5604
rect 17871 5592 17898 5604
rect 17863 5584 17898 5592
rect 17863 5583 17892 5584
rect 17583 5570 17797 5574
rect 17598 5568 17797 5570
rect 17832 5570 17845 5580
rect 17863 5570 17880 5583
rect 17832 5568 17880 5570
rect 17474 5564 17507 5568
rect 17470 5562 17507 5564
rect 17470 5561 17537 5562
rect 17470 5556 17501 5561
rect 17507 5556 17537 5561
rect 17470 5552 17537 5556
rect 17443 5549 17537 5552
rect 17443 5542 17492 5549
rect 17443 5536 17473 5542
rect 17492 5537 17497 5542
rect 17409 5520 17489 5536
rect 17501 5528 17537 5549
rect 17598 5544 17787 5568
rect 17832 5567 17879 5568
rect 17845 5562 17879 5567
rect 17613 5541 17787 5544
rect 17606 5538 17787 5541
rect 17815 5561 17879 5562
rect 17409 5518 17428 5520
rect 17443 5518 17477 5520
rect 17409 5502 17489 5518
rect 17409 5496 17428 5502
rect 17125 5470 17228 5480
rect 17079 5468 17228 5470
rect 17249 5468 17284 5480
rect 16918 5466 17080 5468
rect 16930 5446 16949 5466
rect 16964 5464 16994 5466
rect 16813 5438 16854 5446
rect 16936 5442 16949 5446
rect 17001 5450 17080 5466
rect 17112 5466 17284 5468
rect 17112 5450 17191 5466
rect 17198 5464 17228 5466
rect 16776 5428 16805 5438
rect 16819 5428 16848 5438
rect 16863 5428 16893 5442
rect 16936 5428 16979 5442
rect 17001 5438 17191 5450
rect 17256 5446 17262 5466
rect 16986 5428 17016 5438
rect 17017 5428 17175 5438
rect 17179 5428 17209 5438
rect 17213 5428 17243 5442
rect 17271 5428 17284 5466
rect 17356 5480 17385 5496
rect 17399 5480 17428 5496
rect 17443 5486 17473 5502
rect 17501 5480 17507 5528
rect 17510 5522 17529 5528
rect 17544 5522 17574 5530
rect 17510 5514 17574 5522
rect 17510 5498 17590 5514
rect 17606 5507 17668 5538
rect 17684 5507 17746 5538
rect 17815 5536 17864 5561
rect 17879 5536 17909 5552
rect 17778 5522 17808 5530
rect 17815 5528 17925 5536
rect 17778 5514 17823 5522
rect 17510 5496 17529 5498
rect 17544 5496 17590 5498
rect 17510 5480 17590 5496
rect 17617 5494 17652 5507
rect 17693 5504 17730 5507
rect 17693 5502 17735 5504
rect 17622 5491 17652 5494
rect 17631 5487 17638 5491
rect 17638 5486 17639 5487
rect 17597 5480 17607 5486
rect 17356 5472 17391 5480
rect 17356 5446 17357 5472
rect 17364 5446 17391 5472
rect 17299 5428 17329 5442
rect 17356 5438 17391 5446
rect 17393 5472 17434 5480
rect 17393 5446 17408 5472
rect 17415 5446 17434 5472
rect 17498 5468 17529 5480
rect 17544 5468 17647 5480
rect 17659 5470 17685 5496
rect 17700 5491 17730 5502
rect 17762 5498 17824 5514
rect 17762 5496 17808 5498
rect 17762 5480 17824 5496
rect 17836 5480 17842 5528
rect 17845 5520 17925 5528
rect 17845 5518 17864 5520
rect 17879 5518 17913 5520
rect 17845 5502 17925 5518
rect 17845 5480 17864 5502
rect 17879 5486 17909 5502
rect 17937 5496 17943 5570
rect 17946 5496 17965 5640
rect 17980 5496 17986 5640
rect 17995 5570 18008 5640
rect 18060 5636 18082 5640
rect 18053 5614 18082 5628
rect 18135 5614 18151 5628
rect 18189 5624 18195 5626
rect 18202 5624 18310 5640
rect 18317 5624 18323 5626
rect 18331 5624 18346 5640
rect 18412 5634 18431 5637
rect 18053 5612 18151 5614
rect 18178 5612 18346 5624
rect 18361 5614 18377 5628
rect 18412 5615 18434 5634
rect 18444 5628 18460 5629
rect 18443 5626 18460 5628
rect 18444 5621 18460 5626
rect 18434 5614 18440 5615
rect 18443 5614 18472 5621
rect 18361 5613 18472 5614
rect 18361 5612 18478 5613
rect 18037 5604 18088 5612
rect 18135 5604 18169 5612
rect 18037 5592 18062 5604
rect 18069 5592 18088 5604
rect 18142 5602 18169 5604
rect 18178 5602 18399 5612
rect 18434 5609 18440 5612
rect 18142 5598 18399 5602
rect 18037 5584 18088 5592
rect 18135 5584 18399 5598
rect 18443 5604 18478 5612
rect 17989 5536 18008 5570
rect 18053 5576 18082 5584
rect 18053 5570 18070 5576
rect 18053 5568 18087 5570
rect 18135 5568 18151 5584
rect 18152 5574 18360 5584
rect 18361 5574 18377 5584
rect 18425 5580 18440 5595
rect 18443 5592 18444 5604
rect 18451 5592 18478 5604
rect 18443 5584 18478 5592
rect 18443 5583 18472 5584
rect 18163 5570 18377 5574
rect 18178 5568 18377 5570
rect 18412 5570 18425 5580
rect 18443 5570 18460 5583
rect 18412 5568 18460 5570
rect 18054 5564 18087 5568
rect 18050 5562 18087 5564
rect 18050 5561 18117 5562
rect 18050 5556 18081 5561
rect 18087 5556 18117 5561
rect 18050 5552 18117 5556
rect 18023 5549 18117 5552
rect 18023 5542 18072 5549
rect 18023 5536 18053 5542
rect 18072 5537 18077 5542
rect 17989 5520 18069 5536
rect 18081 5528 18117 5549
rect 18178 5544 18367 5568
rect 18412 5567 18459 5568
rect 18425 5562 18459 5567
rect 18193 5541 18367 5544
rect 18186 5538 18367 5541
rect 18395 5561 18459 5562
rect 17989 5518 18008 5520
rect 18023 5518 18057 5520
rect 17989 5502 18069 5518
rect 17989 5496 18008 5502
rect 17705 5470 17808 5480
rect 17659 5468 17808 5470
rect 17829 5468 17864 5480
rect 17498 5466 17660 5468
rect 17510 5446 17529 5466
rect 17544 5464 17574 5466
rect 17393 5438 17434 5446
rect 17516 5442 17529 5446
rect 17581 5450 17660 5466
rect 17692 5466 17864 5468
rect 17692 5450 17771 5466
rect 17778 5464 17808 5466
rect 17356 5428 17385 5438
rect 17399 5428 17428 5438
rect 17443 5428 17473 5442
rect 17516 5428 17559 5442
rect 17581 5438 17771 5450
rect 17836 5446 17842 5466
rect 17566 5428 17596 5438
rect 17597 5428 17755 5438
rect 17759 5428 17789 5438
rect 17793 5428 17823 5442
rect 17851 5428 17864 5466
rect 17936 5480 17965 5496
rect 17979 5480 18008 5496
rect 18023 5486 18053 5502
rect 18081 5480 18087 5528
rect 18090 5522 18109 5528
rect 18124 5522 18154 5530
rect 18090 5514 18154 5522
rect 18090 5498 18170 5514
rect 18186 5507 18248 5538
rect 18264 5507 18326 5538
rect 18395 5536 18444 5561
rect 18459 5536 18489 5552
rect 18358 5522 18388 5530
rect 18395 5528 18505 5536
rect 18358 5514 18403 5522
rect 18090 5496 18109 5498
rect 18124 5496 18170 5498
rect 18090 5480 18170 5496
rect 18197 5494 18232 5507
rect 18273 5504 18310 5507
rect 18273 5502 18315 5504
rect 18202 5491 18232 5494
rect 18211 5487 18218 5491
rect 18218 5486 18219 5487
rect 18177 5480 18187 5486
rect 17936 5472 17971 5480
rect 17936 5446 17937 5472
rect 17944 5446 17971 5472
rect 17879 5428 17909 5442
rect 17936 5438 17971 5446
rect 17973 5472 18014 5480
rect 17973 5446 17988 5472
rect 17995 5446 18014 5472
rect 18078 5468 18109 5480
rect 18124 5468 18227 5480
rect 18239 5470 18265 5496
rect 18280 5491 18310 5502
rect 18342 5498 18404 5514
rect 18342 5496 18388 5498
rect 18342 5480 18404 5496
rect 18416 5480 18422 5528
rect 18425 5520 18505 5528
rect 18425 5518 18444 5520
rect 18459 5518 18493 5520
rect 18425 5502 18505 5518
rect 18425 5480 18444 5502
rect 18459 5486 18489 5502
rect 18517 5496 18523 5570
rect 18532 5496 18545 5640
rect 18285 5470 18388 5480
rect 18239 5468 18388 5470
rect 18409 5468 18444 5480
rect 18078 5466 18240 5468
rect 18090 5446 18109 5466
rect 18124 5464 18154 5466
rect 17973 5438 18014 5446
rect 18096 5442 18109 5446
rect 18161 5450 18240 5466
rect 18272 5466 18444 5468
rect 18272 5450 18351 5466
rect 18358 5464 18388 5466
rect 17936 5428 17965 5438
rect 17979 5428 18008 5438
rect 18023 5428 18053 5442
rect 18096 5428 18139 5442
rect 18161 5438 18351 5450
rect 18416 5446 18422 5466
rect 18146 5428 18176 5438
rect 18177 5428 18335 5438
rect 18339 5428 18369 5438
rect 18373 5428 18403 5442
rect 18431 5428 18444 5466
rect 18516 5480 18545 5496
rect 18516 5472 18551 5480
rect 18516 5446 18517 5472
rect 18524 5446 18551 5472
rect 18459 5428 18489 5442
rect 18516 5438 18551 5446
rect 18516 5428 18545 5438
rect -1 5422 18545 5428
rect 0 5414 18545 5422
rect 15 5384 28 5414
rect 43 5400 73 5414
rect 116 5400 159 5414
rect 166 5400 386 5414
rect 393 5400 423 5414
rect 83 5386 98 5398
rect 117 5386 130 5400
rect 198 5396 351 5400
rect 80 5384 102 5386
rect 180 5384 372 5396
rect 451 5384 464 5414
rect 479 5400 509 5414
rect 546 5384 565 5414
rect 580 5384 586 5414
rect 595 5384 608 5414
rect 623 5400 653 5414
rect 696 5400 739 5414
rect 746 5400 966 5414
rect 973 5400 1003 5414
rect 663 5386 678 5398
rect 697 5386 710 5400
rect 778 5396 931 5400
rect 660 5384 682 5386
rect 760 5384 952 5396
rect 1031 5384 1044 5414
rect 1059 5400 1089 5414
rect 1126 5384 1145 5414
rect 1160 5384 1166 5414
rect 1175 5384 1188 5414
rect 1203 5400 1233 5414
rect 1276 5400 1319 5414
rect 1326 5400 1546 5414
rect 1553 5400 1583 5414
rect 1243 5386 1258 5398
rect 1277 5386 1290 5400
rect 1358 5396 1511 5400
rect 1240 5384 1262 5386
rect 1340 5384 1532 5396
rect 1611 5384 1624 5414
rect 1639 5400 1669 5414
rect 1706 5384 1725 5414
rect 1740 5384 1746 5414
rect 1755 5384 1768 5414
rect 1783 5400 1813 5414
rect 1856 5400 1899 5414
rect 1906 5400 2126 5414
rect 2133 5400 2163 5414
rect 1823 5386 1838 5398
rect 1857 5386 1870 5400
rect 1938 5396 2091 5400
rect 1820 5384 1842 5386
rect 1920 5384 2112 5396
rect 2191 5384 2204 5414
rect 2219 5400 2249 5414
rect 2286 5384 2305 5414
rect 2320 5384 2326 5414
rect 2335 5384 2348 5414
rect 2363 5400 2393 5414
rect 2436 5400 2479 5414
rect 2486 5400 2706 5414
rect 2713 5400 2743 5414
rect 2403 5386 2418 5398
rect 2437 5386 2450 5400
rect 2518 5396 2671 5400
rect 2400 5384 2422 5386
rect 2500 5384 2692 5396
rect 2771 5384 2784 5414
rect 2799 5400 2829 5414
rect 2866 5384 2885 5414
rect 2900 5384 2906 5414
rect 2915 5384 2928 5414
rect 2943 5400 2973 5414
rect 3016 5400 3059 5414
rect 3066 5400 3286 5414
rect 3293 5400 3323 5414
rect 2983 5386 2998 5398
rect 3017 5386 3030 5400
rect 3098 5396 3251 5400
rect 2980 5384 3002 5386
rect 3080 5384 3272 5396
rect 3351 5384 3364 5414
rect 3379 5400 3409 5414
rect 3446 5384 3465 5414
rect 3480 5384 3486 5414
rect 3495 5384 3508 5414
rect 3523 5400 3553 5414
rect 3596 5400 3639 5414
rect 3646 5400 3866 5414
rect 3873 5400 3903 5414
rect 3563 5386 3578 5398
rect 3597 5386 3610 5400
rect 3678 5396 3831 5400
rect 3560 5384 3582 5386
rect 3660 5384 3852 5396
rect 3931 5384 3944 5414
rect 3959 5400 3989 5414
rect 4026 5384 4045 5414
rect 4060 5384 4066 5414
rect 4075 5384 4088 5414
rect 4103 5400 4133 5414
rect 4176 5400 4219 5414
rect 4226 5400 4446 5414
rect 4453 5400 4483 5414
rect 4143 5386 4158 5398
rect 4177 5386 4190 5400
rect 4258 5396 4411 5400
rect 4140 5384 4162 5386
rect 4240 5384 4432 5396
rect 4511 5384 4524 5414
rect 4539 5400 4569 5414
rect 4606 5384 4625 5414
rect 4640 5384 4646 5414
rect 4655 5384 4668 5414
rect 4683 5400 4713 5414
rect 4756 5400 4799 5414
rect 4806 5400 5026 5414
rect 5033 5400 5063 5414
rect 4723 5386 4738 5398
rect 4757 5386 4770 5400
rect 4838 5396 4991 5400
rect 4720 5384 4742 5386
rect 4820 5384 5012 5396
rect 5091 5384 5104 5414
rect 5119 5400 5149 5414
rect 5186 5384 5205 5414
rect 5220 5384 5226 5414
rect 5235 5384 5248 5414
rect 5263 5400 5293 5414
rect 5336 5400 5379 5414
rect 5386 5400 5606 5414
rect 5613 5400 5643 5414
rect 5303 5386 5318 5398
rect 5337 5386 5350 5400
rect 5418 5396 5571 5400
rect 5300 5384 5322 5386
rect 5400 5384 5592 5396
rect 5671 5384 5684 5414
rect 5699 5400 5729 5414
rect 5766 5384 5785 5414
rect 5800 5384 5806 5414
rect 5815 5384 5828 5414
rect 5843 5400 5873 5414
rect 5916 5400 5959 5414
rect 5966 5400 6186 5414
rect 6193 5400 6223 5414
rect 5883 5386 5898 5398
rect 5917 5386 5930 5400
rect 5998 5396 6151 5400
rect 5880 5384 5902 5386
rect 5980 5384 6172 5396
rect 6251 5384 6264 5414
rect 6279 5400 6309 5414
rect 6346 5384 6365 5414
rect 6380 5384 6386 5414
rect 6395 5384 6408 5414
rect 6423 5400 6453 5414
rect 6496 5400 6539 5414
rect 6546 5400 6766 5414
rect 6773 5400 6803 5414
rect 6463 5386 6478 5398
rect 6497 5386 6510 5400
rect 6578 5396 6731 5400
rect 6460 5384 6482 5386
rect 6560 5384 6752 5396
rect 6831 5384 6844 5414
rect 6859 5400 6889 5414
rect 6926 5384 6945 5414
rect 6960 5384 6966 5414
rect 6975 5384 6988 5414
rect 7003 5400 7033 5414
rect 7076 5400 7119 5414
rect 7126 5400 7346 5414
rect 7353 5400 7383 5414
rect 7043 5386 7058 5398
rect 7077 5386 7090 5400
rect 7158 5396 7311 5400
rect 7040 5384 7062 5386
rect 7140 5384 7332 5396
rect 7411 5384 7424 5414
rect 7439 5400 7469 5414
rect 7506 5384 7525 5414
rect 7540 5384 7546 5414
rect 7555 5384 7568 5414
rect 7583 5400 7613 5414
rect 7656 5400 7699 5414
rect 7706 5400 7926 5414
rect 7933 5400 7963 5414
rect 7623 5386 7638 5398
rect 7657 5386 7670 5400
rect 7738 5396 7891 5400
rect 7620 5384 7642 5386
rect 7720 5384 7912 5396
rect 7991 5384 8004 5414
rect 8019 5400 8049 5414
rect 8086 5384 8105 5414
rect 8120 5384 8126 5414
rect 8135 5384 8148 5414
rect 8163 5400 8193 5414
rect 8236 5400 8279 5414
rect 8286 5400 8506 5414
rect 8513 5400 8543 5414
rect 8203 5386 8218 5398
rect 8237 5386 8250 5400
rect 8318 5396 8471 5400
rect 8200 5384 8222 5386
rect 8300 5384 8492 5396
rect 8571 5384 8584 5414
rect 8599 5400 8629 5414
rect 8666 5384 8685 5414
rect 8700 5384 8706 5414
rect 8715 5384 8728 5414
rect 8743 5400 8773 5414
rect 8816 5400 8859 5414
rect 8866 5400 9086 5414
rect 9093 5400 9123 5414
rect 8783 5386 8798 5398
rect 8817 5386 8830 5400
rect 8898 5396 9051 5400
rect 8780 5384 8802 5386
rect 8880 5384 9072 5396
rect 9151 5384 9164 5414
rect 9179 5400 9209 5414
rect 9246 5384 9265 5414
rect 9280 5384 9286 5414
rect 9295 5384 9308 5414
rect 9323 5400 9353 5414
rect 9396 5400 9439 5414
rect 9446 5400 9666 5414
rect 9673 5400 9703 5414
rect 9363 5386 9378 5398
rect 9397 5386 9410 5400
rect 9478 5396 9631 5400
rect 9360 5384 9382 5386
rect 9460 5384 9652 5396
rect 9731 5384 9744 5414
rect 9759 5400 9789 5414
rect 9826 5384 9845 5414
rect 9860 5384 9866 5414
rect 9875 5384 9888 5414
rect 9903 5400 9933 5414
rect 9976 5400 10019 5414
rect 10026 5400 10246 5414
rect 10253 5400 10283 5414
rect 9943 5386 9958 5398
rect 9977 5386 9990 5400
rect 10058 5396 10211 5400
rect 9940 5384 9962 5386
rect 10040 5384 10232 5396
rect 10311 5384 10324 5414
rect 10339 5400 10369 5414
rect 10406 5384 10425 5414
rect 10440 5384 10446 5414
rect 10455 5384 10468 5414
rect 10483 5400 10513 5414
rect 10556 5400 10599 5414
rect 10606 5400 10826 5414
rect 10833 5400 10863 5414
rect 10523 5386 10538 5398
rect 10557 5386 10570 5400
rect 10638 5396 10791 5400
rect 10520 5384 10542 5386
rect 10620 5384 10812 5396
rect 10891 5384 10904 5414
rect 10919 5400 10949 5414
rect 10986 5384 11005 5414
rect 11020 5384 11026 5414
rect 11035 5384 11048 5414
rect 11063 5400 11093 5414
rect 11136 5400 11179 5414
rect 11186 5400 11406 5414
rect 11413 5400 11443 5414
rect 11103 5386 11118 5398
rect 11137 5386 11150 5400
rect 11218 5396 11371 5400
rect 11100 5384 11122 5386
rect 11200 5384 11392 5396
rect 11471 5384 11484 5414
rect 11499 5400 11529 5414
rect 11566 5384 11585 5414
rect 11600 5384 11606 5414
rect 11615 5384 11628 5414
rect 11643 5400 11673 5414
rect 11716 5400 11759 5414
rect 11766 5400 11986 5414
rect 11993 5400 12023 5414
rect 11683 5386 11698 5398
rect 11717 5386 11730 5400
rect 11798 5396 11951 5400
rect 11680 5384 11702 5386
rect 11780 5384 11972 5396
rect 12051 5384 12064 5414
rect 12079 5400 12109 5414
rect 12146 5384 12165 5414
rect 12180 5384 12186 5414
rect 12195 5384 12208 5414
rect 12223 5400 12253 5414
rect 12296 5400 12339 5414
rect 12346 5400 12566 5414
rect 12573 5400 12603 5414
rect 12263 5386 12278 5398
rect 12297 5386 12310 5400
rect 12378 5396 12531 5400
rect 12260 5384 12282 5386
rect 12360 5384 12552 5396
rect 12631 5384 12644 5414
rect 12659 5400 12689 5414
rect 12726 5384 12745 5414
rect 12760 5384 12766 5414
rect 12775 5384 12788 5414
rect 12803 5400 12833 5414
rect 12876 5400 12919 5414
rect 12926 5400 13146 5414
rect 13153 5400 13183 5414
rect 12843 5386 12858 5398
rect 12877 5386 12890 5400
rect 12958 5396 13111 5400
rect 12840 5384 12862 5386
rect 12940 5384 13132 5396
rect 13211 5384 13224 5414
rect 13239 5400 13269 5414
rect 13306 5384 13325 5414
rect 13340 5384 13346 5414
rect 13355 5384 13368 5414
rect 13383 5400 13413 5414
rect 13456 5400 13499 5414
rect 13506 5400 13726 5414
rect 13733 5400 13763 5414
rect 13423 5386 13438 5398
rect 13457 5386 13470 5400
rect 13538 5396 13691 5400
rect 13420 5384 13442 5386
rect 13520 5384 13712 5396
rect 13791 5384 13804 5414
rect 13819 5400 13849 5414
rect 13886 5384 13905 5414
rect 13920 5384 13926 5414
rect 13935 5384 13948 5414
rect 13963 5400 13993 5414
rect 14036 5400 14079 5414
rect 14086 5400 14306 5414
rect 14313 5400 14343 5414
rect 14003 5386 14018 5398
rect 14037 5386 14050 5400
rect 14118 5396 14271 5400
rect 14000 5384 14022 5386
rect 14100 5384 14292 5396
rect 14371 5384 14384 5414
rect 14399 5400 14429 5414
rect 14466 5384 14485 5414
rect 14500 5384 14506 5414
rect 14515 5384 14528 5414
rect 14543 5400 14573 5414
rect 14616 5400 14659 5414
rect 14666 5400 14886 5414
rect 14893 5400 14923 5414
rect 14583 5386 14598 5398
rect 14617 5386 14630 5400
rect 14698 5396 14851 5400
rect 14580 5384 14602 5386
rect 14680 5384 14872 5396
rect 14951 5384 14964 5414
rect 14979 5400 15009 5414
rect 15046 5384 15065 5414
rect 15080 5384 15086 5414
rect 15095 5384 15108 5414
rect 15123 5400 15153 5414
rect 15196 5400 15239 5414
rect 15246 5400 15466 5414
rect 15473 5400 15503 5414
rect 15163 5386 15178 5398
rect 15197 5386 15210 5400
rect 15278 5396 15431 5400
rect 15160 5384 15182 5386
rect 15260 5384 15452 5396
rect 15531 5384 15544 5414
rect 15559 5400 15589 5414
rect 15626 5384 15645 5414
rect 15660 5384 15666 5414
rect 15675 5384 15688 5414
rect 15703 5400 15733 5414
rect 15776 5400 15819 5414
rect 15826 5400 16046 5414
rect 16053 5400 16083 5414
rect 15743 5386 15758 5398
rect 15777 5386 15790 5400
rect 15858 5396 16011 5400
rect 15740 5384 15762 5386
rect 15840 5384 16032 5396
rect 16111 5384 16124 5414
rect 16139 5400 16169 5414
rect 16206 5384 16225 5414
rect 16240 5384 16246 5414
rect 16255 5384 16268 5414
rect 16283 5400 16313 5414
rect 16356 5400 16399 5414
rect 16406 5400 16626 5414
rect 16633 5400 16663 5414
rect 16323 5386 16338 5398
rect 16357 5386 16370 5400
rect 16438 5396 16591 5400
rect 16320 5384 16342 5386
rect 16420 5384 16612 5396
rect 16691 5384 16704 5414
rect 16719 5400 16749 5414
rect 16786 5384 16805 5414
rect 16820 5384 16826 5414
rect 16835 5384 16848 5414
rect 16863 5400 16893 5414
rect 16936 5400 16979 5414
rect 16986 5400 17206 5414
rect 17213 5400 17243 5414
rect 16903 5386 16918 5398
rect 16937 5386 16950 5400
rect 17018 5396 17171 5400
rect 16900 5384 16922 5386
rect 17000 5384 17192 5396
rect 17271 5384 17284 5414
rect 17299 5400 17329 5414
rect 17366 5384 17385 5414
rect 17400 5384 17406 5414
rect 17415 5384 17428 5414
rect 17443 5400 17473 5414
rect 17516 5400 17559 5414
rect 17566 5400 17786 5414
rect 17793 5400 17823 5414
rect 17483 5386 17498 5398
rect 17517 5386 17530 5400
rect 17598 5396 17751 5400
rect 17480 5384 17502 5386
rect 17580 5384 17772 5396
rect 17851 5384 17864 5414
rect 17879 5400 17909 5414
rect 17946 5384 17965 5414
rect 17980 5384 17986 5414
rect 17995 5384 18008 5414
rect 18023 5400 18053 5414
rect 18096 5400 18139 5414
rect 18146 5400 18366 5414
rect 18373 5400 18403 5414
rect 18063 5386 18078 5398
rect 18097 5386 18110 5400
rect 18178 5396 18331 5400
rect 18060 5384 18082 5386
rect 18160 5384 18352 5396
rect 18431 5384 18444 5414
rect 18459 5400 18489 5414
rect 18532 5384 18545 5414
rect 0 5370 18545 5384
rect 15 5300 28 5370
rect 80 5366 102 5370
rect 73 5344 102 5358
rect 155 5344 171 5358
rect 209 5354 215 5356
rect 222 5354 330 5370
rect 337 5354 343 5356
rect 351 5354 366 5370
rect 432 5364 451 5367
rect 73 5342 171 5344
rect 198 5342 366 5354
rect 381 5344 397 5358
rect 432 5345 454 5364
rect 464 5358 480 5359
rect 463 5356 480 5358
rect 464 5351 480 5356
rect 454 5344 460 5345
rect 463 5344 492 5351
rect 381 5343 492 5344
rect 381 5342 498 5343
rect 57 5334 108 5342
rect 155 5334 189 5342
rect 57 5322 82 5334
rect 89 5322 108 5334
rect 162 5332 189 5334
rect 198 5332 419 5342
rect 454 5339 460 5342
rect 162 5328 419 5332
rect 57 5314 108 5322
rect 155 5314 419 5328
rect 463 5334 498 5342
rect 9 5266 28 5300
rect 73 5306 102 5314
rect 73 5300 90 5306
rect 73 5298 107 5300
rect 155 5298 171 5314
rect 172 5304 380 5314
rect 381 5304 397 5314
rect 445 5310 460 5325
rect 463 5322 464 5334
rect 471 5322 498 5334
rect 463 5314 498 5322
rect 463 5313 492 5314
rect 183 5300 397 5304
rect 198 5298 397 5300
rect 432 5300 445 5310
rect 463 5300 480 5313
rect 432 5298 480 5300
rect 74 5294 107 5298
rect 70 5292 107 5294
rect 70 5291 137 5292
rect 70 5286 101 5291
rect 107 5286 137 5291
rect 70 5282 137 5286
rect 43 5279 137 5282
rect 43 5272 92 5279
rect 43 5266 73 5272
rect 92 5267 97 5272
rect 9 5250 89 5266
rect 101 5258 137 5279
rect 198 5274 387 5298
rect 432 5297 479 5298
rect 445 5292 479 5297
rect 213 5271 387 5274
rect 206 5268 387 5271
rect 415 5291 479 5292
rect 9 5248 28 5250
rect 43 5248 77 5250
rect 9 5232 89 5248
rect 9 5226 28 5232
rect -1 5210 28 5226
rect 43 5216 73 5232
rect 101 5210 107 5258
rect 110 5252 129 5258
rect 144 5252 174 5260
rect 110 5244 174 5252
rect 110 5228 190 5244
rect 206 5237 268 5268
rect 284 5237 346 5268
rect 415 5266 464 5291
rect 479 5266 509 5282
rect 378 5252 408 5260
rect 415 5258 525 5266
rect 378 5244 423 5252
rect 110 5226 129 5228
rect 144 5226 190 5228
rect 110 5210 190 5226
rect 217 5224 252 5237
rect 293 5234 330 5237
rect 293 5232 335 5234
rect 222 5221 252 5224
rect 231 5217 238 5221
rect 238 5216 239 5217
rect 197 5210 207 5216
rect -7 5202 34 5210
rect -7 5176 8 5202
rect 15 5176 34 5202
rect 98 5198 129 5210
rect 144 5198 247 5210
rect 259 5200 285 5226
rect 300 5221 330 5232
rect 362 5228 424 5244
rect 362 5226 408 5228
rect 362 5210 424 5226
rect 436 5210 442 5258
rect 445 5250 525 5258
rect 445 5248 464 5250
rect 479 5248 513 5250
rect 445 5232 525 5248
rect 445 5210 464 5232
rect 479 5216 509 5232
rect 537 5226 543 5300
rect 546 5226 565 5370
rect 580 5226 586 5370
rect 595 5300 608 5370
rect 660 5366 682 5370
rect 653 5344 682 5358
rect 735 5344 751 5358
rect 789 5354 795 5356
rect 802 5354 910 5370
rect 917 5354 923 5356
rect 931 5354 946 5370
rect 1012 5364 1031 5367
rect 653 5342 751 5344
rect 778 5342 946 5354
rect 961 5344 977 5358
rect 1012 5345 1034 5364
rect 1044 5358 1060 5359
rect 1043 5356 1060 5358
rect 1044 5351 1060 5356
rect 1034 5344 1040 5345
rect 1043 5344 1072 5351
rect 961 5343 1072 5344
rect 961 5342 1078 5343
rect 637 5334 688 5342
rect 735 5334 769 5342
rect 637 5322 662 5334
rect 669 5322 688 5334
rect 742 5332 769 5334
rect 778 5332 999 5342
rect 1034 5339 1040 5342
rect 742 5328 999 5332
rect 637 5314 688 5322
rect 735 5314 999 5328
rect 1043 5334 1078 5342
rect 589 5266 608 5300
rect 653 5306 682 5314
rect 653 5300 670 5306
rect 653 5298 687 5300
rect 735 5298 751 5314
rect 752 5304 960 5314
rect 961 5304 977 5314
rect 1025 5310 1040 5325
rect 1043 5322 1044 5334
rect 1051 5322 1078 5334
rect 1043 5314 1078 5322
rect 1043 5313 1072 5314
rect 763 5300 977 5304
rect 778 5298 977 5300
rect 1012 5300 1025 5310
rect 1043 5300 1060 5313
rect 1012 5298 1060 5300
rect 654 5294 687 5298
rect 650 5292 687 5294
rect 650 5291 717 5292
rect 650 5286 681 5291
rect 687 5286 717 5291
rect 650 5282 717 5286
rect 623 5279 717 5282
rect 623 5272 672 5279
rect 623 5266 653 5272
rect 672 5267 677 5272
rect 589 5250 669 5266
rect 681 5258 717 5279
rect 778 5274 967 5298
rect 1012 5297 1059 5298
rect 1025 5292 1059 5297
rect 793 5271 967 5274
rect 786 5268 967 5271
rect 995 5291 1059 5292
rect 589 5248 608 5250
rect 623 5248 657 5250
rect 589 5232 669 5248
rect 589 5226 608 5232
rect 305 5200 408 5210
rect 259 5198 408 5200
rect 429 5198 464 5210
rect 98 5196 260 5198
rect 110 5176 129 5196
rect 144 5194 174 5196
rect -7 5168 34 5176
rect 116 5172 129 5176
rect 181 5180 260 5196
rect 292 5196 464 5198
rect 292 5180 371 5196
rect 378 5194 408 5196
rect -1 5158 28 5168
rect 43 5158 73 5172
rect 116 5158 159 5172
rect 181 5168 371 5180
rect 436 5176 442 5196
rect 166 5158 196 5168
rect 197 5158 355 5168
rect 359 5158 389 5168
rect 393 5158 423 5172
rect 451 5158 464 5196
rect 536 5210 565 5226
rect 579 5210 608 5226
rect 623 5216 653 5232
rect 681 5210 687 5258
rect 690 5252 709 5258
rect 724 5252 754 5260
rect 690 5244 754 5252
rect 690 5228 770 5244
rect 786 5237 848 5268
rect 864 5237 926 5268
rect 995 5266 1044 5291
rect 1059 5266 1089 5282
rect 958 5252 988 5260
rect 995 5258 1105 5266
rect 958 5244 1003 5252
rect 690 5226 709 5228
rect 724 5226 770 5228
rect 690 5210 770 5226
rect 797 5224 832 5237
rect 873 5234 910 5237
rect 873 5232 915 5234
rect 802 5221 832 5224
rect 811 5217 818 5221
rect 818 5216 819 5217
rect 777 5210 787 5216
rect 536 5202 571 5210
rect 536 5176 537 5202
rect 544 5176 571 5202
rect 479 5158 509 5172
rect 536 5168 571 5176
rect 573 5202 614 5210
rect 573 5176 588 5202
rect 595 5176 614 5202
rect 678 5198 709 5210
rect 724 5198 827 5210
rect 839 5200 865 5226
rect 880 5221 910 5232
rect 942 5228 1004 5244
rect 942 5226 988 5228
rect 942 5210 1004 5226
rect 1016 5210 1022 5258
rect 1025 5250 1105 5258
rect 1025 5248 1044 5250
rect 1059 5248 1093 5250
rect 1025 5232 1105 5248
rect 1025 5210 1044 5232
rect 1059 5216 1089 5232
rect 1117 5226 1123 5300
rect 1126 5226 1145 5370
rect 1160 5226 1166 5370
rect 1175 5300 1188 5370
rect 1240 5366 1262 5370
rect 1233 5344 1262 5358
rect 1315 5344 1331 5358
rect 1369 5354 1375 5356
rect 1382 5354 1490 5370
rect 1497 5354 1503 5356
rect 1511 5354 1526 5370
rect 1592 5364 1611 5367
rect 1233 5342 1331 5344
rect 1358 5342 1526 5354
rect 1541 5344 1557 5358
rect 1592 5345 1614 5364
rect 1624 5358 1640 5359
rect 1623 5356 1640 5358
rect 1624 5351 1640 5356
rect 1614 5344 1620 5345
rect 1623 5344 1652 5351
rect 1541 5343 1652 5344
rect 1541 5342 1658 5343
rect 1217 5334 1268 5342
rect 1315 5334 1349 5342
rect 1217 5322 1242 5334
rect 1249 5322 1268 5334
rect 1322 5332 1349 5334
rect 1358 5332 1579 5342
rect 1614 5339 1620 5342
rect 1322 5328 1579 5332
rect 1217 5314 1268 5322
rect 1315 5314 1579 5328
rect 1623 5334 1658 5342
rect 1169 5266 1188 5300
rect 1233 5306 1262 5314
rect 1233 5300 1250 5306
rect 1233 5298 1267 5300
rect 1315 5298 1331 5314
rect 1332 5304 1540 5314
rect 1541 5304 1557 5314
rect 1605 5310 1620 5325
rect 1623 5322 1624 5334
rect 1631 5322 1658 5334
rect 1623 5314 1658 5322
rect 1623 5313 1652 5314
rect 1343 5300 1557 5304
rect 1358 5298 1557 5300
rect 1592 5300 1605 5310
rect 1623 5300 1640 5313
rect 1592 5298 1640 5300
rect 1234 5294 1267 5298
rect 1230 5292 1267 5294
rect 1230 5291 1297 5292
rect 1230 5286 1261 5291
rect 1267 5286 1297 5291
rect 1230 5282 1297 5286
rect 1203 5279 1297 5282
rect 1203 5272 1252 5279
rect 1203 5266 1233 5272
rect 1252 5267 1257 5272
rect 1169 5250 1249 5266
rect 1261 5258 1297 5279
rect 1358 5274 1547 5298
rect 1592 5297 1639 5298
rect 1605 5292 1639 5297
rect 1373 5271 1547 5274
rect 1366 5268 1547 5271
rect 1575 5291 1639 5292
rect 1169 5248 1188 5250
rect 1203 5248 1237 5250
rect 1169 5232 1249 5248
rect 1169 5226 1188 5232
rect 885 5200 988 5210
rect 839 5198 988 5200
rect 1009 5198 1044 5210
rect 678 5196 840 5198
rect 690 5176 709 5196
rect 724 5194 754 5196
rect 573 5168 614 5176
rect 696 5172 709 5176
rect 761 5180 840 5196
rect 872 5196 1044 5198
rect 872 5180 951 5196
rect 958 5194 988 5196
rect 536 5158 565 5168
rect 579 5158 608 5168
rect 623 5158 653 5172
rect 696 5158 739 5172
rect 761 5168 951 5180
rect 1016 5176 1022 5196
rect 746 5158 776 5168
rect 777 5158 935 5168
rect 939 5158 969 5168
rect 973 5158 1003 5172
rect 1031 5158 1044 5196
rect 1116 5210 1145 5226
rect 1159 5210 1188 5226
rect 1203 5216 1233 5232
rect 1261 5210 1267 5258
rect 1270 5252 1289 5258
rect 1304 5252 1334 5260
rect 1270 5244 1334 5252
rect 1270 5228 1350 5244
rect 1366 5237 1428 5268
rect 1444 5237 1506 5268
rect 1575 5266 1624 5291
rect 1639 5266 1669 5282
rect 1538 5252 1568 5260
rect 1575 5258 1685 5266
rect 1538 5244 1583 5252
rect 1270 5226 1289 5228
rect 1304 5226 1350 5228
rect 1270 5210 1350 5226
rect 1377 5224 1412 5237
rect 1453 5234 1490 5237
rect 1453 5232 1495 5234
rect 1382 5221 1412 5224
rect 1391 5217 1398 5221
rect 1398 5216 1399 5217
rect 1357 5210 1367 5216
rect 1116 5202 1151 5210
rect 1116 5176 1117 5202
rect 1124 5176 1151 5202
rect 1059 5158 1089 5172
rect 1116 5168 1151 5176
rect 1153 5202 1194 5210
rect 1153 5176 1168 5202
rect 1175 5176 1194 5202
rect 1258 5198 1289 5210
rect 1304 5198 1407 5210
rect 1419 5200 1445 5226
rect 1460 5221 1490 5232
rect 1522 5228 1584 5244
rect 1522 5226 1568 5228
rect 1522 5210 1584 5226
rect 1596 5210 1602 5258
rect 1605 5250 1685 5258
rect 1605 5248 1624 5250
rect 1639 5248 1673 5250
rect 1605 5232 1685 5248
rect 1605 5210 1624 5232
rect 1639 5216 1669 5232
rect 1697 5226 1703 5300
rect 1706 5226 1725 5370
rect 1740 5226 1746 5370
rect 1755 5300 1768 5370
rect 1820 5366 1842 5370
rect 1813 5344 1842 5358
rect 1895 5344 1911 5358
rect 1949 5354 1955 5356
rect 1962 5354 2070 5370
rect 2077 5354 2083 5356
rect 2091 5354 2106 5370
rect 2172 5364 2191 5367
rect 1813 5342 1911 5344
rect 1938 5342 2106 5354
rect 2121 5344 2137 5358
rect 2172 5345 2194 5364
rect 2204 5358 2220 5359
rect 2203 5356 2220 5358
rect 2204 5351 2220 5356
rect 2194 5344 2200 5345
rect 2203 5344 2232 5351
rect 2121 5343 2232 5344
rect 2121 5342 2238 5343
rect 1797 5334 1848 5342
rect 1895 5334 1929 5342
rect 1797 5322 1822 5334
rect 1829 5322 1848 5334
rect 1902 5332 1929 5334
rect 1938 5332 2159 5342
rect 2194 5339 2200 5342
rect 1902 5328 2159 5332
rect 1797 5314 1848 5322
rect 1895 5314 2159 5328
rect 2203 5334 2238 5342
rect 1749 5266 1768 5300
rect 1813 5306 1842 5314
rect 1813 5300 1830 5306
rect 1813 5298 1847 5300
rect 1895 5298 1911 5314
rect 1912 5304 2120 5314
rect 2121 5304 2137 5314
rect 2185 5310 2200 5325
rect 2203 5322 2204 5334
rect 2211 5322 2238 5334
rect 2203 5314 2238 5322
rect 2203 5313 2232 5314
rect 1923 5300 2137 5304
rect 1938 5298 2137 5300
rect 2172 5300 2185 5310
rect 2203 5300 2220 5313
rect 2172 5298 2220 5300
rect 1814 5294 1847 5298
rect 1810 5292 1847 5294
rect 1810 5291 1877 5292
rect 1810 5286 1841 5291
rect 1847 5286 1877 5291
rect 1810 5282 1877 5286
rect 1783 5279 1877 5282
rect 1783 5272 1832 5279
rect 1783 5266 1813 5272
rect 1832 5267 1837 5272
rect 1749 5250 1829 5266
rect 1841 5258 1877 5279
rect 1938 5274 2127 5298
rect 2172 5297 2219 5298
rect 2185 5292 2219 5297
rect 1953 5271 2127 5274
rect 1946 5268 2127 5271
rect 2155 5291 2219 5292
rect 1749 5248 1768 5250
rect 1783 5248 1817 5250
rect 1749 5232 1829 5248
rect 1749 5226 1768 5232
rect 1465 5200 1568 5210
rect 1419 5198 1568 5200
rect 1589 5198 1624 5210
rect 1258 5196 1420 5198
rect 1270 5176 1289 5196
rect 1304 5194 1334 5196
rect 1153 5168 1194 5176
rect 1276 5172 1289 5176
rect 1341 5180 1420 5196
rect 1452 5196 1624 5198
rect 1452 5180 1531 5196
rect 1538 5194 1568 5196
rect 1116 5158 1145 5168
rect 1159 5158 1188 5168
rect 1203 5158 1233 5172
rect 1276 5158 1319 5172
rect 1341 5168 1531 5180
rect 1596 5176 1602 5196
rect 1326 5158 1356 5168
rect 1357 5158 1515 5168
rect 1519 5158 1549 5168
rect 1553 5158 1583 5172
rect 1611 5158 1624 5196
rect 1696 5210 1725 5226
rect 1739 5210 1768 5226
rect 1783 5216 1813 5232
rect 1841 5210 1847 5258
rect 1850 5252 1869 5258
rect 1884 5252 1914 5260
rect 1850 5244 1914 5252
rect 1850 5228 1930 5244
rect 1946 5237 2008 5268
rect 2024 5237 2086 5268
rect 2155 5266 2204 5291
rect 2219 5266 2249 5282
rect 2118 5252 2148 5260
rect 2155 5258 2265 5266
rect 2118 5244 2163 5252
rect 1850 5226 1869 5228
rect 1884 5226 1930 5228
rect 1850 5210 1930 5226
rect 1957 5224 1992 5237
rect 2033 5234 2070 5237
rect 2033 5232 2075 5234
rect 1962 5221 1992 5224
rect 1971 5217 1978 5221
rect 1978 5216 1979 5217
rect 1937 5210 1947 5216
rect 1696 5202 1731 5210
rect 1696 5176 1697 5202
rect 1704 5176 1731 5202
rect 1639 5158 1669 5172
rect 1696 5168 1731 5176
rect 1733 5202 1774 5210
rect 1733 5176 1748 5202
rect 1755 5176 1774 5202
rect 1838 5198 1869 5210
rect 1884 5198 1987 5210
rect 1999 5200 2025 5226
rect 2040 5221 2070 5232
rect 2102 5228 2164 5244
rect 2102 5226 2148 5228
rect 2102 5210 2164 5226
rect 2176 5210 2182 5258
rect 2185 5250 2265 5258
rect 2185 5248 2204 5250
rect 2219 5248 2253 5250
rect 2185 5232 2265 5248
rect 2185 5210 2204 5232
rect 2219 5216 2249 5232
rect 2277 5226 2283 5300
rect 2286 5226 2305 5370
rect 2320 5226 2326 5370
rect 2335 5300 2348 5370
rect 2400 5366 2422 5370
rect 2393 5344 2422 5358
rect 2475 5344 2491 5358
rect 2529 5354 2535 5356
rect 2542 5354 2650 5370
rect 2657 5354 2663 5356
rect 2671 5354 2686 5370
rect 2752 5364 2771 5367
rect 2393 5342 2491 5344
rect 2518 5342 2686 5354
rect 2701 5344 2717 5358
rect 2752 5345 2774 5364
rect 2784 5358 2800 5359
rect 2783 5356 2800 5358
rect 2784 5351 2800 5356
rect 2774 5344 2780 5345
rect 2783 5344 2812 5351
rect 2701 5343 2812 5344
rect 2701 5342 2818 5343
rect 2377 5334 2428 5342
rect 2475 5334 2509 5342
rect 2377 5322 2402 5334
rect 2409 5322 2428 5334
rect 2482 5332 2509 5334
rect 2518 5332 2739 5342
rect 2774 5339 2780 5342
rect 2482 5328 2739 5332
rect 2377 5314 2428 5322
rect 2475 5314 2739 5328
rect 2783 5334 2818 5342
rect 2329 5266 2348 5300
rect 2393 5306 2422 5314
rect 2393 5300 2410 5306
rect 2393 5298 2427 5300
rect 2475 5298 2491 5314
rect 2492 5304 2700 5314
rect 2701 5304 2717 5314
rect 2765 5310 2780 5325
rect 2783 5322 2784 5334
rect 2791 5322 2818 5334
rect 2783 5314 2818 5322
rect 2783 5313 2812 5314
rect 2503 5300 2717 5304
rect 2518 5298 2717 5300
rect 2752 5300 2765 5310
rect 2783 5300 2800 5313
rect 2752 5298 2800 5300
rect 2394 5294 2427 5298
rect 2390 5292 2427 5294
rect 2390 5291 2457 5292
rect 2390 5286 2421 5291
rect 2427 5286 2457 5291
rect 2390 5282 2457 5286
rect 2363 5279 2457 5282
rect 2363 5272 2412 5279
rect 2363 5266 2393 5272
rect 2412 5267 2417 5272
rect 2329 5250 2409 5266
rect 2421 5258 2457 5279
rect 2518 5274 2707 5298
rect 2752 5297 2799 5298
rect 2765 5292 2799 5297
rect 2533 5271 2707 5274
rect 2526 5268 2707 5271
rect 2735 5291 2799 5292
rect 2329 5248 2348 5250
rect 2363 5248 2397 5250
rect 2329 5232 2409 5248
rect 2329 5226 2348 5232
rect 2045 5200 2148 5210
rect 1999 5198 2148 5200
rect 2169 5198 2204 5210
rect 1838 5196 2000 5198
rect 1850 5176 1869 5196
rect 1884 5194 1914 5196
rect 1733 5168 1774 5176
rect 1856 5172 1869 5176
rect 1921 5180 2000 5196
rect 2032 5196 2204 5198
rect 2032 5180 2111 5196
rect 2118 5194 2148 5196
rect 1696 5158 1725 5168
rect 1739 5158 1768 5168
rect 1783 5158 1813 5172
rect 1856 5158 1899 5172
rect 1921 5168 2111 5180
rect 2176 5176 2182 5196
rect 1906 5158 1936 5168
rect 1937 5158 2095 5168
rect 2099 5158 2129 5168
rect 2133 5158 2163 5172
rect 2191 5158 2204 5196
rect 2276 5210 2305 5226
rect 2319 5210 2348 5226
rect 2363 5216 2393 5232
rect 2421 5210 2427 5258
rect 2430 5252 2449 5258
rect 2464 5252 2494 5260
rect 2430 5244 2494 5252
rect 2430 5228 2510 5244
rect 2526 5237 2588 5268
rect 2604 5237 2666 5268
rect 2735 5266 2784 5291
rect 2799 5266 2829 5282
rect 2698 5252 2728 5260
rect 2735 5258 2845 5266
rect 2698 5244 2743 5252
rect 2430 5226 2449 5228
rect 2464 5226 2510 5228
rect 2430 5210 2510 5226
rect 2537 5224 2572 5237
rect 2613 5234 2650 5237
rect 2613 5232 2655 5234
rect 2542 5221 2572 5224
rect 2551 5217 2558 5221
rect 2558 5216 2559 5217
rect 2517 5210 2527 5216
rect 2276 5202 2311 5210
rect 2276 5176 2277 5202
rect 2284 5176 2311 5202
rect 2219 5158 2249 5172
rect 2276 5168 2311 5176
rect 2313 5202 2354 5210
rect 2313 5176 2328 5202
rect 2335 5176 2354 5202
rect 2418 5198 2449 5210
rect 2464 5198 2567 5210
rect 2579 5200 2605 5226
rect 2620 5221 2650 5232
rect 2682 5228 2744 5244
rect 2682 5226 2728 5228
rect 2682 5210 2744 5226
rect 2756 5210 2762 5258
rect 2765 5250 2845 5258
rect 2765 5248 2784 5250
rect 2799 5248 2833 5250
rect 2765 5232 2845 5248
rect 2765 5210 2784 5232
rect 2799 5216 2829 5232
rect 2857 5226 2863 5300
rect 2866 5226 2885 5370
rect 2900 5226 2906 5370
rect 2915 5300 2928 5370
rect 2980 5366 3002 5370
rect 2973 5344 3002 5358
rect 3055 5344 3071 5358
rect 3109 5354 3115 5356
rect 3122 5354 3230 5370
rect 3237 5354 3243 5356
rect 3251 5354 3266 5370
rect 3332 5364 3351 5367
rect 2973 5342 3071 5344
rect 3098 5342 3266 5354
rect 3281 5344 3297 5358
rect 3332 5345 3354 5364
rect 3364 5358 3380 5359
rect 3363 5356 3380 5358
rect 3364 5351 3380 5356
rect 3354 5344 3360 5345
rect 3363 5344 3392 5351
rect 3281 5343 3392 5344
rect 3281 5342 3398 5343
rect 2957 5334 3008 5342
rect 3055 5334 3089 5342
rect 2957 5322 2982 5334
rect 2989 5322 3008 5334
rect 3062 5332 3089 5334
rect 3098 5332 3319 5342
rect 3354 5339 3360 5342
rect 3062 5328 3319 5332
rect 2957 5314 3008 5322
rect 3055 5314 3319 5328
rect 3363 5334 3398 5342
rect 2909 5266 2928 5300
rect 2973 5306 3002 5314
rect 2973 5300 2990 5306
rect 2973 5298 3007 5300
rect 3055 5298 3071 5314
rect 3072 5304 3280 5314
rect 3281 5304 3297 5314
rect 3345 5310 3360 5325
rect 3363 5322 3364 5334
rect 3371 5322 3398 5334
rect 3363 5314 3398 5322
rect 3363 5313 3392 5314
rect 3083 5300 3297 5304
rect 3098 5298 3297 5300
rect 3332 5300 3345 5310
rect 3363 5300 3380 5313
rect 3332 5298 3380 5300
rect 2974 5294 3007 5298
rect 2970 5292 3007 5294
rect 2970 5291 3037 5292
rect 2970 5286 3001 5291
rect 3007 5286 3037 5291
rect 2970 5282 3037 5286
rect 2943 5279 3037 5282
rect 2943 5272 2992 5279
rect 2943 5266 2973 5272
rect 2992 5267 2997 5272
rect 2909 5250 2989 5266
rect 3001 5258 3037 5279
rect 3098 5274 3287 5298
rect 3332 5297 3379 5298
rect 3345 5292 3379 5297
rect 3113 5271 3287 5274
rect 3106 5268 3287 5271
rect 3315 5291 3379 5292
rect 2909 5248 2928 5250
rect 2943 5248 2977 5250
rect 2909 5232 2989 5248
rect 2909 5226 2928 5232
rect 2625 5200 2728 5210
rect 2579 5198 2728 5200
rect 2749 5198 2784 5210
rect 2418 5196 2580 5198
rect 2430 5176 2449 5196
rect 2464 5194 2494 5196
rect 2313 5168 2354 5176
rect 2436 5172 2449 5176
rect 2501 5180 2580 5196
rect 2612 5196 2784 5198
rect 2612 5180 2691 5196
rect 2698 5194 2728 5196
rect 2276 5158 2305 5168
rect 2319 5158 2348 5168
rect 2363 5158 2393 5172
rect 2436 5158 2479 5172
rect 2501 5168 2691 5180
rect 2756 5176 2762 5196
rect 2486 5158 2516 5168
rect 2517 5158 2675 5168
rect 2679 5158 2709 5168
rect 2713 5158 2743 5172
rect 2771 5158 2784 5196
rect 2856 5210 2885 5226
rect 2899 5210 2928 5226
rect 2943 5216 2973 5232
rect 3001 5210 3007 5258
rect 3010 5252 3029 5258
rect 3044 5252 3074 5260
rect 3010 5244 3074 5252
rect 3010 5228 3090 5244
rect 3106 5237 3168 5268
rect 3184 5237 3246 5268
rect 3315 5266 3364 5291
rect 3379 5266 3409 5282
rect 3278 5252 3308 5260
rect 3315 5258 3425 5266
rect 3278 5244 3323 5252
rect 3010 5226 3029 5228
rect 3044 5226 3090 5228
rect 3010 5210 3090 5226
rect 3117 5224 3152 5237
rect 3193 5234 3230 5237
rect 3193 5232 3235 5234
rect 3122 5221 3152 5224
rect 3131 5217 3138 5221
rect 3138 5216 3139 5217
rect 3097 5210 3107 5216
rect 2856 5202 2891 5210
rect 2856 5176 2857 5202
rect 2864 5176 2891 5202
rect 2799 5158 2829 5172
rect 2856 5168 2891 5176
rect 2893 5202 2934 5210
rect 2893 5176 2908 5202
rect 2915 5176 2934 5202
rect 2998 5198 3029 5210
rect 3044 5198 3147 5210
rect 3159 5200 3185 5226
rect 3200 5221 3230 5232
rect 3262 5228 3324 5244
rect 3262 5226 3308 5228
rect 3262 5210 3324 5226
rect 3336 5210 3342 5258
rect 3345 5250 3425 5258
rect 3345 5248 3364 5250
rect 3379 5248 3413 5250
rect 3345 5232 3425 5248
rect 3345 5210 3364 5232
rect 3379 5216 3409 5232
rect 3437 5226 3443 5300
rect 3446 5226 3465 5370
rect 3480 5226 3486 5370
rect 3495 5300 3508 5370
rect 3560 5366 3582 5370
rect 3553 5344 3582 5358
rect 3635 5344 3651 5358
rect 3689 5354 3695 5356
rect 3702 5354 3810 5370
rect 3817 5354 3823 5356
rect 3831 5354 3846 5370
rect 3912 5364 3931 5367
rect 3553 5342 3651 5344
rect 3678 5342 3846 5354
rect 3861 5344 3877 5358
rect 3912 5345 3934 5364
rect 3944 5358 3960 5359
rect 3943 5356 3960 5358
rect 3944 5351 3960 5356
rect 3934 5344 3940 5345
rect 3943 5344 3972 5351
rect 3861 5343 3972 5344
rect 3861 5342 3978 5343
rect 3537 5334 3588 5342
rect 3635 5334 3669 5342
rect 3537 5322 3562 5334
rect 3569 5322 3588 5334
rect 3642 5332 3669 5334
rect 3678 5332 3899 5342
rect 3934 5339 3940 5342
rect 3642 5328 3899 5332
rect 3537 5314 3588 5322
rect 3635 5314 3899 5328
rect 3943 5334 3978 5342
rect 3489 5266 3508 5300
rect 3553 5306 3582 5314
rect 3553 5300 3570 5306
rect 3553 5298 3587 5300
rect 3635 5298 3651 5314
rect 3652 5304 3860 5314
rect 3861 5304 3877 5314
rect 3925 5310 3940 5325
rect 3943 5322 3944 5334
rect 3951 5322 3978 5334
rect 3943 5314 3978 5322
rect 3943 5313 3972 5314
rect 3663 5300 3877 5304
rect 3678 5298 3877 5300
rect 3912 5300 3925 5310
rect 3943 5300 3960 5313
rect 3912 5298 3960 5300
rect 3554 5294 3587 5298
rect 3550 5292 3587 5294
rect 3550 5291 3617 5292
rect 3550 5286 3581 5291
rect 3587 5286 3617 5291
rect 3550 5282 3617 5286
rect 3523 5279 3617 5282
rect 3523 5272 3572 5279
rect 3523 5266 3553 5272
rect 3572 5267 3577 5272
rect 3489 5250 3569 5266
rect 3581 5258 3617 5279
rect 3678 5274 3867 5298
rect 3912 5297 3959 5298
rect 3925 5292 3959 5297
rect 3693 5271 3867 5274
rect 3686 5268 3867 5271
rect 3895 5291 3959 5292
rect 3489 5248 3508 5250
rect 3523 5248 3557 5250
rect 3489 5232 3569 5248
rect 3489 5226 3508 5232
rect 3205 5200 3308 5210
rect 3159 5198 3308 5200
rect 3329 5198 3364 5210
rect 2998 5196 3160 5198
rect 3010 5176 3029 5196
rect 3044 5194 3074 5196
rect 2893 5168 2934 5176
rect 3016 5172 3029 5176
rect 3081 5180 3160 5196
rect 3192 5196 3364 5198
rect 3192 5180 3271 5196
rect 3278 5194 3308 5196
rect 2856 5158 2885 5168
rect 2899 5158 2928 5168
rect 2943 5158 2973 5172
rect 3016 5158 3059 5172
rect 3081 5168 3271 5180
rect 3336 5176 3342 5196
rect 3066 5158 3096 5168
rect 3097 5158 3255 5168
rect 3259 5158 3289 5168
rect 3293 5158 3323 5172
rect 3351 5158 3364 5196
rect 3436 5210 3465 5226
rect 3479 5210 3508 5226
rect 3523 5216 3553 5232
rect 3581 5210 3587 5258
rect 3590 5252 3609 5258
rect 3624 5252 3654 5260
rect 3590 5244 3654 5252
rect 3590 5228 3670 5244
rect 3686 5237 3748 5268
rect 3764 5237 3826 5268
rect 3895 5266 3944 5291
rect 3959 5266 3989 5282
rect 3858 5252 3888 5260
rect 3895 5258 4005 5266
rect 3858 5244 3903 5252
rect 3590 5226 3609 5228
rect 3624 5226 3670 5228
rect 3590 5210 3670 5226
rect 3697 5224 3732 5237
rect 3773 5234 3810 5237
rect 3773 5232 3815 5234
rect 3702 5221 3732 5224
rect 3711 5217 3718 5221
rect 3718 5216 3719 5217
rect 3677 5210 3687 5216
rect 3436 5202 3471 5210
rect 3436 5176 3437 5202
rect 3444 5176 3471 5202
rect 3379 5158 3409 5172
rect 3436 5168 3471 5176
rect 3473 5202 3514 5210
rect 3473 5176 3488 5202
rect 3495 5176 3514 5202
rect 3578 5198 3609 5210
rect 3624 5198 3727 5210
rect 3739 5200 3765 5226
rect 3780 5221 3810 5232
rect 3842 5228 3904 5244
rect 3842 5226 3888 5228
rect 3842 5210 3904 5226
rect 3916 5210 3922 5258
rect 3925 5250 4005 5258
rect 3925 5248 3944 5250
rect 3959 5248 3993 5250
rect 3925 5232 4005 5248
rect 3925 5210 3944 5232
rect 3959 5216 3989 5232
rect 4017 5226 4023 5300
rect 4026 5226 4045 5370
rect 4060 5226 4066 5370
rect 4075 5300 4088 5370
rect 4140 5366 4162 5370
rect 4133 5344 4162 5358
rect 4215 5344 4231 5358
rect 4269 5354 4275 5356
rect 4282 5354 4390 5370
rect 4397 5354 4403 5356
rect 4411 5354 4426 5370
rect 4492 5364 4511 5367
rect 4133 5342 4231 5344
rect 4258 5342 4426 5354
rect 4441 5344 4457 5358
rect 4492 5345 4514 5364
rect 4524 5358 4540 5359
rect 4523 5356 4540 5358
rect 4524 5351 4540 5356
rect 4514 5344 4520 5345
rect 4523 5344 4552 5351
rect 4441 5343 4552 5344
rect 4441 5342 4558 5343
rect 4117 5334 4168 5342
rect 4215 5334 4249 5342
rect 4117 5322 4142 5334
rect 4149 5322 4168 5334
rect 4222 5332 4249 5334
rect 4258 5332 4479 5342
rect 4514 5339 4520 5342
rect 4222 5328 4479 5332
rect 4117 5314 4168 5322
rect 4215 5314 4479 5328
rect 4523 5334 4558 5342
rect 4069 5266 4088 5300
rect 4133 5306 4162 5314
rect 4133 5300 4150 5306
rect 4133 5298 4167 5300
rect 4215 5298 4231 5314
rect 4232 5304 4440 5314
rect 4441 5304 4457 5314
rect 4505 5310 4520 5325
rect 4523 5322 4524 5334
rect 4531 5322 4558 5334
rect 4523 5314 4558 5322
rect 4523 5313 4552 5314
rect 4243 5300 4457 5304
rect 4258 5298 4457 5300
rect 4492 5300 4505 5310
rect 4523 5300 4540 5313
rect 4492 5298 4540 5300
rect 4134 5294 4167 5298
rect 4130 5292 4167 5294
rect 4130 5291 4197 5292
rect 4130 5286 4161 5291
rect 4167 5286 4197 5291
rect 4130 5282 4197 5286
rect 4103 5279 4197 5282
rect 4103 5272 4152 5279
rect 4103 5266 4133 5272
rect 4152 5267 4157 5272
rect 4069 5250 4149 5266
rect 4161 5258 4197 5279
rect 4258 5274 4447 5298
rect 4492 5297 4539 5298
rect 4505 5292 4539 5297
rect 4273 5271 4447 5274
rect 4266 5268 4447 5271
rect 4475 5291 4539 5292
rect 4069 5248 4088 5250
rect 4103 5248 4137 5250
rect 4069 5232 4149 5248
rect 4069 5226 4088 5232
rect 3785 5200 3888 5210
rect 3739 5198 3888 5200
rect 3909 5198 3944 5210
rect 3578 5196 3740 5198
rect 3590 5176 3609 5196
rect 3624 5194 3654 5196
rect 3473 5168 3514 5176
rect 3596 5172 3609 5176
rect 3661 5180 3740 5196
rect 3772 5196 3944 5198
rect 3772 5180 3851 5196
rect 3858 5194 3888 5196
rect 3436 5158 3465 5168
rect 3479 5158 3508 5168
rect 3523 5158 3553 5172
rect 3596 5158 3639 5172
rect 3661 5168 3851 5180
rect 3916 5176 3922 5196
rect 3646 5158 3676 5168
rect 3677 5158 3835 5168
rect 3839 5158 3869 5168
rect 3873 5158 3903 5172
rect 3931 5158 3944 5196
rect 4016 5210 4045 5226
rect 4059 5210 4088 5226
rect 4103 5216 4133 5232
rect 4161 5210 4167 5258
rect 4170 5252 4189 5258
rect 4204 5252 4234 5260
rect 4170 5244 4234 5252
rect 4170 5228 4250 5244
rect 4266 5237 4328 5268
rect 4344 5237 4406 5268
rect 4475 5266 4524 5291
rect 4539 5266 4569 5282
rect 4438 5252 4468 5260
rect 4475 5258 4585 5266
rect 4438 5244 4483 5252
rect 4170 5226 4189 5228
rect 4204 5226 4250 5228
rect 4170 5210 4250 5226
rect 4277 5224 4312 5237
rect 4353 5234 4390 5237
rect 4353 5232 4395 5234
rect 4282 5221 4312 5224
rect 4291 5217 4298 5221
rect 4298 5216 4299 5217
rect 4257 5210 4267 5216
rect 4016 5202 4051 5210
rect 4016 5176 4017 5202
rect 4024 5176 4051 5202
rect 3959 5158 3989 5172
rect 4016 5168 4051 5176
rect 4053 5202 4094 5210
rect 4053 5176 4068 5202
rect 4075 5176 4094 5202
rect 4158 5198 4189 5210
rect 4204 5198 4307 5210
rect 4319 5200 4345 5226
rect 4360 5221 4390 5232
rect 4422 5228 4484 5244
rect 4422 5226 4468 5228
rect 4422 5210 4484 5226
rect 4496 5210 4502 5258
rect 4505 5250 4585 5258
rect 4505 5248 4524 5250
rect 4539 5248 4573 5250
rect 4505 5232 4585 5248
rect 4505 5210 4524 5232
rect 4539 5216 4569 5232
rect 4597 5226 4603 5300
rect 4606 5226 4625 5370
rect 4640 5226 4646 5370
rect 4655 5300 4668 5370
rect 4720 5366 4742 5370
rect 4713 5344 4742 5358
rect 4795 5344 4811 5358
rect 4849 5354 4855 5356
rect 4862 5354 4970 5370
rect 4977 5354 4983 5356
rect 4991 5354 5006 5370
rect 5072 5364 5091 5367
rect 4713 5342 4811 5344
rect 4838 5342 5006 5354
rect 5021 5344 5037 5358
rect 5072 5345 5094 5364
rect 5104 5358 5120 5359
rect 5103 5356 5120 5358
rect 5104 5351 5120 5356
rect 5094 5344 5100 5345
rect 5103 5344 5132 5351
rect 5021 5343 5132 5344
rect 5021 5342 5138 5343
rect 4697 5334 4748 5342
rect 4795 5334 4829 5342
rect 4697 5322 4722 5334
rect 4729 5322 4748 5334
rect 4802 5332 4829 5334
rect 4838 5332 5059 5342
rect 5094 5339 5100 5342
rect 4802 5328 5059 5332
rect 4697 5314 4748 5322
rect 4795 5314 5059 5328
rect 5103 5334 5138 5342
rect 4649 5266 4668 5300
rect 4713 5306 4742 5314
rect 4713 5300 4730 5306
rect 4713 5298 4747 5300
rect 4795 5298 4811 5314
rect 4812 5304 5020 5314
rect 5021 5304 5037 5314
rect 5085 5310 5100 5325
rect 5103 5322 5104 5334
rect 5111 5322 5138 5334
rect 5103 5314 5138 5322
rect 5103 5313 5132 5314
rect 4823 5300 5037 5304
rect 4838 5298 5037 5300
rect 5072 5300 5085 5310
rect 5103 5300 5120 5313
rect 5072 5298 5120 5300
rect 4714 5294 4747 5298
rect 4710 5292 4747 5294
rect 4710 5291 4777 5292
rect 4710 5286 4741 5291
rect 4747 5286 4777 5291
rect 4710 5282 4777 5286
rect 4683 5279 4777 5282
rect 4683 5272 4732 5279
rect 4683 5266 4713 5272
rect 4732 5267 4737 5272
rect 4649 5250 4729 5266
rect 4741 5258 4777 5279
rect 4838 5274 5027 5298
rect 5072 5297 5119 5298
rect 5085 5292 5119 5297
rect 4853 5271 5027 5274
rect 4846 5268 5027 5271
rect 5055 5291 5119 5292
rect 4649 5248 4668 5250
rect 4683 5248 4717 5250
rect 4649 5232 4729 5248
rect 4649 5226 4668 5232
rect 4365 5200 4468 5210
rect 4319 5198 4468 5200
rect 4489 5198 4524 5210
rect 4158 5196 4320 5198
rect 4170 5176 4189 5196
rect 4204 5194 4234 5196
rect 4053 5168 4094 5176
rect 4176 5172 4189 5176
rect 4241 5180 4320 5196
rect 4352 5196 4524 5198
rect 4352 5180 4431 5196
rect 4438 5194 4468 5196
rect 4016 5158 4045 5168
rect 4059 5158 4088 5168
rect 4103 5158 4133 5172
rect 4176 5158 4219 5172
rect 4241 5168 4431 5180
rect 4496 5176 4502 5196
rect 4226 5158 4256 5168
rect 4257 5158 4415 5168
rect 4419 5158 4449 5168
rect 4453 5158 4483 5172
rect 4511 5158 4524 5196
rect 4596 5210 4625 5226
rect 4639 5210 4668 5226
rect 4683 5216 4713 5232
rect 4741 5210 4747 5258
rect 4750 5252 4769 5258
rect 4784 5252 4814 5260
rect 4750 5244 4814 5252
rect 4750 5228 4830 5244
rect 4846 5237 4908 5268
rect 4924 5237 4986 5268
rect 5055 5266 5104 5291
rect 5119 5266 5149 5282
rect 5018 5252 5048 5260
rect 5055 5258 5165 5266
rect 5018 5244 5063 5252
rect 4750 5226 4769 5228
rect 4784 5226 4830 5228
rect 4750 5210 4830 5226
rect 4857 5224 4892 5237
rect 4933 5234 4970 5237
rect 4933 5232 4975 5234
rect 4862 5221 4892 5224
rect 4871 5217 4878 5221
rect 4878 5216 4879 5217
rect 4837 5210 4847 5216
rect 4596 5202 4631 5210
rect 4596 5176 4597 5202
rect 4604 5176 4631 5202
rect 4539 5158 4569 5172
rect 4596 5168 4631 5176
rect 4633 5202 4674 5210
rect 4633 5176 4648 5202
rect 4655 5176 4674 5202
rect 4738 5198 4769 5210
rect 4784 5198 4887 5210
rect 4899 5200 4925 5226
rect 4940 5221 4970 5232
rect 5002 5228 5064 5244
rect 5002 5226 5048 5228
rect 5002 5210 5064 5226
rect 5076 5210 5082 5258
rect 5085 5250 5165 5258
rect 5085 5248 5104 5250
rect 5119 5248 5153 5250
rect 5085 5232 5165 5248
rect 5085 5210 5104 5232
rect 5119 5216 5149 5232
rect 5177 5226 5183 5300
rect 5186 5226 5205 5370
rect 5220 5226 5226 5370
rect 5235 5300 5248 5370
rect 5300 5366 5322 5370
rect 5293 5344 5322 5358
rect 5375 5344 5391 5358
rect 5429 5354 5435 5356
rect 5442 5354 5550 5370
rect 5557 5354 5563 5356
rect 5571 5354 5586 5370
rect 5652 5364 5671 5367
rect 5293 5342 5391 5344
rect 5418 5342 5586 5354
rect 5601 5344 5617 5358
rect 5652 5345 5674 5364
rect 5684 5358 5700 5359
rect 5683 5356 5700 5358
rect 5684 5351 5700 5356
rect 5674 5344 5680 5345
rect 5683 5344 5712 5351
rect 5601 5343 5712 5344
rect 5601 5342 5718 5343
rect 5277 5334 5328 5342
rect 5375 5334 5409 5342
rect 5277 5322 5302 5334
rect 5309 5322 5328 5334
rect 5382 5332 5409 5334
rect 5418 5332 5639 5342
rect 5674 5339 5680 5342
rect 5382 5328 5639 5332
rect 5277 5314 5328 5322
rect 5375 5314 5639 5328
rect 5683 5334 5718 5342
rect 5229 5266 5248 5300
rect 5293 5306 5322 5314
rect 5293 5300 5310 5306
rect 5293 5298 5327 5300
rect 5375 5298 5391 5314
rect 5392 5304 5600 5314
rect 5601 5304 5617 5314
rect 5665 5310 5680 5325
rect 5683 5322 5684 5334
rect 5691 5322 5718 5334
rect 5683 5314 5718 5322
rect 5683 5313 5712 5314
rect 5403 5300 5617 5304
rect 5418 5298 5617 5300
rect 5652 5300 5665 5310
rect 5683 5300 5700 5313
rect 5652 5298 5700 5300
rect 5294 5294 5327 5298
rect 5290 5292 5327 5294
rect 5290 5291 5357 5292
rect 5290 5286 5321 5291
rect 5327 5286 5357 5291
rect 5290 5282 5357 5286
rect 5263 5279 5357 5282
rect 5263 5272 5312 5279
rect 5263 5266 5293 5272
rect 5312 5267 5317 5272
rect 5229 5250 5309 5266
rect 5321 5258 5357 5279
rect 5418 5274 5607 5298
rect 5652 5297 5699 5298
rect 5665 5292 5699 5297
rect 5433 5271 5607 5274
rect 5426 5268 5607 5271
rect 5635 5291 5699 5292
rect 5229 5248 5248 5250
rect 5263 5248 5297 5250
rect 5229 5232 5309 5248
rect 5229 5226 5248 5232
rect 4945 5200 5048 5210
rect 4899 5198 5048 5200
rect 5069 5198 5104 5210
rect 4738 5196 4900 5198
rect 4750 5176 4769 5196
rect 4784 5194 4814 5196
rect 4633 5168 4674 5176
rect 4756 5172 4769 5176
rect 4821 5180 4900 5196
rect 4932 5196 5104 5198
rect 4932 5180 5011 5196
rect 5018 5194 5048 5196
rect 4596 5158 4625 5168
rect 4639 5158 4668 5168
rect 4683 5158 4713 5172
rect 4756 5158 4799 5172
rect 4821 5168 5011 5180
rect 5076 5176 5082 5196
rect 4806 5158 4836 5168
rect 4837 5158 4995 5168
rect 4999 5158 5029 5168
rect 5033 5158 5063 5172
rect 5091 5158 5104 5196
rect 5176 5210 5205 5226
rect 5219 5210 5248 5226
rect 5263 5216 5293 5232
rect 5321 5210 5327 5258
rect 5330 5252 5349 5258
rect 5364 5252 5394 5260
rect 5330 5244 5394 5252
rect 5330 5228 5410 5244
rect 5426 5237 5488 5268
rect 5504 5237 5566 5268
rect 5635 5266 5684 5291
rect 5699 5266 5729 5282
rect 5598 5252 5628 5260
rect 5635 5258 5745 5266
rect 5598 5244 5643 5252
rect 5330 5226 5349 5228
rect 5364 5226 5410 5228
rect 5330 5210 5410 5226
rect 5437 5224 5472 5237
rect 5513 5234 5550 5237
rect 5513 5232 5555 5234
rect 5442 5221 5472 5224
rect 5451 5217 5458 5221
rect 5458 5216 5459 5217
rect 5417 5210 5427 5216
rect 5176 5202 5211 5210
rect 5176 5176 5177 5202
rect 5184 5176 5211 5202
rect 5119 5158 5149 5172
rect 5176 5168 5211 5176
rect 5213 5202 5254 5210
rect 5213 5176 5228 5202
rect 5235 5176 5254 5202
rect 5318 5198 5349 5210
rect 5364 5198 5467 5210
rect 5479 5200 5505 5226
rect 5520 5221 5550 5232
rect 5582 5228 5644 5244
rect 5582 5226 5628 5228
rect 5582 5210 5644 5226
rect 5656 5210 5662 5258
rect 5665 5250 5745 5258
rect 5665 5248 5684 5250
rect 5699 5248 5733 5250
rect 5665 5232 5745 5248
rect 5665 5210 5684 5232
rect 5699 5216 5729 5232
rect 5757 5226 5763 5300
rect 5766 5226 5785 5370
rect 5800 5226 5806 5370
rect 5815 5300 5828 5370
rect 5880 5366 5902 5370
rect 5873 5344 5902 5358
rect 5955 5344 5971 5358
rect 6009 5354 6015 5356
rect 6022 5354 6130 5370
rect 6137 5354 6143 5356
rect 6151 5354 6166 5370
rect 6232 5364 6251 5367
rect 5873 5342 5971 5344
rect 5998 5342 6166 5354
rect 6181 5344 6197 5358
rect 6232 5345 6254 5364
rect 6264 5358 6280 5359
rect 6263 5356 6280 5358
rect 6264 5351 6280 5356
rect 6254 5344 6260 5345
rect 6263 5344 6292 5351
rect 6181 5343 6292 5344
rect 6181 5342 6298 5343
rect 5857 5334 5908 5342
rect 5955 5334 5989 5342
rect 5857 5322 5882 5334
rect 5889 5322 5908 5334
rect 5962 5332 5989 5334
rect 5998 5332 6219 5342
rect 6254 5339 6260 5342
rect 5962 5328 6219 5332
rect 5857 5314 5908 5322
rect 5955 5314 6219 5328
rect 6263 5334 6298 5342
rect 5809 5266 5828 5300
rect 5873 5306 5902 5314
rect 5873 5300 5890 5306
rect 5873 5298 5907 5300
rect 5955 5298 5971 5314
rect 5972 5304 6180 5314
rect 6181 5304 6197 5314
rect 6245 5310 6260 5325
rect 6263 5322 6264 5334
rect 6271 5322 6298 5334
rect 6263 5314 6298 5322
rect 6263 5313 6292 5314
rect 5983 5300 6197 5304
rect 5998 5298 6197 5300
rect 6232 5300 6245 5310
rect 6263 5300 6280 5313
rect 6232 5298 6280 5300
rect 5874 5294 5907 5298
rect 5870 5292 5907 5294
rect 5870 5291 5937 5292
rect 5870 5286 5901 5291
rect 5907 5286 5937 5291
rect 5870 5282 5937 5286
rect 5843 5279 5937 5282
rect 5843 5272 5892 5279
rect 5843 5266 5873 5272
rect 5892 5267 5897 5272
rect 5809 5250 5889 5266
rect 5901 5258 5937 5279
rect 5998 5274 6187 5298
rect 6232 5297 6279 5298
rect 6245 5292 6279 5297
rect 6013 5271 6187 5274
rect 6006 5268 6187 5271
rect 6215 5291 6279 5292
rect 5809 5248 5828 5250
rect 5843 5248 5877 5250
rect 5809 5232 5889 5248
rect 5809 5226 5828 5232
rect 5525 5200 5628 5210
rect 5479 5198 5628 5200
rect 5649 5198 5684 5210
rect 5318 5196 5480 5198
rect 5330 5176 5349 5196
rect 5364 5194 5394 5196
rect 5213 5168 5254 5176
rect 5336 5172 5349 5176
rect 5401 5180 5480 5196
rect 5512 5196 5684 5198
rect 5512 5180 5591 5196
rect 5598 5194 5628 5196
rect 5176 5158 5205 5168
rect 5219 5158 5248 5168
rect 5263 5158 5293 5172
rect 5336 5158 5379 5172
rect 5401 5168 5591 5180
rect 5656 5176 5662 5196
rect 5386 5158 5416 5168
rect 5417 5158 5575 5168
rect 5579 5158 5609 5168
rect 5613 5158 5643 5172
rect 5671 5158 5684 5196
rect 5756 5210 5785 5226
rect 5799 5210 5828 5226
rect 5843 5216 5873 5232
rect 5901 5210 5907 5258
rect 5910 5252 5929 5258
rect 5944 5252 5974 5260
rect 5910 5244 5974 5252
rect 5910 5228 5990 5244
rect 6006 5237 6068 5268
rect 6084 5237 6146 5268
rect 6215 5266 6264 5291
rect 6279 5266 6309 5282
rect 6178 5252 6208 5260
rect 6215 5258 6325 5266
rect 6178 5244 6223 5252
rect 5910 5226 5929 5228
rect 5944 5226 5990 5228
rect 5910 5210 5990 5226
rect 6017 5224 6052 5237
rect 6093 5234 6130 5237
rect 6093 5232 6135 5234
rect 6022 5221 6052 5224
rect 6031 5217 6038 5221
rect 6038 5216 6039 5217
rect 5997 5210 6007 5216
rect 5756 5202 5791 5210
rect 5756 5176 5757 5202
rect 5764 5176 5791 5202
rect 5699 5158 5729 5172
rect 5756 5168 5791 5176
rect 5793 5202 5834 5210
rect 5793 5176 5808 5202
rect 5815 5176 5834 5202
rect 5898 5198 5929 5210
rect 5944 5198 6047 5210
rect 6059 5200 6085 5226
rect 6100 5221 6130 5232
rect 6162 5228 6224 5244
rect 6162 5226 6208 5228
rect 6162 5210 6224 5226
rect 6236 5210 6242 5258
rect 6245 5250 6325 5258
rect 6245 5248 6264 5250
rect 6279 5248 6313 5250
rect 6245 5232 6325 5248
rect 6245 5210 6264 5232
rect 6279 5216 6309 5232
rect 6337 5226 6343 5300
rect 6346 5226 6365 5370
rect 6380 5226 6386 5370
rect 6395 5300 6408 5370
rect 6460 5366 6482 5370
rect 6453 5344 6482 5358
rect 6535 5344 6551 5358
rect 6589 5354 6595 5356
rect 6602 5354 6710 5370
rect 6717 5354 6723 5356
rect 6731 5354 6746 5370
rect 6812 5364 6831 5367
rect 6453 5342 6551 5344
rect 6578 5342 6746 5354
rect 6761 5344 6777 5358
rect 6812 5345 6834 5364
rect 6844 5358 6860 5359
rect 6843 5356 6860 5358
rect 6844 5351 6860 5356
rect 6834 5344 6840 5345
rect 6843 5344 6872 5351
rect 6761 5343 6872 5344
rect 6761 5342 6878 5343
rect 6437 5334 6488 5342
rect 6535 5334 6569 5342
rect 6437 5322 6462 5334
rect 6469 5322 6488 5334
rect 6542 5332 6569 5334
rect 6578 5332 6799 5342
rect 6834 5339 6840 5342
rect 6542 5328 6799 5332
rect 6437 5314 6488 5322
rect 6535 5314 6799 5328
rect 6843 5334 6878 5342
rect 6389 5266 6408 5300
rect 6453 5306 6482 5314
rect 6453 5300 6470 5306
rect 6453 5298 6487 5300
rect 6535 5298 6551 5314
rect 6552 5304 6760 5314
rect 6761 5304 6777 5314
rect 6825 5310 6840 5325
rect 6843 5322 6844 5334
rect 6851 5322 6878 5334
rect 6843 5314 6878 5322
rect 6843 5313 6872 5314
rect 6563 5300 6777 5304
rect 6578 5298 6777 5300
rect 6812 5300 6825 5310
rect 6843 5300 6860 5313
rect 6812 5298 6860 5300
rect 6454 5294 6487 5298
rect 6450 5292 6487 5294
rect 6450 5291 6517 5292
rect 6450 5286 6481 5291
rect 6487 5286 6517 5291
rect 6450 5282 6517 5286
rect 6423 5279 6517 5282
rect 6423 5272 6472 5279
rect 6423 5266 6453 5272
rect 6472 5267 6477 5272
rect 6389 5250 6469 5266
rect 6481 5258 6517 5279
rect 6578 5274 6767 5298
rect 6812 5297 6859 5298
rect 6825 5292 6859 5297
rect 6593 5271 6767 5274
rect 6586 5268 6767 5271
rect 6795 5291 6859 5292
rect 6389 5248 6408 5250
rect 6423 5248 6457 5250
rect 6389 5232 6469 5248
rect 6389 5226 6408 5232
rect 6105 5200 6208 5210
rect 6059 5198 6208 5200
rect 6229 5198 6264 5210
rect 5898 5196 6060 5198
rect 5910 5176 5929 5196
rect 5944 5194 5974 5196
rect 5793 5168 5834 5176
rect 5916 5172 5929 5176
rect 5981 5180 6060 5196
rect 6092 5196 6264 5198
rect 6092 5180 6171 5196
rect 6178 5194 6208 5196
rect 5756 5158 5785 5168
rect 5799 5158 5828 5168
rect 5843 5158 5873 5172
rect 5916 5158 5959 5172
rect 5981 5168 6171 5180
rect 6236 5176 6242 5196
rect 5966 5158 5996 5168
rect 5997 5158 6155 5168
rect 6159 5158 6189 5168
rect 6193 5158 6223 5172
rect 6251 5158 6264 5196
rect 6336 5210 6365 5226
rect 6379 5210 6408 5226
rect 6423 5216 6453 5232
rect 6481 5210 6487 5258
rect 6490 5252 6509 5258
rect 6524 5252 6554 5260
rect 6490 5244 6554 5252
rect 6490 5228 6570 5244
rect 6586 5237 6648 5268
rect 6664 5237 6726 5268
rect 6795 5266 6844 5291
rect 6859 5266 6889 5282
rect 6758 5252 6788 5260
rect 6795 5258 6905 5266
rect 6758 5244 6803 5252
rect 6490 5226 6509 5228
rect 6524 5226 6570 5228
rect 6490 5210 6570 5226
rect 6597 5224 6632 5237
rect 6673 5234 6710 5237
rect 6673 5232 6715 5234
rect 6602 5221 6632 5224
rect 6611 5217 6618 5221
rect 6618 5216 6619 5217
rect 6577 5210 6587 5216
rect 6336 5202 6371 5210
rect 6336 5176 6337 5202
rect 6344 5176 6371 5202
rect 6279 5158 6309 5172
rect 6336 5168 6371 5176
rect 6373 5202 6414 5210
rect 6373 5176 6388 5202
rect 6395 5176 6414 5202
rect 6478 5198 6509 5210
rect 6524 5198 6627 5210
rect 6639 5200 6665 5226
rect 6680 5221 6710 5232
rect 6742 5228 6804 5244
rect 6742 5226 6788 5228
rect 6742 5210 6804 5226
rect 6816 5210 6822 5258
rect 6825 5250 6905 5258
rect 6825 5248 6844 5250
rect 6859 5248 6893 5250
rect 6825 5232 6905 5248
rect 6825 5210 6844 5232
rect 6859 5216 6889 5232
rect 6917 5226 6923 5300
rect 6926 5226 6945 5370
rect 6960 5226 6966 5370
rect 6975 5300 6988 5370
rect 7040 5366 7062 5370
rect 7033 5344 7062 5358
rect 7115 5344 7131 5358
rect 7169 5354 7175 5356
rect 7182 5354 7290 5370
rect 7297 5354 7303 5356
rect 7311 5354 7326 5370
rect 7392 5364 7411 5367
rect 7033 5342 7131 5344
rect 7158 5342 7326 5354
rect 7341 5344 7357 5358
rect 7392 5345 7414 5364
rect 7424 5358 7440 5359
rect 7423 5356 7440 5358
rect 7424 5351 7440 5356
rect 7414 5344 7420 5345
rect 7423 5344 7452 5351
rect 7341 5343 7452 5344
rect 7341 5342 7458 5343
rect 7017 5334 7068 5342
rect 7115 5334 7149 5342
rect 7017 5322 7042 5334
rect 7049 5322 7068 5334
rect 7122 5332 7149 5334
rect 7158 5332 7379 5342
rect 7414 5339 7420 5342
rect 7122 5328 7379 5332
rect 7017 5314 7068 5322
rect 7115 5314 7379 5328
rect 7423 5334 7458 5342
rect 6969 5266 6988 5300
rect 7033 5306 7062 5314
rect 7033 5300 7050 5306
rect 7033 5298 7067 5300
rect 7115 5298 7131 5314
rect 7132 5304 7340 5314
rect 7341 5304 7357 5314
rect 7405 5310 7420 5325
rect 7423 5322 7424 5334
rect 7431 5322 7458 5334
rect 7423 5314 7458 5322
rect 7423 5313 7452 5314
rect 7143 5300 7357 5304
rect 7158 5298 7357 5300
rect 7392 5300 7405 5310
rect 7423 5300 7440 5313
rect 7392 5298 7440 5300
rect 7034 5294 7067 5298
rect 7030 5292 7067 5294
rect 7030 5291 7097 5292
rect 7030 5286 7061 5291
rect 7067 5286 7097 5291
rect 7030 5282 7097 5286
rect 7003 5279 7097 5282
rect 7003 5272 7052 5279
rect 7003 5266 7033 5272
rect 7052 5267 7057 5272
rect 6969 5250 7049 5266
rect 7061 5258 7097 5279
rect 7158 5274 7347 5298
rect 7392 5297 7439 5298
rect 7405 5292 7439 5297
rect 7173 5271 7347 5274
rect 7166 5268 7347 5271
rect 7375 5291 7439 5292
rect 6969 5248 6988 5250
rect 7003 5248 7037 5250
rect 6969 5232 7049 5248
rect 6969 5226 6988 5232
rect 6685 5200 6788 5210
rect 6639 5198 6788 5200
rect 6809 5198 6844 5210
rect 6478 5196 6640 5198
rect 6490 5176 6509 5196
rect 6524 5194 6554 5196
rect 6373 5168 6414 5176
rect 6496 5172 6509 5176
rect 6561 5180 6640 5196
rect 6672 5196 6844 5198
rect 6672 5180 6751 5196
rect 6758 5194 6788 5196
rect 6336 5158 6365 5168
rect 6379 5158 6408 5168
rect 6423 5158 6453 5172
rect 6496 5158 6539 5172
rect 6561 5168 6751 5180
rect 6816 5176 6822 5196
rect 6546 5158 6576 5168
rect 6577 5158 6735 5168
rect 6739 5158 6769 5168
rect 6773 5158 6803 5172
rect 6831 5158 6844 5196
rect 6916 5210 6945 5226
rect 6959 5210 6988 5226
rect 7003 5216 7033 5232
rect 7061 5210 7067 5258
rect 7070 5252 7089 5258
rect 7104 5252 7134 5260
rect 7070 5244 7134 5252
rect 7070 5228 7150 5244
rect 7166 5237 7228 5268
rect 7244 5237 7306 5268
rect 7375 5266 7424 5291
rect 7439 5266 7469 5282
rect 7338 5252 7368 5260
rect 7375 5258 7485 5266
rect 7338 5244 7383 5252
rect 7070 5226 7089 5228
rect 7104 5226 7150 5228
rect 7070 5210 7150 5226
rect 7177 5224 7212 5237
rect 7253 5234 7290 5237
rect 7253 5232 7295 5234
rect 7182 5221 7212 5224
rect 7191 5217 7198 5221
rect 7198 5216 7199 5217
rect 7157 5210 7167 5216
rect 6916 5202 6951 5210
rect 6916 5176 6917 5202
rect 6924 5176 6951 5202
rect 6859 5158 6889 5172
rect 6916 5168 6951 5176
rect 6953 5202 6994 5210
rect 6953 5176 6968 5202
rect 6975 5176 6994 5202
rect 7058 5198 7089 5210
rect 7104 5198 7207 5210
rect 7219 5200 7245 5226
rect 7260 5221 7290 5232
rect 7322 5228 7384 5244
rect 7322 5226 7368 5228
rect 7322 5210 7384 5226
rect 7396 5210 7402 5258
rect 7405 5250 7485 5258
rect 7405 5248 7424 5250
rect 7439 5248 7473 5250
rect 7405 5232 7485 5248
rect 7405 5210 7424 5232
rect 7439 5216 7469 5232
rect 7497 5226 7503 5300
rect 7506 5226 7525 5370
rect 7540 5226 7546 5370
rect 7555 5300 7568 5370
rect 7620 5366 7642 5370
rect 7613 5344 7642 5358
rect 7695 5344 7711 5358
rect 7749 5354 7755 5356
rect 7762 5354 7870 5370
rect 7877 5354 7883 5356
rect 7891 5354 7906 5370
rect 7972 5364 7991 5367
rect 7613 5342 7711 5344
rect 7738 5342 7906 5354
rect 7921 5344 7937 5358
rect 7972 5345 7994 5364
rect 8004 5358 8020 5359
rect 8003 5356 8020 5358
rect 8004 5351 8020 5356
rect 7994 5344 8000 5345
rect 8003 5344 8032 5351
rect 7921 5343 8032 5344
rect 7921 5342 8038 5343
rect 7597 5334 7648 5342
rect 7695 5334 7729 5342
rect 7597 5322 7622 5334
rect 7629 5322 7648 5334
rect 7702 5332 7729 5334
rect 7738 5332 7959 5342
rect 7994 5339 8000 5342
rect 7702 5328 7959 5332
rect 7597 5314 7648 5322
rect 7695 5314 7959 5328
rect 8003 5334 8038 5342
rect 7549 5266 7568 5300
rect 7613 5306 7642 5314
rect 7613 5300 7630 5306
rect 7613 5298 7647 5300
rect 7695 5298 7711 5314
rect 7712 5304 7920 5314
rect 7921 5304 7937 5314
rect 7985 5310 8000 5325
rect 8003 5322 8004 5334
rect 8011 5322 8038 5334
rect 8003 5314 8038 5322
rect 8003 5313 8032 5314
rect 7723 5300 7937 5304
rect 7738 5298 7937 5300
rect 7972 5300 7985 5310
rect 8003 5300 8020 5313
rect 7972 5298 8020 5300
rect 7614 5294 7647 5298
rect 7610 5292 7647 5294
rect 7610 5291 7677 5292
rect 7610 5286 7641 5291
rect 7647 5286 7677 5291
rect 7610 5282 7677 5286
rect 7583 5279 7677 5282
rect 7583 5272 7632 5279
rect 7583 5266 7613 5272
rect 7632 5267 7637 5272
rect 7549 5250 7629 5266
rect 7641 5258 7677 5279
rect 7738 5274 7927 5298
rect 7972 5297 8019 5298
rect 7985 5292 8019 5297
rect 7753 5271 7927 5274
rect 7746 5268 7927 5271
rect 7955 5291 8019 5292
rect 7549 5248 7568 5250
rect 7583 5248 7617 5250
rect 7549 5232 7629 5248
rect 7549 5226 7568 5232
rect 7265 5200 7368 5210
rect 7219 5198 7368 5200
rect 7389 5198 7424 5210
rect 7058 5196 7220 5198
rect 7070 5176 7089 5196
rect 7104 5194 7134 5196
rect 6953 5168 6994 5176
rect 7076 5172 7089 5176
rect 7141 5180 7220 5196
rect 7252 5196 7424 5198
rect 7252 5180 7331 5196
rect 7338 5194 7368 5196
rect 6916 5158 6945 5168
rect 6959 5158 6988 5168
rect 7003 5158 7033 5172
rect 7076 5158 7119 5172
rect 7141 5168 7331 5180
rect 7396 5176 7402 5196
rect 7126 5158 7156 5168
rect 7157 5158 7315 5168
rect 7319 5158 7349 5168
rect 7353 5158 7383 5172
rect 7411 5158 7424 5196
rect 7496 5210 7525 5226
rect 7539 5210 7568 5226
rect 7583 5216 7613 5232
rect 7641 5210 7647 5258
rect 7650 5252 7669 5258
rect 7684 5252 7714 5260
rect 7650 5244 7714 5252
rect 7650 5228 7730 5244
rect 7746 5237 7808 5268
rect 7824 5237 7886 5268
rect 7955 5266 8004 5291
rect 8019 5266 8049 5282
rect 7918 5252 7948 5260
rect 7955 5258 8065 5266
rect 7918 5244 7963 5252
rect 7650 5226 7669 5228
rect 7684 5226 7730 5228
rect 7650 5210 7730 5226
rect 7757 5224 7792 5237
rect 7833 5234 7870 5237
rect 7833 5232 7875 5234
rect 7762 5221 7792 5224
rect 7771 5217 7778 5221
rect 7778 5216 7779 5217
rect 7737 5210 7747 5216
rect 7496 5202 7531 5210
rect 7496 5176 7497 5202
rect 7504 5176 7531 5202
rect 7439 5158 7469 5172
rect 7496 5168 7531 5176
rect 7533 5202 7574 5210
rect 7533 5176 7548 5202
rect 7555 5176 7574 5202
rect 7638 5198 7669 5210
rect 7684 5198 7787 5210
rect 7799 5200 7825 5226
rect 7840 5221 7870 5232
rect 7902 5228 7964 5244
rect 7902 5226 7948 5228
rect 7902 5210 7964 5226
rect 7976 5210 7982 5258
rect 7985 5250 8065 5258
rect 7985 5248 8004 5250
rect 8019 5248 8053 5250
rect 7985 5232 8065 5248
rect 7985 5210 8004 5232
rect 8019 5216 8049 5232
rect 8077 5226 8083 5300
rect 8086 5226 8105 5370
rect 8120 5226 8126 5370
rect 8135 5300 8148 5370
rect 8200 5366 8222 5370
rect 8193 5344 8222 5358
rect 8275 5344 8291 5358
rect 8329 5354 8335 5356
rect 8342 5354 8450 5370
rect 8457 5354 8463 5356
rect 8471 5354 8486 5370
rect 8552 5364 8571 5367
rect 8193 5342 8291 5344
rect 8318 5342 8486 5354
rect 8501 5344 8517 5358
rect 8552 5345 8574 5364
rect 8584 5358 8600 5359
rect 8583 5356 8600 5358
rect 8584 5351 8600 5356
rect 8574 5344 8580 5345
rect 8583 5344 8612 5351
rect 8501 5343 8612 5344
rect 8501 5342 8618 5343
rect 8177 5334 8228 5342
rect 8275 5334 8309 5342
rect 8177 5322 8202 5334
rect 8209 5322 8228 5334
rect 8282 5332 8309 5334
rect 8318 5332 8539 5342
rect 8574 5339 8580 5342
rect 8282 5328 8539 5332
rect 8177 5314 8228 5322
rect 8275 5314 8539 5328
rect 8583 5334 8618 5342
rect 8129 5266 8148 5300
rect 8193 5306 8222 5314
rect 8193 5300 8210 5306
rect 8193 5298 8227 5300
rect 8275 5298 8291 5314
rect 8292 5304 8500 5314
rect 8501 5304 8517 5314
rect 8565 5310 8580 5325
rect 8583 5322 8584 5334
rect 8591 5322 8618 5334
rect 8583 5314 8618 5322
rect 8583 5313 8612 5314
rect 8303 5300 8517 5304
rect 8318 5298 8517 5300
rect 8552 5300 8565 5310
rect 8583 5300 8600 5313
rect 8552 5298 8600 5300
rect 8194 5294 8227 5298
rect 8190 5292 8227 5294
rect 8190 5291 8257 5292
rect 8190 5286 8221 5291
rect 8227 5286 8257 5291
rect 8190 5282 8257 5286
rect 8163 5279 8257 5282
rect 8163 5272 8212 5279
rect 8163 5266 8193 5272
rect 8212 5267 8217 5272
rect 8129 5250 8209 5266
rect 8221 5258 8257 5279
rect 8318 5274 8507 5298
rect 8552 5297 8599 5298
rect 8565 5292 8599 5297
rect 8333 5271 8507 5274
rect 8326 5268 8507 5271
rect 8535 5291 8599 5292
rect 8129 5248 8148 5250
rect 8163 5248 8197 5250
rect 8129 5232 8209 5248
rect 8129 5226 8148 5232
rect 7845 5200 7948 5210
rect 7799 5198 7948 5200
rect 7969 5198 8004 5210
rect 7638 5196 7800 5198
rect 7650 5176 7669 5196
rect 7684 5194 7714 5196
rect 7533 5168 7574 5176
rect 7656 5172 7669 5176
rect 7721 5180 7800 5196
rect 7832 5196 8004 5198
rect 7832 5180 7911 5196
rect 7918 5194 7948 5196
rect 7496 5158 7525 5168
rect 7539 5158 7568 5168
rect 7583 5158 7613 5172
rect 7656 5158 7699 5172
rect 7721 5168 7911 5180
rect 7976 5176 7982 5196
rect 7706 5158 7736 5168
rect 7737 5158 7895 5168
rect 7899 5158 7929 5168
rect 7933 5158 7963 5172
rect 7991 5158 8004 5196
rect 8076 5210 8105 5226
rect 8119 5210 8148 5226
rect 8163 5216 8193 5232
rect 8221 5210 8227 5258
rect 8230 5252 8249 5258
rect 8264 5252 8294 5260
rect 8230 5244 8294 5252
rect 8230 5228 8310 5244
rect 8326 5237 8388 5268
rect 8404 5237 8466 5268
rect 8535 5266 8584 5291
rect 8599 5266 8629 5282
rect 8498 5252 8528 5260
rect 8535 5258 8645 5266
rect 8498 5244 8543 5252
rect 8230 5226 8249 5228
rect 8264 5226 8310 5228
rect 8230 5210 8310 5226
rect 8337 5224 8372 5237
rect 8413 5234 8450 5237
rect 8413 5232 8455 5234
rect 8342 5221 8372 5224
rect 8351 5217 8358 5221
rect 8358 5216 8359 5217
rect 8317 5210 8327 5216
rect 8076 5202 8111 5210
rect 8076 5176 8077 5202
rect 8084 5176 8111 5202
rect 8019 5158 8049 5172
rect 8076 5168 8111 5176
rect 8113 5202 8154 5210
rect 8113 5176 8128 5202
rect 8135 5176 8154 5202
rect 8218 5198 8249 5210
rect 8264 5198 8367 5210
rect 8379 5200 8405 5226
rect 8420 5221 8450 5232
rect 8482 5228 8544 5244
rect 8482 5226 8528 5228
rect 8482 5210 8544 5226
rect 8556 5210 8562 5258
rect 8565 5250 8645 5258
rect 8565 5248 8584 5250
rect 8599 5248 8633 5250
rect 8565 5232 8645 5248
rect 8565 5210 8584 5232
rect 8599 5216 8629 5232
rect 8657 5226 8663 5300
rect 8666 5226 8685 5370
rect 8700 5226 8706 5370
rect 8715 5300 8728 5370
rect 8780 5366 8802 5370
rect 8773 5344 8802 5358
rect 8855 5344 8871 5358
rect 8909 5354 8915 5356
rect 8922 5354 9030 5370
rect 9037 5354 9043 5356
rect 9051 5354 9066 5370
rect 9132 5364 9151 5367
rect 8773 5342 8871 5344
rect 8898 5342 9066 5354
rect 9081 5344 9097 5358
rect 9132 5345 9154 5364
rect 9164 5358 9180 5359
rect 9163 5356 9180 5358
rect 9164 5351 9180 5356
rect 9154 5344 9160 5345
rect 9163 5344 9192 5351
rect 9081 5343 9192 5344
rect 9081 5342 9198 5343
rect 8757 5334 8808 5342
rect 8855 5334 8889 5342
rect 8757 5322 8782 5334
rect 8789 5322 8808 5334
rect 8862 5332 8889 5334
rect 8898 5332 9119 5342
rect 9154 5339 9160 5342
rect 8862 5328 9119 5332
rect 8757 5314 8808 5322
rect 8855 5314 9119 5328
rect 9163 5334 9198 5342
rect 8709 5266 8728 5300
rect 8773 5306 8802 5314
rect 8773 5300 8790 5306
rect 8773 5298 8807 5300
rect 8855 5298 8871 5314
rect 8872 5304 9080 5314
rect 9081 5304 9097 5314
rect 9145 5310 9160 5325
rect 9163 5322 9164 5334
rect 9171 5322 9198 5334
rect 9163 5314 9198 5322
rect 9163 5313 9192 5314
rect 8883 5300 9097 5304
rect 8898 5298 9097 5300
rect 9132 5300 9145 5310
rect 9163 5300 9180 5313
rect 9132 5298 9180 5300
rect 8774 5294 8807 5298
rect 8770 5292 8807 5294
rect 8770 5291 8837 5292
rect 8770 5286 8801 5291
rect 8807 5286 8837 5291
rect 8770 5282 8837 5286
rect 8743 5279 8837 5282
rect 8743 5272 8792 5279
rect 8743 5266 8773 5272
rect 8792 5267 8797 5272
rect 8709 5250 8789 5266
rect 8801 5258 8837 5279
rect 8898 5274 9087 5298
rect 9132 5297 9179 5298
rect 9145 5292 9179 5297
rect 8913 5271 9087 5274
rect 8906 5268 9087 5271
rect 9115 5291 9179 5292
rect 8709 5248 8728 5250
rect 8743 5248 8777 5250
rect 8709 5232 8789 5248
rect 8709 5226 8728 5232
rect 8425 5200 8528 5210
rect 8379 5198 8528 5200
rect 8549 5198 8584 5210
rect 8218 5196 8380 5198
rect 8230 5176 8249 5196
rect 8264 5194 8294 5196
rect 8113 5168 8154 5176
rect 8236 5172 8249 5176
rect 8301 5180 8380 5196
rect 8412 5196 8584 5198
rect 8412 5180 8491 5196
rect 8498 5194 8528 5196
rect 8076 5158 8105 5168
rect 8119 5158 8148 5168
rect 8163 5158 8193 5172
rect 8236 5158 8279 5172
rect 8301 5168 8491 5180
rect 8556 5176 8562 5196
rect 8286 5158 8316 5168
rect 8317 5158 8475 5168
rect 8479 5158 8509 5168
rect 8513 5158 8543 5172
rect 8571 5158 8584 5196
rect 8656 5210 8685 5226
rect 8699 5210 8728 5226
rect 8743 5216 8773 5232
rect 8801 5210 8807 5258
rect 8810 5252 8829 5258
rect 8844 5252 8874 5260
rect 8810 5244 8874 5252
rect 8810 5228 8890 5244
rect 8906 5237 8968 5268
rect 8984 5237 9046 5268
rect 9115 5266 9164 5291
rect 9179 5266 9209 5282
rect 9078 5252 9108 5260
rect 9115 5258 9225 5266
rect 9078 5244 9123 5252
rect 8810 5226 8829 5228
rect 8844 5226 8890 5228
rect 8810 5210 8890 5226
rect 8917 5224 8952 5237
rect 8993 5234 9030 5237
rect 8993 5232 9035 5234
rect 8922 5221 8952 5224
rect 8931 5217 8938 5221
rect 8938 5216 8939 5217
rect 8897 5210 8907 5216
rect 8656 5202 8691 5210
rect 8656 5176 8657 5202
rect 8664 5176 8691 5202
rect 8599 5158 8629 5172
rect 8656 5168 8691 5176
rect 8693 5202 8734 5210
rect 8693 5176 8708 5202
rect 8715 5176 8734 5202
rect 8798 5198 8829 5210
rect 8844 5198 8947 5210
rect 8959 5200 8985 5226
rect 9000 5221 9030 5232
rect 9062 5228 9124 5244
rect 9062 5226 9108 5228
rect 9062 5210 9124 5226
rect 9136 5210 9142 5258
rect 9145 5250 9225 5258
rect 9145 5248 9164 5250
rect 9179 5248 9213 5250
rect 9145 5232 9225 5248
rect 9145 5210 9164 5232
rect 9179 5216 9209 5232
rect 9237 5226 9243 5300
rect 9246 5226 9265 5370
rect 9280 5226 9286 5370
rect 9295 5300 9308 5370
rect 9360 5366 9382 5370
rect 9353 5344 9382 5358
rect 9435 5344 9451 5358
rect 9489 5354 9495 5356
rect 9502 5354 9610 5370
rect 9617 5354 9623 5356
rect 9631 5354 9646 5370
rect 9712 5364 9731 5367
rect 9353 5342 9451 5344
rect 9478 5342 9646 5354
rect 9661 5344 9677 5358
rect 9712 5345 9734 5364
rect 9744 5358 9760 5359
rect 9743 5356 9760 5358
rect 9744 5351 9760 5356
rect 9734 5344 9740 5345
rect 9743 5344 9772 5351
rect 9661 5343 9772 5344
rect 9661 5342 9778 5343
rect 9337 5334 9388 5342
rect 9435 5334 9469 5342
rect 9337 5322 9362 5334
rect 9369 5322 9388 5334
rect 9442 5332 9469 5334
rect 9478 5332 9699 5342
rect 9734 5339 9740 5342
rect 9442 5328 9699 5332
rect 9337 5314 9388 5322
rect 9435 5314 9699 5328
rect 9743 5334 9778 5342
rect 9289 5266 9308 5300
rect 9353 5306 9382 5314
rect 9353 5300 9370 5306
rect 9353 5298 9387 5300
rect 9435 5298 9451 5314
rect 9452 5304 9660 5314
rect 9661 5304 9677 5314
rect 9725 5310 9740 5325
rect 9743 5322 9744 5334
rect 9751 5322 9778 5334
rect 9743 5314 9778 5322
rect 9743 5313 9772 5314
rect 9463 5300 9677 5304
rect 9478 5298 9677 5300
rect 9712 5300 9725 5310
rect 9743 5300 9760 5313
rect 9712 5298 9760 5300
rect 9354 5294 9387 5298
rect 9350 5292 9387 5294
rect 9350 5291 9417 5292
rect 9350 5286 9381 5291
rect 9387 5286 9417 5291
rect 9350 5282 9417 5286
rect 9323 5279 9417 5282
rect 9323 5272 9372 5279
rect 9323 5266 9353 5272
rect 9372 5267 9377 5272
rect 9289 5250 9369 5266
rect 9381 5258 9417 5279
rect 9478 5274 9667 5298
rect 9712 5297 9759 5298
rect 9725 5292 9759 5297
rect 9493 5271 9667 5274
rect 9486 5268 9667 5271
rect 9695 5291 9759 5292
rect 9289 5248 9308 5250
rect 9323 5248 9357 5250
rect 9289 5232 9369 5248
rect 9289 5226 9308 5232
rect 9005 5200 9108 5210
rect 8959 5198 9108 5200
rect 9129 5198 9164 5210
rect 8798 5196 8960 5198
rect 8810 5176 8829 5196
rect 8844 5194 8874 5196
rect 8693 5168 8734 5176
rect 8816 5172 8829 5176
rect 8881 5180 8960 5196
rect 8992 5196 9164 5198
rect 8992 5180 9071 5196
rect 9078 5194 9108 5196
rect 8656 5158 8685 5168
rect 8699 5158 8728 5168
rect 8743 5158 8773 5172
rect 8816 5158 8859 5172
rect 8881 5168 9071 5180
rect 9136 5176 9142 5196
rect 8866 5158 8896 5168
rect 8897 5158 9055 5168
rect 9059 5158 9089 5168
rect 9093 5158 9123 5172
rect 9151 5158 9164 5196
rect 9236 5210 9265 5226
rect 9279 5210 9308 5226
rect 9323 5216 9353 5232
rect 9381 5210 9387 5258
rect 9390 5252 9409 5258
rect 9424 5252 9454 5260
rect 9390 5244 9454 5252
rect 9390 5228 9470 5244
rect 9486 5237 9548 5268
rect 9564 5237 9626 5268
rect 9695 5266 9744 5291
rect 9759 5266 9789 5282
rect 9658 5252 9688 5260
rect 9695 5258 9805 5266
rect 9658 5244 9703 5252
rect 9390 5226 9409 5228
rect 9424 5226 9470 5228
rect 9390 5210 9470 5226
rect 9497 5224 9532 5237
rect 9573 5234 9610 5237
rect 9573 5232 9615 5234
rect 9502 5221 9532 5224
rect 9511 5217 9518 5221
rect 9518 5216 9519 5217
rect 9477 5210 9487 5216
rect 9236 5202 9271 5210
rect 9236 5176 9237 5202
rect 9244 5176 9271 5202
rect 9179 5158 9209 5172
rect 9236 5168 9271 5176
rect 9273 5202 9314 5210
rect 9273 5176 9288 5202
rect 9295 5176 9314 5202
rect 9378 5198 9409 5210
rect 9424 5198 9527 5210
rect 9539 5200 9565 5226
rect 9580 5221 9610 5232
rect 9642 5228 9704 5244
rect 9642 5226 9688 5228
rect 9642 5210 9704 5226
rect 9716 5210 9722 5258
rect 9725 5250 9805 5258
rect 9725 5248 9744 5250
rect 9759 5248 9793 5250
rect 9725 5232 9805 5248
rect 9725 5210 9744 5232
rect 9759 5216 9789 5232
rect 9817 5226 9823 5300
rect 9826 5226 9845 5370
rect 9860 5226 9866 5370
rect 9875 5300 9888 5370
rect 9940 5366 9962 5370
rect 9933 5344 9962 5358
rect 10015 5344 10031 5358
rect 10069 5354 10075 5356
rect 10082 5354 10190 5370
rect 10197 5354 10203 5356
rect 10211 5354 10226 5370
rect 10292 5364 10311 5367
rect 9933 5342 10031 5344
rect 10058 5342 10226 5354
rect 10241 5344 10257 5358
rect 10292 5345 10314 5364
rect 10324 5358 10340 5359
rect 10323 5356 10340 5358
rect 10324 5351 10340 5356
rect 10314 5344 10320 5345
rect 10323 5344 10352 5351
rect 10241 5343 10352 5344
rect 10241 5342 10358 5343
rect 9917 5334 9968 5342
rect 10015 5334 10049 5342
rect 9917 5322 9942 5334
rect 9949 5322 9968 5334
rect 10022 5332 10049 5334
rect 10058 5332 10279 5342
rect 10314 5339 10320 5342
rect 10022 5328 10279 5332
rect 9917 5314 9968 5322
rect 10015 5314 10279 5328
rect 10323 5334 10358 5342
rect 9869 5266 9888 5300
rect 9933 5306 9962 5314
rect 9933 5300 9950 5306
rect 9933 5298 9967 5300
rect 10015 5298 10031 5314
rect 10032 5304 10240 5314
rect 10241 5304 10257 5314
rect 10305 5310 10320 5325
rect 10323 5322 10324 5334
rect 10331 5322 10358 5334
rect 10323 5314 10358 5322
rect 10323 5313 10352 5314
rect 10043 5300 10257 5304
rect 10058 5298 10257 5300
rect 10292 5300 10305 5310
rect 10323 5300 10340 5313
rect 10292 5298 10340 5300
rect 9934 5294 9967 5298
rect 9930 5292 9967 5294
rect 9930 5291 9997 5292
rect 9930 5286 9961 5291
rect 9967 5286 9997 5291
rect 9930 5282 9997 5286
rect 9903 5279 9997 5282
rect 9903 5272 9952 5279
rect 9903 5266 9933 5272
rect 9952 5267 9957 5272
rect 9869 5250 9949 5266
rect 9961 5258 9997 5279
rect 10058 5274 10247 5298
rect 10292 5297 10339 5298
rect 10305 5292 10339 5297
rect 10073 5271 10247 5274
rect 10066 5268 10247 5271
rect 10275 5291 10339 5292
rect 9869 5248 9888 5250
rect 9903 5248 9937 5250
rect 9869 5232 9949 5248
rect 9869 5226 9888 5232
rect 9585 5200 9688 5210
rect 9539 5198 9688 5200
rect 9709 5198 9744 5210
rect 9378 5196 9540 5198
rect 9390 5176 9409 5196
rect 9424 5194 9454 5196
rect 9273 5168 9314 5176
rect 9396 5172 9409 5176
rect 9461 5180 9540 5196
rect 9572 5196 9744 5198
rect 9572 5180 9651 5196
rect 9658 5194 9688 5196
rect 9236 5158 9265 5168
rect 9279 5158 9308 5168
rect 9323 5158 9353 5172
rect 9396 5158 9439 5172
rect 9461 5168 9651 5180
rect 9716 5176 9722 5196
rect 9446 5158 9476 5168
rect 9477 5158 9635 5168
rect 9639 5158 9669 5168
rect 9673 5158 9703 5172
rect 9731 5158 9744 5196
rect 9816 5210 9845 5226
rect 9859 5210 9888 5226
rect 9903 5216 9933 5232
rect 9961 5210 9967 5258
rect 9970 5252 9989 5258
rect 10004 5252 10034 5260
rect 9970 5244 10034 5252
rect 9970 5228 10050 5244
rect 10066 5237 10128 5268
rect 10144 5237 10206 5268
rect 10275 5266 10324 5291
rect 10339 5266 10369 5282
rect 10238 5252 10268 5260
rect 10275 5258 10385 5266
rect 10238 5244 10283 5252
rect 9970 5226 9989 5228
rect 10004 5226 10050 5228
rect 9970 5210 10050 5226
rect 10077 5224 10112 5237
rect 10153 5234 10190 5237
rect 10153 5232 10195 5234
rect 10082 5221 10112 5224
rect 10091 5217 10098 5221
rect 10098 5216 10099 5217
rect 10057 5210 10067 5216
rect 9816 5202 9851 5210
rect 9816 5176 9817 5202
rect 9824 5176 9851 5202
rect 9759 5158 9789 5172
rect 9816 5168 9851 5176
rect 9853 5202 9894 5210
rect 9853 5176 9868 5202
rect 9875 5176 9894 5202
rect 9958 5198 9989 5210
rect 10004 5198 10107 5210
rect 10119 5200 10145 5226
rect 10160 5221 10190 5232
rect 10222 5228 10284 5244
rect 10222 5226 10268 5228
rect 10222 5210 10284 5226
rect 10296 5210 10302 5258
rect 10305 5250 10385 5258
rect 10305 5248 10324 5250
rect 10339 5248 10373 5250
rect 10305 5232 10385 5248
rect 10305 5210 10324 5232
rect 10339 5216 10369 5232
rect 10397 5226 10403 5300
rect 10406 5226 10425 5370
rect 10440 5226 10446 5370
rect 10455 5300 10468 5370
rect 10520 5366 10542 5370
rect 10513 5344 10542 5358
rect 10595 5344 10611 5358
rect 10649 5354 10655 5356
rect 10662 5354 10770 5370
rect 10777 5354 10783 5356
rect 10791 5354 10806 5370
rect 10872 5364 10891 5367
rect 10513 5342 10611 5344
rect 10638 5342 10806 5354
rect 10821 5344 10837 5358
rect 10872 5345 10894 5364
rect 10904 5358 10920 5359
rect 10903 5356 10920 5358
rect 10904 5351 10920 5356
rect 10894 5344 10900 5345
rect 10903 5344 10932 5351
rect 10821 5343 10932 5344
rect 10821 5342 10938 5343
rect 10497 5334 10548 5342
rect 10595 5334 10629 5342
rect 10497 5322 10522 5334
rect 10529 5322 10548 5334
rect 10602 5332 10629 5334
rect 10638 5332 10859 5342
rect 10894 5339 10900 5342
rect 10602 5328 10859 5332
rect 10497 5314 10548 5322
rect 10595 5314 10859 5328
rect 10903 5334 10938 5342
rect 10449 5266 10468 5300
rect 10513 5306 10542 5314
rect 10513 5300 10530 5306
rect 10513 5298 10547 5300
rect 10595 5298 10611 5314
rect 10612 5304 10820 5314
rect 10821 5304 10837 5314
rect 10885 5310 10900 5325
rect 10903 5322 10904 5334
rect 10911 5322 10938 5334
rect 10903 5314 10938 5322
rect 10903 5313 10932 5314
rect 10623 5300 10837 5304
rect 10638 5298 10837 5300
rect 10872 5300 10885 5310
rect 10903 5300 10920 5313
rect 10872 5298 10920 5300
rect 10514 5294 10547 5298
rect 10510 5292 10547 5294
rect 10510 5291 10577 5292
rect 10510 5286 10541 5291
rect 10547 5286 10577 5291
rect 10510 5282 10577 5286
rect 10483 5279 10577 5282
rect 10483 5272 10532 5279
rect 10483 5266 10513 5272
rect 10532 5267 10537 5272
rect 10449 5250 10529 5266
rect 10541 5258 10577 5279
rect 10638 5274 10827 5298
rect 10872 5297 10919 5298
rect 10885 5292 10919 5297
rect 10653 5271 10827 5274
rect 10646 5268 10827 5271
rect 10855 5291 10919 5292
rect 10449 5248 10468 5250
rect 10483 5248 10517 5250
rect 10449 5232 10529 5248
rect 10449 5226 10468 5232
rect 10165 5200 10268 5210
rect 10119 5198 10268 5200
rect 10289 5198 10324 5210
rect 9958 5196 10120 5198
rect 9970 5176 9989 5196
rect 10004 5194 10034 5196
rect 9853 5168 9894 5176
rect 9976 5172 9989 5176
rect 10041 5180 10120 5196
rect 10152 5196 10324 5198
rect 10152 5180 10231 5196
rect 10238 5194 10268 5196
rect 9816 5158 9845 5168
rect 9859 5158 9888 5168
rect 9903 5158 9933 5172
rect 9976 5158 10019 5172
rect 10041 5168 10231 5180
rect 10296 5176 10302 5196
rect 10026 5158 10056 5168
rect 10057 5158 10215 5168
rect 10219 5158 10249 5168
rect 10253 5158 10283 5172
rect 10311 5158 10324 5196
rect 10396 5210 10425 5226
rect 10439 5210 10468 5226
rect 10483 5216 10513 5232
rect 10541 5210 10547 5258
rect 10550 5252 10569 5258
rect 10584 5252 10614 5260
rect 10550 5244 10614 5252
rect 10550 5228 10630 5244
rect 10646 5237 10708 5268
rect 10724 5237 10786 5268
rect 10855 5266 10904 5291
rect 10919 5266 10949 5282
rect 10818 5252 10848 5260
rect 10855 5258 10965 5266
rect 10818 5244 10863 5252
rect 10550 5226 10569 5228
rect 10584 5226 10630 5228
rect 10550 5210 10630 5226
rect 10657 5224 10692 5237
rect 10733 5234 10770 5237
rect 10733 5232 10775 5234
rect 10662 5221 10692 5224
rect 10671 5217 10678 5221
rect 10678 5216 10679 5217
rect 10637 5210 10647 5216
rect 10396 5202 10431 5210
rect 10396 5176 10397 5202
rect 10404 5176 10431 5202
rect 10339 5158 10369 5172
rect 10396 5168 10431 5176
rect 10433 5202 10474 5210
rect 10433 5176 10448 5202
rect 10455 5176 10474 5202
rect 10538 5198 10569 5210
rect 10584 5198 10687 5210
rect 10699 5200 10725 5226
rect 10740 5221 10770 5232
rect 10802 5228 10864 5244
rect 10802 5226 10848 5228
rect 10802 5210 10864 5226
rect 10876 5210 10882 5258
rect 10885 5250 10965 5258
rect 10885 5248 10904 5250
rect 10919 5248 10953 5250
rect 10885 5232 10965 5248
rect 10885 5210 10904 5232
rect 10919 5216 10949 5232
rect 10977 5226 10983 5300
rect 10986 5226 11005 5370
rect 11020 5226 11026 5370
rect 11035 5300 11048 5370
rect 11100 5366 11122 5370
rect 11093 5344 11122 5358
rect 11175 5344 11191 5358
rect 11229 5354 11235 5356
rect 11242 5354 11350 5370
rect 11357 5354 11363 5356
rect 11371 5354 11386 5370
rect 11452 5364 11471 5367
rect 11093 5342 11191 5344
rect 11218 5342 11386 5354
rect 11401 5344 11417 5358
rect 11452 5345 11474 5364
rect 11484 5358 11500 5359
rect 11483 5356 11500 5358
rect 11484 5351 11500 5356
rect 11474 5344 11480 5345
rect 11483 5344 11512 5351
rect 11401 5343 11512 5344
rect 11401 5342 11518 5343
rect 11077 5334 11128 5342
rect 11175 5334 11209 5342
rect 11077 5322 11102 5334
rect 11109 5322 11128 5334
rect 11182 5332 11209 5334
rect 11218 5332 11439 5342
rect 11474 5339 11480 5342
rect 11182 5328 11439 5332
rect 11077 5314 11128 5322
rect 11175 5314 11439 5328
rect 11483 5334 11518 5342
rect 11029 5266 11048 5300
rect 11093 5306 11122 5314
rect 11093 5300 11110 5306
rect 11093 5298 11127 5300
rect 11175 5298 11191 5314
rect 11192 5304 11400 5314
rect 11401 5304 11417 5314
rect 11465 5310 11480 5325
rect 11483 5322 11484 5334
rect 11491 5322 11518 5334
rect 11483 5314 11518 5322
rect 11483 5313 11512 5314
rect 11203 5300 11417 5304
rect 11218 5298 11417 5300
rect 11452 5300 11465 5310
rect 11483 5300 11500 5313
rect 11452 5298 11500 5300
rect 11094 5294 11127 5298
rect 11090 5292 11127 5294
rect 11090 5291 11157 5292
rect 11090 5286 11121 5291
rect 11127 5286 11157 5291
rect 11090 5282 11157 5286
rect 11063 5279 11157 5282
rect 11063 5272 11112 5279
rect 11063 5266 11093 5272
rect 11112 5267 11117 5272
rect 11029 5250 11109 5266
rect 11121 5258 11157 5279
rect 11218 5274 11407 5298
rect 11452 5297 11499 5298
rect 11465 5292 11499 5297
rect 11233 5271 11407 5274
rect 11226 5268 11407 5271
rect 11435 5291 11499 5292
rect 11029 5248 11048 5250
rect 11063 5248 11097 5250
rect 11029 5232 11109 5248
rect 11029 5226 11048 5232
rect 10745 5200 10848 5210
rect 10699 5198 10848 5200
rect 10869 5198 10904 5210
rect 10538 5196 10700 5198
rect 10550 5176 10569 5196
rect 10584 5194 10614 5196
rect 10433 5168 10474 5176
rect 10556 5172 10569 5176
rect 10621 5180 10700 5196
rect 10732 5196 10904 5198
rect 10732 5180 10811 5196
rect 10818 5194 10848 5196
rect 10396 5158 10425 5168
rect 10439 5158 10468 5168
rect 10483 5158 10513 5172
rect 10556 5158 10599 5172
rect 10621 5168 10811 5180
rect 10876 5176 10882 5196
rect 10606 5158 10636 5168
rect 10637 5158 10795 5168
rect 10799 5158 10829 5168
rect 10833 5158 10863 5172
rect 10891 5158 10904 5196
rect 10976 5210 11005 5226
rect 11019 5210 11048 5226
rect 11063 5216 11093 5232
rect 11121 5210 11127 5258
rect 11130 5252 11149 5258
rect 11164 5252 11194 5260
rect 11130 5244 11194 5252
rect 11130 5228 11210 5244
rect 11226 5237 11288 5268
rect 11304 5237 11366 5268
rect 11435 5266 11484 5291
rect 11499 5266 11529 5282
rect 11398 5252 11428 5260
rect 11435 5258 11545 5266
rect 11398 5244 11443 5252
rect 11130 5226 11149 5228
rect 11164 5226 11210 5228
rect 11130 5210 11210 5226
rect 11237 5224 11272 5237
rect 11313 5234 11350 5237
rect 11313 5232 11355 5234
rect 11242 5221 11272 5224
rect 11251 5217 11258 5221
rect 11258 5216 11259 5217
rect 11217 5210 11227 5216
rect 10976 5202 11011 5210
rect 10976 5176 10977 5202
rect 10984 5176 11011 5202
rect 10919 5158 10949 5172
rect 10976 5168 11011 5176
rect 11013 5202 11054 5210
rect 11013 5176 11028 5202
rect 11035 5176 11054 5202
rect 11118 5198 11149 5210
rect 11164 5198 11267 5210
rect 11279 5200 11305 5226
rect 11320 5221 11350 5232
rect 11382 5228 11444 5244
rect 11382 5226 11428 5228
rect 11382 5210 11444 5226
rect 11456 5210 11462 5258
rect 11465 5250 11545 5258
rect 11465 5248 11484 5250
rect 11499 5248 11533 5250
rect 11465 5232 11545 5248
rect 11465 5210 11484 5232
rect 11499 5216 11529 5232
rect 11557 5226 11563 5300
rect 11566 5226 11585 5370
rect 11600 5226 11606 5370
rect 11615 5300 11628 5370
rect 11680 5366 11702 5370
rect 11673 5344 11702 5358
rect 11755 5344 11771 5358
rect 11809 5354 11815 5356
rect 11822 5354 11930 5370
rect 11937 5354 11943 5356
rect 11951 5354 11966 5370
rect 12032 5364 12051 5367
rect 11673 5342 11771 5344
rect 11798 5342 11966 5354
rect 11981 5344 11997 5358
rect 12032 5345 12054 5364
rect 12064 5358 12080 5359
rect 12063 5356 12080 5358
rect 12064 5351 12080 5356
rect 12054 5344 12060 5345
rect 12063 5344 12092 5351
rect 11981 5343 12092 5344
rect 11981 5342 12098 5343
rect 11657 5334 11708 5342
rect 11755 5334 11789 5342
rect 11657 5322 11682 5334
rect 11689 5322 11708 5334
rect 11762 5332 11789 5334
rect 11798 5332 12019 5342
rect 12054 5339 12060 5342
rect 11762 5328 12019 5332
rect 11657 5314 11708 5322
rect 11755 5314 12019 5328
rect 12063 5334 12098 5342
rect 11609 5266 11628 5300
rect 11673 5306 11702 5314
rect 11673 5300 11690 5306
rect 11673 5298 11707 5300
rect 11755 5298 11771 5314
rect 11772 5304 11980 5314
rect 11981 5304 11997 5314
rect 12045 5310 12060 5325
rect 12063 5322 12064 5334
rect 12071 5322 12098 5334
rect 12063 5314 12098 5322
rect 12063 5313 12092 5314
rect 11783 5300 11997 5304
rect 11798 5298 11997 5300
rect 12032 5300 12045 5310
rect 12063 5300 12080 5313
rect 12032 5298 12080 5300
rect 11674 5294 11707 5298
rect 11670 5292 11707 5294
rect 11670 5291 11737 5292
rect 11670 5286 11701 5291
rect 11707 5286 11737 5291
rect 11670 5282 11737 5286
rect 11643 5279 11737 5282
rect 11643 5272 11692 5279
rect 11643 5266 11673 5272
rect 11692 5267 11697 5272
rect 11609 5250 11689 5266
rect 11701 5258 11737 5279
rect 11798 5274 11987 5298
rect 12032 5297 12079 5298
rect 12045 5292 12079 5297
rect 11813 5271 11987 5274
rect 11806 5268 11987 5271
rect 12015 5291 12079 5292
rect 11609 5248 11628 5250
rect 11643 5248 11677 5250
rect 11609 5232 11689 5248
rect 11609 5226 11628 5232
rect 11325 5200 11428 5210
rect 11279 5198 11428 5200
rect 11449 5198 11484 5210
rect 11118 5196 11280 5198
rect 11130 5176 11149 5196
rect 11164 5194 11194 5196
rect 11013 5168 11054 5176
rect 11136 5172 11149 5176
rect 11201 5180 11280 5196
rect 11312 5196 11484 5198
rect 11312 5180 11391 5196
rect 11398 5194 11428 5196
rect 10976 5158 11005 5168
rect 11019 5158 11048 5168
rect 11063 5158 11093 5172
rect 11136 5158 11179 5172
rect 11201 5168 11391 5180
rect 11456 5176 11462 5196
rect 11186 5158 11216 5168
rect 11217 5158 11375 5168
rect 11379 5158 11409 5168
rect 11413 5158 11443 5172
rect 11471 5158 11484 5196
rect 11556 5210 11585 5226
rect 11599 5210 11628 5226
rect 11643 5216 11673 5232
rect 11701 5210 11707 5258
rect 11710 5252 11729 5258
rect 11744 5252 11774 5260
rect 11710 5244 11774 5252
rect 11710 5228 11790 5244
rect 11806 5237 11868 5268
rect 11884 5237 11946 5268
rect 12015 5266 12064 5291
rect 12079 5266 12109 5282
rect 11978 5252 12008 5260
rect 12015 5258 12125 5266
rect 11978 5244 12023 5252
rect 11710 5226 11729 5228
rect 11744 5226 11790 5228
rect 11710 5210 11790 5226
rect 11817 5224 11852 5237
rect 11893 5234 11930 5237
rect 11893 5232 11935 5234
rect 11822 5221 11852 5224
rect 11831 5217 11838 5221
rect 11838 5216 11839 5217
rect 11797 5210 11807 5216
rect 11556 5202 11591 5210
rect 11556 5176 11557 5202
rect 11564 5176 11591 5202
rect 11499 5158 11529 5172
rect 11556 5168 11591 5176
rect 11593 5202 11634 5210
rect 11593 5176 11608 5202
rect 11615 5176 11634 5202
rect 11698 5198 11729 5210
rect 11744 5198 11847 5210
rect 11859 5200 11885 5226
rect 11900 5221 11930 5232
rect 11962 5228 12024 5244
rect 11962 5226 12008 5228
rect 11962 5210 12024 5226
rect 12036 5210 12042 5258
rect 12045 5250 12125 5258
rect 12045 5248 12064 5250
rect 12079 5248 12113 5250
rect 12045 5232 12125 5248
rect 12045 5210 12064 5232
rect 12079 5216 12109 5232
rect 12137 5226 12143 5300
rect 12146 5226 12165 5370
rect 12180 5226 12186 5370
rect 12195 5300 12208 5370
rect 12260 5366 12282 5370
rect 12253 5344 12282 5358
rect 12335 5344 12351 5358
rect 12389 5354 12395 5356
rect 12402 5354 12510 5370
rect 12517 5354 12523 5356
rect 12531 5354 12546 5370
rect 12612 5364 12631 5367
rect 12253 5342 12351 5344
rect 12378 5342 12546 5354
rect 12561 5344 12577 5358
rect 12612 5345 12634 5364
rect 12644 5358 12660 5359
rect 12643 5356 12660 5358
rect 12644 5351 12660 5356
rect 12634 5344 12640 5345
rect 12643 5344 12672 5351
rect 12561 5343 12672 5344
rect 12561 5342 12678 5343
rect 12237 5334 12288 5342
rect 12335 5334 12369 5342
rect 12237 5322 12262 5334
rect 12269 5322 12288 5334
rect 12342 5332 12369 5334
rect 12378 5332 12599 5342
rect 12634 5339 12640 5342
rect 12342 5328 12599 5332
rect 12237 5314 12288 5322
rect 12335 5314 12599 5328
rect 12643 5334 12678 5342
rect 12189 5266 12208 5300
rect 12253 5306 12282 5314
rect 12253 5300 12270 5306
rect 12253 5298 12287 5300
rect 12335 5298 12351 5314
rect 12352 5304 12560 5314
rect 12561 5304 12577 5314
rect 12625 5310 12640 5325
rect 12643 5322 12644 5334
rect 12651 5322 12678 5334
rect 12643 5314 12678 5322
rect 12643 5313 12672 5314
rect 12363 5300 12577 5304
rect 12378 5298 12577 5300
rect 12612 5300 12625 5310
rect 12643 5300 12660 5313
rect 12612 5298 12660 5300
rect 12254 5294 12287 5298
rect 12250 5292 12287 5294
rect 12250 5291 12317 5292
rect 12250 5286 12281 5291
rect 12287 5286 12317 5291
rect 12250 5282 12317 5286
rect 12223 5279 12317 5282
rect 12223 5272 12272 5279
rect 12223 5266 12253 5272
rect 12272 5267 12277 5272
rect 12189 5250 12269 5266
rect 12281 5258 12317 5279
rect 12378 5274 12567 5298
rect 12612 5297 12659 5298
rect 12625 5292 12659 5297
rect 12393 5271 12567 5274
rect 12386 5268 12567 5271
rect 12595 5291 12659 5292
rect 12189 5248 12208 5250
rect 12223 5248 12257 5250
rect 12189 5232 12269 5248
rect 12189 5226 12208 5232
rect 11905 5200 12008 5210
rect 11859 5198 12008 5200
rect 12029 5198 12064 5210
rect 11698 5196 11860 5198
rect 11710 5176 11729 5196
rect 11744 5194 11774 5196
rect 11593 5168 11634 5176
rect 11716 5172 11729 5176
rect 11781 5180 11860 5196
rect 11892 5196 12064 5198
rect 11892 5180 11971 5196
rect 11978 5194 12008 5196
rect 11556 5158 11585 5168
rect 11599 5158 11628 5168
rect 11643 5158 11673 5172
rect 11716 5158 11759 5172
rect 11781 5168 11971 5180
rect 12036 5176 12042 5196
rect 11766 5158 11796 5168
rect 11797 5158 11955 5168
rect 11959 5158 11989 5168
rect 11993 5158 12023 5172
rect 12051 5158 12064 5196
rect 12136 5210 12165 5226
rect 12179 5210 12208 5226
rect 12223 5216 12253 5232
rect 12281 5210 12287 5258
rect 12290 5252 12309 5258
rect 12324 5252 12354 5260
rect 12290 5244 12354 5252
rect 12290 5228 12370 5244
rect 12386 5237 12448 5268
rect 12464 5237 12526 5268
rect 12595 5266 12644 5291
rect 12659 5266 12689 5282
rect 12558 5252 12588 5260
rect 12595 5258 12705 5266
rect 12558 5244 12603 5252
rect 12290 5226 12309 5228
rect 12324 5226 12370 5228
rect 12290 5210 12370 5226
rect 12397 5224 12432 5237
rect 12473 5234 12510 5237
rect 12473 5232 12515 5234
rect 12402 5221 12432 5224
rect 12411 5217 12418 5221
rect 12418 5216 12419 5217
rect 12377 5210 12387 5216
rect 12136 5202 12171 5210
rect 12136 5176 12137 5202
rect 12144 5176 12171 5202
rect 12079 5158 12109 5172
rect 12136 5168 12171 5176
rect 12173 5202 12214 5210
rect 12173 5176 12188 5202
rect 12195 5176 12214 5202
rect 12278 5198 12309 5210
rect 12324 5198 12427 5210
rect 12439 5200 12465 5226
rect 12480 5221 12510 5232
rect 12542 5228 12604 5244
rect 12542 5226 12588 5228
rect 12542 5210 12604 5226
rect 12616 5210 12622 5258
rect 12625 5250 12705 5258
rect 12625 5248 12644 5250
rect 12659 5248 12693 5250
rect 12625 5232 12705 5248
rect 12625 5210 12644 5232
rect 12659 5216 12689 5232
rect 12717 5226 12723 5300
rect 12726 5226 12745 5370
rect 12760 5226 12766 5370
rect 12775 5300 12788 5370
rect 12840 5366 12862 5370
rect 12833 5344 12862 5358
rect 12915 5344 12931 5358
rect 12969 5354 12975 5356
rect 12982 5354 13090 5370
rect 13097 5354 13103 5356
rect 13111 5354 13126 5370
rect 13192 5364 13211 5367
rect 12833 5342 12931 5344
rect 12958 5342 13126 5354
rect 13141 5344 13157 5358
rect 13192 5345 13214 5364
rect 13224 5358 13240 5359
rect 13223 5356 13240 5358
rect 13224 5351 13240 5356
rect 13214 5344 13220 5345
rect 13223 5344 13252 5351
rect 13141 5343 13252 5344
rect 13141 5342 13258 5343
rect 12817 5334 12868 5342
rect 12915 5334 12949 5342
rect 12817 5322 12842 5334
rect 12849 5322 12868 5334
rect 12922 5332 12949 5334
rect 12958 5332 13179 5342
rect 13214 5339 13220 5342
rect 12922 5328 13179 5332
rect 12817 5314 12868 5322
rect 12915 5314 13179 5328
rect 13223 5334 13258 5342
rect 12769 5266 12788 5300
rect 12833 5306 12862 5314
rect 12833 5300 12850 5306
rect 12833 5298 12867 5300
rect 12915 5298 12931 5314
rect 12932 5304 13140 5314
rect 13141 5304 13157 5314
rect 13205 5310 13220 5325
rect 13223 5322 13224 5334
rect 13231 5322 13258 5334
rect 13223 5314 13258 5322
rect 13223 5313 13252 5314
rect 12943 5300 13157 5304
rect 12958 5298 13157 5300
rect 13192 5300 13205 5310
rect 13223 5300 13240 5313
rect 13192 5298 13240 5300
rect 12834 5294 12867 5298
rect 12830 5292 12867 5294
rect 12830 5291 12897 5292
rect 12830 5286 12861 5291
rect 12867 5286 12897 5291
rect 12830 5282 12897 5286
rect 12803 5279 12897 5282
rect 12803 5272 12852 5279
rect 12803 5266 12833 5272
rect 12852 5267 12857 5272
rect 12769 5250 12849 5266
rect 12861 5258 12897 5279
rect 12958 5274 13147 5298
rect 13192 5297 13239 5298
rect 13205 5292 13239 5297
rect 12973 5271 13147 5274
rect 12966 5268 13147 5271
rect 13175 5291 13239 5292
rect 12769 5248 12788 5250
rect 12803 5248 12837 5250
rect 12769 5232 12849 5248
rect 12769 5226 12788 5232
rect 12485 5200 12588 5210
rect 12439 5198 12588 5200
rect 12609 5198 12644 5210
rect 12278 5196 12440 5198
rect 12290 5176 12309 5196
rect 12324 5194 12354 5196
rect 12173 5168 12214 5176
rect 12296 5172 12309 5176
rect 12361 5180 12440 5196
rect 12472 5196 12644 5198
rect 12472 5180 12551 5196
rect 12558 5194 12588 5196
rect 12136 5158 12165 5168
rect 12179 5158 12208 5168
rect 12223 5158 12253 5172
rect 12296 5158 12339 5172
rect 12361 5168 12551 5180
rect 12616 5176 12622 5196
rect 12346 5158 12376 5168
rect 12377 5158 12535 5168
rect 12539 5158 12569 5168
rect 12573 5158 12603 5172
rect 12631 5158 12644 5196
rect 12716 5210 12745 5226
rect 12759 5210 12788 5226
rect 12803 5216 12833 5232
rect 12861 5210 12867 5258
rect 12870 5252 12889 5258
rect 12904 5252 12934 5260
rect 12870 5244 12934 5252
rect 12870 5228 12950 5244
rect 12966 5237 13028 5268
rect 13044 5237 13106 5268
rect 13175 5266 13224 5291
rect 13239 5266 13269 5282
rect 13138 5252 13168 5260
rect 13175 5258 13285 5266
rect 13138 5244 13183 5252
rect 12870 5226 12889 5228
rect 12904 5226 12950 5228
rect 12870 5210 12950 5226
rect 12977 5224 13012 5237
rect 13053 5234 13090 5237
rect 13053 5232 13095 5234
rect 12982 5221 13012 5224
rect 12991 5217 12998 5221
rect 12998 5216 12999 5217
rect 12957 5210 12967 5216
rect 12716 5202 12751 5210
rect 12716 5176 12717 5202
rect 12724 5176 12751 5202
rect 12659 5158 12689 5172
rect 12716 5168 12751 5176
rect 12753 5202 12794 5210
rect 12753 5176 12768 5202
rect 12775 5176 12794 5202
rect 12858 5198 12889 5210
rect 12904 5198 13007 5210
rect 13019 5200 13045 5226
rect 13060 5221 13090 5232
rect 13122 5228 13184 5244
rect 13122 5226 13168 5228
rect 13122 5210 13184 5226
rect 13196 5210 13202 5258
rect 13205 5250 13285 5258
rect 13205 5248 13224 5250
rect 13239 5248 13273 5250
rect 13205 5232 13285 5248
rect 13205 5210 13224 5232
rect 13239 5216 13269 5232
rect 13297 5226 13303 5300
rect 13306 5226 13325 5370
rect 13340 5226 13346 5370
rect 13355 5300 13368 5370
rect 13420 5366 13442 5370
rect 13413 5344 13442 5358
rect 13495 5344 13511 5358
rect 13549 5354 13555 5356
rect 13562 5354 13670 5370
rect 13677 5354 13683 5356
rect 13691 5354 13706 5370
rect 13772 5364 13791 5367
rect 13413 5342 13511 5344
rect 13538 5342 13706 5354
rect 13721 5344 13737 5358
rect 13772 5345 13794 5364
rect 13804 5358 13820 5359
rect 13803 5356 13820 5358
rect 13804 5351 13820 5356
rect 13794 5344 13800 5345
rect 13803 5344 13832 5351
rect 13721 5343 13832 5344
rect 13721 5342 13838 5343
rect 13397 5334 13448 5342
rect 13495 5334 13529 5342
rect 13397 5322 13422 5334
rect 13429 5322 13448 5334
rect 13502 5332 13529 5334
rect 13538 5332 13759 5342
rect 13794 5339 13800 5342
rect 13502 5328 13759 5332
rect 13397 5314 13448 5322
rect 13495 5314 13759 5328
rect 13803 5334 13838 5342
rect 13349 5266 13368 5300
rect 13413 5306 13442 5314
rect 13413 5300 13430 5306
rect 13413 5298 13447 5300
rect 13495 5298 13511 5314
rect 13512 5304 13720 5314
rect 13721 5304 13737 5314
rect 13785 5310 13800 5325
rect 13803 5322 13804 5334
rect 13811 5322 13838 5334
rect 13803 5314 13838 5322
rect 13803 5313 13832 5314
rect 13523 5300 13737 5304
rect 13538 5298 13737 5300
rect 13772 5300 13785 5310
rect 13803 5300 13820 5313
rect 13772 5298 13820 5300
rect 13414 5294 13447 5298
rect 13410 5292 13447 5294
rect 13410 5291 13477 5292
rect 13410 5286 13441 5291
rect 13447 5286 13477 5291
rect 13410 5282 13477 5286
rect 13383 5279 13477 5282
rect 13383 5272 13432 5279
rect 13383 5266 13413 5272
rect 13432 5267 13437 5272
rect 13349 5250 13429 5266
rect 13441 5258 13477 5279
rect 13538 5274 13727 5298
rect 13772 5297 13819 5298
rect 13785 5292 13819 5297
rect 13553 5271 13727 5274
rect 13546 5268 13727 5271
rect 13755 5291 13819 5292
rect 13349 5248 13368 5250
rect 13383 5248 13417 5250
rect 13349 5232 13429 5248
rect 13349 5226 13368 5232
rect 13065 5200 13168 5210
rect 13019 5198 13168 5200
rect 13189 5198 13224 5210
rect 12858 5196 13020 5198
rect 12870 5176 12889 5196
rect 12904 5194 12934 5196
rect 12753 5168 12794 5176
rect 12876 5172 12889 5176
rect 12941 5180 13020 5196
rect 13052 5196 13224 5198
rect 13052 5180 13131 5196
rect 13138 5194 13168 5196
rect 12716 5158 12745 5168
rect 12759 5158 12788 5168
rect 12803 5158 12833 5172
rect 12876 5158 12919 5172
rect 12941 5168 13131 5180
rect 13196 5176 13202 5196
rect 12926 5158 12956 5168
rect 12957 5158 13115 5168
rect 13119 5158 13149 5168
rect 13153 5158 13183 5172
rect 13211 5158 13224 5196
rect 13296 5210 13325 5226
rect 13339 5210 13368 5226
rect 13383 5216 13413 5232
rect 13441 5210 13447 5258
rect 13450 5252 13469 5258
rect 13484 5252 13514 5260
rect 13450 5244 13514 5252
rect 13450 5228 13530 5244
rect 13546 5237 13608 5268
rect 13624 5237 13686 5268
rect 13755 5266 13804 5291
rect 13819 5266 13849 5282
rect 13718 5252 13748 5260
rect 13755 5258 13865 5266
rect 13718 5244 13763 5252
rect 13450 5226 13469 5228
rect 13484 5226 13530 5228
rect 13450 5210 13530 5226
rect 13557 5224 13592 5237
rect 13633 5234 13670 5237
rect 13633 5232 13675 5234
rect 13562 5221 13592 5224
rect 13571 5217 13578 5221
rect 13578 5216 13579 5217
rect 13537 5210 13547 5216
rect 13296 5202 13331 5210
rect 13296 5176 13297 5202
rect 13304 5176 13331 5202
rect 13239 5158 13269 5172
rect 13296 5168 13331 5176
rect 13333 5202 13374 5210
rect 13333 5176 13348 5202
rect 13355 5176 13374 5202
rect 13438 5198 13469 5210
rect 13484 5198 13587 5210
rect 13599 5200 13625 5226
rect 13640 5221 13670 5232
rect 13702 5228 13764 5244
rect 13702 5226 13748 5228
rect 13702 5210 13764 5226
rect 13776 5210 13782 5258
rect 13785 5250 13865 5258
rect 13785 5248 13804 5250
rect 13819 5248 13853 5250
rect 13785 5232 13865 5248
rect 13785 5210 13804 5232
rect 13819 5216 13849 5232
rect 13877 5226 13883 5300
rect 13886 5226 13905 5370
rect 13920 5226 13926 5370
rect 13935 5300 13948 5370
rect 14000 5366 14022 5370
rect 13993 5344 14022 5358
rect 14075 5344 14091 5358
rect 14129 5354 14135 5356
rect 14142 5354 14250 5370
rect 14257 5354 14263 5356
rect 14271 5354 14286 5370
rect 14352 5364 14371 5367
rect 13993 5342 14091 5344
rect 14118 5342 14286 5354
rect 14301 5344 14317 5358
rect 14352 5345 14374 5364
rect 14384 5358 14400 5359
rect 14383 5356 14400 5358
rect 14384 5351 14400 5356
rect 14374 5344 14380 5345
rect 14383 5344 14412 5351
rect 14301 5343 14412 5344
rect 14301 5342 14418 5343
rect 13977 5334 14028 5342
rect 14075 5334 14109 5342
rect 13977 5322 14002 5334
rect 14009 5322 14028 5334
rect 14082 5332 14109 5334
rect 14118 5332 14339 5342
rect 14374 5339 14380 5342
rect 14082 5328 14339 5332
rect 13977 5314 14028 5322
rect 14075 5314 14339 5328
rect 14383 5334 14418 5342
rect 13929 5266 13948 5300
rect 13993 5306 14022 5314
rect 13993 5300 14010 5306
rect 13993 5298 14027 5300
rect 14075 5298 14091 5314
rect 14092 5304 14300 5314
rect 14301 5304 14317 5314
rect 14365 5310 14380 5325
rect 14383 5322 14384 5334
rect 14391 5322 14418 5334
rect 14383 5314 14418 5322
rect 14383 5313 14412 5314
rect 14103 5300 14317 5304
rect 14118 5298 14317 5300
rect 14352 5300 14365 5310
rect 14383 5300 14400 5313
rect 14352 5298 14400 5300
rect 13994 5294 14027 5298
rect 13990 5292 14027 5294
rect 13990 5291 14057 5292
rect 13990 5286 14021 5291
rect 14027 5286 14057 5291
rect 13990 5282 14057 5286
rect 13963 5279 14057 5282
rect 13963 5272 14012 5279
rect 13963 5266 13993 5272
rect 14012 5267 14017 5272
rect 13929 5250 14009 5266
rect 14021 5258 14057 5279
rect 14118 5274 14307 5298
rect 14352 5297 14399 5298
rect 14365 5292 14399 5297
rect 14133 5271 14307 5274
rect 14126 5268 14307 5271
rect 14335 5291 14399 5292
rect 13929 5248 13948 5250
rect 13963 5248 13997 5250
rect 13929 5232 14009 5248
rect 13929 5226 13948 5232
rect 13645 5200 13748 5210
rect 13599 5198 13748 5200
rect 13769 5198 13804 5210
rect 13438 5196 13600 5198
rect 13450 5176 13469 5196
rect 13484 5194 13514 5196
rect 13333 5168 13374 5176
rect 13456 5172 13469 5176
rect 13521 5180 13600 5196
rect 13632 5196 13804 5198
rect 13632 5180 13711 5196
rect 13718 5194 13748 5196
rect 13296 5158 13325 5168
rect 13339 5158 13368 5168
rect 13383 5158 13413 5172
rect 13456 5158 13499 5172
rect 13521 5168 13711 5180
rect 13776 5176 13782 5196
rect 13506 5158 13536 5168
rect 13537 5158 13695 5168
rect 13699 5158 13729 5168
rect 13733 5158 13763 5172
rect 13791 5158 13804 5196
rect 13876 5210 13905 5226
rect 13919 5210 13948 5226
rect 13963 5216 13993 5232
rect 14021 5210 14027 5258
rect 14030 5252 14049 5258
rect 14064 5252 14094 5260
rect 14030 5244 14094 5252
rect 14030 5228 14110 5244
rect 14126 5237 14188 5268
rect 14204 5237 14266 5268
rect 14335 5266 14384 5291
rect 14399 5266 14429 5282
rect 14298 5252 14328 5260
rect 14335 5258 14445 5266
rect 14298 5244 14343 5252
rect 14030 5226 14049 5228
rect 14064 5226 14110 5228
rect 14030 5210 14110 5226
rect 14137 5224 14172 5237
rect 14213 5234 14250 5237
rect 14213 5232 14255 5234
rect 14142 5221 14172 5224
rect 14151 5217 14158 5221
rect 14158 5216 14159 5217
rect 14117 5210 14127 5216
rect 13876 5202 13911 5210
rect 13876 5176 13877 5202
rect 13884 5176 13911 5202
rect 13819 5158 13849 5172
rect 13876 5168 13911 5176
rect 13913 5202 13954 5210
rect 13913 5176 13928 5202
rect 13935 5176 13954 5202
rect 14018 5198 14049 5210
rect 14064 5198 14167 5210
rect 14179 5200 14205 5226
rect 14220 5221 14250 5232
rect 14282 5228 14344 5244
rect 14282 5226 14328 5228
rect 14282 5210 14344 5226
rect 14356 5210 14362 5258
rect 14365 5250 14445 5258
rect 14365 5248 14384 5250
rect 14399 5248 14433 5250
rect 14365 5232 14445 5248
rect 14365 5210 14384 5232
rect 14399 5216 14429 5232
rect 14457 5226 14463 5300
rect 14466 5226 14485 5370
rect 14500 5226 14506 5370
rect 14515 5300 14528 5370
rect 14580 5366 14602 5370
rect 14573 5344 14602 5358
rect 14655 5344 14671 5358
rect 14709 5354 14715 5356
rect 14722 5354 14830 5370
rect 14837 5354 14843 5356
rect 14851 5354 14866 5370
rect 14932 5364 14951 5367
rect 14573 5342 14671 5344
rect 14698 5342 14866 5354
rect 14881 5344 14897 5358
rect 14932 5345 14954 5364
rect 14964 5358 14980 5359
rect 14963 5356 14980 5358
rect 14964 5351 14980 5356
rect 14954 5344 14960 5345
rect 14963 5344 14992 5351
rect 14881 5343 14992 5344
rect 14881 5342 14998 5343
rect 14557 5334 14608 5342
rect 14655 5334 14689 5342
rect 14557 5322 14582 5334
rect 14589 5322 14608 5334
rect 14662 5332 14689 5334
rect 14698 5332 14919 5342
rect 14954 5339 14960 5342
rect 14662 5328 14919 5332
rect 14557 5314 14608 5322
rect 14655 5314 14919 5328
rect 14963 5334 14998 5342
rect 14509 5266 14528 5300
rect 14573 5306 14602 5314
rect 14573 5300 14590 5306
rect 14573 5298 14607 5300
rect 14655 5298 14671 5314
rect 14672 5304 14880 5314
rect 14881 5304 14897 5314
rect 14945 5310 14960 5325
rect 14963 5322 14964 5334
rect 14971 5322 14998 5334
rect 14963 5314 14998 5322
rect 14963 5313 14992 5314
rect 14683 5300 14897 5304
rect 14698 5298 14897 5300
rect 14932 5300 14945 5310
rect 14963 5300 14980 5313
rect 14932 5298 14980 5300
rect 14574 5294 14607 5298
rect 14570 5292 14607 5294
rect 14570 5291 14637 5292
rect 14570 5286 14601 5291
rect 14607 5286 14637 5291
rect 14570 5282 14637 5286
rect 14543 5279 14637 5282
rect 14543 5272 14592 5279
rect 14543 5266 14573 5272
rect 14592 5267 14597 5272
rect 14509 5250 14589 5266
rect 14601 5258 14637 5279
rect 14698 5274 14887 5298
rect 14932 5297 14979 5298
rect 14945 5292 14979 5297
rect 14713 5271 14887 5274
rect 14706 5268 14887 5271
rect 14915 5291 14979 5292
rect 14509 5248 14528 5250
rect 14543 5248 14577 5250
rect 14509 5232 14589 5248
rect 14509 5226 14528 5232
rect 14225 5200 14328 5210
rect 14179 5198 14328 5200
rect 14349 5198 14384 5210
rect 14018 5196 14180 5198
rect 14030 5176 14049 5196
rect 14064 5194 14094 5196
rect 13913 5168 13954 5176
rect 14036 5172 14049 5176
rect 14101 5180 14180 5196
rect 14212 5196 14384 5198
rect 14212 5180 14291 5196
rect 14298 5194 14328 5196
rect 13876 5158 13905 5168
rect 13919 5158 13948 5168
rect 13963 5158 13993 5172
rect 14036 5158 14079 5172
rect 14101 5168 14291 5180
rect 14356 5176 14362 5196
rect 14086 5158 14116 5168
rect 14117 5158 14275 5168
rect 14279 5158 14309 5168
rect 14313 5158 14343 5172
rect 14371 5158 14384 5196
rect 14456 5210 14485 5226
rect 14499 5210 14528 5226
rect 14543 5216 14573 5232
rect 14601 5210 14607 5258
rect 14610 5252 14629 5258
rect 14644 5252 14674 5260
rect 14610 5244 14674 5252
rect 14610 5228 14690 5244
rect 14706 5237 14768 5268
rect 14784 5237 14846 5268
rect 14915 5266 14964 5291
rect 14979 5266 15009 5282
rect 14878 5252 14908 5260
rect 14915 5258 15025 5266
rect 14878 5244 14923 5252
rect 14610 5226 14629 5228
rect 14644 5226 14690 5228
rect 14610 5210 14690 5226
rect 14717 5224 14752 5237
rect 14793 5234 14830 5237
rect 14793 5232 14835 5234
rect 14722 5221 14752 5224
rect 14731 5217 14738 5221
rect 14738 5216 14739 5217
rect 14697 5210 14707 5216
rect 14456 5202 14491 5210
rect 14456 5176 14457 5202
rect 14464 5176 14491 5202
rect 14399 5158 14429 5172
rect 14456 5168 14491 5176
rect 14493 5202 14534 5210
rect 14493 5176 14508 5202
rect 14515 5176 14534 5202
rect 14598 5198 14629 5210
rect 14644 5198 14747 5210
rect 14759 5200 14785 5226
rect 14800 5221 14830 5232
rect 14862 5228 14924 5244
rect 14862 5226 14908 5228
rect 14862 5210 14924 5226
rect 14936 5210 14942 5258
rect 14945 5250 15025 5258
rect 14945 5248 14964 5250
rect 14979 5248 15013 5250
rect 14945 5232 15025 5248
rect 14945 5210 14964 5232
rect 14979 5216 15009 5232
rect 15037 5226 15043 5300
rect 15046 5226 15065 5370
rect 15080 5226 15086 5370
rect 15095 5300 15108 5370
rect 15160 5366 15182 5370
rect 15153 5344 15182 5358
rect 15235 5344 15251 5358
rect 15289 5354 15295 5356
rect 15302 5354 15410 5370
rect 15417 5354 15423 5356
rect 15431 5354 15446 5370
rect 15512 5364 15531 5367
rect 15153 5342 15251 5344
rect 15278 5342 15446 5354
rect 15461 5344 15477 5358
rect 15512 5345 15534 5364
rect 15544 5358 15560 5359
rect 15543 5356 15560 5358
rect 15544 5351 15560 5356
rect 15534 5344 15540 5345
rect 15543 5344 15572 5351
rect 15461 5343 15572 5344
rect 15461 5342 15578 5343
rect 15137 5334 15188 5342
rect 15235 5334 15269 5342
rect 15137 5322 15162 5334
rect 15169 5322 15188 5334
rect 15242 5332 15269 5334
rect 15278 5332 15499 5342
rect 15534 5339 15540 5342
rect 15242 5328 15499 5332
rect 15137 5314 15188 5322
rect 15235 5314 15499 5328
rect 15543 5334 15578 5342
rect 15089 5266 15108 5300
rect 15153 5306 15182 5314
rect 15153 5300 15170 5306
rect 15153 5298 15187 5300
rect 15235 5298 15251 5314
rect 15252 5304 15460 5314
rect 15461 5304 15477 5314
rect 15525 5310 15540 5325
rect 15543 5322 15544 5334
rect 15551 5322 15578 5334
rect 15543 5314 15578 5322
rect 15543 5313 15572 5314
rect 15263 5300 15477 5304
rect 15278 5298 15477 5300
rect 15512 5300 15525 5310
rect 15543 5300 15560 5313
rect 15512 5298 15560 5300
rect 15154 5294 15187 5298
rect 15150 5292 15187 5294
rect 15150 5291 15217 5292
rect 15150 5286 15181 5291
rect 15187 5286 15217 5291
rect 15150 5282 15217 5286
rect 15123 5279 15217 5282
rect 15123 5272 15172 5279
rect 15123 5266 15153 5272
rect 15172 5267 15177 5272
rect 15089 5250 15169 5266
rect 15181 5258 15217 5279
rect 15278 5274 15467 5298
rect 15512 5297 15559 5298
rect 15525 5292 15559 5297
rect 15293 5271 15467 5274
rect 15286 5268 15467 5271
rect 15495 5291 15559 5292
rect 15089 5248 15108 5250
rect 15123 5248 15157 5250
rect 15089 5232 15169 5248
rect 15089 5226 15108 5232
rect 14805 5200 14908 5210
rect 14759 5198 14908 5200
rect 14929 5198 14964 5210
rect 14598 5196 14760 5198
rect 14610 5176 14629 5196
rect 14644 5194 14674 5196
rect 14493 5168 14534 5176
rect 14616 5172 14629 5176
rect 14681 5180 14760 5196
rect 14792 5196 14964 5198
rect 14792 5180 14871 5196
rect 14878 5194 14908 5196
rect 14456 5158 14485 5168
rect 14499 5158 14528 5168
rect 14543 5158 14573 5172
rect 14616 5158 14659 5172
rect 14681 5168 14871 5180
rect 14936 5176 14942 5196
rect 14666 5158 14696 5168
rect 14697 5158 14855 5168
rect 14859 5158 14889 5168
rect 14893 5158 14923 5172
rect 14951 5158 14964 5196
rect 15036 5210 15065 5226
rect 15079 5210 15108 5226
rect 15123 5216 15153 5232
rect 15181 5210 15187 5258
rect 15190 5252 15209 5258
rect 15224 5252 15254 5260
rect 15190 5244 15254 5252
rect 15190 5228 15270 5244
rect 15286 5237 15348 5268
rect 15364 5237 15426 5268
rect 15495 5266 15544 5291
rect 15559 5266 15589 5282
rect 15458 5252 15488 5260
rect 15495 5258 15605 5266
rect 15458 5244 15503 5252
rect 15190 5226 15209 5228
rect 15224 5226 15270 5228
rect 15190 5210 15270 5226
rect 15297 5224 15332 5237
rect 15373 5234 15410 5237
rect 15373 5232 15415 5234
rect 15302 5221 15332 5224
rect 15311 5217 15318 5221
rect 15318 5216 15319 5217
rect 15277 5210 15287 5216
rect 15036 5202 15071 5210
rect 15036 5176 15037 5202
rect 15044 5176 15071 5202
rect 14979 5158 15009 5172
rect 15036 5168 15071 5176
rect 15073 5202 15114 5210
rect 15073 5176 15088 5202
rect 15095 5176 15114 5202
rect 15178 5198 15209 5210
rect 15224 5198 15327 5210
rect 15339 5200 15365 5226
rect 15380 5221 15410 5232
rect 15442 5228 15504 5244
rect 15442 5226 15488 5228
rect 15442 5210 15504 5226
rect 15516 5210 15522 5258
rect 15525 5250 15605 5258
rect 15525 5248 15544 5250
rect 15559 5248 15593 5250
rect 15525 5232 15605 5248
rect 15525 5210 15544 5232
rect 15559 5216 15589 5232
rect 15617 5226 15623 5300
rect 15626 5226 15645 5370
rect 15660 5226 15666 5370
rect 15675 5300 15688 5370
rect 15740 5366 15762 5370
rect 15733 5344 15762 5358
rect 15815 5344 15831 5358
rect 15869 5354 15875 5356
rect 15882 5354 15990 5370
rect 15997 5354 16003 5356
rect 16011 5354 16026 5370
rect 16092 5364 16111 5367
rect 15733 5342 15831 5344
rect 15858 5342 16026 5354
rect 16041 5344 16057 5358
rect 16092 5345 16114 5364
rect 16124 5358 16140 5359
rect 16123 5356 16140 5358
rect 16124 5351 16140 5356
rect 16114 5344 16120 5345
rect 16123 5344 16152 5351
rect 16041 5343 16152 5344
rect 16041 5342 16158 5343
rect 15717 5334 15768 5342
rect 15815 5334 15849 5342
rect 15717 5322 15742 5334
rect 15749 5322 15768 5334
rect 15822 5332 15849 5334
rect 15858 5332 16079 5342
rect 16114 5339 16120 5342
rect 15822 5328 16079 5332
rect 15717 5314 15768 5322
rect 15815 5314 16079 5328
rect 16123 5334 16158 5342
rect 15669 5266 15688 5300
rect 15733 5306 15762 5314
rect 15733 5300 15750 5306
rect 15733 5298 15767 5300
rect 15815 5298 15831 5314
rect 15832 5304 16040 5314
rect 16041 5304 16057 5314
rect 16105 5310 16120 5325
rect 16123 5322 16124 5334
rect 16131 5322 16158 5334
rect 16123 5314 16158 5322
rect 16123 5313 16152 5314
rect 15843 5300 16057 5304
rect 15858 5298 16057 5300
rect 16092 5300 16105 5310
rect 16123 5300 16140 5313
rect 16092 5298 16140 5300
rect 15734 5294 15767 5298
rect 15730 5292 15767 5294
rect 15730 5291 15797 5292
rect 15730 5286 15761 5291
rect 15767 5286 15797 5291
rect 15730 5282 15797 5286
rect 15703 5279 15797 5282
rect 15703 5272 15752 5279
rect 15703 5266 15733 5272
rect 15752 5267 15757 5272
rect 15669 5250 15749 5266
rect 15761 5258 15797 5279
rect 15858 5274 16047 5298
rect 16092 5297 16139 5298
rect 16105 5292 16139 5297
rect 15873 5271 16047 5274
rect 15866 5268 16047 5271
rect 16075 5291 16139 5292
rect 15669 5248 15688 5250
rect 15703 5248 15737 5250
rect 15669 5232 15749 5248
rect 15669 5226 15688 5232
rect 15385 5200 15488 5210
rect 15339 5198 15488 5200
rect 15509 5198 15544 5210
rect 15178 5196 15340 5198
rect 15190 5176 15209 5196
rect 15224 5194 15254 5196
rect 15073 5168 15114 5176
rect 15196 5172 15209 5176
rect 15261 5180 15340 5196
rect 15372 5196 15544 5198
rect 15372 5180 15451 5196
rect 15458 5194 15488 5196
rect 15036 5158 15065 5168
rect 15079 5158 15108 5168
rect 15123 5158 15153 5172
rect 15196 5158 15239 5172
rect 15261 5168 15451 5180
rect 15516 5176 15522 5196
rect 15246 5158 15276 5168
rect 15277 5158 15435 5168
rect 15439 5158 15469 5168
rect 15473 5158 15503 5172
rect 15531 5158 15544 5196
rect 15616 5210 15645 5226
rect 15659 5210 15688 5226
rect 15703 5216 15733 5232
rect 15761 5210 15767 5258
rect 15770 5252 15789 5258
rect 15804 5252 15834 5260
rect 15770 5244 15834 5252
rect 15770 5228 15850 5244
rect 15866 5237 15928 5268
rect 15944 5237 16006 5268
rect 16075 5266 16124 5291
rect 16139 5266 16169 5282
rect 16038 5252 16068 5260
rect 16075 5258 16185 5266
rect 16038 5244 16083 5252
rect 15770 5226 15789 5228
rect 15804 5226 15850 5228
rect 15770 5210 15850 5226
rect 15877 5224 15912 5237
rect 15953 5234 15990 5237
rect 15953 5232 15995 5234
rect 15882 5221 15912 5224
rect 15891 5217 15898 5221
rect 15898 5216 15899 5217
rect 15857 5210 15867 5216
rect 15616 5202 15651 5210
rect 15616 5176 15617 5202
rect 15624 5176 15651 5202
rect 15559 5158 15589 5172
rect 15616 5168 15651 5176
rect 15653 5202 15694 5210
rect 15653 5176 15668 5202
rect 15675 5176 15694 5202
rect 15758 5198 15789 5210
rect 15804 5198 15907 5210
rect 15919 5200 15945 5226
rect 15960 5221 15990 5232
rect 16022 5228 16084 5244
rect 16022 5226 16068 5228
rect 16022 5210 16084 5226
rect 16096 5210 16102 5258
rect 16105 5250 16185 5258
rect 16105 5248 16124 5250
rect 16139 5248 16173 5250
rect 16105 5232 16185 5248
rect 16105 5210 16124 5232
rect 16139 5216 16169 5232
rect 16197 5226 16203 5300
rect 16206 5226 16225 5370
rect 16240 5226 16246 5370
rect 16255 5300 16268 5370
rect 16320 5366 16342 5370
rect 16313 5344 16342 5358
rect 16395 5344 16411 5358
rect 16449 5354 16455 5356
rect 16462 5354 16570 5370
rect 16577 5354 16583 5356
rect 16591 5354 16606 5370
rect 16672 5364 16691 5367
rect 16313 5342 16411 5344
rect 16438 5342 16606 5354
rect 16621 5344 16637 5358
rect 16672 5345 16694 5364
rect 16704 5358 16720 5359
rect 16703 5356 16720 5358
rect 16704 5351 16720 5356
rect 16694 5344 16700 5345
rect 16703 5344 16732 5351
rect 16621 5343 16732 5344
rect 16621 5342 16738 5343
rect 16297 5334 16348 5342
rect 16395 5334 16429 5342
rect 16297 5322 16322 5334
rect 16329 5322 16348 5334
rect 16402 5332 16429 5334
rect 16438 5332 16659 5342
rect 16694 5339 16700 5342
rect 16402 5328 16659 5332
rect 16297 5314 16348 5322
rect 16395 5314 16659 5328
rect 16703 5334 16738 5342
rect 16249 5266 16268 5300
rect 16313 5306 16342 5314
rect 16313 5300 16330 5306
rect 16313 5298 16347 5300
rect 16395 5298 16411 5314
rect 16412 5304 16620 5314
rect 16621 5304 16637 5314
rect 16685 5310 16700 5325
rect 16703 5322 16704 5334
rect 16711 5322 16738 5334
rect 16703 5314 16738 5322
rect 16703 5313 16732 5314
rect 16423 5300 16637 5304
rect 16438 5298 16637 5300
rect 16672 5300 16685 5310
rect 16703 5300 16720 5313
rect 16672 5298 16720 5300
rect 16314 5294 16347 5298
rect 16310 5292 16347 5294
rect 16310 5291 16377 5292
rect 16310 5286 16341 5291
rect 16347 5286 16377 5291
rect 16310 5282 16377 5286
rect 16283 5279 16377 5282
rect 16283 5272 16332 5279
rect 16283 5266 16313 5272
rect 16332 5267 16337 5272
rect 16249 5250 16329 5266
rect 16341 5258 16377 5279
rect 16438 5274 16627 5298
rect 16672 5297 16719 5298
rect 16685 5292 16719 5297
rect 16453 5271 16627 5274
rect 16446 5268 16627 5271
rect 16655 5291 16719 5292
rect 16249 5248 16268 5250
rect 16283 5248 16317 5250
rect 16249 5232 16329 5248
rect 16249 5226 16268 5232
rect 15965 5200 16068 5210
rect 15919 5198 16068 5200
rect 16089 5198 16124 5210
rect 15758 5196 15920 5198
rect 15770 5176 15789 5196
rect 15804 5194 15834 5196
rect 15653 5168 15694 5176
rect 15776 5172 15789 5176
rect 15841 5180 15920 5196
rect 15952 5196 16124 5198
rect 15952 5180 16031 5196
rect 16038 5194 16068 5196
rect 15616 5158 15645 5168
rect 15659 5158 15688 5168
rect 15703 5158 15733 5172
rect 15776 5158 15819 5172
rect 15841 5168 16031 5180
rect 16096 5176 16102 5196
rect 15826 5158 15856 5168
rect 15857 5158 16015 5168
rect 16019 5158 16049 5168
rect 16053 5158 16083 5172
rect 16111 5158 16124 5196
rect 16196 5210 16225 5226
rect 16239 5210 16268 5226
rect 16283 5216 16313 5232
rect 16341 5210 16347 5258
rect 16350 5252 16369 5258
rect 16384 5252 16414 5260
rect 16350 5244 16414 5252
rect 16350 5228 16430 5244
rect 16446 5237 16508 5268
rect 16524 5237 16586 5268
rect 16655 5266 16704 5291
rect 16719 5266 16749 5282
rect 16618 5252 16648 5260
rect 16655 5258 16765 5266
rect 16618 5244 16663 5252
rect 16350 5226 16369 5228
rect 16384 5226 16430 5228
rect 16350 5210 16430 5226
rect 16457 5224 16492 5237
rect 16533 5234 16570 5237
rect 16533 5232 16575 5234
rect 16462 5221 16492 5224
rect 16471 5217 16478 5221
rect 16478 5216 16479 5217
rect 16437 5210 16447 5216
rect 16196 5202 16231 5210
rect 16196 5176 16197 5202
rect 16204 5176 16231 5202
rect 16139 5158 16169 5172
rect 16196 5168 16231 5176
rect 16233 5202 16274 5210
rect 16233 5176 16248 5202
rect 16255 5176 16274 5202
rect 16338 5198 16369 5210
rect 16384 5198 16487 5210
rect 16499 5200 16525 5226
rect 16540 5221 16570 5232
rect 16602 5228 16664 5244
rect 16602 5226 16648 5228
rect 16602 5210 16664 5226
rect 16676 5210 16682 5258
rect 16685 5250 16765 5258
rect 16685 5248 16704 5250
rect 16719 5248 16753 5250
rect 16685 5232 16765 5248
rect 16685 5210 16704 5232
rect 16719 5216 16749 5232
rect 16777 5226 16783 5300
rect 16786 5226 16805 5370
rect 16820 5226 16826 5370
rect 16835 5300 16848 5370
rect 16900 5366 16922 5370
rect 16893 5344 16922 5358
rect 16975 5344 16991 5358
rect 17029 5354 17035 5356
rect 17042 5354 17150 5370
rect 17157 5354 17163 5356
rect 17171 5354 17186 5370
rect 17252 5364 17271 5367
rect 16893 5342 16991 5344
rect 17018 5342 17186 5354
rect 17201 5344 17217 5358
rect 17252 5345 17274 5364
rect 17284 5358 17300 5359
rect 17283 5356 17300 5358
rect 17284 5351 17300 5356
rect 17274 5344 17280 5345
rect 17283 5344 17312 5351
rect 17201 5343 17312 5344
rect 17201 5342 17318 5343
rect 16877 5334 16928 5342
rect 16975 5334 17009 5342
rect 16877 5322 16902 5334
rect 16909 5322 16928 5334
rect 16982 5332 17009 5334
rect 17018 5332 17239 5342
rect 17274 5339 17280 5342
rect 16982 5328 17239 5332
rect 16877 5314 16928 5322
rect 16975 5314 17239 5328
rect 17283 5334 17318 5342
rect 16829 5266 16848 5300
rect 16893 5306 16922 5314
rect 16893 5300 16910 5306
rect 16893 5298 16927 5300
rect 16975 5298 16991 5314
rect 16992 5304 17200 5314
rect 17201 5304 17217 5314
rect 17265 5310 17280 5325
rect 17283 5322 17284 5334
rect 17291 5322 17318 5334
rect 17283 5314 17318 5322
rect 17283 5313 17312 5314
rect 17003 5300 17217 5304
rect 17018 5298 17217 5300
rect 17252 5300 17265 5310
rect 17283 5300 17300 5313
rect 17252 5298 17300 5300
rect 16894 5294 16927 5298
rect 16890 5292 16927 5294
rect 16890 5291 16957 5292
rect 16890 5286 16921 5291
rect 16927 5286 16957 5291
rect 16890 5282 16957 5286
rect 16863 5279 16957 5282
rect 16863 5272 16912 5279
rect 16863 5266 16893 5272
rect 16912 5267 16917 5272
rect 16829 5250 16909 5266
rect 16921 5258 16957 5279
rect 17018 5274 17207 5298
rect 17252 5297 17299 5298
rect 17265 5292 17299 5297
rect 17033 5271 17207 5274
rect 17026 5268 17207 5271
rect 17235 5291 17299 5292
rect 16829 5248 16848 5250
rect 16863 5248 16897 5250
rect 16829 5232 16909 5248
rect 16829 5226 16848 5232
rect 16545 5200 16648 5210
rect 16499 5198 16648 5200
rect 16669 5198 16704 5210
rect 16338 5196 16500 5198
rect 16350 5176 16369 5196
rect 16384 5194 16414 5196
rect 16233 5168 16274 5176
rect 16356 5172 16369 5176
rect 16421 5180 16500 5196
rect 16532 5196 16704 5198
rect 16532 5180 16611 5196
rect 16618 5194 16648 5196
rect 16196 5158 16225 5168
rect 16239 5158 16268 5168
rect 16283 5158 16313 5172
rect 16356 5158 16399 5172
rect 16421 5168 16611 5180
rect 16676 5176 16682 5196
rect 16406 5158 16436 5168
rect 16437 5158 16595 5168
rect 16599 5158 16629 5168
rect 16633 5158 16663 5172
rect 16691 5158 16704 5196
rect 16776 5210 16805 5226
rect 16819 5210 16848 5226
rect 16863 5216 16893 5232
rect 16921 5210 16927 5258
rect 16930 5252 16949 5258
rect 16964 5252 16994 5260
rect 16930 5244 16994 5252
rect 16930 5228 17010 5244
rect 17026 5237 17088 5268
rect 17104 5237 17166 5268
rect 17235 5266 17284 5291
rect 17299 5266 17329 5282
rect 17198 5252 17228 5260
rect 17235 5258 17345 5266
rect 17198 5244 17243 5252
rect 16930 5226 16949 5228
rect 16964 5226 17010 5228
rect 16930 5210 17010 5226
rect 17037 5224 17072 5237
rect 17113 5234 17150 5237
rect 17113 5232 17155 5234
rect 17042 5221 17072 5224
rect 17051 5217 17058 5221
rect 17058 5216 17059 5217
rect 17017 5210 17027 5216
rect 16776 5202 16811 5210
rect 16776 5176 16777 5202
rect 16784 5176 16811 5202
rect 16719 5158 16749 5172
rect 16776 5168 16811 5176
rect 16813 5202 16854 5210
rect 16813 5176 16828 5202
rect 16835 5176 16854 5202
rect 16918 5198 16949 5210
rect 16964 5198 17067 5210
rect 17079 5200 17105 5226
rect 17120 5221 17150 5232
rect 17182 5228 17244 5244
rect 17182 5226 17228 5228
rect 17182 5210 17244 5226
rect 17256 5210 17262 5258
rect 17265 5250 17345 5258
rect 17265 5248 17284 5250
rect 17299 5248 17333 5250
rect 17265 5232 17345 5248
rect 17265 5210 17284 5232
rect 17299 5216 17329 5232
rect 17357 5226 17363 5300
rect 17366 5226 17385 5370
rect 17400 5226 17406 5370
rect 17415 5300 17428 5370
rect 17480 5366 17502 5370
rect 17473 5344 17502 5358
rect 17555 5344 17571 5358
rect 17609 5354 17615 5356
rect 17622 5354 17730 5370
rect 17737 5354 17743 5356
rect 17751 5354 17766 5370
rect 17832 5364 17851 5367
rect 17473 5342 17571 5344
rect 17598 5342 17766 5354
rect 17781 5344 17797 5358
rect 17832 5345 17854 5364
rect 17864 5358 17880 5359
rect 17863 5356 17880 5358
rect 17864 5351 17880 5356
rect 17854 5344 17860 5345
rect 17863 5344 17892 5351
rect 17781 5343 17892 5344
rect 17781 5342 17898 5343
rect 17457 5334 17508 5342
rect 17555 5334 17589 5342
rect 17457 5322 17482 5334
rect 17489 5322 17508 5334
rect 17562 5332 17589 5334
rect 17598 5332 17819 5342
rect 17854 5339 17860 5342
rect 17562 5328 17819 5332
rect 17457 5314 17508 5322
rect 17555 5314 17819 5328
rect 17863 5334 17898 5342
rect 17409 5266 17428 5300
rect 17473 5306 17502 5314
rect 17473 5300 17490 5306
rect 17473 5298 17507 5300
rect 17555 5298 17571 5314
rect 17572 5304 17780 5314
rect 17781 5304 17797 5314
rect 17845 5310 17860 5325
rect 17863 5322 17864 5334
rect 17871 5322 17898 5334
rect 17863 5314 17898 5322
rect 17863 5313 17892 5314
rect 17583 5300 17797 5304
rect 17598 5298 17797 5300
rect 17832 5300 17845 5310
rect 17863 5300 17880 5313
rect 17832 5298 17880 5300
rect 17474 5294 17507 5298
rect 17470 5292 17507 5294
rect 17470 5291 17537 5292
rect 17470 5286 17501 5291
rect 17507 5286 17537 5291
rect 17470 5282 17537 5286
rect 17443 5279 17537 5282
rect 17443 5272 17492 5279
rect 17443 5266 17473 5272
rect 17492 5267 17497 5272
rect 17409 5250 17489 5266
rect 17501 5258 17537 5279
rect 17598 5274 17787 5298
rect 17832 5297 17879 5298
rect 17845 5292 17879 5297
rect 17613 5271 17787 5274
rect 17606 5268 17787 5271
rect 17815 5291 17879 5292
rect 17409 5248 17428 5250
rect 17443 5248 17477 5250
rect 17409 5232 17489 5248
rect 17409 5226 17428 5232
rect 17125 5200 17228 5210
rect 17079 5198 17228 5200
rect 17249 5198 17284 5210
rect 16918 5196 17080 5198
rect 16930 5176 16949 5196
rect 16964 5194 16994 5196
rect 16813 5168 16854 5176
rect 16936 5172 16949 5176
rect 17001 5180 17080 5196
rect 17112 5196 17284 5198
rect 17112 5180 17191 5196
rect 17198 5194 17228 5196
rect 16776 5158 16805 5168
rect 16819 5158 16848 5168
rect 16863 5158 16893 5172
rect 16936 5158 16979 5172
rect 17001 5168 17191 5180
rect 17256 5176 17262 5196
rect 16986 5158 17016 5168
rect 17017 5158 17175 5168
rect 17179 5158 17209 5168
rect 17213 5158 17243 5172
rect 17271 5158 17284 5196
rect 17356 5210 17385 5226
rect 17399 5210 17428 5226
rect 17443 5216 17473 5232
rect 17501 5210 17507 5258
rect 17510 5252 17529 5258
rect 17544 5252 17574 5260
rect 17510 5244 17574 5252
rect 17510 5228 17590 5244
rect 17606 5237 17668 5268
rect 17684 5237 17746 5268
rect 17815 5266 17864 5291
rect 17879 5266 17909 5282
rect 17778 5252 17808 5260
rect 17815 5258 17925 5266
rect 17778 5244 17823 5252
rect 17510 5226 17529 5228
rect 17544 5226 17590 5228
rect 17510 5210 17590 5226
rect 17617 5224 17652 5237
rect 17693 5234 17730 5237
rect 17693 5232 17735 5234
rect 17622 5221 17652 5224
rect 17631 5217 17638 5221
rect 17638 5216 17639 5217
rect 17597 5210 17607 5216
rect 17356 5202 17391 5210
rect 17356 5176 17357 5202
rect 17364 5176 17391 5202
rect 17299 5158 17329 5172
rect 17356 5168 17391 5176
rect 17393 5202 17434 5210
rect 17393 5176 17408 5202
rect 17415 5176 17434 5202
rect 17498 5198 17529 5210
rect 17544 5198 17647 5210
rect 17659 5200 17685 5226
rect 17700 5221 17730 5232
rect 17762 5228 17824 5244
rect 17762 5226 17808 5228
rect 17762 5210 17824 5226
rect 17836 5210 17842 5258
rect 17845 5250 17925 5258
rect 17845 5248 17864 5250
rect 17879 5248 17913 5250
rect 17845 5232 17925 5248
rect 17845 5210 17864 5232
rect 17879 5216 17909 5232
rect 17937 5226 17943 5300
rect 17946 5226 17965 5370
rect 17980 5226 17986 5370
rect 17995 5300 18008 5370
rect 18060 5366 18082 5370
rect 18053 5344 18082 5358
rect 18135 5344 18151 5358
rect 18189 5354 18195 5356
rect 18202 5354 18310 5370
rect 18317 5354 18323 5356
rect 18331 5354 18346 5370
rect 18412 5364 18431 5367
rect 18053 5342 18151 5344
rect 18178 5342 18346 5354
rect 18361 5344 18377 5358
rect 18412 5345 18434 5364
rect 18444 5358 18460 5359
rect 18443 5356 18460 5358
rect 18444 5351 18460 5356
rect 18434 5344 18440 5345
rect 18443 5344 18472 5351
rect 18361 5343 18472 5344
rect 18361 5342 18478 5343
rect 18037 5334 18088 5342
rect 18135 5334 18169 5342
rect 18037 5322 18062 5334
rect 18069 5322 18088 5334
rect 18142 5332 18169 5334
rect 18178 5332 18399 5342
rect 18434 5339 18440 5342
rect 18142 5328 18399 5332
rect 18037 5314 18088 5322
rect 18135 5314 18399 5328
rect 18443 5334 18478 5342
rect 17989 5266 18008 5300
rect 18053 5306 18082 5314
rect 18053 5300 18070 5306
rect 18053 5298 18087 5300
rect 18135 5298 18151 5314
rect 18152 5304 18360 5314
rect 18361 5304 18377 5314
rect 18425 5310 18440 5325
rect 18443 5322 18444 5334
rect 18451 5322 18478 5334
rect 18443 5314 18478 5322
rect 18443 5313 18472 5314
rect 18163 5300 18377 5304
rect 18178 5298 18377 5300
rect 18412 5300 18425 5310
rect 18443 5300 18460 5313
rect 18412 5298 18460 5300
rect 18054 5294 18087 5298
rect 18050 5292 18087 5294
rect 18050 5291 18117 5292
rect 18050 5286 18081 5291
rect 18087 5286 18117 5291
rect 18050 5282 18117 5286
rect 18023 5279 18117 5282
rect 18023 5272 18072 5279
rect 18023 5266 18053 5272
rect 18072 5267 18077 5272
rect 17989 5250 18069 5266
rect 18081 5258 18117 5279
rect 18178 5274 18367 5298
rect 18412 5297 18459 5298
rect 18425 5292 18459 5297
rect 18193 5271 18367 5274
rect 18186 5268 18367 5271
rect 18395 5291 18459 5292
rect 17989 5248 18008 5250
rect 18023 5248 18057 5250
rect 17989 5232 18069 5248
rect 17989 5226 18008 5232
rect 17705 5200 17808 5210
rect 17659 5198 17808 5200
rect 17829 5198 17864 5210
rect 17498 5196 17660 5198
rect 17510 5176 17529 5196
rect 17544 5194 17574 5196
rect 17393 5168 17434 5176
rect 17516 5172 17529 5176
rect 17581 5180 17660 5196
rect 17692 5196 17864 5198
rect 17692 5180 17771 5196
rect 17778 5194 17808 5196
rect 17356 5158 17385 5168
rect 17399 5158 17428 5168
rect 17443 5158 17473 5172
rect 17516 5158 17559 5172
rect 17581 5168 17771 5180
rect 17836 5176 17842 5196
rect 17566 5158 17596 5168
rect 17597 5158 17755 5168
rect 17759 5158 17789 5168
rect 17793 5158 17823 5172
rect 17851 5158 17864 5196
rect 17936 5210 17965 5226
rect 17979 5210 18008 5226
rect 18023 5216 18053 5232
rect 18081 5210 18087 5258
rect 18090 5252 18109 5258
rect 18124 5252 18154 5260
rect 18090 5244 18154 5252
rect 18090 5228 18170 5244
rect 18186 5237 18248 5268
rect 18264 5237 18326 5268
rect 18395 5266 18444 5291
rect 18459 5266 18489 5282
rect 18358 5252 18388 5260
rect 18395 5258 18505 5266
rect 18358 5244 18403 5252
rect 18090 5226 18109 5228
rect 18124 5226 18170 5228
rect 18090 5210 18170 5226
rect 18197 5224 18232 5237
rect 18273 5234 18310 5237
rect 18273 5232 18315 5234
rect 18202 5221 18232 5224
rect 18211 5217 18218 5221
rect 18218 5216 18219 5217
rect 18177 5210 18187 5216
rect 17936 5202 17971 5210
rect 17936 5176 17937 5202
rect 17944 5176 17971 5202
rect 17879 5158 17909 5172
rect 17936 5168 17971 5176
rect 17973 5202 18014 5210
rect 17973 5176 17988 5202
rect 17995 5176 18014 5202
rect 18078 5198 18109 5210
rect 18124 5198 18227 5210
rect 18239 5200 18265 5226
rect 18280 5221 18310 5232
rect 18342 5228 18404 5244
rect 18342 5226 18388 5228
rect 18342 5210 18404 5226
rect 18416 5210 18422 5258
rect 18425 5250 18505 5258
rect 18425 5248 18444 5250
rect 18459 5248 18493 5250
rect 18425 5232 18505 5248
rect 18425 5210 18444 5232
rect 18459 5216 18489 5232
rect 18517 5226 18523 5300
rect 18532 5226 18545 5370
rect 18285 5200 18388 5210
rect 18239 5198 18388 5200
rect 18409 5198 18444 5210
rect 18078 5196 18240 5198
rect 18090 5176 18109 5196
rect 18124 5194 18154 5196
rect 17973 5168 18014 5176
rect 18096 5172 18109 5176
rect 18161 5180 18240 5196
rect 18272 5196 18444 5198
rect 18272 5180 18351 5196
rect 18358 5194 18388 5196
rect 17936 5158 17965 5168
rect 17979 5158 18008 5168
rect 18023 5158 18053 5172
rect 18096 5158 18139 5172
rect 18161 5168 18351 5180
rect 18416 5176 18422 5196
rect 18146 5158 18176 5168
rect 18177 5158 18335 5168
rect 18339 5158 18369 5168
rect 18373 5158 18403 5172
rect 18431 5158 18444 5196
rect 18516 5210 18545 5226
rect 18516 5202 18551 5210
rect 18516 5176 18517 5202
rect 18524 5176 18551 5202
rect 18459 5158 18489 5172
rect 18516 5168 18551 5176
rect 18516 5158 18545 5168
rect -1 5152 18545 5158
rect 0 5144 18545 5152
rect 15 5114 28 5144
rect 43 5130 73 5144
rect 116 5130 159 5144
rect 166 5130 386 5144
rect 393 5130 423 5144
rect 83 5116 98 5128
rect 117 5116 130 5130
rect 198 5126 351 5130
rect 80 5114 102 5116
rect 180 5114 372 5126
rect 451 5114 464 5144
rect 479 5130 509 5144
rect 546 5114 565 5144
rect 580 5114 586 5144
rect 595 5114 608 5144
rect 623 5130 653 5144
rect 696 5130 739 5144
rect 746 5130 966 5144
rect 973 5130 1003 5144
rect 663 5116 678 5128
rect 697 5116 710 5130
rect 778 5126 931 5130
rect 660 5114 682 5116
rect 760 5114 952 5126
rect 1031 5114 1044 5144
rect 1059 5130 1089 5144
rect 1126 5114 1145 5144
rect 1160 5114 1166 5144
rect 1175 5114 1188 5144
rect 1203 5130 1233 5144
rect 1276 5130 1319 5144
rect 1326 5130 1546 5144
rect 1553 5130 1583 5144
rect 1243 5116 1258 5128
rect 1277 5116 1290 5130
rect 1358 5126 1511 5130
rect 1240 5114 1262 5116
rect 1340 5114 1532 5126
rect 1611 5114 1624 5144
rect 1639 5130 1669 5144
rect 1706 5114 1725 5144
rect 1740 5114 1746 5144
rect 1755 5114 1768 5144
rect 1783 5130 1813 5144
rect 1856 5130 1899 5144
rect 1906 5130 2126 5144
rect 2133 5130 2163 5144
rect 1823 5116 1838 5128
rect 1857 5116 1870 5130
rect 1938 5126 2091 5130
rect 1820 5114 1842 5116
rect 1920 5114 2112 5126
rect 2191 5114 2204 5144
rect 2219 5130 2249 5144
rect 2286 5114 2305 5144
rect 2320 5114 2326 5144
rect 2335 5114 2348 5144
rect 2363 5130 2393 5144
rect 2436 5130 2479 5144
rect 2486 5130 2706 5144
rect 2713 5130 2743 5144
rect 2403 5116 2418 5128
rect 2437 5116 2450 5130
rect 2518 5126 2671 5130
rect 2400 5114 2422 5116
rect 2500 5114 2692 5126
rect 2771 5114 2784 5144
rect 2799 5130 2829 5144
rect 2866 5114 2885 5144
rect 2900 5114 2906 5144
rect 2915 5114 2928 5144
rect 2943 5130 2973 5144
rect 3016 5130 3059 5144
rect 3066 5130 3286 5144
rect 3293 5130 3323 5144
rect 2983 5116 2998 5128
rect 3017 5116 3030 5130
rect 3098 5126 3251 5130
rect 2980 5114 3002 5116
rect 3080 5114 3272 5126
rect 3351 5114 3364 5144
rect 3379 5130 3409 5144
rect 3446 5114 3465 5144
rect 3480 5114 3486 5144
rect 3495 5114 3508 5144
rect 3523 5130 3553 5144
rect 3596 5130 3639 5144
rect 3646 5130 3866 5144
rect 3873 5130 3903 5144
rect 3563 5116 3578 5128
rect 3597 5116 3610 5130
rect 3678 5126 3831 5130
rect 3560 5114 3582 5116
rect 3660 5114 3852 5126
rect 3931 5114 3944 5144
rect 3959 5130 3989 5144
rect 4026 5114 4045 5144
rect 4060 5114 4066 5144
rect 4075 5114 4088 5144
rect 4103 5130 4133 5144
rect 4176 5130 4219 5144
rect 4226 5130 4446 5144
rect 4453 5130 4483 5144
rect 4143 5116 4158 5128
rect 4177 5116 4190 5130
rect 4258 5126 4411 5130
rect 4140 5114 4162 5116
rect 4240 5114 4432 5126
rect 4511 5114 4524 5144
rect 4539 5130 4569 5144
rect 4606 5114 4625 5144
rect 4640 5114 4646 5144
rect 4655 5114 4668 5144
rect 4683 5130 4713 5144
rect 4756 5130 4799 5144
rect 4806 5130 5026 5144
rect 5033 5130 5063 5144
rect 4723 5116 4738 5128
rect 4757 5116 4770 5130
rect 4838 5126 4991 5130
rect 4720 5114 4742 5116
rect 4820 5114 5012 5126
rect 5091 5114 5104 5144
rect 5119 5130 5149 5144
rect 5186 5114 5205 5144
rect 5220 5114 5226 5144
rect 5235 5114 5248 5144
rect 5263 5130 5293 5144
rect 5336 5130 5379 5144
rect 5386 5130 5606 5144
rect 5613 5130 5643 5144
rect 5303 5116 5318 5128
rect 5337 5116 5350 5130
rect 5418 5126 5571 5130
rect 5300 5114 5322 5116
rect 5400 5114 5592 5126
rect 5671 5114 5684 5144
rect 5699 5130 5729 5144
rect 5766 5114 5785 5144
rect 5800 5114 5806 5144
rect 5815 5114 5828 5144
rect 5843 5130 5873 5144
rect 5916 5130 5959 5144
rect 5966 5130 6186 5144
rect 6193 5130 6223 5144
rect 5883 5116 5898 5128
rect 5917 5116 5930 5130
rect 5998 5126 6151 5130
rect 5880 5114 5902 5116
rect 5980 5114 6172 5126
rect 6251 5114 6264 5144
rect 6279 5130 6309 5144
rect 6346 5114 6365 5144
rect 6380 5114 6386 5144
rect 6395 5114 6408 5144
rect 6423 5130 6453 5144
rect 6496 5130 6539 5144
rect 6546 5130 6766 5144
rect 6773 5130 6803 5144
rect 6463 5116 6478 5128
rect 6497 5116 6510 5130
rect 6578 5126 6731 5130
rect 6460 5114 6482 5116
rect 6560 5114 6752 5126
rect 6831 5114 6844 5144
rect 6859 5130 6889 5144
rect 6926 5114 6945 5144
rect 6960 5114 6966 5144
rect 6975 5114 6988 5144
rect 7003 5130 7033 5144
rect 7076 5130 7119 5144
rect 7126 5130 7346 5144
rect 7353 5130 7383 5144
rect 7043 5116 7058 5128
rect 7077 5116 7090 5130
rect 7158 5126 7311 5130
rect 7040 5114 7062 5116
rect 7140 5114 7332 5126
rect 7411 5114 7424 5144
rect 7439 5130 7469 5144
rect 7506 5114 7525 5144
rect 7540 5114 7546 5144
rect 7555 5114 7568 5144
rect 7583 5130 7613 5144
rect 7656 5130 7699 5144
rect 7706 5130 7926 5144
rect 7933 5130 7963 5144
rect 7623 5116 7638 5128
rect 7657 5116 7670 5130
rect 7738 5126 7891 5130
rect 7620 5114 7642 5116
rect 7720 5114 7912 5126
rect 7991 5114 8004 5144
rect 8019 5130 8049 5144
rect 8086 5114 8105 5144
rect 8120 5114 8126 5144
rect 8135 5114 8148 5144
rect 8163 5130 8193 5144
rect 8236 5130 8279 5144
rect 8286 5130 8506 5144
rect 8513 5130 8543 5144
rect 8203 5116 8218 5128
rect 8237 5116 8250 5130
rect 8318 5126 8471 5130
rect 8200 5114 8222 5116
rect 8300 5114 8492 5126
rect 8571 5114 8584 5144
rect 8599 5130 8629 5144
rect 8666 5114 8685 5144
rect 8700 5114 8706 5144
rect 8715 5114 8728 5144
rect 8743 5130 8773 5144
rect 8816 5130 8859 5144
rect 8866 5130 9086 5144
rect 9093 5130 9123 5144
rect 8783 5116 8798 5128
rect 8817 5116 8830 5130
rect 8898 5126 9051 5130
rect 8780 5114 8802 5116
rect 8880 5114 9072 5126
rect 9151 5114 9164 5144
rect 9179 5130 9209 5144
rect 9246 5114 9265 5144
rect 9280 5114 9286 5144
rect 9295 5114 9308 5144
rect 9323 5130 9353 5144
rect 9396 5130 9439 5144
rect 9446 5130 9666 5144
rect 9673 5130 9703 5144
rect 9363 5116 9378 5128
rect 9397 5116 9410 5130
rect 9478 5126 9631 5130
rect 9360 5114 9382 5116
rect 9460 5114 9652 5126
rect 9731 5114 9744 5144
rect 9759 5130 9789 5144
rect 9826 5114 9845 5144
rect 9860 5114 9866 5144
rect 9875 5114 9888 5144
rect 9903 5130 9933 5144
rect 9976 5130 10019 5144
rect 10026 5130 10246 5144
rect 10253 5130 10283 5144
rect 9943 5116 9958 5128
rect 9977 5116 9990 5130
rect 10058 5126 10211 5130
rect 9940 5114 9962 5116
rect 10040 5114 10232 5126
rect 10311 5114 10324 5144
rect 10339 5130 10369 5144
rect 10406 5114 10425 5144
rect 10440 5114 10446 5144
rect 10455 5114 10468 5144
rect 10483 5130 10513 5144
rect 10556 5130 10599 5144
rect 10606 5130 10826 5144
rect 10833 5130 10863 5144
rect 10523 5116 10538 5128
rect 10557 5116 10570 5130
rect 10638 5126 10791 5130
rect 10520 5114 10542 5116
rect 10620 5114 10812 5126
rect 10891 5114 10904 5144
rect 10919 5130 10949 5144
rect 10986 5114 11005 5144
rect 11020 5114 11026 5144
rect 11035 5114 11048 5144
rect 11063 5130 11093 5144
rect 11136 5130 11179 5144
rect 11186 5130 11406 5144
rect 11413 5130 11443 5144
rect 11103 5116 11118 5128
rect 11137 5116 11150 5130
rect 11218 5126 11371 5130
rect 11100 5114 11122 5116
rect 11200 5114 11392 5126
rect 11471 5114 11484 5144
rect 11499 5130 11529 5144
rect 11566 5114 11585 5144
rect 11600 5114 11606 5144
rect 11615 5114 11628 5144
rect 11643 5130 11673 5144
rect 11716 5130 11759 5144
rect 11766 5130 11986 5144
rect 11993 5130 12023 5144
rect 11683 5116 11698 5128
rect 11717 5116 11730 5130
rect 11798 5126 11951 5130
rect 11680 5114 11702 5116
rect 11780 5114 11972 5126
rect 12051 5114 12064 5144
rect 12079 5130 12109 5144
rect 12146 5114 12165 5144
rect 12180 5114 12186 5144
rect 12195 5114 12208 5144
rect 12223 5130 12253 5144
rect 12296 5130 12339 5144
rect 12346 5130 12566 5144
rect 12573 5130 12603 5144
rect 12263 5116 12278 5128
rect 12297 5116 12310 5130
rect 12378 5126 12531 5130
rect 12260 5114 12282 5116
rect 12360 5114 12552 5126
rect 12631 5114 12644 5144
rect 12659 5130 12689 5144
rect 12726 5114 12745 5144
rect 12760 5114 12766 5144
rect 12775 5114 12788 5144
rect 12803 5130 12833 5144
rect 12876 5130 12919 5144
rect 12926 5130 13146 5144
rect 13153 5130 13183 5144
rect 12843 5116 12858 5128
rect 12877 5116 12890 5130
rect 12958 5126 13111 5130
rect 12840 5114 12862 5116
rect 12940 5114 13132 5126
rect 13211 5114 13224 5144
rect 13239 5130 13269 5144
rect 13306 5114 13325 5144
rect 13340 5114 13346 5144
rect 13355 5114 13368 5144
rect 13383 5130 13413 5144
rect 13456 5130 13499 5144
rect 13506 5130 13726 5144
rect 13733 5130 13763 5144
rect 13423 5116 13438 5128
rect 13457 5116 13470 5130
rect 13538 5126 13691 5130
rect 13420 5114 13442 5116
rect 13520 5114 13712 5126
rect 13791 5114 13804 5144
rect 13819 5130 13849 5144
rect 13886 5114 13905 5144
rect 13920 5114 13926 5144
rect 13935 5114 13948 5144
rect 13963 5130 13993 5144
rect 14036 5130 14079 5144
rect 14086 5130 14306 5144
rect 14313 5130 14343 5144
rect 14003 5116 14018 5128
rect 14037 5116 14050 5130
rect 14118 5126 14271 5130
rect 14000 5114 14022 5116
rect 14100 5114 14292 5126
rect 14371 5114 14384 5144
rect 14399 5130 14429 5144
rect 14466 5114 14485 5144
rect 14500 5114 14506 5144
rect 14515 5114 14528 5144
rect 14543 5130 14573 5144
rect 14616 5130 14659 5144
rect 14666 5130 14886 5144
rect 14893 5130 14923 5144
rect 14583 5116 14598 5128
rect 14617 5116 14630 5130
rect 14698 5126 14851 5130
rect 14580 5114 14602 5116
rect 14680 5114 14872 5126
rect 14951 5114 14964 5144
rect 14979 5130 15009 5144
rect 15046 5114 15065 5144
rect 15080 5114 15086 5144
rect 15095 5114 15108 5144
rect 15123 5130 15153 5144
rect 15196 5130 15239 5144
rect 15246 5130 15466 5144
rect 15473 5130 15503 5144
rect 15163 5116 15178 5128
rect 15197 5116 15210 5130
rect 15278 5126 15431 5130
rect 15160 5114 15182 5116
rect 15260 5114 15452 5126
rect 15531 5114 15544 5144
rect 15559 5130 15589 5144
rect 15626 5114 15645 5144
rect 15660 5114 15666 5144
rect 15675 5114 15688 5144
rect 15703 5130 15733 5144
rect 15776 5130 15819 5144
rect 15826 5130 16046 5144
rect 16053 5130 16083 5144
rect 15743 5116 15758 5128
rect 15777 5116 15790 5130
rect 15858 5126 16011 5130
rect 15740 5114 15762 5116
rect 15840 5114 16032 5126
rect 16111 5114 16124 5144
rect 16139 5130 16169 5144
rect 16206 5114 16225 5144
rect 16240 5114 16246 5144
rect 16255 5114 16268 5144
rect 16283 5130 16313 5144
rect 16356 5130 16399 5144
rect 16406 5130 16626 5144
rect 16633 5130 16663 5144
rect 16323 5116 16338 5128
rect 16357 5116 16370 5130
rect 16438 5126 16591 5130
rect 16320 5114 16342 5116
rect 16420 5114 16612 5126
rect 16691 5114 16704 5144
rect 16719 5130 16749 5144
rect 16786 5114 16805 5144
rect 16820 5114 16826 5144
rect 16835 5114 16848 5144
rect 16863 5130 16893 5144
rect 16936 5130 16979 5144
rect 16986 5130 17206 5144
rect 17213 5130 17243 5144
rect 16903 5116 16918 5128
rect 16937 5116 16950 5130
rect 17018 5126 17171 5130
rect 16900 5114 16922 5116
rect 17000 5114 17192 5126
rect 17271 5114 17284 5144
rect 17299 5130 17329 5144
rect 17366 5114 17385 5144
rect 17400 5114 17406 5144
rect 17415 5114 17428 5144
rect 17443 5130 17473 5144
rect 17516 5130 17559 5144
rect 17566 5130 17786 5144
rect 17793 5130 17823 5144
rect 17483 5116 17498 5128
rect 17517 5116 17530 5130
rect 17598 5126 17751 5130
rect 17480 5114 17502 5116
rect 17580 5114 17772 5126
rect 17851 5114 17864 5144
rect 17879 5130 17909 5144
rect 17946 5114 17965 5144
rect 17980 5114 17986 5144
rect 17995 5114 18008 5144
rect 18023 5130 18053 5144
rect 18096 5130 18139 5144
rect 18146 5130 18366 5144
rect 18373 5130 18403 5144
rect 18063 5116 18078 5128
rect 18097 5116 18110 5130
rect 18178 5126 18331 5130
rect 18060 5114 18082 5116
rect 18160 5114 18352 5126
rect 18431 5114 18444 5144
rect 18459 5130 18489 5144
rect 18532 5114 18545 5144
rect 0 5100 18545 5114
rect 15 5030 28 5100
rect 80 5096 102 5100
rect 73 5074 102 5088
rect 155 5074 171 5088
rect 209 5084 215 5086
rect 222 5084 330 5100
rect 337 5084 343 5086
rect 351 5084 366 5100
rect 432 5094 451 5097
rect 73 5072 171 5074
rect 198 5072 366 5084
rect 381 5074 397 5088
rect 432 5075 454 5094
rect 464 5088 480 5089
rect 463 5086 480 5088
rect 464 5081 480 5086
rect 454 5074 460 5075
rect 463 5074 492 5081
rect 381 5073 492 5074
rect 381 5072 498 5073
rect 57 5064 108 5072
rect 155 5064 189 5072
rect 57 5052 82 5064
rect 89 5052 108 5064
rect 162 5062 189 5064
rect 198 5062 419 5072
rect 454 5069 460 5072
rect 162 5058 419 5062
rect 57 5044 108 5052
rect 155 5044 419 5058
rect 463 5064 498 5072
rect 9 4996 28 5030
rect 73 5036 102 5044
rect 73 5030 90 5036
rect 73 5028 107 5030
rect 155 5028 171 5044
rect 172 5034 380 5044
rect 381 5034 397 5044
rect 445 5040 460 5055
rect 463 5052 464 5064
rect 471 5052 498 5064
rect 463 5044 498 5052
rect 463 5043 492 5044
rect 183 5030 397 5034
rect 198 5028 397 5030
rect 432 5030 445 5040
rect 463 5030 480 5043
rect 432 5028 480 5030
rect 74 5024 107 5028
rect 70 5022 107 5024
rect 70 5021 137 5022
rect 70 5016 101 5021
rect 107 5016 137 5021
rect 70 5012 137 5016
rect 43 5009 137 5012
rect 43 5002 92 5009
rect 43 4996 73 5002
rect 92 4997 97 5002
rect 9 4980 89 4996
rect 101 4988 137 5009
rect 198 5004 387 5028
rect 432 5027 479 5028
rect 445 5022 479 5027
rect 213 5001 387 5004
rect 206 4998 387 5001
rect 415 5021 479 5022
rect 9 4978 28 4980
rect 43 4978 77 4980
rect 9 4962 89 4978
rect 9 4956 28 4962
rect -1 4940 28 4956
rect 43 4946 73 4962
rect 101 4940 107 4988
rect 110 4982 129 4988
rect 144 4982 174 4990
rect 110 4974 174 4982
rect 110 4958 190 4974
rect 206 4967 268 4998
rect 284 4967 346 4998
rect 415 4996 464 5021
rect 479 4996 509 5012
rect 378 4982 408 4990
rect 415 4988 525 4996
rect 378 4974 423 4982
rect 110 4956 129 4958
rect 144 4956 190 4958
rect 110 4940 190 4956
rect 217 4954 252 4967
rect 293 4964 330 4967
rect 293 4962 335 4964
rect 222 4951 252 4954
rect 231 4947 238 4951
rect 238 4946 239 4947
rect 197 4940 207 4946
rect -7 4932 34 4940
rect -7 4906 8 4932
rect 15 4906 34 4932
rect 98 4928 129 4940
rect 144 4928 247 4940
rect 259 4930 285 4956
rect 300 4951 330 4962
rect 362 4958 424 4974
rect 362 4956 408 4958
rect 362 4940 424 4956
rect 436 4940 442 4988
rect 445 4980 525 4988
rect 445 4978 464 4980
rect 479 4978 513 4980
rect 445 4962 525 4978
rect 445 4940 464 4962
rect 479 4946 509 4962
rect 537 4956 543 5030
rect 546 4956 565 5100
rect 580 4956 586 5100
rect 595 5030 608 5100
rect 660 5096 682 5100
rect 653 5074 682 5088
rect 735 5074 751 5088
rect 789 5084 795 5086
rect 802 5084 910 5100
rect 917 5084 923 5086
rect 931 5084 946 5100
rect 1012 5094 1031 5097
rect 653 5072 751 5074
rect 778 5072 946 5084
rect 961 5074 977 5088
rect 1012 5075 1034 5094
rect 1044 5088 1060 5089
rect 1043 5086 1060 5088
rect 1044 5081 1060 5086
rect 1034 5074 1040 5075
rect 1043 5074 1072 5081
rect 961 5073 1072 5074
rect 961 5072 1078 5073
rect 637 5064 688 5072
rect 735 5064 769 5072
rect 637 5052 662 5064
rect 669 5052 688 5064
rect 742 5062 769 5064
rect 778 5062 999 5072
rect 1034 5069 1040 5072
rect 742 5058 999 5062
rect 637 5044 688 5052
rect 735 5044 999 5058
rect 1043 5064 1078 5072
rect 589 4996 608 5030
rect 653 5036 682 5044
rect 653 5030 670 5036
rect 653 5028 687 5030
rect 735 5028 751 5044
rect 752 5034 960 5044
rect 961 5034 977 5044
rect 1025 5040 1040 5055
rect 1043 5052 1044 5064
rect 1051 5052 1078 5064
rect 1043 5044 1078 5052
rect 1043 5043 1072 5044
rect 763 5030 977 5034
rect 778 5028 977 5030
rect 1012 5030 1025 5040
rect 1043 5030 1060 5043
rect 1012 5028 1060 5030
rect 654 5024 687 5028
rect 650 5022 687 5024
rect 650 5021 717 5022
rect 650 5016 681 5021
rect 687 5016 717 5021
rect 650 5012 717 5016
rect 623 5009 717 5012
rect 623 5002 672 5009
rect 623 4996 653 5002
rect 672 4997 677 5002
rect 589 4980 669 4996
rect 681 4988 717 5009
rect 778 5004 967 5028
rect 1012 5027 1059 5028
rect 1025 5022 1059 5027
rect 793 5001 967 5004
rect 786 4998 967 5001
rect 995 5021 1059 5022
rect 589 4978 608 4980
rect 623 4978 657 4980
rect 589 4962 669 4978
rect 589 4956 608 4962
rect 305 4930 408 4940
rect 259 4928 408 4930
rect 429 4928 464 4940
rect 98 4926 260 4928
rect 110 4906 129 4926
rect 144 4924 174 4926
rect -7 4898 34 4906
rect 116 4902 129 4906
rect 181 4910 260 4926
rect 292 4926 464 4928
rect 292 4910 371 4926
rect 378 4924 408 4926
rect -1 4888 28 4898
rect 43 4888 73 4902
rect 116 4888 159 4902
rect 181 4898 371 4910
rect 436 4906 442 4926
rect 166 4888 196 4898
rect 197 4888 355 4898
rect 359 4888 389 4898
rect 393 4888 423 4902
rect 451 4888 464 4926
rect 536 4940 565 4956
rect 579 4940 608 4956
rect 623 4946 653 4962
rect 681 4940 687 4988
rect 690 4982 709 4988
rect 724 4982 754 4990
rect 690 4974 754 4982
rect 690 4958 770 4974
rect 786 4967 848 4998
rect 864 4967 926 4998
rect 995 4996 1044 5021
rect 1059 4996 1089 5012
rect 958 4982 988 4990
rect 995 4988 1105 4996
rect 958 4974 1003 4982
rect 690 4956 709 4958
rect 724 4956 770 4958
rect 690 4940 770 4956
rect 797 4954 832 4967
rect 873 4964 910 4967
rect 873 4962 915 4964
rect 802 4951 832 4954
rect 811 4947 818 4951
rect 818 4946 819 4947
rect 777 4940 787 4946
rect 536 4932 571 4940
rect 536 4906 537 4932
rect 544 4906 571 4932
rect 479 4888 509 4902
rect 536 4898 571 4906
rect 573 4932 614 4940
rect 573 4906 588 4932
rect 595 4906 614 4932
rect 678 4928 709 4940
rect 724 4928 827 4940
rect 839 4930 865 4956
rect 880 4951 910 4962
rect 942 4958 1004 4974
rect 942 4956 988 4958
rect 942 4940 1004 4956
rect 1016 4940 1022 4988
rect 1025 4980 1105 4988
rect 1025 4978 1044 4980
rect 1059 4978 1093 4980
rect 1025 4962 1105 4978
rect 1025 4940 1044 4962
rect 1059 4946 1089 4962
rect 1117 4956 1123 5030
rect 1126 4956 1145 5100
rect 1160 4956 1166 5100
rect 1175 5030 1188 5100
rect 1240 5096 1262 5100
rect 1233 5074 1262 5088
rect 1315 5074 1331 5088
rect 1369 5084 1375 5086
rect 1382 5084 1490 5100
rect 1497 5084 1503 5086
rect 1511 5084 1526 5100
rect 1592 5094 1611 5097
rect 1233 5072 1331 5074
rect 1358 5072 1526 5084
rect 1541 5074 1557 5088
rect 1592 5075 1614 5094
rect 1624 5088 1640 5089
rect 1623 5086 1640 5088
rect 1624 5081 1640 5086
rect 1614 5074 1620 5075
rect 1623 5074 1652 5081
rect 1541 5073 1652 5074
rect 1541 5072 1658 5073
rect 1217 5064 1268 5072
rect 1315 5064 1349 5072
rect 1217 5052 1242 5064
rect 1249 5052 1268 5064
rect 1322 5062 1349 5064
rect 1358 5062 1579 5072
rect 1614 5069 1620 5072
rect 1322 5058 1579 5062
rect 1217 5044 1268 5052
rect 1315 5044 1579 5058
rect 1623 5064 1658 5072
rect 1169 4996 1188 5030
rect 1233 5036 1262 5044
rect 1233 5030 1250 5036
rect 1233 5028 1267 5030
rect 1315 5028 1331 5044
rect 1332 5034 1540 5044
rect 1541 5034 1557 5044
rect 1605 5040 1620 5055
rect 1623 5052 1624 5064
rect 1631 5052 1658 5064
rect 1623 5044 1658 5052
rect 1623 5043 1652 5044
rect 1343 5030 1557 5034
rect 1358 5028 1557 5030
rect 1592 5030 1605 5040
rect 1623 5030 1640 5043
rect 1592 5028 1640 5030
rect 1234 5024 1267 5028
rect 1230 5022 1267 5024
rect 1230 5021 1297 5022
rect 1230 5016 1261 5021
rect 1267 5016 1297 5021
rect 1230 5012 1297 5016
rect 1203 5009 1297 5012
rect 1203 5002 1252 5009
rect 1203 4996 1233 5002
rect 1252 4997 1257 5002
rect 1169 4980 1249 4996
rect 1261 4988 1297 5009
rect 1358 5004 1547 5028
rect 1592 5027 1639 5028
rect 1605 5022 1639 5027
rect 1373 5001 1547 5004
rect 1366 4998 1547 5001
rect 1575 5021 1639 5022
rect 1169 4978 1188 4980
rect 1203 4978 1237 4980
rect 1169 4962 1249 4978
rect 1169 4956 1188 4962
rect 885 4930 988 4940
rect 839 4928 988 4930
rect 1009 4928 1044 4940
rect 678 4926 840 4928
rect 690 4906 709 4926
rect 724 4924 754 4926
rect 573 4898 614 4906
rect 696 4902 709 4906
rect 761 4910 840 4926
rect 872 4926 1044 4928
rect 872 4910 951 4926
rect 958 4924 988 4926
rect 536 4888 565 4898
rect 579 4888 608 4898
rect 623 4888 653 4902
rect 696 4888 739 4902
rect 761 4898 951 4910
rect 1016 4906 1022 4926
rect 746 4888 776 4898
rect 777 4888 935 4898
rect 939 4888 969 4898
rect 973 4888 1003 4902
rect 1031 4888 1044 4926
rect 1116 4940 1145 4956
rect 1159 4940 1188 4956
rect 1203 4946 1233 4962
rect 1261 4940 1267 4988
rect 1270 4982 1289 4988
rect 1304 4982 1334 4990
rect 1270 4974 1334 4982
rect 1270 4958 1350 4974
rect 1366 4967 1428 4998
rect 1444 4967 1506 4998
rect 1575 4996 1624 5021
rect 1639 4996 1669 5012
rect 1538 4982 1568 4990
rect 1575 4988 1685 4996
rect 1538 4974 1583 4982
rect 1270 4956 1289 4958
rect 1304 4956 1350 4958
rect 1270 4940 1350 4956
rect 1377 4954 1412 4967
rect 1453 4964 1490 4967
rect 1453 4962 1495 4964
rect 1382 4951 1412 4954
rect 1391 4947 1398 4951
rect 1398 4946 1399 4947
rect 1357 4940 1367 4946
rect 1116 4932 1151 4940
rect 1116 4906 1117 4932
rect 1124 4906 1151 4932
rect 1059 4888 1089 4902
rect 1116 4898 1151 4906
rect 1153 4932 1194 4940
rect 1153 4906 1168 4932
rect 1175 4906 1194 4932
rect 1258 4928 1289 4940
rect 1304 4928 1407 4940
rect 1419 4930 1445 4956
rect 1460 4951 1490 4962
rect 1522 4958 1584 4974
rect 1522 4956 1568 4958
rect 1522 4940 1584 4956
rect 1596 4940 1602 4988
rect 1605 4980 1685 4988
rect 1605 4978 1624 4980
rect 1639 4978 1673 4980
rect 1605 4962 1685 4978
rect 1605 4940 1624 4962
rect 1639 4946 1669 4962
rect 1697 4956 1703 5030
rect 1706 4956 1725 5100
rect 1740 4956 1746 5100
rect 1755 5030 1768 5100
rect 1820 5096 1842 5100
rect 1813 5074 1842 5088
rect 1895 5074 1911 5088
rect 1949 5084 1955 5086
rect 1962 5084 2070 5100
rect 2077 5084 2083 5086
rect 2091 5084 2106 5100
rect 2172 5094 2191 5097
rect 1813 5072 1911 5074
rect 1938 5072 2106 5084
rect 2121 5074 2137 5088
rect 2172 5075 2194 5094
rect 2204 5088 2220 5089
rect 2203 5086 2220 5088
rect 2204 5081 2220 5086
rect 2194 5074 2200 5075
rect 2203 5074 2232 5081
rect 2121 5073 2232 5074
rect 2121 5072 2238 5073
rect 1797 5064 1848 5072
rect 1895 5064 1929 5072
rect 1797 5052 1822 5064
rect 1829 5052 1848 5064
rect 1902 5062 1929 5064
rect 1938 5062 2159 5072
rect 2194 5069 2200 5072
rect 1902 5058 2159 5062
rect 1797 5044 1848 5052
rect 1895 5044 2159 5058
rect 2203 5064 2238 5072
rect 1749 4996 1768 5030
rect 1813 5036 1842 5044
rect 1813 5030 1830 5036
rect 1813 5028 1847 5030
rect 1895 5028 1911 5044
rect 1912 5034 2120 5044
rect 2121 5034 2137 5044
rect 2185 5040 2200 5055
rect 2203 5052 2204 5064
rect 2211 5052 2238 5064
rect 2203 5044 2238 5052
rect 2203 5043 2232 5044
rect 1923 5030 2137 5034
rect 1938 5028 2137 5030
rect 2172 5030 2185 5040
rect 2203 5030 2220 5043
rect 2172 5028 2220 5030
rect 1814 5024 1847 5028
rect 1810 5022 1847 5024
rect 1810 5021 1877 5022
rect 1810 5016 1841 5021
rect 1847 5016 1877 5021
rect 1810 5012 1877 5016
rect 1783 5009 1877 5012
rect 1783 5002 1832 5009
rect 1783 4996 1813 5002
rect 1832 4997 1837 5002
rect 1749 4980 1829 4996
rect 1841 4988 1877 5009
rect 1938 5004 2127 5028
rect 2172 5027 2219 5028
rect 2185 5022 2219 5027
rect 1953 5001 2127 5004
rect 1946 4998 2127 5001
rect 2155 5021 2219 5022
rect 1749 4978 1768 4980
rect 1783 4978 1817 4980
rect 1749 4962 1829 4978
rect 1749 4956 1768 4962
rect 1465 4930 1568 4940
rect 1419 4928 1568 4930
rect 1589 4928 1624 4940
rect 1258 4926 1420 4928
rect 1270 4906 1289 4926
rect 1304 4924 1334 4926
rect 1153 4898 1194 4906
rect 1276 4902 1289 4906
rect 1341 4910 1420 4926
rect 1452 4926 1624 4928
rect 1452 4910 1531 4926
rect 1538 4924 1568 4926
rect 1116 4888 1145 4898
rect 1159 4888 1188 4898
rect 1203 4888 1233 4902
rect 1276 4888 1319 4902
rect 1341 4898 1531 4910
rect 1596 4906 1602 4926
rect 1326 4888 1356 4898
rect 1357 4888 1515 4898
rect 1519 4888 1549 4898
rect 1553 4888 1583 4902
rect 1611 4888 1624 4926
rect 1696 4940 1725 4956
rect 1739 4940 1768 4956
rect 1783 4946 1813 4962
rect 1841 4940 1847 4988
rect 1850 4982 1869 4988
rect 1884 4982 1914 4990
rect 1850 4974 1914 4982
rect 1850 4958 1930 4974
rect 1946 4967 2008 4998
rect 2024 4967 2086 4998
rect 2155 4996 2204 5021
rect 2219 4996 2249 5012
rect 2118 4982 2148 4990
rect 2155 4988 2265 4996
rect 2118 4974 2163 4982
rect 1850 4956 1869 4958
rect 1884 4956 1930 4958
rect 1850 4940 1930 4956
rect 1957 4954 1992 4967
rect 2033 4964 2070 4967
rect 2033 4962 2075 4964
rect 1962 4951 1992 4954
rect 1971 4947 1978 4951
rect 1978 4946 1979 4947
rect 1937 4940 1947 4946
rect 1696 4932 1731 4940
rect 1696 4906 1697 4932
rect 1704 4906 1731 4932
rect 1639 4888 1669 4902
rect 1696 4898 1731 4906
rect 1733 4932 1774 4940
rect 1733 4906 1748 4932
rect 1755 4906 1774 4932
rect 1838 4928 1869 4940
rect 1884 4928 1987 4940
rect 1999 4930 2025 4956
rect 2040 4951 2070 4962
rect 2102 4958 2164 4974
rect 2102 4956 2148 4958
rect 2102 4940 2164 4956
rect 2176 4940 2182 4988
rect 2185 4980 2265 4988
rect 2185 4978 2204 4980
rect 2219 4978 2253 4980
rect 2185 4962 2265 4978
rect 2185 4940 2204 4962
rect 2219 4946 2249 4962
rect 2277 4956 2283 5030
rect 2286 4956 2305 5100
rect 2320 4956 2326 5100
rect 2335 5030 2348 5100
rect 2400 5096 2422 5100
rect 2393 5074 2422 5088
rect 2475 5074 2491 5088
rect 2529 5084 2535 5086
rect 2542 5084 2650 5100
rect 2657 5084 2663 5086
rect 2671 5084 2686 5100
rect 2752 5094 2771 5097
rect 2393 5072 2491 5074
rect 2518 5072 2686 5084
rect 2701 5074 2717 5088
rect 2752 5075 2774 5094
rect 2784 5088 2800 5089
rect 2783 5086 2800 5088
rect 2784 5081 2800 5086
rect 2774 5074 2780 5075
rect 2783 5074 2812 5081
rect 2701 5073 2812 5074
rect 2701 5072 2818 5073
rect 2377 5064 2428 5072
rect 2475 5064 2509 5072
rect 2377 5052 2402 5064
rect 2409 5052 2428 5064
rect 2482 5062 2509 5064
rect 2518 5062 2739 5072
rect 2774 5069 2780 5072
rect 2482 5058 2739 5062
rect 2377 5044 2428 5052
rect 2475 5044 2739 5058
rect 2783 5064 2818 5072
rect 2329 4996 2348 5030
rect 2393 5036 2422 5044
rect 2393 5030 2410 5036
rect 2393 5028 2427 5030
rect 2475 5028 2491 5044
rect 2492 5034 2700 5044
rect 2701 5034 2717 5044
rect 2765 5040 2780 5055
rect 2783 5052 2784 5064
rect 2791 5052 2818 5064
rect 2783 5044 2818 5052
rect 2783 5043 2812 5044
rect 2503 5030 2717 5034
rect 2518 5028 2717 5030
rect 2752 5030 2765 5040
rect 2783 5030 2800 5043
rect 2752 5028 2800 5030
rect 2394 5024 2427 5028
rect 2390 5022 2427 5024
rect 2390 5021 2457 5022
rect 2390 5016 2421 5021
rect 2427 5016 2457 5021
rect 2390 5012 2457 5016
rect 2363 5009 2457 5012
rect 2363 5002 2412 5009
rect 2363 4996 2393 5002
rect 2412 4997 2417 5002
rect 2329 4980 2409 4996
rect 2421 4988 2457 5009
rect 2518 5004 2707 5028
rect 2752 5027 2799 5028
rect 2765 5022 2799 5027
rect 2533 5001 2707 5004
rect 2526 4998 2707 5001
rect 2735 5021 2799 5022
rect 2329 4978 2348 4980
rect 2363 4978 2397 4980
rect 2329 4962 2409 4978
rect 2329 4956 2348 4962
rect 2045 4930 2148 4940
rect 1999 4928 2148 4930
rect 2169 4928 2204 4940
rect 1838 4926 2000 4928
rect 1850 4906 1869 4926
rect 1884 4924 1914 4926
rect 1733 4898 1774 4906
rect 1856 4902 1869 4906
rect 1921 4910 2000 4926
rect 2032 4926 2204 4928
rect 2032 4910 2111 4926
rect 2118 4924 2148 4926
rect 1696 4888 1725 4898
rect 1739 4888 1768 4898
rect 1783 4888 1813 4902
rect 1856 4888 1899 4902
rect 1921 4898 2111 4910
rect 2176 4906 2182 4926
rect 1906 4888 1936 4898
rect 1937 4888 2095 4898
rect 2099 4888 2129 4898
rect 2133 4888 2163 4902
rect 2191 4888 2204 4926
rect 2276 4940 2305 4956
rect 2319 4940 2348 4956
rect 2363 4946 2393 4962
rect 2421 4940 2427 4988
rect 2430 4982 2449 4988
rect 2464 4982 2494 4990
rect 2430 4974 2494 4982
rect 2430 4958 2510 4974
rect 2526 4967 2588 4998
rect 2604 4967 2666 4998
rect 2735 4996 2784 5021
rect 2799 4996 2829 5012
rect 2698 4982 2728 4990
rect 2735 4988 2845 4996
rect 2698 4974 2743 4982
rect 2430 4956 2449 4958
rect 2464 4956 2510 4958
rect 2430 4940 2510 4956
rect 2537 4954 2572 4967
rect 2613 4964 2650 4967
rect 2613 4962 2655 4964
rect 2542 4951 2572 4954
rect 2551 4947 2558 4951
rect 2558 4946 2559 4947
rect 2517 4940 2527 4946
rect 2276 4932 2311 4940
rect 2276 4906 2277 4932
rect 2284 4906 2311 4932
rect 2219 4888 2249 4902
rect 2276 4898 2311 4906
rect 2313 4932 2354 4940
rect 2313 4906 2328 4932
rect 2335 4906 2354 4932
rect 2418 4928 2449 4940
rect 2464 4928 2567 4940
rect 2579 4930 2605 4956
rect 2620 4951 2650 4962
rect 2682 4958 2744 4974
rect 2682 4956 2728 4958
rect 2682 4940 2744 4956
rect 2756 4940 2762 4988
rect 2765 4980 2845 4988
rect 2765 4978 2784 4980
rect 2799 4978 2833 4980
rect 2765 4962 2845 4978
rect 2765 4940 2784 4962
rect 2799 4946 2829 4962
rect 2857 4956 2863 5030
rect 2866 4956 2885 5100
rect 2900 4956 2906 5100
rect 2915 5030 2928 5100
rect 2980 5096 3002 5100
rect 2973 5074 3002 5088
rect 3055 5074 3071 5088
rect 3109 5084 3115 5086
rect 3122 5084 3230 5100
rect 3237 5084 3243 5086
rect 3251 5084 3266 5100
rect 3332 5094 3351 5097
rect 2973 5072 3071 5074
rect 3098 5072 3266 5084
rect 3281 5074 3297 5088
rect 3332 5075 3354 5094
rect 3364 5088 3380 5089
rect 3363 5086 3380 5088
rect 3364 5081 3380 5086
rect 3354 5074 3360 5075
rect 3363 5074 3392 5081
rect 3281 5073 3392 5074
rect 3281 5072 3398 5073
rect 2957 5064 3008 5072
rect 3055 5064 3089 5072
rect 2957 5052 2982 5064
rect 2989 5052 3008 5064
rect 3062 5062 3089 5064
rect 3098 5062 3319 5072
rect 3354 5069 3360 5072
rect 3062 5058 3319 5062
rect 2957 5044 3008 5052
rect 3055 5044 3319 5058
rect 3363 5064 3398 5072
rect 2909 4996 2928 5030
rect 2973 5036 3002 5044
rect 2973 5030 2990 5036
rect 2973 5028 3007 5030
rect 3055 5028 3071 5044
rect 3072 5034 3280 5044
rect 3281 5034 3297 5044
rect 3345 5040 3360 5055
rect 3363 5052 3364 5064
rect 3371 5052 3398 5064
rect 3363 5044 3398 5052
rect 3363 5043 3392 5044
rect 3083 5030 3297 5034
rect 3098 5028 3297 5030
rect 3332 5030 3345 5040
rect 3363 5030 3380 5043
rect 3332 5028 3380 5030
rect 2974 5024 3007 5028
rect 2970 5022 3007 5024
rect 2970 5021 3037 5022
rect 2970 5016 3001 5021
rect 3007 5016 3037 5021
rect 2970 5012 3037 5016
rect 2943 5009 3037 5012
rect 2943 5002 2992 5009
rect 2943 4996 2973 5002
rect 2992 4997 2997 5002
rect 2909 4980 2989 4996
rect 3001 4988 3037 5009
rect 3098 5004 3287 5028
rect 3332 5027 3379 5028
rect 3345 5022 3379 5027
rect 3113 5001 3287 5004
rect 3106 4998 3287 5001
rect 3315 5021 3379 5022
rect 2909 4978 2928 4980
rect 2943 4978 2977 4980
rect 2909 4962 2989 4978
rect 2909 4956 2928 4962
rect 2625 4930 2728 4940
rect 2579 4928 2728 4930
rect 2749 4928 2784 4940
rect 2418 4926 2580 4928
rect 2430 4906 2449 4926
rect 2464 4924 2494 4926
rect 2313 4898 2354 4906
rect 2436 4902 2449 4906
rect 2501 4910 2580 4926
rect 2612 4926 2784 4928
rect 2612 4910 2691 4926
rect 2698 4924 2728 4926
rect 2276 4888 2305 4898
rect 2319 4888 2348 4898
rect 2363 4888 2393 4902
rect 2436 4888 2479 4902
rect 2501 4898 2691 4910
rect 2756 4906 2762 4926
rect 2486 4888 2516 4898
rect 2517 4888 2675 4898
rect 2679 4888 2709 4898
rect 2713 4888 2743 4902
rect 2771 4888 2784 4926
rect 2856 4940 2885 4956
rect 2899 4940 2928 4956
rect 2943 4946 2973 4962
rect 3001 4940 3007 4988
rect 3010 4982 3029 4988
rect 3044 4982 3074 4990
rect 3010 4974 3074 4982
rect 3010 4958 3090 4974
rect 3106 4967 3168 4998
rect 3184 4967 3246 4998
rect 3315 4996 3364 5021
rect 3379 4996 3409 5012
rect 3278 4982 3308 4990
rect 3315 4988 3425 4996
rect 3278 4974 3323 4982
rect 3010 4956 3029 4958
rect 3044 4956 3090 4958
rect 3010 4940 3090 4956
rect 3117 4954 3152 4967
rect 3193 4964 3230 4967
rect 3193 4962 3235 4964
rect 3122 4951 3152 4954
rect 3131 4947 3138 4951
rect 3138 4946 3139 4947
rect 3097 4940 3107 4946
rect 2856 4932 2891 4940
rect 2856 4906 2857 4932
rect 2864 4906 2891 4932
rect 2799 4888 2829 4902
rect 2856 4898 2891 4906
rect 2893 4932 2934 4940
rect 2893 4906 2908 4932
rect 2915 4906 2934 4932
rect 2998 4928 3029 4940
rect 3044 4928 3147 4940
rect 3159 4930 3185 4956
rect 3200 4951 3230 4962
rect 3262 4958 3324 4974
rect 3262 4956 3308 4958
rect 3262 4940 3324 4956
rect 3336 4940 3342 4988
rect 3345 4980 3425 4988
rect 3345 4978 3364 4980
rect 3379 4978 3413 4980
rect 3345 4962 3425 4978
rect 3345 4940 3364 4962
rect 3379 4946 3409 4962
rect 3437 4956 3443 5030
rect 3446 4956 3465 5100
rect 3480 4956 3486 5100
rect 3495 5030 3508 5100
rect 3560 5096 3582 5100
rect 3553 5074 3582 5088
rect 3635 5074 3651 5088
rect 3689 5084 3695 5086
rect 3702 5084 3810 5100
rect 3817 5084 3823 5086
rect 3831 5084 3846 5100
rect 3912 5094 3931 5097
rect 3553 5072 3651 5074
rect 3678 5072 3846 5084
rect 3861 5074 3877 5088
rect 3912 5075 3934 5094
rect 3944 5088 3960 5089
rect 3943 5086 3960 5088
rect 3944 5081 3960 5086
rect 3934 5074 3940 5075
rect 3943 5074 3972 5081
rect 3861 5073 3972 5074
rect 3861 5072 3978 5073
rect 3537 5064 3588 5072
rect 3635 5064 3669 5072
rect 3537 5052 3562 5064
rect 3569 5052 3588 5064
rect 3642 5062 3669 5064
rect 3678 5062 3899 5072
rect 3934 5069 3940 5072
rect 3642 5058 3899 5062
rect 3537 5044 3588 5052
rect 3635 5044 3899 5058
rect 3943 5064 3978 5072
rect 3489 4996 3508 5030
rect 3553 5036 3582 5044
rect 3553 5030 3570 5036
rect 3553 5028 3587 5030
rect 3635 5028 3651 5044
rect 3652 5034 3860 5044
rect 3861 5034 3877 5044
rect 3925 5040 3940 5055
rect 3943 5052 3944 5064
rect 3951 5052 3978 5064
rect 3943 5044 3978 5052
rect 3943 5043 3972 5044
rect 3663 5030 3877 5034
rect 3678 5028 3877 5030
rect 3912 5030 3925 5040
rect 3943 5030 3960 5043
rect 3912 5028 3960 5030
rect 3554 5024 3587 5028
rect 3550 5022 3587 5024
rect 3550 5021 3617 5022
rect 3550 5016 3581 5021
rect 3587 5016 3617 5021
rect 3550 5012 3617 5016
rect 3523 5009 3617 5012
rect 3523 5002 3572 5009
rect 3523 4996 3553 5002
rect 3572 4997 3577 5002
rect 3489 4980 3569 4996
rect 3581 4988 3617 5009
rect 3678 5004 3867 5028
rect 3912 5027 3959 5028
rect 3925 5022 3959 5027
rect 3693 5001 3867 5004
rect 3686 4998 3867 5001
rect 3895 5021 3959 5022
rect 3489 4978 3508 4980
rect 3523 4978 3557 4980
rect 3489 4962 3569 4978
rect 3489 4956 3508 4962
rect 3205 4930 3308 4940
rect 3159 4928 3308 4930
rect 3329 4928 3364 4940
rect 2998 4926 3160 4928
rect 3010 4906 3029 4926
rect 3044 4924 3074 4926
rect 2893 4898 2934 4906
rect 3016 4902 3029 4906
rect 3081 4910 3160 4926
rect 3192 4926 3364 4928
rect 3192 4910 3271 4926
rect 3278 4924 3308 4926
rect 2856 4888 2885 4898
rect 2899 4888 2928 4898
rect 2943 4888 2973 4902
rect 3016 4888 3059 4902
rect 3081 4898 3271 4910
rect 3336 4906 3342 4926
rect 3066 4888 3096 4898
rect 3097 4888 3255 4898
rect 3259 4888 3289 4898
rect 3293 4888 3323 4902
rect 3351 4888 3364 4926
rect 3436 4940 3465 4956
rect 3479 4940 3508 4956
rect 3523 4946 3553 4962
rect 3581 4940 3587 4988
rect 3590 4982 3609 4988
rect 3624 4982 3654 4990
rect 3590 4974 3654 4982
rect 3590 4958 3670 4974
rect 3686 4967 3748 4998
rect 3764 4967 3826 4998
rect 3895 4996 3944 5021
rect 3959 4996 3989 5012
rect 3858 4982 3888 4990
rect 3895 4988 4005 4996
rect 3858 4974 3903 4982
rect 3590 4956 3609 4958
rect 3624 4956 3670 4958
rect 3590 4940 3670 4956
rect 3697 4954 3732 4967
rect 3773 4964 3810 4967
rect 3773 4962 3815 4964
rect 3702 4951 3732 4954
rect 3711 4947 3718 4951
rect 3718 4946 3719 4947
rect 3677 4940 3687 4946
rect 3436 4932 3471 4940
rect 3436 4906 3437 4932
rect 3444 4906 3471 4932
rect 3379 4888 3409 4902
rect 3436 4898 3471 4906
rect 3473 4932 3514 4940
rect 3473 4906 3488 4932
rect 3495 4906 3514 4932
rect 3578 4928 3609 4940
rect 3624 4928 3727 4940
rect 3739 4930 3765 4956
rect 3780 4951 3810 4962
rect 3842 4958 3904 4974
rect 3842 4956 3888 4958
rect 3842 4940 3904 4956
rect 3916 4940 3922 4988
rect 3925 4980 4005 4988
rect 3925 4978 3944 4980
rect 3959 4978 3993 4980
rect 3925 4962 4005 4978
rect 3925 4940 3944 4962
rect 3959 4946 3989 4962
rect 4017 4956 4023 5030
rect 4026 4956 4045 5100
rect 4060 4956 4066 5100
rect 4075 5030 4088 5100
rect 4140 5096 4162 5100
rect 4133 5074 4162 5088
rect 4215 5074 4231 5088
rect 4269 5084 4275 5086
rect 4282 5084 4390 5100
rect 4397 5084 4403 5086
rect 4411 5084 4426 5100
rect 4492 5094 4511 5097
rect 4133 5072 4231 5074
rect 4258 5072 4426 5084
rect 4441 5074 4457 5088
rect 4492 5075 4514 5094
rect 4524 5088 4540 5089
rect 4523 5086 4540 5088
rect 4524 5081 4540 5086
rect 4514 5074 4520 5075
rect 4523 5074 4552 5081
rect 4441 5073 4552 5074
rect 4441 5072 4558 5073
rect 4117 5064 4168 5072
rect 4215 5064 4249 5072
rect 4117 5052 4142 5064
rect 4149 5052 4168 5064
rect 4222 5062 4249 5064
rect 4258 5062 4479 5072
rect 4514 5069 4520 5072
rect 4222 5058 4479 5062
rect 4117 5044 4168 5052
rect 4215 5044 4479 5058
rect 4523 5064 4558 5072
rect 4069 4996 4088 5030
rect 4133 5036 4162 5044
rect 4133 5030 4150 5036
rect 4133 5028 4167 5030
rect 4215 5028 4231 5044
rect 4232 5034 4440 5044
rect 4441 5034 4457 5044
rect 4505 5040 4520 5055
rect 4523 5052 4524 5064
rect 4531 5052 4558 5064
rect 4523 5044 4558 5052
rect 4523 5043 4552 5044
rect 4243 5030 4457 5034
rect 4258 5028 4457 5030
rect 4492 5030 4505 5040
rect 4523 5030 4540 5043
rect 4492 5028 4540 5030
rect 4134 5024 4167 5028
rect 4130 5022 4167 5024
rect 4130 5021 4197 5022
rect 4130 5016 4161 5021
rect 4167 5016 4197 5021
rect 4130 5012 4197 5016
rect 4103 5009 4197 5012
rect 4103 5002 4152 5009
rect 4103 4996 4133 5002
rect 4152 4997 4157 5002
rect 4069 4980 4149 4996
rect 4161 4988 4197 5009
rect 4258 5004 4447 5028
rect 4492 5027 4539 5028
rect 4505 5022 4539 5027
rect 4273 5001 4447 5004
rect 4266 4998 4447 5001
rect 4475 5021 4539 5022
rect 4069 4978 4088 4980
rect 4103 4978 4137 4980
rect 4069 4962 4149 4978
rect 4069 4956 4088 4962
rect 3785 4930 3888 4940
rect 3739 4928 3888 4930
rect 3909 4928 3944 4940
rect 3578 4926 3740 4928
rect 3590 4906 3609 4926
rect 3624 4924 3654 4926
rect 3473 4898 3514 4906
rect 3596 4902 3609 4906
rect 3661 4910 3740 4926
rect 3772 4926 3944 4928
rect 3772 4910 3851 4926
rect 3858 4924 3888 4926
rect 3436 4888 3465 4898
rect 3479 4888 3508 4898
rect 3523 4888 3553 4902
rect 3596 4888 3639 4902
rect 3661 4898 3851 4910
rect 3916 4906 3922 4926
rect 3646 4888 3676 4898
rect 3677 4888 3835 4898
rect 3839 4888 3869 4898
rect 3873 4888 3903 4902
rect 3931 4888 3944 4926
rect 4016 4940 4045 4956
rect 4059 4940 4088 4956
rect 4103 4946 4133 4962
rect 4161 4940 4167 4988
rect 4170 4982 4189 4988
rect 4204 4982 4234 4990
rect 4170 4974 4234 4982
rect 4170 4958 4250 4974
rect 4266 4967 4328 4998
rect 4344 4967 4406 4998
rect 4475 4996 4524 5021
rect 4539 4996 4569 5012
rect 4438 4982 4468 4990
rect 4475 4988 4585 4996
rect 4438 4974 4483 4982
rect 4170 4956 4189 4958
rect 4204 4956 4250 4958
rect 4170 4940 4250 4956
rect 4277 4954 4312 4967
rect 4353 4964 4390 4967
rect 4353 4962 4395 4964
rect 4282 4951 4312 4954
rect 4291 4947 4298 4951
rect 4298 4946 4299 4947
rect 4257 4940 4267 4946
rect 4016 4932 4051 4940
rect 4016 4906 4017 4932
rect 4024 4906 4051 4932
rect 3959 4888 3989 4902
rect 4016 4898 4051 4906
rect 4053 4932 4094 4940
rect 4053 4906 4068 4932
rect 4075 4906 4094 4932
rect 4158 4928 4189 4940
rect 4204 4928 4307 4940
rect 4319 4930 4345 4956
rect 4360 4951 4390 4962
rect 4422 4958 4484 4974
rect 4422 4956 4468 4958
rect 4422 4940 4484 4956
rect 4496 4940 4502 4988
rect 4505 4980 4585 4988
rect 4505 4978 4524 4980
rect 4539 4978 4573 4980
rect 4505 4962 4585 4978
rect 4505 4940 4524 4962
rect 4539 4946 4569 4962
rect 4597 4956 4603 5030
rect 4606 4956 4625 5100
rect 4640 4956 4646 5100
rect 4655 5030 4668 5100
rect 4720 5096 4742 5100
rect 4713 5074 4742 5088
rect 4795 5074 4811 5088
rect 4849 5084 4855 5086
rect 4862 5084 4970 5100
rect 4977 5084 4983 5086
rect 4991 5084 5006 5100
rect 5072 5094 5091 5097
rect 4713 5072 4811 5074
rect 4838 5072 5006 5084
rect 5021 5074 5037 5088
rect 5072 5075 5094 5094
rect 5104 5088 5120 5089
rect 5103 5086 5120 5088
rect 5104 5081 5120 5086
rect 5094 5074 5100 5075
rect 5103 5074 5132 5081
rect 5021 5073 5132 5074
rect 5021 5072 5138 5073
rect 4697 5064 4748 5072
rect 4795 5064 4829 5072
rect 4697 5052 4722 5064
rect 4729 5052 4748 5064
rect 4802 5062 4829 5064
rect 4838 5062 5059 5072
rect 5094 5069 5100 5072
rect 4802 5058 5059 5062
rect 4697 5044 4748 5052
rect 4795 5044 5059 5058
rect 5103 5064 5138 5072
rect 4649 4996 4668 5030
rect 4713 5036 4742 5044
rect 4713 5030 4730 5036
rect 4713 5028 4747 5030
rect 4795 5028 4811 5044
rect 4812 5034 5020 5044
rect 5021 5034 5037 5044
rect 5085 5040 5100 5055
rect 5103 5052 5104 5064
rect 5111 5052 5138 5064
rect 5103 5044 5138 5052
rect 5103 5043 5132 5044
rect 4823 5030 5037 5034
rect 4838 5028 5037 5030
rect 5072 5030 5085 5040
rect 5103 5030 5120 5043
rect 5072 5028 5120 5030
rect 4714 5024 4747 5028
rect 4710 5022 4747 5024
rect 4710 5021 4777 5022
rect 4710 5016 4741 5021
rect 4747 5016 4777 5021
rect 4710 5012 4777 5016
rect 4683 5009 4777 5012
rect 4683 5002 4732 5009
rect 4683 4996 4713 5002
rect 4732 4997 4737 5002
rect 4649 4980 4729 4996
rect 4741 4988 4777 5009
rect 4838 5004 5027 5028
rect 5072 5027 5119 5028
rect 5085 5022 5119 5027
rect 4853 5001 5027 5004
rect 4846 4998 5027 5001
rect 5055 5021 5119 5022
rect 4649 4978 4668 4980
rect 4683 4978 4717 4980
rect 4649 4962 4729 4978
rect 4649 4956 4668 4962
rect 4365 4930 4468 4940
rect 4319 4928 4468 4930
rect 4489 4928 4524 4940
rect 4158 4926 4320 4928
rect 4170 4906 4189 4926
rect 4204 4924 4234 4926
rect 4053 4898 4094 4906
rect 4176 4902 4189 4906
rect 4241 4910 4320 4926
rect 4352 4926 4524 4928
rect 4352 4910 4431 4926
rect 4438 4924 4468 4926
rect 4016 4888 4045 4898
rect 4059 4888 4088 4898
rect 4103 4888 4133 4902
rect 4176 4888 4219 4902
rect 4241 4898 4431 4910
rect 4496 4906 4502 4926
rect 4226 4888 4256 4898
rect 4257 4888 4415 4898
rect 4419 4888 4449 4898
rect 4453 4888 4483 4902
rect 4511 4888 4524 4926
rect 4596 4940 4625 4956
rect 4639 4940 4668 4956
rect 4683 4946 4713 4962
rect 4741 4940 4747 4988
rect 4750 4982 4769 4988
rect 4784 4982 4814 4990
rect 4750 4974 4814 4982
rect 4750 4958 4830 4974
rect 4846 4967 4908 4998
rect 4924 4967 4986 4998
rect 5055 4996 5104 5021
rect 5119 4996 5149 5012
rect 5018 4982 5048 4990
rect 5055 4988 5165 4996
rect 5018 4974 5063 4982
rect 4750 4956 4769 4958
rect 4784 4956 4830 4958
rect 4750 4940 4830 4956
rect 4857 4954 4892 4967
rect 4933 4964 4970 4967
rect 4933 4962 4975 4964
rect 4862 4951 4892 4954
rect 4871 4947 4878 4951
rect 4878 4946 4879 4947
rect 4837 4940 4847 4946
rect 4596 4932 4631 4940
rect 4596 4906 4597 4932
rect 4604 4906 4631 4932
rect 4539 4888 4569 4902
rect 4596 4898 4631 4906
rect 4633 4932 4674 4940
rect 4633 4906 4648 4932
rect 4655 4906 4674 4932
rect 4738 4928 4769 4940
rect 4784 4928 4887 4940
rect 4899 4930 4925 4956
rect 4940 4951 4970 4962
rect 5002 4958 5064 4974
rect 5002 4956 5048 4958
rect 5002 4940 5064 4956
rect 5076 4940 5082 4988
rect 5085 4980 5165 4988
rect 5085 4978 5104 4980
rect 5119 4978 5153 4980
rect 5085 4962 5165 4978
rect 5085 4940 5104 4962
rect 5119 4946 5149 4962
rect 5177 4956 5183 5030
rect 5186 4956 5205 5100
rect 5220 4956 5226 5100
rect 5235 5030 5248 5100
rect 5300 5096 5322 5100
rect 5293 5074 5322 5088
rect 5375 5074 5391 5088
rect 5429 5084 5435 5086
rect 5442 5084 5550 5100
rect 5557 5084 5563 5086
rect 5571 5084 5586 5100
rect 5652 5094 5671 5097
rect 5293 5072 5391 5074
rect 5418 5072 5586 5084
rect 5601 5074 5617 5088
rect 5652 5075 5674 5094
rect 5684 5088 5700 5089
rect 5683 5086 5700 5088
rect 5684 5081 5700 5086
rect 5674 5074 5680 5075
rect 5683 5074 5712 5081
rect 5601 5073 5712 5074
rect 5601 5072 5718 5073
rect 5277 5064 5328 5072
rect 5375 5064 5409 5072
rect 5277 5052 5302 5064
rect 5309 5052 5328 5064
rect 5382 5062 5409 5064
rect 5418 5062 5639 5072
rect 5674 5069 5680 5072
rect 5382 5058 5639 5062
rect 5277 5044 5328 5052
rect 5375 5044 5639 5058
rect 5683 5064 5718 5072
rect 5229 4996 5248 5030
rect 5293 5036 5322 5044
rect 5293 5030 5310 5036
rect 5293 5028 5327 5030
rect 5375 5028 5391 5044
rect 5392 5034 5600 5044
rect 5601 5034 5617 5044
rect 5665 5040 5680 5055
rect 5683 5052 5684 5064
rect 5691 5052 5718 5064
rect 5683 5044 5718 5052
rect 5683 5043 5712 5044
rect 5403 5030 5617 5034
rect 5418 5028 5617 5030
rect 5652 5030 5665 5040
rect 5683 5030 5700 5043
rect 5652 5028 5700 5030
rect 5294 5024 5327 5028
rect 5290 5022 5327 5024
rect 5290 5021 5357 5022
rect 5290 5016 5321 5021
rect 5327 5016 5357 5021
rect 5290 5012 5357 5016
rect 5263 5009 5357 5012
rect 5263 5002 5312 5009
rect 5263 4996 5293 5002
rect 5312 4997 5317 5002
rect 5229 4980 5309 4996
rect 5321 4988 5357 5009
rect 5418 5004 5607 5028
rect 5652 5027 5699 5028
rect 5665 5022 5699 5027
rect 5433 5001 5607 5004
rect 5426 4998 5607 5001
rect 5635 5021 5699 5022
rect 5229 4978 5248 4980
rect 5263 4978 5297 4980
rect 5229 4962 5309 4978
rect 5229 4956 5248 4962
rect 4945 4930 5048 4940
rect 4899 4928 5048 4930
rect 5069 4928 5104 4940
rect 4738 4926 4900 4928
rect 4750 4906 4769 4926
rect 4784 4924 4814 4926
rect 4633 4898 4674 4906
rect 4756 4902 4769 4906
rect 4821 4910 4900 4926
rect 4932 4926 5104 4928
rect 4932 4910 5011 4926
rect 5018 4924 5048 4926
rect 4596 4888 4625 4898
rect 4639 4888 4668 4898
rect 4683 4888 4713 4902
rect 4756 4888 4799 4902
rect 4821 4898 5011 4910
rect 5076 4906 5082 4926
rect 4806 4888 4836 4898
rect 4837 4888 4995 4898
rect 4999 4888 5029 4898
rect 5033 4888 5063 4902
rect 5091 4888 5104 4926
rect 5176 4940 5205 4956
rect 5219 4940 5248 4956
rect 5263 4946 5293 4962
rect 5321 4940 5327 4988
rect 5330 4982 5349 4988
rect 5364 4982 5394 4990
rect 5330 4974 5394 4982
rect 5330 4958 5410 4974
rect 5426 4967 5488 4998
rect 5504 4967 5566 4998
rect 5635 4996 5684 5021
rect 5699 4996 5729 5012
rect 5598 4982 5628 4990
rect 5635 4988 5745 4996
rect 5598 4974 5643 4982
rect 5330 4956 5349 4958
rect 5364 4956 5410 4958
rect 5330 4940 5410 4956
rect 5437 4954 5472 4967
rect 5513 4964 5550 4967
rect 5513 4962 5555 4964
rect 5442 4951 5472 4954
rect 5451 4947 5458 4951
rect 5458 4946 5459 4947
rect 5417 4940 5427 4946
rect 5176 4932 5211 4940
rect 5176 4906 5177 4932
rect 5184 4906 5211 4932
rect 5119 4888 5149 4902
rect 5176 4898 5211 4906
rect 5213 4932 5254 4940
rect 5213 4906 5228 4932
rect 5235 4906 5254 4932
rect 5318 4928 5349 4940
rect 5364 4928 5467 4940
rect 5479 4930 5505 4956
rect 5520 4951 5550 4962
rect 5582 4958 5644 4974
rect 5582 4956 5628 4958
rect 5582 4940 5644 4956
rect 5656 4940 5662 4988
rect 5665 4980 5745 4988
rect 5665 4978 5684 4980
rect 5699 4978 5733 4980
rect 5665 4962 5745 4978
rect 5665 4940 5684 4962
rect 5699 4946 5729 4962
rect 5757 4956 5763 5030
rect 5766 4956 5785 5100
rect 5800 4956 5806 5100
rect 5815 5030 5828 5100
rect 5880 5096 5902 5100
rect 5873 5074 5902 5088
rect 5955 5074 5971 5088
rect 6009 5084 6015 5086
rect 6022 5084 6130 5100
rect 6137 5084 6143 5086
rect 6151 5084 6166 5100
rect 6232 5094 6251 5097
rect 5873 5072 5971 5074
rect 5998 5072 6166 5084
rect 6181 5074 6197 5088
rect 6232 5075 6254 5094
rect 6264 5088 6280 5089
rect 6263 5086 6280 5088
rect 6264 5081 6280 5086
rect 6254 5074 6260 5075
rect 6263 5074 6292 5081
rect 6181 5073 6292 5074
rect 6181 5072 6298 5073
rect 5857 5064 5908 5072
rect 5955 5064 5989 5072
rect 5857 5052 5882 5064
rect 5889 5052 5908 5064
rect 5962 5062 5989 5064
rect 5998 5062 6219 5072
rect 6254 5069 6260 5072
rect 5962 5058 6219 5062
rect 5857 5044 5908 5052
rect 5955 5044 6219 5058
rect 6263 5064 6298 5072
rect 5809 4996 5828 5030
rect 5873 5036 5902 5044
rect 5873 5030 5890 5036
rect 5873 5028 5907 5030
rect 5955 5028 5971 5044
rect 5972 5034 6180 5044
rect 6181 5034 6197 5044
rect 6245 5040 6260 5055
rect 6263 5052 6264 5064
rect 6271 5052 6298 5064
rect 6263 5044 6298 5052
rect 6263 5043 6292 5044
rect 5983 5030 6197 5034
rect 5998 5028 6197 5030
rect 6232 5030 6245 5040
rect 6263 5030 6280 5043
rect 6232 5028 6280 5030
rect 5874 5024 5907 5028
rect 5870 5022 5907 5024
rect 5870 5021 5937 5022
rect 5870 5016 5901 5021
rect 5907 5016 5937 5021
rect 5870 5012 5937 5016
rect 5843 5009 5937 5012
rect 5843 5002 5892 5009
rect 5843 4996 5873 5002
rect 5892 4997 5897 5002
rect 5809 4980 5889 4996
rect 5901 4988 5937 5009
rect 5998 5004 6187 5028
rect 6232 5027 6279 5028
rect 6245 5022 6279 5027
rect 6013 5001 6187 5004
rect 6006 4998 6187 5001
rect 6215 5021 6279 5022
rect 5809 4978 5828 4980
rect 5843 4978 5877 4980
rect 5809 4962 5889 4978
rect 5809 4956 5828 4962
rect 5525 4930 5628 4940
rect 5479 4928 5628 4930
rect 5649 4928 5684 4940
rect 5318 4926 5480 4928
rect 5330 4906 5349 4926
rect 5364 4924 5394 4926
rect 5213 4898 5254 4906
rect 5336 4902 5349 4906
rect 5401 4910 5480 4926
rect 5512 4926 5684 4928
rect 5512 4910 5591 4926
rect 5598 4924 5628 4926
rect 5176 4888 5205 4898
rect 5219 4888 5248 4898
rect 5263 4888 5293 4902
rect 5336 4888 5379 4902
rect 5401 4898 5591 4910
rect 5656 4906 5662 4926
rect 5386 4888 5416 4898
rect 5417 4888 5575 4898
rect 5579 4888 5609 4898
rect 5613 4888 5643 4902
rect 5671 4888 5684 4926
rect 5756 4940 5785 4956
rect 5799 4940 5828 4956
rect 5843 4946 5873 4962
rect 5901 4940 5907 4988
rect 5910 4982 5929 4988
rect 5944 4982 5974 4990
rect 5910 4974 5974 4982
rect 5910 4958 5990 4974
rect 6006 4967 6068 4998
rect 6084 4967 6146 4998
rect 6215 4996 6264 5021
rect 6279 4996 6309 5012
rect 6178 4982 6208 4990
rect 6215 4988 6325 4996
rect 6178 4974 6223 4982
rect 5910 4956 5929 4958
rect 5944 4956 5990 4958
rect 5910 4940 5990 4956
rect 6017 4954 6052 4967
rect 6093 4964 6130 4967
rect 6093 4962 6135 4964
rect 6022 4951 6052 4954
rect 6031 4947 6038 4951
rect 6038 4946 6039 4947
rect 5997 4940 6007 4946
rect 5756 4932 5791 4940
rect 5756 4906 5757 4932
rect 5764 4906 5791 4932
rect 5699 4888 5729 4902
rect 5756 4898 5791 4906
rect 5793 4932 5834 4940
rect 5793 4906 5808 4932
rect 5815 4906 5834 4932
rect 5898 4928 5929 4940
rect 5944 4928 6047 4940
rect 6059 4930 6085 4956
rect 6100 4951 6130 4962
rect 6162 4958 6224 4974
rect 6162 4956 6208 4958
rect 6162 4940 6224 4956
rect 6236 4940 6242 4988
rect 6245 4980 6325 4988
rect 6245 4978 6264 4980
rect 6279 4978 6313 4980
rect 6245 4962 6325 4978
rect 6245 4940 6264 4962
rect 6279 4946 6309 4962
rect 6337 4956 6343 5030
rect 6346 4956 6365 5100
rect 6380 4956 6386 5100
rect 6395 5030 6408 5100
rect 6460 5096 6482 5100
rect 6453 5074 6482 5088
rect 6535 5074 6551 5088
rect 6589 5084 6595 5086
rect 6602 5084 6710 5100
rect 6717 5084 6723 5086
rect 6731 5084 6746 5100
rect 6812 5094 6831 5097
rect 6453 5072 6551 5074
rect 6578 5072 6746 5084
rect 6761 5074 6777 5088
rect 6812 5075 6834 5094
rect 6844 5088 6860 5089
rect 6843 5086 6860 5088
rect 6844 5081 6860 5086
rect 6834 5074 6840 5075
rect 6843 5074 6872 5081
rect 6761 5073 6872 5074
rect 6761 5072 6878 5073
rect 6437 5064 6488 5072
rect 6535 5064 6569 5072
rect 6437 5052 6462 5064
rect 6469 5052 6488 5064
rect 6542 5062 6569 5064
rect 6578 5062 6799 5072
rect 6834 5069 6840 5072
rect 6542 5058 6799 5062
rect 6437 5044 6488 5052
rect 6535 5044 6799 5058
rect 6843 5064 6878 5072
rect 6389 4996 6408 5030
rect 6453 5036 6482 5044
rect 6453 5030 6470 5036
rect 6453 5028 6487 5030
rect 6535 5028 6551 5044
rect 6552 5034 6760 5044
rect 6761 5034 6777 5044
rect 6825 5040 6840 5055
rect 6843 5052 6844 5064
rect 6851 5052 6878 5064
rect 6843 5044 6878 5052
rect 6843 5043 6872 5044
rect 6563 5030 6777 5034
rect 6578 5028 6777 5030
rect 6812 5030 6825 5040
rect 6843 5030 6860 5043
rect 6812 5028 6860 5030
rect 6454 5024 6487 5028
rect 6450 5022 6487 5024
rect 6450 5021 6517 5022
rect 6450 5016 6481 5021
rect 6487 5016 6517 5021
rect 6450 5012 6517 5016
rect 6423 5009 6517 5012
rect 6423 5002 6472 5009
rect 6423 4996 6453 5002
rect 6472 4997 6477 5002
rect 6389 4980 6469 4996
rect 6481 4988 6517 5009
rect 6578 5004 6767 5028
rect 6812 5027 6859 5028
rect 6825 5022 6859 5027
rect 6593 5001 6767 5004
rect 6586 4998 6767 5001
rect 6795 5021 6859 5022
rect 6389 4978 6408 4980
rect 6423 4978 6457 4980
rect 6389 4962 6469 4978
rect 6389 4956 6408 4962
rect 6105 4930 6208 4940
rect 6059 4928 6208 4930
rect 6229 4928 6264 4940
rect 5898 4926 6060 4928
rect 5910 4906 5929 4926
rect 5944 4924 5974 4926
rect 5793 4898 5834 4906
rect 5916 4902 5929 4906
rect 5981 4910 6060 4926
rect 6092 4926 6264 4928
rect 6092 4910 6171 4926
rect 6178 4924 6208 4926
rect 5756 4888 5785 4898
rect 5799 4888 5828 4898
rect 5843 4888 5873 4902
rect 5916 4888 5959 4902
rect 5981 4898 6171 4910
rect 6236 4906 6242 4926
rect 5966 4888 5996 4898
rect 5997 4888 6155 4898
rect 6159 4888 6189 4898
rect 6193 4888 6223 4902
rect 6251 4888 6264 4926
rect 6336 4940 6365 4956
rect 6379 4940 6408 4956
rect 6423 4946 6453 4962
rect 6481 4940 6487 4988
rect 6490 4982 6509 4988
rect 6524 4982 6554 4990
rect 6490 4974 6554 4982
rect 6490 4958 6570 4974
rect 6586 4967 6648 4998
rect 6664 4967 6726 4998
rect 6795 4996 6844 5021
rect 6859 4996 6889 5012
rect 6758 4982 6788 4990
rect 6795 4988 6905 4996
rect 6758 4974 6803 4982
rect 6490 4956 6509 4958
rect 6524 4956 6570 4958
rect 6490 4940 6570 4956
rect 6597 4954 6632 4967
rect 6673 4964 6710 4967
rect 6673 4962 6715 4964
rect 6602 4951 6632 4954
rect 6611 4947 6618 4951
rect 6618 4946 6619 4947
rect 6577 4940 6587 4946
rect 6336 4932 6371 4940
rect 6336 4906 6337 4932
rect 6344 4906 6371 4932
rect 6279 4888 6309 4902
rect 6336 4898 6371 4906
rect 6373 4932 6414 4940
rect 6373 4906 6388 4932
rect 6395 4906 6414 4932
rect 6478 4928 6509 4940
rect 6524 4928 6627 4940
rect 6639 4930 6665 4956
rect 6680 4951 6710 4962
rect 6742 4958 6804 4974
rect 6742 4956 6788 4958
rect 6742 4940 6804 4956
rect 6816 4940 6822 4988
rect 6825 4980 6905 4988
rect 6825 4978 6844 4980
rect 6859 4978 6893 4980
rect 6825 4962 6905 4978
rect 6825 4940 6844 4962
rect 6859 4946 6889 4962
rect 6917 4956 6923 5030
rect 6926 4956 6945 5100
rect 6960 4956 6966 5100
rect 6975 5030 6988 5100
rect 7040 5096 7062 5100
rect 7033 5074 7062 5088
rect 7115 5074 7131 5088
rect 7169 5084 7175 5086
rect 7182 5084 7290 5100
rect 7297 5084 7303 5086
rect 7311 5084 7326 5100
rect 7392 5094 7411 5097
rect 7033 5072 7131 5074
rect 7158 5072 7326 5084
rect 7341 5074 7357 5088
rect 7392 5075 7414 5094
rect 7424 5088 7440 5089
rect 7423 5086 7440 5088
rect 7424 5081 7440 5086
rect 7414 5074 7420 5075
rect 7423 5074 7452 5081
rect 7341 5073 7452 5074
rect 7341 5072 7458 5073
rect 7017 5064 7068 5072
rect 7115 5064 7149 5072
rect 7017 5052 7042 5064
rect 7049 5052 7068 5064
rect 7122 5062 7149 5064
rect 7158 5062 7379 5072
rect 7414 5069 7420 5072
rect 7122 5058 7379 5062
rect 7017 5044 7068 5052
rect 7115 5044 7379 5058
rect 7423 5064 7458 5072
rect 6969 4996 6988 5030
rect 7033 5036 7062 5044
rect 7033 5030 7050 5036
rect 7033 5028 7067 5030
rect 7115 5028 7131 5044
rect 7132 5034 7340 5044
rect 7341 5034 7357 5044
rect 7405 5040 7420 5055
rect 7423 5052 7424 5064
rect 7431 5052 7458 5064
rect 7423 5044 7458 5052
rect 7423 5043 7452 5044
rect 7143 5030 7357 5034
rect 7158 5028 7357 5030
rect 7392 5030 7405 5040
rect 7423 5030 7440 5043
rect 7392 5028 7440 5030
rect 7034 5024 7067 5028
rect 7030 5022 7067 5024
rect 7030 5021 7097 5022
rect 7030 5016 7061 5021
rect 7067 5016 7097 5021
rect 7030 5012 7097 5016
rect 7003 5009 7097 5012
rect 7003 5002 7052 5009
rect 7003 4996 7033 5002
rect 7052 4997 7057 5002
rect 6969 4980 7049 4996
rect 7061 4988 7097 5009
rect 7158 5004 7347 5028
rect 7392 5027 7439 5028
rect 7405 5022 7439 5027
rect 7173 5001 7347 5004
rect 7166 4998 7347 5001
rect 7375 5021 7439 5022
rect 6969 4978 6988 4980
rect 7003 4978 7037 4980
rect 6969 4962 7049 4978
rect 6969 4956 6988 4962
rect 6685 4930 6788 4940
rect 6639 4928 6788 4930
rect 6809 4928 6844 4940
rect 6478 4926 6640 4928
rect 6490 4906 6509 4926
rect 6524 4924 6554 4926
rect 6373 4898 6414 4906
rect 6496 4902 6509 4906
rect 6561 4910 6640 4926
rect 6672 4926 6844 4928
rect 6672 4910 6751 4926
rect 6758 4924 6788 4926
rect 6336 4888 6365 4898
rect 6379 4888 6408 4898
rect 6423 4888 6453 4902
rect 6496 4888 6539 4902
rect 6561 4898 6751 4910
rect 6816 4906 6822 4926
rect 6546 4888 6576 4898
rect 6577 4888 6735 4898
rect 6739 4888 6769 4898
rect 6773 4888 6803 4902
rect 6831 4888 6844 4926
rect 6916 4940 6945 4956
rect 6959 4940 6988 4956
rect 7003 4946 7033 4962
rect 7061 4940 7067 4988
rect 7070 4982 7089 4988
rect 7104 4982 7134 4990
rect 7070 4974 7134 4982
rect 7070 4958 7150 4974
rect 7166 4967 7228 4998
rect 7244 4967 7306 4998
rect 7375 4996 7424 5021
rect 7439 4996 7469 5012
rect 7338 4982 7368 4990
rect 7375 4988 7485 4996
rect 7338 4974 7383 4982
rect 7070 4956 7089 4958
rect 7104 4956 7150 4958
rect 7070 4940 7150 4956
rect 7177 4954 7212 4967
rect 7253 4964 7290 4967
rect 7253 4962 7295 4964
rect 7182 4951 7212 4954
rect 7191 4947 7198 4951
rect 7198 4946 7199 4947
rect 7157 4940 7167 4946
rect 6916 4932 6951 4940
rect 6916 4906 6917 4932
rect 6924 4906 6951 4932
rect 6859 4888 6889 4902
rect 6916 4898 6951 4906
rect 6953 4932 6994 4940
rect 6953 4906 6968 4932
rect 6975 4906 6994 4932
rect 7058 4928 7089 4940
rect 7104 4928 7207 4940
rect 7219 4930 7245 4956
rect 7260 4951 7290 4962
rect 7322 4958 7384 4974
rect 7322 4956 7368 4958
rect 7322 4940 7384 4956
rect 7396 4940 7402 4988
rect 7405 4980 7485 4988
rect 7405 4978 7424 4980
rect 7439 4978 7473 4980
rect 7405 4962 7485 4978
rect 7405 4940 7424 4962
rect 7439 4946 7469 4962
rect 7497 4956 7503 5030
rect 7506 4956 7525 5100
rect 7540 4956 7546 5100
rect 7555 5030 7568 5100
rect 7620 5096 7642 5100
rect 7613 5074 7642 5088
rect 7695 5074 7711 5088
rect 7749 5084 7755 5086
rect 7762 5084 7870 5100
rect 7877 5084 7883 5086
rect 7891 5084 7906 5100
rect 7972 5094 7991 5097
rect 7613 5072 7711 5074
rect 7738 5072 7906 5084
rect 7921 5074 7937 5088
rect 7972 5075 7994 5094
rect 8004 5088 8020 5089
rect 8003 5086 8020 5088
rect 8004 5081 8020 5086
rect 7994 5074 8000 5075
rect 8003 5074 8032 5081
rect 7921 5073 8032 5074
rect 7921 5072 8038 5073
rect 7597 5064 7648 5072
rect 7695 5064 7729 5072
rect 7597 5052 7622 5064
rect 7629 5052 7648 5064
rect 7702 5062 7729 5064
rect 7738 5062 7959 5072
rect 7994 5069 8000 5072
rect 7702 5058 7959 5062
rect 7597 5044 7648 5052
rect 7695 5044 7959 5058
rect 8003 5064 8038 5072
rect 7549 4996 7568 5030
rect 7613 5036 7642 5044
rect 7613 5030 7630 5036
rect 7613 5028 7647 5030
rect 7695 5028 7711 5044
rect 7712 5034 7920 5044
rect 7921 5034 7937 5044
rect 7985 5040 8000 5055
rect 8003 5052 8004 5064
rect 8011 5052 8038 5064
rect 8003 5044 8038 5052
rect 8003 5043 8032 5044
rect 7723 5030 7937 5034
rect 7738 5028 7937 5030
rect 7972 5030 7985 5040
rect 8003 5030 8020 5043
rect 7972 5028 8020 5030
rect 7614 5024 7647 5028
rect 7610 5022 7647 5024
rect 7610 5021 7677 5022
rect 7610 5016 7641 5021
rect 7647 5016 7677 5021
rect 7610 5012 7677 5016
rect 7583 5009 7677 5012
rect 7583 5002 7632 5009
rect 7583 4996 7613 5002
rect 7632 4997 7637 5002
rect 7549 4980 7629 4996
rect 7641 4988 7677 5009
rect 7738 5004 7927 5028
rect 7972 5027 8019 5028
rect 7985 5022 8019 5027
rect 7753 5001 7927 5004
rect 7746 4998 7927 5001
rect 7955 5021 8019 5022
rect 7549 4978 7568 4980
rect 7583 4978 7617 4980
rect 7549 4962 7629 4978
rect 7549 4956 7568 4962
rect 7265 4930 7368 4940
rect 7219 4928 7368 4930
rect 7389 4928 7424 4940
rect 7058 4926 7220 4928
rect 7070 4906 7089 4926
rect 7104 4924 7134 4926
rect 6953 4898 6994 4906
rect 7076 4902 7089 4906
rect 7141 4910 7220 4926
rect 7252 4926 7424 4928
rect 7252 4910 7331 4926
rect 7338 4924 7368 4926
rect 6916 4888 6945 4898
rect 6959 4888 6988 4898
rect 7003 4888 7033 4902
rect 7076 4888 7119 4902
rect 7141 4898 7331 4910
rect 7396 4906 7402 4926
rect 7126 4888 7156 4898
rect 7157 4888 7315 4898
rect 7319 4888 7349 4898
rect 7353 4888 7383 4902
rect 7411 4888 7424 4926
rect 7496 4940 7525 4956
rect 7539 4940 7568 4956
rect 7583 4946 7613 4962
rect 7641 4940 7647 4988
rect 7650 4982 7669 4988
rect 7684 4982 7714 4990
rect 7650 4974 7714 4982
rect 7650 4958 7730 4974
rect 7746 4967 7808 4998
rect 7824 4967 7886 4998
rect 7955 4996 8004 5021
rect 8019 4996 8049 5012
rect 7918 4982 7948 4990
rect 7955 4988 8065 4996
rect 7918 4974 7963 4982
rect 7650 4956 7669 4958
rect 7684 4956 7730 4958
rect 7650 4940 7730 4956
rect 7757 4954 7792 4967
rect 7833 4964 7870 4967
rect 7833 4962 7875 4964
rect 7762 4951 7792 4954
rect 7771 4947 7778 4951
rect 7778 4946 7779 4947
rect 7737 4940 7747 4946
rect 7496 4932 7531 4940
rect 7496 4906 7497 4932
rect 7504 4906 7531 4932
rect 7439 4888 7469 4902
rect 7496 4898 7531 4906
rect 7533 4932 7574 4940
rect 7533 4906 7548 4932
rect 7555 4906 7574 4932
rect 7638 4928 7669 4940
rect 7684 4928 7787 4940
rect 7799 4930 7825 4956
rect 7840 4951 7870 4962
rect 7902 4958 7964 4974
rect 7902 4956 7948 4958
rect 7902 4940 7964 4956
rect 7976 4940 7982 4988
rect 7985 4980 8065 4988
rect 7985 4978 8004 4980
rect 8019 4978 8053 4980
rect 7985 4962 8065 4978
rect 7985 4940 8004 4962
rect 8019 4946 8049 4962
rect 8077 4956 8083 5030
rect 8086 4956 8105 5100
rect 8120 4956 8126 5100
rect 8135 5030 8148 5100
rect 8200 5096 8222 5100
rect 8193 5074 8222 5088
rect 8275 5074 8291 5088
rect 8329 5084 8335 5086
rect 8342 5084 8450 5100
rect 8457 5084 8463 5086
rect 8471 5084 8486 5100
rect 8552 5094 8571 5097
rect 8193 5072 8291 5074
rect 8318 5072 8486 5084
rect 8501 5074 8517 5088
rect 8552 5075 8574 5094
rect 8584 5088 8600 5089
rect 8583 5086 8600 5088
rect 8584 5081 8600 5086
rect 8574 5074 8580 5075
rect 8583 5074 8612 5081
rect 8501 5073 8612 5074
rect 8501 5072 8618 5073
rect 8177 5064 8228 5072
rect 8275 5064 8309 5072
rect 8177 5052 8202 5064
rect 8209 5052 8228 5064
rect 8282 5062 8309 5064
rect 8318 5062 8539 5072
rect 8574 5069 8580 5072
rect 8282 5058 8539 5062
rect 8177 5044 8228 5052
rect 8275 5044 8539 5058
rect 8583 5064 8618 5072
rect 8129 4996 8148 5030
rect 8193 5036 8222 5044
rect 8193 5030 8210 5036
rect 8193 5028 8227 5030
rect 8275 5028 8291 5044
rect 8292 5034 8500 5044
rect 8501 5034 8517 5044
rect 8565 5040 8580 5055
rect 8583 5052 8584 5064
rect 8591 5052 8618 5064
rect 8583 5044 8618 5052
rect 8583 5043 8612 5044
rect 8303 5030 8517 5034
rect 8318 5028 8517 5030
rect 8552 5030 8565 5040
rect 8583 5030 8600 5043
rect 8552 5028 8600 5030
rect 8194 5024 8227 5028
rect 8190 5022 8227 5024
rect 8190 5021 8257 5022
rect 8190 5016 8221 5021
rect 8227 5016 8257 5021
rect 8190 5012 8257 5016
rect 8163 5009 8257 5012
rect 8163 5002 8212 5009
rect 8163 4996 8193 5002
rect 8212 4997 8217 5002
rect 8129 4980 8209 4996
rect 8221 4988 8257 5009
rect 8318 5004 8507 5028
rect 8552 5027 8599 5028
rect 8565 5022 8599 5027
rect 8333 5001 8507 5004
rect 8326 4998 8507 5001
rect 8535 5021 8599 5022
rect 8129 4978 8148 4980
rect 8163 4978 8197 4980
rect 8129 4962 8209 4978
rect 8129 4956 8148 4962
rect 7845 4930 7948 4940
rect 7799 4928 7948 4930
rect 7969 4928 8004 4940
rect 7638 4926 7800 4928
rect 7650 4906 7669 4926
rect 7684 4924 7714 4926
rect 7533 4898 7574 4906
rect 7656 4902 7669 4906
rect 7721 4910 7800 4926
rect 7832 4926 8004 4928
rect 7832 4910 7911 4926
rect 7918 4924 7948 4926
rect 7496 4888 7525 4898
rect 7539 4888 7568 4898
rect 7583 4888 7613 4902
rect 7656 4888 7699 4902
rect 7721 4898 7911 4910
rect 7976 4906 7982 4926
rect 7706 4888 7736 4898
rect 7737 4888 7895 4898
rect 7899 4888 7929 4898
rect 7933 4888 7963 4902
rect 7991 4888 8004 4926
rect 8076 4940 8105 4956
rect 8119 4940 8148 4956
rect 8163 4946 8193 4962
rect 8221 4940 8227 4988
rect 8230 4982 8249 4988
rect 8264 4982 8294 4990
rect 8230 4974 8294 4982
rect 8230 4958 8310 4974
rect 8326 4967 8388 4998
rect 8404 4967 8466 4998
rect 8535 4996 8584 5021
rect 8599 4996 8629 5012
rect 8498 4982 8528 4990
rect 8535 4988 8645 4996
rect 8498 4974 8543 4982
rect 8230 4956 8249 4958
rect 8264 4956 8310 4958
rect 8230 4940 8310 4956
rect 8337 4954 8372 4967
rect 8413 4964 8450 4967
rect 8413 4962 8455 4964
rect 8342 4951 8372 4954
rect 8351 4947 8358 4951
rect 8358 4946 8359 4947
rect 8317 4940 8327 4946
rect 8076 4932 8111 4940
rect 8076 4906 8077 4932
rect 8084 4906 8111 4932
rect 8019 4888 8049 4902
rect 8076 4898 8111 4906
rect 8113 4932 8154 4940
rect 8113 4906 8128 4932
rect 8135 4906 8154 4932
rect 8218 4928 8249 4940
rect 8264 4928 8367 4940
rect 8379 4930 8405 4956
rect 8420 4951 8450 4962
rect 8482 4958 8544 4974
rect 8482 4956 8528 4958
rect 8482 4940 8544 4956
rect 8556 4940 8562 4988
rect 8565 4980 8645 4988
rect 8565 4978 8584 4980
rect 8599 4978 8633 4980
rect 8565 4962 8645 4978
rect 8565 4940 8584 4962
rect 8599 4946 8629 4962
rect 8657 4956 8663 5030
rect 8666 4956 8685 5100
rect 8700 4956 8706 5100
rect 8715 5030 8728 5100
rect 8780 5096 8802 5100
rect 8773 5074 8802 5088
rect 8855 5074 8871 5088
rect 8909 5084 8915 5086
rect 8922 5084 9030 5100
rect 9037 5084 9043 5086
rect 9051 5084 9066 5100
rect 9132 5094 9151 5097
rect 8773 5072 8871 5074
rect 8898 5072 9066 5084
rect 9081 5074 9097 5088
rect 9132 5075 9154 5094
rect 9164 5088 9180 5089
rect 9163 5086 9180 5088
rect 9164 5081 9180 5086
rect 9154 5074 9160 5075
rect 9163 5074 9192 5081
rect 9081 5073 9192 5074
rect 9081 5072 9198 5073
rect 8757 5064 8808 5072
rect 8855 5064 8889 5072
rect 8757 5052 8782 5064
rect 8789 5052 8808 5064
rect 8862 5062 8889 5064
rect 8898 5062 9119 5072
rect 9154 5069 9160 5072
rect 8862 5058 9119 5062
rect 8757 5044 8808 5052
rect 8855 5044 9119 5058
rect 9163 5064 9198 5072
rect 8709 4996 8728 5030
rect 8773 5036 8802 5044
rect 8773 5030 8790 5036
rect 8773 5028 8807 5030
rect 8855 5028 8871 5044
rect 8872 5034 9080 5044
rect 9081 5034 9097 5044
rect 9145 5040 9160 5055
rect 9163 5052 9164 5064
rect 9171 5052 9198 5064
rect 9163 5044 9198 5052
rect 9163 5043 9192 5044
rect 8883 5030 9097 5034
rect 8898 5028 9097 5030
rect 9132 5030 9145 5040
rect 9163 5030 9180 5043
rect 9132 5028 9180 5030
rect 8774 5024 8807 5028
rect 8770 5022 8807 5024
rect 8770 5021 8837 5022
rect 8770 5016 8801 5021
rect 8807 5016 8837 5021
rect 8770 5012 8837 5016
rect 8743 5009 8837 5012
rect 8743 5002 8792 5009
rect 8743 4996 8773 5002
rect 8792 4997 8797 5002
rect 8709 4980 8789 4996
rect 8801 4988 8837 5009
rect 8898 5004 9087 5028
rect 9132 5027 9179 5028
rect 9145 5022 9179 5027
rect 8913 5001 9087 5004
rect 8906 4998 9087 5001
rect 9115 5021 9179 5022
rect 8709 4978 8728 4980
rect 8743 4978 8777 4980
rect 8709 4962 8789 4978
rect 8709 4956 8728 4962
rect 8425 4930 8528 4940
rect 8379 4928 8528 4930
rect 8549 4928 8584 4940
rect 8218 4926 8380 4928
rect 8230 4906 8249 4926
rect 8264 4924 8294 4926
rect 8113 4898 8154 4906
rect 8236 4902 8249 4906
rect 8301 4910 8380 4926
rect 8412 4926 8584 4928
rect 8412 4910 8491 4926
rect 8498 4924 8528 4926
rect 8076 4888 8105 4898
rect 8119 4888 8148 4898
rect 8163 4888 8193 4902
rect 8236 4888 8279 4902
rect 8301 4898 8491 4910
rect 8556 4906 8562 4926
rect 8286 4888 8316 4898
rect 8317 4888 8475 4898
rect 8479 4888 8509 4898
rect 8513 4888 8543 4902
rect 8571 4888 8584 4926
rect 8656 4940 8685 4956
rect 8699 4940 8728 4956
rect 8743 4946 8773 4962
rect 8801 4940 8807 4988
rect 8810 4982 8829 4988
rect 8844 4982 8874 4990
rect 8810 4974 8874 4982
rect 8810 4958 8890 4974
rect 8906 4967 8968 4998
rect 8984 4967 9046 4998
rect 9115 4996 9164 5021
rect 9179 4996 9209 5012
rect 9078 4982 9108 4990
rect 9115 4988 9225 4996
rect 9078 4974 9123 4982
rect 8810 4956 8829 4958
rect 8844 4956 8890 4958
rect 8810 4940 8890 4956
rect 8917 4954 8952 4967
rect 8993 4964 9030 4967
rect 8993 4962 9035 4964
rect 8922 4951 8952 4954
rect 8931 4947 8938 4951
rect 8938 4946 8939 4947
rect 8897 4940 8907 4946
rect 8656 4932 8691 4940
rect 8656 4906 8657 4932
rect 8664 4906 8691 4932
rect 8599 4888 8629 4902
rect 8656 4898 8691 4906
rect 8693 4932 8734 4940
rect 8693 4906 8708 4932
rect 8715 4906 8734 4932
rect 8798 4928 8829 4940
rect 8844 4928 8947 4940
rect 8959 4930 8985 4956
rect 9000 4951 9030 4962
rect 9062 4958 9124 4974
rect 9062 4956 9108 4958
rect 9062 4940 9124 4956
rect 9136 4940 9142 4988
rect 9145 4980 9225 4988
rect 9145 4978 9164 4980
rect 9179 4978 9213 4980
rect 9145 4962 9225 4978
rect 9145 4940 9164 4962
rect 9179 4946 9209 4962
rect 9237 4956 9243 5030
rect 9246 4956 9265 5100
rect 9280 4956 9286 5100
rect 9295 5030 9308 5100
rect 9360 5096 9382 5100
rect 9353 5074 9382 5088
rect 9435 5074 9451 5088
rect 9489 5084 9495 5086
rect 9502 5084 9610 5100
rect 9617 5084 9623 5086
rect 9631 5084 9646 5100
rect 9712 5094 9731 5097
rect 9353 5072 9451 5074
rect 9478 5072 9646 5084
rect 9661 5074 9677 5088
rect 9712 5075 9734 5094
rect 9744 5088 9760 5089
rect 9743 5086 9760 5088
rect 9744 5081 9760 5086
rect 9734 5074 9740 5075
rect 9743 5074 9772 5081
rect 9661 5073 9772 5074
rect 9661 5072 9778 5073
rect 9337 5064 9388 5072
rect 9435 5064 9469 5072
rect 9337 5052 9362 5064
rect 9369 5052 9388 5064
rect 9442 5062 9469 5064
rect 9478 5062 9699 5072
rect 9734 5069 9740 5072
rect 9442 5058 9699 5062
rect 9337 5044 9388 5052
rect 9435 5044 9699 5058
rect 9743 5064 9778 5072
rect 9289 4996 9308 5030
rect 9353 5036 9382 5044
rect 9353 5030 9370 5036
rect 9353 5028 9387 5030
rect 9435 5028 9451 5044
rect 9452 5034 9660 5044
rect 9661 5034 9677 5044
rect 9725 5040 9740 5055
rect 9743 5052 9744 5064
rect 9751 5052 9778 5064
rect 9743 5044 9778 5052
rect 9743 5043 9772 5044
rect 9463 5030 9677 5034
rect 9478 5028 9677 5030
rect 9712 5030 9725 5040
rect 9743 5030 9760 5043
rect 9712 5028 9760 5030
rect 9354 5024 9387 5028
rect 9350 5022 9387 5024
rect 9350 5021 9417 5022
rect 9350 5016 9381 5021
rect 9387 5016 9417 5021
rect 9350 5012 9417 5016
rect 9323 5009 9417 5012
rect 9323 5002 9372 5009
rect 9323 4996 9353 5002
rect 9372 4997 9377 5002
rect 9289 4980 9369 4996
rect 9381 4988 9417 5009
rect 9478 5004 9667 5028
rect 9712 5027 9759 5028
rect 9725 5022 9759 5027
rect 9493 5001 9667 5004
rect 9486 4998 9667 5001
rect 9695 5021 9759 5022
rect 9289 4978 9308 4980
rect 9323 4978 9357 4980
rect 9289 4962 9369 4978
rect 9289 4956 9308 4962
rect 9005 4930 9108 4940
rect 8959 4928 9108 4930
rect 9129 4928 9164 4940
rect 8798 4926 8960 4928
rect 8810 4906 8829 4926
rect 8844 4924 8874 4926
rect 8693 4898 8734 4906
rect 8816 4902 8829 4906
rect 8881 4910 8960 4926
rect 8992 4926 9164 4928
rect 8992 4910 9071 4926
rect 9078 4924 9108 4926
rect 8656 4888 8685 4898
rect 8699 4888 8728 4898
rect 8743 4888 8773 4902
rect 8816 4888 8859 4902
rect 8881 4898 9071 4910
rect 9136 4906 9142 4926
rect 8866 4888 8896 4898
rect 8897 4888 9055 4898
rect 9059 4888 9089 4898
rect 9093 4888 9123 4902
rect 9151 4888 9164 4926
rect 9236 4940 9265 4956
rect 9279 4940 9308 4956
rect 9323 4946 9353 4962
rect 9381 4940 9387 4988
rect 9390 4982 9409 4988
rect 9424 4982 9454 4990
rect 9390 4974 9454 4982
rect 9390 4958 9470 4974
rect 9486 4967 9548 4998
rect 9564 4967 9626 4998
rect 9695 4996 9744 5021
rect 9759 4996 9789 5012
rect 9658 4982 9688 4990
rect 9695 4988 9805 4996
rect 9658 4974 9703 4982
rect 9390 4956 9409 4958
rect 9424 4956 9470 4958
rect 9390 4940 9470 4956
rect 9497 4954 9532 4967
rect 9573 4964 9610 4967
rect 9573 4962 9615 4964
rect 9502 4951 9532 4954
rect 9511 4947 9518 4951
rect 9518 4946 9519 4947
rect 9477 4940 9487 4946
rect 9236 4932 9271 4940
rect 9236 4906 9237 4932
rect 9244 4906 9271 4932
rect 9179 4888 9209 4902
rect 9236 4898 9271 4906
rect 9273 4932 9314 4940
rect 9273 4906 9288 4932
rect 9295 4906 9314 4932
rect 9378 4928 9409 4940
rect 9424 4928 9527 4940
rect 9539 4930 9565 4956
rect 9580 4951 9610 4962
rect 9642 4958 9704 4974
rect 9642 4956 9688 4958
rect 9642 4940 9704 4956
rect 9716 4940 9722 4988
rect 9725 4980 9805 4988
rect 9725 4978 9744 4980
rect 9759 4978 9793 4980
rect 9725 4962 9805 4978
rect 9725 4940 9744 4962
rect 9759 4946 9789 4962
rect 9817 4956 9823 5030
rect 9826 4956 9845 5100
rect 9860 4956 9866 5100
rect 9875 5030 9888 5100
rect 9940 5096 9962 5100
rect 9933 5074 9962 5088
rect 10015 5074 10031 5088
rect 10069 5084 10075 5086
rect 10082 5084 10190 5100
rect 10197 5084 10203 5086
rect 10211 5084 10226 5100
rect 10292 5094 10311 5097
rect 9933 5072 10031 5074
rect 10058 5072 10226 5084
rect 10241 5074 10257 5088
rect 10292 5075 10314 5094
rect 10324 5088 10340 5089
rect 10323 5086 10340 5088
rect 10324 5081 10340 5086
rect 10314 5074 10320 5075
rect 10323 5074 10352 5081
rect 10241 5073 10352 5074
rect 10241 5072 10358 5073
rect 9917 5064 9968 5072
rect 10015 5064 10049 5072
rect 9917 5052 9942 5064
rect 9949 5052 9968 5064
rect 10022 5062 10049 5064
rect 10058 5062 10279 5072
rect 10314 5069 10320 5072
rect 10022 5058 10279 5062
rect 9917 5044 9968 5052
rect 10015 5044 10279 5058
rect 10323 5064 10358 5072
rect 9869 4996 9888 5030
rect 9933 5036 9962 5044
rect 9933 5030 9950 5036
rect 9933 5028 9967 5030
rect 10015 5028 10031 5044
rect 10032 5034 10240 5044
rect 10241 5034 10257 5044
rect 10305 5040 10320 5055
rect 10323 5052 10324 5064
rect 10331 5052 10358 5064
rect 10323 5044 10358 5052
rect 10323 5043 10352 5044
rect 10043 5030 10257 5034
rect 10058 5028 10257 5030
rect 10292 5030 10305 5040
rect 10323 5030 10340 5043
rect 10292 5028 10340 5030
rect 9934 5024 9967 5028
rect 9930 5022 9967 5024
rect 9930 5021 9997 5022
rect 9930 5016 9961 5021
rect 9967 5016 9997 5021
rect 9930 5012 9997 5016
rect 9903 5009 9997 5012
rect 9903 5002 9952 5009
rect 9903 4996 9933 5002
rect 9952 4997 9957 5002
rect 9869 4980 9949 4996
rect 9961 4988 9997 5009
rect 10058 5004 10247 5028
rect 10292 5027 10339 5028
rect 10305 5022 10339 5027
rect 10073 5001 10247 5004
rect 10066 4998 10247 5001
rect 10275 5021 10339 5022
rect 9869 4978 9888 4980
rect 9903 4978 9937 4980
rect 9869 4962 9949 4978
rect 9869 4956 9888 4962
rect 9585 4930 9688 4940
rect 9539 4928 9688 4930
rect 9709 4928 9744 4940
rect 9378 4926 9540 4928
rect 9390 4906 9409 4926
rect 9424 4924 9454 4926
rect 9273 4898 9314 4906
rect 9396 4902 9409 4906
rect 9461 4910 9540 4926
rect 9572 4926 9744 4928
rect 9572 4910 9651 4926
rect 9658 4924 9688 4926
rect 9236 4888 9265 4898
rect 9279 4888 9308 4898
rect 9323 4888 9353 4902
rect 9396 4888 9439 4902
rect 9461 4898 9651 4910
rect 9716 4906 9722 4926
rect 9446 4888 9476 4898
rect 9477 4888 9635 4898
rect 9639 4888 9669 4898
rect 9673 4888 9703 4902
rect 9731 4888 9744 4926
rect 9816 4940 9845 4956
rect 9859 4940 9888 4956
rect 9903 4946 9933 4962
rect 9961 4940 9967 4988
rect 9970 4982 9989 4988
rect 10004 4982 10034 4990
rect 9970 4974 10034 4982
rect 9970 4958 10050 4974
rect 10066 4967 10128 4998
rect 10144 4967 10206 4998
rect 10275 4996 10324 5021
rect 10339 4996 10369 5012
rect 10238 4982 10268 4990
rect 10275 4988 10385 4996
rect 10238 4974 10283 4982
rect 9970 4956 9989 4958
rect 10004 4956 10050 4958
rect 9970 4940 10050 4956
rect 10077 4954 10112 4967
rect 10153 4964 10190 4967
rect 10153 4962 10195 4964
rect 10082 4951 10112 4954
rect 10091 4947 10098 4951
rect 10098 4946 10099 4947
rect 10057 4940 10067 4946
rect 9816 4932 9851 4940
rect 9816 4906 9817 4932
rect 9824 4906 9851 4932
rect 9759 4888 9789 4902
rect 9816 4898 9851 4906
rect 9853 4932 9894 4940
rect 9853 4906 9868 4932
rect 9875 4906 9894 4932
rect 9958 4928 9989 4940
rect 10004 4928 10107 4940
rect 10119 4930 10145 4956
rect 10160 4951 10190 4962
rect 10222 4958 10284 4974
rect 10222 4956 10268 4958
rect 10222 4940 10284 4956
rect 10296 4940 10302 4988
rect 10305 4980 10385 4988
rect 10305 4978 10324 4980
rect 10339 4978 10373 4980
rect 10305 4962 10385 4978
rect 10305 4940 10324 4962
rect 10339 4946 10369 4962
rect 10397 4956 10403 5030
rect 10406 4956 10425 5100
rect 10440 4956 10446 5100
rect 10455 5030 10468 5100
rect 10520 5096 10542 5100
rect 10513 5074 10542 5088
rect 10595 5074 10611 5088
rect 10649 5084 10655 5086
rect 10662 5084 10770 5100
rect 10777 5084 10783 5086
rect 10791 5084 10806 5100
rect 10872 5094 10891 5097
rect 10513 5072 10611 5074
rect 10638 5072 10806 5084
rect 10821 5074 10837 5088
rect 10872 5075 10894 5094
rect 10904 5088 10920 5089
rect 10903 5086 10920 5088
rect 10904 5081 10920 5086
rect 10894 5074 10900 5075
rect 10903 5074 10932 5081
rect 10821 5073 10932 5074
rect 10821 5072 10938 5073
rect 10497 5064 10548 5072
rect 10595 5064 10629 5072
rect 10497 5052 10522 5064
rect 10529 5052 10548 5064
rect 10602 5062 10629 5064
rect 10638 5062 10859 5072
rect 10894 5069 10900 5072
rect 10602 5058 10859 5062
rect 10497 5044 10548 5052
rect 10595 5044 10859 5058
rect 10903 5064 10938 5072
rect 10449 4996 10468 5030
rect 10513 5036 10542 5044
rect 10513 5030 10530 5036
rect 10513 5028 10547 5030
rect 10595 5028 10611 5044
rect 10612 5034 10820 5044
rect 10821 5034 10837 5044
rect 10885 5040 10900 5055
rect 10903 5052 10904 5064
rect 10911 5052 10938 5064
rect 10903 5044 10938 5052
rect 10903 5043 10932 5044
rect 10623 5030 10837 5034
rect 10638 5028 10837 5030
rect 10872 5030 10885 5040
rect 10903 5030 10920 5043
rect 10872 5028 10920 5030
rect 10514 5024 10547 5028
rect 10510 5022 10547 5024
rect 10510 5021 10577 5022
rect 10510 5016 10541 5021
rect 10547 5016 10577 5021
rect 10510 5012 10577 5016
rect 10483 5009 10577 5012
rect 10483 5002 10532 5009
rect 10483 4996 10513 5002
rect 10532 4997 10537 5002
rect 10449 4980 10529 4996
rect 10541 4988 10577 5009
rect 10638 5004 10827 5028
rect 10872 5027 10919 5028
rect 10885 5022 10919 5027
rect 10653 5001 10827 5004
rect 10646 4998 10827 5001
rect 10855 5021 10919 5022
rect 10449 4978 10468 4980
rect 10483 4978 10517 4980
rect 10449 4962 10529 4978
rect 10449 4956 10468 4962
rect 10165 4930 10268 4940
rect 10119 4928 10268 4930
rect 10289 4928 10324 4940
rect 9958 4926 10120 4928
rect 9970 4906 9989 4926
rect 10004 4924 10034 4926
rect 9853 4898 9894 4906
rect 9976 4902 9989 4906
rect 10041 4910 10120 4926
rect 10152 4926 10324 4928
rect 10152 4910 10231 4926
rect 10238 4924 10268 4926
rect 9816 4888 9845 4898
rect 9859 4888 9888 4898
rect 9903 4888 9933 4902
rect 9976 4888 10019 4902
rect 10041 4898 10231 4910
rect 10296 4906 10302 4926
rect 10026 4888 10056 4898
rect 10057 4888 10215 4898
rect 10219 4888 10249 4898
rect 10253 4888 10283 4902
rect 10311 4888 10324 4926
rect 10396 4940 10425 4956
rect 10439 4940 10468 4956
rect 10483 4946 10513 4962
rect 10541 4940 10547 4988
rect 10550 4982 10569 4988
rect 10584 4982 10614 4990
rect 10550 4974 10614 4982
rect 10550 4958 10630 4974
rect 10646 4967 10708 4998
rect 10724 4967 10786 4998
rect 10855 4996 10904 5021
rect 10919 4996 10949 5012
rect 10818 4982 10848 4990
rect 10855 4988 10965 4996
rect 10818 4974 10863 4982
rect 10550 4956 10569 4958
rect 10584 4956 10630 4958
rect 10550 4940 10630 4956
rect 10657 4954 10692 4967
rect 10733 4964 10770 4967
rect 10733 4962 10775 4964
rect 10662 4951 10692 4954
rect 10671 4947 10678 4951
rect 10678 4946 10679 4947
rect 10637 4940 10647 4946
rect 10396 4932 10431 4940
rect 10396 4906 10397 4932
rect 10404 4906 10431 4932
rect 10339 4888 10369 4902
rect 10396 4898 10431 4906
rect 10433 4932 10474 4940
rect 10433 4906 10448 4932
rect 10455 4906 10474 4932
rect 10538 4928 10569 4940
rect 10584 4928 10687 4940
rect 10699 4930 10725 4956
rect 10740 4951 10770 4962
rect 10802 4958 10864 4974
rect 10802 4956 10848 4958
rect 10802 4940 10864 4956
rect 10876 4940 10882 4988
rect 10885 4980 10965 4988
rect 10885 4978 10904 4980
rect 10919 4978 10953 4980
rect 10885 4962 10965 4978
rect 10885 4940 10904 4962
rect 10919 4946 10949 4962
rect 10977 4956 10983 5030
rect 10986 4956 11005 5100
rect 11020 4956 11026 5100
rect 11035 5030 11048 5100
rect 11100 5096 11122 5100
rect 11093 5074 11122 5088
rect 11175 5074 11191 5088
rect 11229 5084 11235 5086
rect 11242 5084 11350 5100
rect 11357 5084 11363 5086
rect 11371 5084 11386 5100
rect 11452 5094 11471 5097
rect 11093 5072 11191 5074
rect 11218 5072 11386 5084
rect 11401 5074 11417 5088
rect 11452 5075 11474 5094
rect 11484 5088 11500 5089
rect 11483 5086 11500 5088
rect 11484 5081 11500 5086
rect 11474 5074 11480 5075
rect 11483 5074 11512 5081
rect 11401 5073 11512 5074
rect 11401 5072 11518 5073
rect 11077 5064 11128 5072
rect 11175 5064 11209 5072
rect 11077 5052 11102 5064
rect 11109 5052 11128 5064
rect 11182 5062 11209 5064
rect 11218 5062 11439 5072
rect 11474 5069 11480 5072
rect 11182 5058 11439 5062
rect 11077 5044 11128 5052
rect 11175 5044 11439 5058
rect 11483 5064 11518 5072
rect 11029 4996 11048 5030
rect 11093 5036 11122 5044
rect 11093 5030 11110 5036
rect 11093 5028 11127 5030
rect 11175 5028 11191 5044
rect 11192 5034 11400 5044
rect 11401 5034 11417 5044
rect 11465 5040 11480 5055
rect 11483 5052 11484 5064
rect 11491 5052 11518 5064
rect 11483 5044 11518 5052
rect 11483 5043 11512 5044
rect 11203 5030 11417 5034
rect 11218 5028 11417 5030
rect 11452 5030 11465 5040
rect 11483 5030 11500 5043
rect 11452 5028 11500 5030
rect 11094 5024 11127 5028
rect 11090 5022 11127 5024
rect 11090 5021 11157 5022
rect 11090 5016 11121 5021
rect 11127 5016 11157 5021
rect 11090 5012 11157 5016
rect 11063 5009 11157 5012
rect 11063 5002 11112 5009
rect 11063 4996 11093 5002
rect 11112 4997 11117 5002
rect 11029 4980 11109 4996
rect 11121 4988 11157 5009
rect 11218 5004 11407 5028
rect 11452 5027 11499 5028
rect 11465 5022 11499 5027
rect 11233 5001 11407 5004
rect 11226 4998 11407 5001
rect 11435 5021 11499 5022
rect 11029 4978 11048 4980
rect 11063 4978 11097 4980
rect 11029 4962 11109 4978
rect 11029 4956 11048 4962
rect 10745 4930 10848 4940
rect 10699 4928 10848 4930
rect 10869 4928 10904 4940
rect 10538 4926 10700 4928
rect 10550 4906 10569 4926
rect 10584 4924 10614 4926
rect 10433 4898 10474 4906
rect 10556 4902 10569 4906
rect 10621 4910 10700 4926
rect 10732 4926 10904 4928
rect 10732 4910 10811 4926
rect 10818 4924 10848 4926
rect 10396 4888 10425 4898
rect 10439 4888 10468 4898
rect 10483 4888 10513 4902
rect 10556 4888 10599 4902
rect 10621 4898 10811 4910
rect 10876 4906 10882 4926
rect 10606 4888 10636 4898
rect 10637 4888 10795 4898
rect 10799 4888 10829 4898
rect 10833 4888 10863 4902
rect 10891 4888 10904 4926
rect 10976 4940 11005 4956
rect 11019 4940 11048 4956
rect 11063 4946 11093 4962
rect 11121 4940 11127 4988
rect 11130 4982 11149 4988
rect 11164 4982 11194 4990
rect 11130 4974 11194 4982
rect 11130 4958 11210 4974
rect 11226 4967 11288 4998
rect 11304 4967 11366 4998
rect 11435 4996 11484 5021
rect 11499 4996 11529 5012
rect 11398 4982 11428 4990
rect 11435 4988 11545 4996
rect 11398 4974 11443 4982
rect 11130 4956 11149 4958
rect 11164 4956 11210 4958
rect 11130 4940 11210 4956
rect 11237 4954 11272 4967
rect 11313 4964 11350 4967
rect 11313 4962 11355 4964
rect 11242 4951 11272 4954
rect 11251 4947 11258 4951
rect 11258 4946 11259 4947
rect 11217 4940 11227 4946
rect 10976 4932 11011 4940
rect 10976 4906 10977 4932
rect 10984 4906 11011 4932
rect 10919 4888 10949 4902
rect 10976 4898 11011 4906
rect 11013 4932 11054 4940
rect 11013 4906 11028 4932
rect 11035 4906 11054 4932
rect 11118 4928 11149 4940
rect 11164 4928 11267 4940
rect 11279 4930 11305 4956
rect 11320 4951 11350 4962
rect 11382 4958 11444 4974
rect 11382 4956 11428 4958
rect 11382 4940 11444 4956
rect 11456 4940 11462 4988
rect 11465 4980 11545 4988
rect 11465 4978 11484 4980
rect 11499 4978 11533 4980
rect 11465 4962 11545 4978
rect 11465 4940 11484 4962
rect 11499 4946 11529 4962
rect 11557 4956 11563 5030
rect 11566 4956 11585 5100
rect 11600 4956 11606 5100
rect 11615 5030 11628 5100
rect 11680 5096 11702 5100
rect 11673 5074 11702 5088
rect 11755 5074 11771 5088
rect 11809 5084 11815 5086
rect 11822 5084 11930 5100
rect 11937 5084 11943 5086
rect 11951 5084 11966 5100
rect 12032 5094 12051 5097
rect 11673 5072 11771 5074
rect 11798 5072 11966 5084
rect 11981 5074 11997 5088
rect 12032 5075 12054 5094
rect 12064 5088 12080 5089
rect 12063 5086 12080 5088
rect 12064 5081 12080 5086
rect 12054 5074 12060 5075
rect 12063 5074 12092 5081
rect 11981 5073 12092 5074
rect 11981 5072 12098 5073
rect 11657 5064 11708 5072
rect 11755 5064 11789 5072
rect 11657 5052 11682 5064
rect 11689 5052 11708 5064
rect 11762 5062 11789 5064
rect 11798 5062 12019 5072
rect 12054 5069 12060 5072
rect 11762 5058 12019 5062
rect 11657 5044 11708 5052
rect 11755 5044 12019 5058
rect 12063 5064 12098 5072
rect 11609 4996 11628 5030
rect 11673 5036 11702 5044
rect 11673 5030 11690 5036
rect 11673 5028 11707 5030
rect 11755 5028 11771 5044
rect 11772 5034 11980 5044
rect 11981 5034 11997 5044
rect 12045 5040 12060 5055
rect 12063 5052 12064 5064
rect 12071 5052 12098 5064
rect 12063 5044 12098 5052
rect 12063 5043 12092 5044
rect 11783 5030 11997 5034
rect 11798 5028 11997 5030
rect 12032 5030 12045 5040
rect 12063 5030 12080 5043
rect 12032 5028 12080 5030
rect 11674 5024 11707 5028
rect 11670 5022 11707 5024
rect 11670 5021 11737 5022
rect 11670 5016 11701 5021
rect 11707 5016 11737 5021
rect 11670 5012 11737 5016
rect 11643 5009 11737 5012
rect 11643 5002 11692 5009
rect 11643 4996 11673 5002
rect 11692 4997 11697 5002
rect 11609 4980 11689 4996
rect 11701 4988 11737 5009
rect 11798 5004 11987 5028
rect 12032 5027 12079 5028
rect 12045 5022 12079 5027
rect 11813 5001 11987 5004
rect 11806 4998 11987 5001
rect 12015 5021 12079 5022
rect 11609 4978 11628 4980
rect 11643 4978 11677 4980
rect 11609 4962 11689 4978
rect 11609 4956 11628 4962
rect 11325 4930 11428 4940
rect 11279 4928 11428 4930
rect 11449 4928 11484 4940
rect 11118 4926 11280 4928
rect 11130 4906 11149 4926
rect 11164 4924 11194 4926
rect 11013 4898 11054 4906
rect 11136 4902 11149 4906
rect 11201 4910 11280 4926
rect 11312 4926 11484 4928
rect 11312 4910 11391 4926
rect 11398 4924 11428 4926
rect 10976 4888 11005 4898
rect 11019 4888 11048 4898
rect 11063 4888 11093 4902
rect 11136 4888 11179 4902
rect 11201 4898 11391 4910
rect 11456 4906 11462 4926
rect 11186 4888 11216 4898
rect 11217 4888 11375 4898
rect 11379 4888 11409 4898
rect 11413 4888 11443 4902
rect 11471 4888 11484 4926
rect 11556 4940 11585 4956
rect 11599 4940 11628 4956
rect 11643 4946 11673 4962
rect 11701 4940 11707 4988
rect 11710 4982 11729 4988
rect 11744 4982 11774 4990
rect 11710 4974 11774 4982
rect 11710 4958 11790 4974
rect 11806 4967 11868 4998
rect 11884 4967 11946 4998
rect 12015 4996 12064 5021
rect 12079 4996 12109 5012
rect 11978 4982 12008 4990
rect 12015 4988 12125 4996
rect 11978 4974 12023 4982
rect 11710 4956 11729 4958
rect 11744 4956 11790 4958
rect 11710 4940 11790 4956
rect 11817 4954 11852 4967
rect 11893 4964 11930 4967
rect 11893 4962 11935 4964
rect 11822 4951 11852 4954
rect 11831 4947 11838 4951
rect 11838 4946 11839 4947
rect 11797 4940 11807 4946
rect 11556 4932 11591 4940
rect 11556 4906 11557 4932
rect 11564 4906 11591 4932
rect 11499 4888 11529 4902
rect 11556 4898 11591 4906
rect 11593 4932 11634 4940
rect 11593 4906 11608 4932
rect 11615 4906 11634 4932
rect 11698 4928 11729 4940
rect 11744 4928 11847 4940
rect 11859 4930 11885 4956
rect 11900 4951 11930 4962
rect 11962 4958 12024 4974
rect 11962 4956 12008 4958
rect 11962 4940 12024 4956
rect 12036 4940 12042 4988
rect 12045 4980 12125 4988
rect 12045 4978 12064 4980
rect 12079 4978 12113 4980
rect 12045 4962 12125 4978
rect 12045 4940 12064 4962
rect 12079 4946 12109 4962
rect 12137 4956 12143 5030
rect 12146 4956 12165 5100
rect 12180 4956 12186 5100
rect 12195 5030 12208 5100
rect 12260 5096 12282 5100
rect 12253 5074 12282 5088
rect 12335 5074 12351 5088
rect 12389 5084 12395 5086
rect 12402 5084 12510 5100
rect 12517 5084 12523 5086
rect 12531 5084 12546 5100
rect 12612 5094 12631 5097
rect 12253 5072 12351 5074
rect 12378 5072 12546 5084
rect 12561 5074 12577 5088
rect 12612 5075 12634 5094
rect 12644 5088 12660 5089
rect 12643 5086 12660 5088
rect 12644 5081 12660 5086
rect 12634 5074 12640 5075
rect 12643 5074 12672 5081
rect 12561 5073 12672 5074
rect 12561 5072 12678 5073
rect 12237 5064 12288 5072
rect 12335 5064 12369 5072
rect 12237 5052 12262 5064
rect 12269 5052 12288 5064
rect 12342 5062 12369 5064
rect 12378 5062 12599 5072
rect 12634 5069 12640 5072
rect 12342 5058 12599 5062
rect 12237 5044 12288 5052
rect 12335 5044 12599 5058
rect 12643 5064 12678 5072
rect 12189 4996 12208 5030
rect 12253 5036 12282 5044
rect 12253 5030 12270 5036
rect 12253 5028 12287 5030
rect 12335 5028 12351 5044
rect 12352 5034 12560 5044
rect 12561 5034 12577 5044
rect 12625 5040 12640 5055
rect 12643 5052 12644 5064
rect 12651 5052 12678 5064
rect 12643 5044 12678 5052
rect 12643 5043 12672 5044
rect 12363 5030 12577 5034
rect 12378 5028 12577 5030
rect 12612 5030 12625 5040
rect 12643 5030 12660 5043
rect 12612 5028 12660 5030
rect 12254 5024 12287 5028
rect 12250 5022 12287 5024
rect 12250 5021 12317 5022
rect 12250 5016 12281 5021
rect 12287 5016 12317 5021
rect 12250 5012 12317 5016
rect 12223 5009 12317 5012
rect 12223 5002 12272 5009
rect 12223 4996 12253 5002
rect 12272 4997 12277 5002
rect 12189 4980 12269 4996
rect 12281 4988 12317 5009
rect 12378 5004 12567 5028
rect 12612 5027 12659 5028
rect 12625 5022 12659 5027
rect 12393 5001 12567 5004
rect 12386 4998 12567 5001
rect 12595 5021 12659 5022
rect 12189 4978 12208 4980
rect 12223 4978 12257 4980
rect 12189 4962 12269 4978
rect 12189 4956 12208 4962
rect 11905 4930 12008 4940
rect 11859 4928 12008 4930
rect 12029 4928 12064 4940
rect 11698 4926 11860 4928
rect 11710 4906 11729 4926
rect 11744 4924 11774 4926
rect 11593 4898 11634 4906
rect 11716 4902 11729 4906
rect 11781 4910 11860 4926
rect 11892 4926 12064 4928
rect 11892 4910 11971 4926
rect 11978 4924 12008 4926
rect 11556 4888 11585 4898
rect 11599 4888 11628 4898
rect 11643 4888 11673 4902
rect 11716 4888 11759 4902
rect 11781 4898 11971 4910
rect 12036 4906 12042 4926
rect 11766 4888 11796 4898
rect 11797 4888 11955 4898
rect 11959 4888 11989 4898
rect 11993 4888 12023 4902
rect 12051 4888 12064 4926
rect 12136 4940 12165 4956
rect 12179 4940 12208 4956
rect 12223 4946 12253 4962
rect 12281 4940 12287 4988
rect 12290 4982 12309 4988
rect 12324 4982 12354 4990
rect 12290 4974 12354 4982
rect 12290 4958 12370 4974
rect 12386 4967 12448 4998
rect 12464 4967 12526 4998
rect 12595 4996 12644 5021
rect 12659 4996 12689 5012
rect 12558 4982 12588 4990
rect 12595 4988 12705 4996
rect 12558 4974 12603 4982
rect 12290 4956 12309 4958
rect 12324 4956 12370 4958
rect 12290 4940 12370 4956
rect 12397 4954 12432 4967
rect 12473 4964 12510 4967
rect 12473 4962 12515 4964
rect 12402 4951 12432 4954
rect 12411 4947 12418 4951
rect 12418 4946 12419 4947
rect 12377 4940 12387 4946
rect 12136 4932 12171 4940
rect 12136 4906 12137 4932
rect 12144 4906 12171 4932
rect 12079 4888 12109 4902
rect 12136 4898 12171 4906
rect 12173 4932 12214 4940
rect 12173 4906 12188 4932
rect 12195 4906 12214 4932
rect 12278 4928 12309 4940
rect 12324 4928 12427 4940
rect 12439 4930 12465 4956
rect 12480 4951 12510 4962
rect 12542 4958 12604 4974
rect 12542 4956 12588 4958
rect 12542 4940 12604 4956
rect 12616 4940 12622 4988
rect 12625 4980 12705 4988
rect 12625 4978 12644 4980
rect 12659 4978 12693 4980
rect 12625 4962 12705 4978
rect 12625 4940 12644 4962
rect 12659 4946 12689 4962
rect 12717 4956 12723 5030
rect 12726 4956 12745 5100
rect 12760 4956 12766 5100
rect 12775 5030 12788 5100
rect 12840 5096 12862 5100
rect 12833 5074 12862 5088
rect 12915 5074 12931 5088
rect 12969 5084 12975 5086
rect 12982 5084 13090 5100
rect 13097 5084 13103 5086
rect 13111 5084 13126 5100
rect 13192 5094 13211 5097
rect 12833 5072 12931 5074
rect 12958 5072 13126 5084
rect 13141 5074 13157 5088
rect 13192 5075 13214 5094
rect 13224 5088 13240 5089
rect 13223 5086 13240 5088
rect 13224 5081 13240 5086
rect 13214 5074 13220 5075
rect 13223 5074 13252 5081
rect 13141 5073 13252 5074
rect 13141 5072 13258 5073
rect 12817 5064 12868 5072
rect 12915 5064 12949 5072
rect 12817 5052 12842 5064
rect 12849 5052 12868 5064
rect 12922 5062 12949 5064
rect 12958 5062 13179 5072
rect 13214 5069 13220 5072
rect 12922 5058 13179 5062
rect 12817 5044 12868 5052
rect 12915 5044 13179 5058
rect 13223 5064 13258 5072
rect 12769 4996 12788 5030
rect 12833 5036 12862 5044
rect 12833 5030 12850 5036
rect 12833 5028 12867 5030
rect 12915 5028 12931 5044
rect 12932 5034 13140 5044
rect 13141 5034 13157 5044
rect 13205 5040 13220 5055
rect 13223 5052 13224 5064
rect 13231 5052 13258 5064
rect 13223 5044 13258 5052
rect 13223 5043 13252 5044
rect 12943 5030 13157 5034
rect 12958 5028 13157 5030
rect 13192 5030 13205 5040
rect 13223 5030 13240 5043
rect 13192 5028 13240 5030
rect 12834 5024 12867 5028
rect 12830 5022 12867 5024
rect 12830 5021 12897 5022
rect 12830 5016 12861 5021
rect 12867 5016 12897 5021
rect 12830 5012 12897 5016
rect 12803 5009 12897 5012
rect 12803 5002 12852 5009
rect 12803 4996 12833 5002
rect 12852 4997 12857 5002
rect 12769 4980 12849 4996
rect 12861 4988 12897 5009
rect 12958 5004 13147 5028
rect 13192 5027 13239 5028
rect 13205 5022 13239 5027
rect 12973 5001 13147 5004
rect 12966 4998 13147 5001
rect 13175 5021 13239 5022
rect 12769 4978 12788 4980
rect 12803 4978 12837 4980
rect 12769 4962 12849 4978
rect 12769 4956 12788 4962
rect 12485 4930 12588 4940
rect 12439 4928 12588 4930
rect 12609 4928 12644 4940
rect 12278 4926 12440 4928
rect 12290 4906 12309 4926
rect 12324 4924 12354 4926
rect 12173 4898 12214 4906
rect 12296 4902 12309 4906
rect 12361 4910 12440 4926
rect 12472 4926 12644 4928
rect 12472 4910 12551 4926
rect 12558 4924 12588 4926
rect 12136 4888 12165 4898
rect 12179 4888 12208 4898
rect 12223 4888 12253 4902
rect 12296 4888 12339 4902
rect 12361 4898 12551 4910
rect 12616 4906 12622 4926
rect 12346 4888 12376 4898
rect 12377 4888 12535 4898
rect 12539 4888 12569 4898
rect 12573 4888 12603 4902
rect 12631 4888 12644 4926
rect 12716 4940 12745 4956
rect 12759 4940 12788 4956
rect 12803 4946 12833 4962
rect 12861 4940 12867 4988
rect 12870 4982 12889 4988
rect 12904 4982 12934 4990
rect 12870 4974 12934 4982
rect 12870 4958 12950 4974
rect 12966 4967 13028 4998
rect 13044 4967 13106 4998
rect 13175 4996 13224 5021
rect 13239 4996 13269 5012
rect 13138 4982 13168 4990
rect 13175 4988 13285 4996
rect 13138 4974 13183 4982
rect 12870 4956 12889 4958
rect 12904 4956 12950 4958
rect 12870 4940 12950 4956
rect 12977 4954 13012 4967
rect 13053 4964 13090 4967
rect 13053 4962 13095 4964
rect 12982 4951 13012 4954
rect 12991 4947 12998 4951
rect 12998 4946 12999 4947
rect 12957 4940 12967 4946
rect 12716 4932 12751 4940
rect 12716 4906 12717 4932
rect 12724 4906 12751 4932
rect 12659 4888 12689 4902
rect 12716 4898 12751 4906
rect 12753 4932 12794 4940
rect 12753 4906 12768 4932
rect 12775 4906 12794 4932
rect 12858 4928 12889 4940
rect 12904 4928 13007 4940
rect 13019 4930 13045 4956
rect 13060 4951 13090 4962
rect 13122 4958 13184 4974
rect 13122 4956 13168 4958
rect 13122 4940 13184 4956
rect 13196 4940 13202 4988
rect 13205 4980 13285 4988
rect 13205 4978 13224 4980
rect 13239 4978 13273 4980
rect 13205 4962 13285 4978
rect 13205 4940 13224 4962
rect 13239 4946 13269 4962
rect 13297 4956 13303 5030
rect 13306 4956 13325 5100
rect 13340 4956 13346 5100
rect 13355 5030 13368 5100
rect 13420 5096 13442 5100
rect 13413 5074 13442 5088
rect 13495 5074 13511 5088
rect 13549 5084 13555 5086
rect 13562 5084 13670 5100
rect 13677 5084 13683 5086
rect 13691 5084 13706 5100
rect 13772 5094 13791 5097
rect 13413 5072 13511 5074
rect 13538 5072 13706 5084
rect 13721 5074 13737 5088
rect 13772 5075 13794 5094
rect 13804 5088 13820 5089
rect 13803 5086 13820 5088
rect 13804 5081 13820 5086
rect 13794 5074 13800 5075
rect 13803 5074 13832 5081
rect 13721 5073 13832 5074
rect 13721 5072 13838 5073
rect 13397 5064 13448 5072
rect 13495 5064 13529 5072
rect 13397 5052 13422 5064
rect 13429 5052 13448 5064
rect 13502 5062 13529 5064
rect 13538 5062 13759 5072
rect 13794 5069 13800 5072
rect 13502 5058 13759 5062
rect 13397 5044 13448 5052
rect 13495 5044 13759 5058
rect 13803 5064 13838 5072
rect 13349 4996 13368 5030
rect 13413 5036 13442 5044
rect 13413 5030 13430 5036
rect 13413 5028 13447 5030
rect 13495 5028 13511 5044
rect 13512 5034 13720 5044
rect 13721 5034 13737 5044
rect 13785 5040 13800 5055
rect 13803 5052 13804 5064
rect 13811 5052 13838 5064
rect 13803 5044 13838 5052
rect 13803 5043 13832 5044
rect 13523 5030 13737 5034
rect 13538 5028 13737 5030
rect 13772 5030 13785 5040
rect 13803 5030 13820 5043
rect 13772 5028 13820 5030
rect 13414 5024 13447 5028
rect 13410 5022 13447 5024
rect 13410 5021 13477 5022
rect 13410 5016 13441 5021
rect 13447 5016 13477 5021
rect 13410 5012 13477 5016
rect 13383 5009 13477 5012
rect 13383 5002 13432 5009
rect 13383 4996 13413 5002
rect 13432 4997 13437 5002
rect 13349 4980 13429 4996
rect 13441 4988 13477 5009
rect 13538 5004 13727 5028
rect 13772 5027 13819 5028
rect 13785 5022 13819 5027
rect 13553 5001 13727 5004
rect 13546 4998 13727 5001
rect 13755 5021 13819 5022
rect 13349 4978 13368 4980
rect 13383 4978 13417 4980
rect 13349 4962 13429 4978
rect 13349 4956 13368 4962
rect 13065 4930 13168 4940
rect 13019 4928 13168 4930
rect 13189 4928 13224 4940
rect 12858 4926 13020 4928
rect 12870 4906 12889 4926
rect 12904 4924 12934 4926
rect 12753 4898 12794 4906
rect 12876 4902 12889 4906
rect 12941 4910 13020 4926
rect 13052 4926 13224 4928
rect 13052 4910 13131 4926
rect 13138 4924 13168 4926
rect 12716 4888 12745 4898
rect 12759 4888 12788 4898
rect 12803 4888 12833 4902
rect 12876 4888 12919 4902
rect 12941 4898 13131 4910
rect 13196 4906 13202 4926
rect 12926 4888 12956 4898
rect 12957 4888 13115 4898
rect 13119 4888 13149 4898
rect 13153 4888 13183 4902
rect 13211 4888 13224 4926
rect 13296 4940 13325 4956
rect 13339 4940 13368 4956
rect 13383 4946 13413 4962
rect 13441 4940 13447 4988
rect 13450 4982 13469 4988
rect 13484 4982 13514 4990
rect 13450 4974 13514 4982
rect 13450 4958 13530 4974
rect 13546 4967 13608 4998
rect 13624 4967 13686 4998
rect 13755 4996 13804 5021
rect 13819 4996 13849 5012
rect 13718 4982 13748 4990
rect 13755 4988 13865 4996
rect 13718 4974 13763 4982
rect 13450 4956 13469 4958
rect 13484 4956 13530 4958
rect 13450 4940 13530 4956
rect 13557 4954 13592 4967
rect 13633 4964 13670 4967
rect 13633 4962 13675 4964
rect 13562 4951 13592 4954
rect 13571 4947 13578 4951
rect 13578 4946 13579 4947
rect 13537 4940 13547 4946
rect 13296 4932 13331 4940
rect 13296 4906 13297 4932
rect 13304 4906 13331 4932
rect 13239 4888 13269 4902
rect 13296 4898 13331 4906
rect 13333 4932 13374 4940
rect 13333 4906 13348 4932
rect 13355 4906 13374 4932
rect 13438 4928 13469 4940
rect 13484 4928 13587 4940
rect 13599 4930 13625 4956
rect 13640 4951 13670 4962
rect 13702 4958 13764 4974
rect 13702 4956 13748 4958
rect 13702 4940 13764 4956
rect 13776 4940 13782 4988
rect 13785 4980 13865 4988
rect 13785 4978 13804 4980
rect 13819 4978 13853 4980
rect 13785 4962 13865 4978
rect 13785 4940 13804 4962
rect 13819 4946 13849 4962
rect 13877 4956 13883 5030
rect 13886 4956 13905 5100
rect 13920 4956 13926 5100
rect 13935 5030 13948 5100
rect 14000 5096 14022 5100
rect 13993 5074 14022 5088
rect 14075 5074 14091 5088
rect 14129 5084 14135 5086
rect 14142 5084 14250 5100
rect 14257 5084 14263 5086
rect 14271 5084 14286 5100
rect 14352 5094 14371 5097
rect 13993 5072 14091 5074
rect 14118 5072 14286 5084
rect 14301 5074 14317 5088
rect 14352 5075 14374 5094
rect 14384 5088 14400 5089
rect 14383 5086 14400 5088
rect 14384 5081 14400 5086
rect 14374 5074 14380 5075
rect 14383 5074 14412 5081
rect 14301 5073 14412 5074
rect 14301 5072 14418 5073
rect 13977 5064 14028 5072
rect 14075 5064 14109 5072
rect 13977 5052 14002 5064
rect 14009 5052 14028 5064
rect 14082 5062 14109 5064
rect 14118 5062 14339 5072
rect 14374 5069 14380 5072
rect 14082 5058 14339 5062
rect 13977 5044 14028 5052
rect 14075 5044 14339 5058
rect 14383 5064 14418 5072
rect 13929 4996 13948 5030
rect 13993 5036 14022 5044
rect 13993 5030 14010 5036
rect 13993 5028 14027 5030
rect 14075 5028 14091 5044
rect 14092 5034 14300 5044
rect 14301 5034 14317 5044
rect 14365 5040 14380 5055
rect 14383 5052 14384 5064
rect 14391 5052 14418 5064
rect 14383 5044 14418 5052
rect 14383 5043 14412 5044
rect 14103 5030 14317 5034
rect 14118 5028 14317 5030
rect 14352 5030 14365 5040
rect 14383 5030 14400 5043
rect 14352 5028 14400 5030
rect 13994 5024 14027 5028
rect 13990 5022 14027 5024
rect 13990 5021 14057 5022
rect 13990 5016 14021 5021
rect 14027 5016 14057 5021
rect 13990 5012 14057 5016
rect 13963 5009 14057 5012
rect 13963 5002 14012 5009
rect 13963 4996 13993 5002
rect 14012 4997 14017 5002
rect 13929 4980 14009 4996
rect 14021 4988 14057 5009
rect 14118 5004 14307 5028
rect 14352 5027 14399 5028
rect 14365 5022 14399 5027
rect 14133 5001 14307 5004
rect 14126 4998 14307 5001
rect 14335 5021 14399 5022
rect 13929 4978 13948 4980
rect 13963 4978 13997 4980
rect 13929 4962 14009 4978
rect 13929 4956 13948 4962
rect 13645 4930 13748 4940
rect 13599 4928 13748 4930
rect 13769 4928 13804 4940
rect 13438 4926 13600 4928
rect 13450 4906 13469 4926
rect 13484 4924 13514 4926
rect 13333 4898 13374 4906
rect 13456 4902 13469 4906
rect 13521 4910 13600 4926
rect 13632 4926 13804 4928
rect 13632 4910 13711 4926
rect 13718 4924 13748 4926
rect 13296 4888 13325 4898
rect 13339 4888 13368 4898
rect 13383 4888 13413 4902
rect 13456 4888 13499 4902
rect 13521 4898 13711 4910
rect 13776 4906 13782 4926
rect 13506 4888 13536 4898
rect 13537 4888 13695 4898
rect 13699 4888 13729 4898
rect 13733 4888 13763 4902
rect 13791 4888 13804 4926
rect 13876 4940 13905 4956
rect 13919 4940 13948 4956
rect 13963 4946 13993 4962
rect 14021 4940 14027 4988
rect 14030 4982 14049 4988
rect 14064 4982 14094 4990
rect 14030 4974 14094 4982
rect 14030 4958 14110 4974
rect 14126 4967 14188 4998
rect 14204 4967 14266 4998
rect 14335 4996 14384 5021
rect 14399 4996 14429 5012
rect 14298 4982 14328 4990
rect 14335 4988 14445 4996
rect 14298 4974 14343 4982
rect 14030 4956 14049 4958
rect 14064 4956 14110 4958
rect 14030 4940 14110 4956
rect 14137 4954 14172 4967
rect 14213 4964 14250 4967
rect 14213 4962 14255 4964
rect 14142 4951 14172 4954
rect 14151 4947 14158 4951
rect 14158 4946 14159 4947
rect 14117 4940 14127 4946
rect 13876 4932 13911 4940
rect 13876 4906 13877 4932
rect 13884 4906 13911 4932
rect 13819 4888 13849 4902
rect 13876 4898 13911 4906
rect 13913 4932 13954 4940
rect 13913 4906 13928 4932
rect 13935 4906 13954 4932
rect 14018 4928 14049 4940
rect 14064 4928 14167 4940
rect 14179 4930 14205 4956
rect 14220 4951 14250 4962
rect 14282 4958 14344 4974
rect 14282 4956 14328 4958
rect 14282 4940 14344 4956
rect 14356 4940 14362 4988
rect 14365 4980 14445 4988
rect 14365 4978 14384 4980
rect 14399 4978 14433 4980
rect 14365 4962 14445 4978
rect 14365 4940 14384 4962
rect 14399 4946 14429 4962
rect 14457 4956 14463 5030
rect 14466 4956 14485 5100
rect 14500 4956 14506 5100
rect 14515 5030 14528 5100
rect 14580 5096 14602 5100
rect 14573 5074 14602 5088
rect 14655 5074 14671 5088
rect 14709 5084 14715 5086
rect 14722 5084 14830 5100
rect 14837 5084 14843 5086
rect 14851 5084 14866 5100
rect 14932 5094 14951 5097
rect 14573 5072 14671 5074
rect 14698 5072 14866 5084
rect 14881 5074 14897 5088
rect 14932 5075 14954 5094
rect 14964 5088 14980 5089
rect 14963 5086 14980 5088
rect 14964 5081 14980 5086
rect 14954 5074 14960 5075
rect 14963 5074 14992 5081
rect 14881 5073 14992 5074
rect 14881 5072 14998 5073
rect 14557 5064 14608 5072
rect 14655 5064 14689 5072
rect 14557 5052 14582 5064
rect 14589 5052 14608 5064
rect 14662 5062 14689 5064
rect 14698 5062 14919 5072
rect 14954 5069 14960 5072
rect 14662 5058 14919 5062
rect 14557 5044 14608 5052
rect 14655 5044 14919 5058
rect 14963 5064 14998 5072
rect 14509 4996 14528 5030
rect 14573 5036 14602 5044
rect 14573 5030 14590 5036
rect 14573 5028 14607 5030
rect 14655 5028 14671 5044
rect 14672 5034 14880 5044
rect 14881 5034 14897 5044
rect 14945 5040 14960 5055
rect 14963 5052 14964 5064
rect 14971 5052 14998 5064
rect 14963 5044 14998 5052
rect 14963 5043 14992 5044
rect 14683 5030 14897 5034
rect 14698 5028 14897 5030
rect 14932 5030 14945 5040
rect 14963 5030 14980 5043
rect 14932 5028 14980 5030
rect 14574 5024 14607 5028
rect 14570 5022 14607 5024
rect 14570 5021 14637 5022
rect 14570 5016 14601 5021
rect 14607 5016 14637 5021
rect 14570 5012 14637 5016
rect 14543 5009 14637 5012
rect 14543 5002 14592 5009
rect 14543 4996 14573 5002
rect 14592 4997 14597 5002
rect 14509 4980 14589 4996
rect 14601 4988 14637 5009
rect 14698 5004 14887 5028
rect 14932 5027 14979 5028
rect 14945 5022 14979 5027
rect 14713 5001 14887 5004
rect 14706 4998 14887 5001
rect 14915 5021 14979 5022
rect 14509 4978 14528 4980
rect 14543 4978 14577 4980
rect 14509 4962 14589 4978
rect 14509 4956 14528 4962
rect 14225 4930 14328 4940
rect 14179 4928 14328 4930
rect 14349 4928 14384 4940
rect 14018 4926 14180 4928
rect 14030 4906 14049 4926
rect 14064 4924 14094 4926
rect 13913 4898 13954 4906
rect 14036 4902 14049 4906
rect 14101 4910 14180 4926
rect 14212 4926 14384 4928
rect 14212 4910 14291 4926
rect 14298 4924 14328 4926
rect 13876 4888 13905 4898
rect 13919 4888 13948 4898
rect 13963 4888 13993 4902
rect 14036 4888 14079 4902
rect 14101 4898 14291 4910
rect 14356 4906 14362 4926
rect 14086 4888 14116 4898
rect 14117 4888 14275 4898
rect 14279 4888 14309 4898
rect 14313 4888 14343 4902
rect 14371 4888 14384 4926
rect 14456 4940 14485 4956
rect 14499 4940 14528 4956
rect 14543 4946 14573 4962
rect 14601 4940 14607 4988
rect 14610 4982 14629 4988
rect 14644 4982 14674 4990
rect 14610 4974 14674 4982
rect 14610 4958 14690 4974
rect 14706 4967 14768 4998
rect 14784 4967 14846 4998
rect 14915 4996 14964 5021
rect 14979 4996 15009 5012
rect 14878 4982 14908 4990
rect 14915 4988 15025 4996
rect 14878 4974 14923 4982
rect 14610 4956 14629 4958
rect 14644 4956 14690 4958
rect 14610 4940 14690 4956
rect 14717 4954 14752 4967
rect 14793 4964 14830 4967
rect 14793 4962 14835 4964
rect 14722 4951 14752 4954
rect 14731 4947 14738 4951
rect 14738 4946 14739 4947
rect 14697 4940 14707 4946
rect 14456 4932 14491 4940
rect 14456 4906 14457 4932
rect 14464 4906 14491 4932
rect 14399 4888 14429 4902
rect 14456 4898 14491 4906
rect 14493 4932 14534 4940
rect 14493 4906 14508 4932
rect 14515 4906 14534 4932
rect 14598 4928 14629 4940
rect 14644 4928 14747 4940
rect 14759 4930 14785 4956
rect 14800 4951 14830 4962
rect 14862 4958 14924 4974
rect 14862 4956 14908 4958
rect 14862 4940 14924 4956
rect 14936 4940 14942 4988
rect 14945 4980 15025 4988
rect 14945 4978 14964 4980
rect 14979 4978 15013 4980
rect 14945 4962 15025 4978
rect 14945 4940 14964 4962
rect 14979 4946 15009 4962
rect 15037 4956 15043 5030
rect 15046 4956 15065 5100
rect 15080 4956 15086 5100
rect 15095 5030 15108 5100
rect 15160 5096 15182 5100
rect 15153 5074 15182 5088
rect 15235 5074 15251 5088
rect 15289 5084 15295 5086
rect 15302 5084 15410 5100
rect 15417 5084 15423 5086
rect 15431 5084 15446 5100
rect 15512 5094 15531 5097
rect 15153 5072 15251 5074
rect 15278 5072 15446 5084
rect 15461 5074 15477 5088
rect 15512 5075 15534 5094
rect 15544 5088 15560 5089
rect 15543 5086 15560 5088
rect 15544 5081 15560 5086
rect 15534 5074 15540 5075
rect 15543 5074 15572 5081
rect 15461 5073 15572 5074
rect 15461 5072 15578 5073
rect 15137 5064 15188 5072
rect 15235 5064 15269 5072
rect 15137 5052 15162 5064
rect 15169 5052 15188 5064
rect 15242 5062 15269 5064
rect 15278 5062 15499 5072
rect 15534 5069 15540 5072
rect 15242 5058 15499 5062
rect 15137 5044 15188 5052
rect 15235 5044 15499 5058
rect 15543 5064 15578 5072
rect 15089 4996 15108 5030
rect 15153 5036 15182 5044
rect 15153 5030 15170 5036
rect 15153 5028 15187 5030
rect 15235 5028 15251 5044
rect 15252 5034 15460 5044
rect 15461 5034 15477 5044
rect 15525 5040 15540 5055
rect 15543 5052 15544 5064
rect 15551 5052 15578 5064
rect 15543 5044 15578 5052
rect 15543 5043 15572 5044
rect 15263 5030 15477 5034
rect 15278 5028 15477 5030
rect 15512 5030 15525 5040
rect 15543 5030 15560 5043
rect 15512 5028 15560 5030
rect 15154 5024 15187 5028
rect 15150 5022 15187 5024
rect 15150 5021 15217 5022
rect 15150 5016 15181 5021
rect 15187 5016 15217 5021
rect 15150 5012 15217 5016
rect 15123 5009 15217 5012
rect 15123 5002 15172 5009
rect 15123 4996 15153 5002
rect 15172 4997 15177 5002
rect 15089 4980 15169 4996
rect 15181 4988 15217 5009
rect 15278 5004 15467 5028
rect 15512 5027 15559 5028
rect 15525 5022 15559 5027
rect 15293 5001 15467 5004
rect 15286 4998 15467 5001
rect 15495 5021 15559 5022
rect 15089 4978 15108 4980
rect 15123 4978 15157 4980
rect 15089 4962 15169 4978
rect 15089 4956 15108 4962
rect 14805 4930 14908 4940
rect 14759 4928 14908 4930
rect 14929 4928 14964 4940
rect 14598 4926 14760 4928
rect 14610 4906 14629 4926
rect 14644 4924 14674 4926
rect 14493 4898 14534 4906
rect 14616 4902 14629 4906
rect 14681 4910 14760 4926
rect 14792 4926 14964 4928
rect 14792 4910 14871 4926
rect 14878 4924 14908 4926
rect 14456 4888 14485 4898
rect 14499 4888 14528 4898
rect 14543 4888 14573 4902
rect 14616 4888 14659 4902
rect 14681 4898 14871 4910
rect 14936 4906 14942 4926
rect 14666 4888 14696 4898
rect 14697 4888 14855 4898
rect 14859 4888 14889 4898
rect 14893 4888 14923 4902
rect 14951 4888 14964 4926
rect 15036 4940 15065 4956
rect 15079 4940 15108 4956
rect 15123 4946 15153 4962
rect 15181 4940 15187 4988
rect 15190 4982 15209 4988
rect 15224 4982 15254 4990
rect 15190 4974 15254 4982
rect 15190 4958 15270 4974
rect 15286 4967 15348 4998
rect 15364 4967 15426 4998
rect 15495 4996 15544 5021
rect 15559 4996 15589 5012
rect 15458 4982 15488 4990
rect 15495 4988 15605 4996
rect 15458 4974 15503 4982
rect 15190 4956 15209 4958
rect 15224 4956 15270 4958
rect 15190 4940 15270 4956
rect 15297 4954 15332 4967
rect 15373 4964 15410 4967
rect 15373 4962 15415 4964
rect 15302 4951 15332 4954
rect 15311 4947 15318 4951
rect 15318 4946 15319 4947
rect 15277 4940 15287 4946
rect 15036 4932 15071 4940
rect 15036 4906 15037 4932
rect 15044 4906 15071 4932
rect 14979 4888 15009 4902
rect 15036 4898 15071 4906
rect 15073 4932 15114 4940
rect 15073 4906 15088 4932
rect 15095 4906 15114 4932
rect 15178 4928 15209 4940
rect 15224 4928 15327 4940
rect 15339 4930 15365 4956
rect 15380 4951 15410 4962
rect 15442 4958 15504 4974
rect 15442 4956 15488 4958
rect 15442 4940 15504 4956
rect 15516 4940 15522 4988
rect 15525 4980 15605 4988
rect 15525 4978 15544 4980
rect 15559 4978 15593 4980
rect 15525 4962 15605 4978
rect 15525 4940 15544 4962
rect 15559 4946 15589 4962
rect 15617 4956 15623 5030
rect 15626 4956 15645 5100
rect 15660 4956 15666 5100
rect 15675 5030 15688 5100
rect 15740 5096 15762 5100
rect 15733 5074 15762 5088
rect 15815 5074 15831 5088
rect 15869 5084 15875 5086
rect 15882 5084 15990 5100
rect 15997 5084 16003 5086
rect 16011 5084 16026 5100
rect 16092 5094 16111 5097
rect 15733 5072 15831 5074
rect 15858 5072 16026 5084
rect 16041 5074 16057 5088
rect 16092 5075 16114 5094
rect 16124 5088 16140 5089
rect 16123 5086 16140 5088
rect 16124 5081 16140 5086
rect 16114 5074 16120 5075
rect 16123 5074 16152 5081
rect 16041 5073 16152 5074
rect 16041 5072 16158 5073
rect 15717 5064 15768 5072
rect 15815 5064 15849 5072
rect 15717 5052 15742 5064
rect 15749 5052 15768 5064
rect 15822 5062 15849 5064
rect 15858 5062 16079 5072
rect 16114 5069 16120 5072
rect 15822 5058 16079 5062
rect 15717 5044 15768 5052
rect 15815 5044 16079 5058
rect 16123 5064 16158 5072
rect 15669 4996 15688 5030
rect 15733 5036 15762 5044
rect 15733 5030 15750 5036
rect 15733 5028 15767 5030
rect 15815 5028 15831 5044
rect 15832 5034 16040 5044
rect 16041 5034 16057 5044
rect 16105 5040 16120 5055
rect 16123 5052 16124 5064
rect 16131 5052 16158 5064
rect 16123 5044 16158 5052
rect 16123 5043 16152 5044
rect 15843 5030 16057 5034
rect 15858 5028 16057 5030
rect 16092 5030 16105 5040
rect 16123 5030 16140 5043
rect 16092 5028 16140 5030
rect 15734 5024 15767 5028
rect 15730 5022 15767 5024
rect 15730 5021 15797 5022
rect 15730 5016 15761 5021
rect 15767 5016 15797 5021
rect 15730 5012 15797 5016
rect 15703 5009 15797 5012
rect 15703 5002 15752 5009
rect 15703 4996 15733 5002
rect 15752 4997 15757 5002
rect 15669 4980 15749 4996
rect 15761 4988 15797 5009
rect 15858 5004 16047 5028
rect 16092 5027 16139 5028
rect 16105 5022 16139 5027
rect 15873 5001 16047 5004
rect 15866 4998 16047 5001
rect 16075 5021 16139 5022
rect 15669 4978 15688 4980
rect 15703 4978 15737 4980
rect 15669 4962 15749 4978
rect 15669 4956 15688 4962
rect 15385 4930 15488 4940
rect 15339 4928 15488 4930
rect 15509 4928 15544 4940
rect 15178 4926 15340 4928
rect 15190 4906 15209 4926
rect 15224 4924 15254 4926
rect 15073 4898 15114 4906
rect 15196 4902 15209 4906
rect 15261 4910 15340 4926
rect 15372 4926 15544 4928
rect 15372 4910 15451 4926
rect 15458 4924 15488 4926
rect 15036 4888 15065 4898
rect 15079 4888 15108 4898
rect 15123 4888 15153 4902
rect 15196 4888 15239 4902
rect 15261 4898 15451 4910
rect 15516 4906 15522 4926
rect 15246 4888 15276 4898
rect 15277 4888 15435 4898
rect 15439 4888 15469 4898
rect 15473 4888 15503 4902
rect 15531 4888 15544 4926
rect 15616 4940 15645 4956
rect 15659 4940 15688 4956
rect 15703 4946 15733 4962
rect 15761 4940 15767 4988
rect 15770 4982 15789 4988
rect 15804 4982 15834 4990
rect 15770 4974 15834 4982
rect 15770 4958 15850 4974
rect 15866 4967 15928 4998
rect 15944 4967 16006 4998
rect 16075 4996 16124 5021
rect 16139 4996 16169 5012
rect 16038 4982 16068 4990
rect 16075 4988 16185 4996
rect 16038 4974 16083 4982
rect 15770 4956 15789 4958
rect 15804 4956 15850 4958
rect 15770 4940 15850 4956
rect 15877 4954 15912 4967
rect 15953 4964 15990 4967
rect 15953 4962 15995 4964
rect 15882 4951 15912 4954
rect 15891 4947 15898 4951
rect 15898 4946 15899 4947
rect 15857 4940 15867 4946
rect 15616 4932 15651 4940
rect 15616 4906 15617 4932
rect 15624 4906 15651 4932
rect 15559 4888 15589 4902
rect 15616 4898 15651 4906
rect 15653 4932 15694 4940
rect 15653 4906 15668 4932
rect 15675 4906 15694 4932
rect 15758 4928 15789 4940
rect 15804 4928 15907 4940
rect 15919 4930 15945 4956
rect 15960 4951 15990 4962
rect 16022 4958 16084 4974
rect 16022 4956 16068 4958
rect 16022 4940 16084 4956
rect 16096 4940 16102 4988
rect 16105 4980 16185 4988
rect 16105 4978 16124 4980
rect 16139 4978 16173 4980
rect 16105 4962 16185 4978
rect 16105 4940 16124 4962
rect 16139 4946 16169 4962
rect 16197 4956 16203 5030
rect 16206 4956 16225 5100
rect 16240 4956 16246 5100
rect 16255 5030 16268 5100
rect 16320 5096 16342 5100
rect 16313 5074 16342 5088
rect 16395 5074 16411 5088
rect 16449 5084 16455 5086
rect 16462 5084 16570 5100
rect 16577 5084 16583 5086
rect 16591 5084 16606 5100
rect 16672 5094 16691 5097
rect 16313 5072 16411 5074
rect 16438 5072 16606 5084
rect 16621 5074 16637 5088
rect 16672 5075 16694 5094
rect 16704 5088 16720 5089
rect 16703 5086 16720 5088
rect 16704 5081 16720 5086
rect 16694 5074 16700 5075
rect 16703 5074 16732 5081
rect 16621 5073 16732 5074
rect 16621 5072 16738 5073
rect 16297 5064 16348 5072
rect 16395 5064 16429 5072
rect 16297 5052 16322 5064
rect 16329 5052 16348 5064
rect 16402 5062 16429 5064
rect 16438 5062 16659 5072
rect 16694 5069 16700 5072
rect 16402 5058 16659 5062
rect 16297 5044 16348 5052
rect 16395 5044 16659 5058
rect 16703 5064 16738 5072
rect 16249 4996 16268 5030
rect 16313 5036 16342 5044
rect 16313 5030 16330 5036
rect 16313 5028 16347 5030
rect 16395 5028 16411 5044
rect 16412 5034 16620 5044
rect 16621 5034 16637 5044
rect 16685 5040 16700 5055
rect 16703 5052 16704 5064
rect 16711 5052 16738 5064
rect 16703 5044 16738 5052
rect 16703 5043 16732 5044
rect 16423 5030 16637 5034
rect 16438 5028 16637 5030
rect 16672 5030 16685 5040
rect 16703 5030 16720 5043
rect 16672 5028 16720 5030
rect 16314 5024 16347 5028
rect 16310 5022 16347 5024
rect 16310 5021 16377 5022
rect 16310 5016 16341 5021
rect 16347 5016 16377 5021
rect 16310 5012 16377 5016
rect 16283 5009 16377 5012
rect 16283 5002 16332 5009
rect 16283 4996 16313 5002
rect 16332 4997 16337 5002
rect 16249 4980 16329 4996
rect 16341 4988 16377 5009
rect 16438 5004 16627 5028
rect 16672 5027 16719 5028
rect 16685 5022 16719 5027
rect 16453 5001 16627 5004
rect 16446 4998 16627 5001
rect 16655 5021 16719 5022
rect 16249 4978 16268 4980
rect 16283 4978 16317 4980
rect 16249 4962 16329 4978
rect 16249 4956 16268 4962
rect 15965 4930 16068 4940
rect 15919 4928 16068 4930
rect 16089 4928 16124 4940
rect 15758 4926 15920 4928
rect 15770 4906 15789 4926
rect 15804 4924 15834 4926
rect 15653 4898 15694 4906
rect 15776 4902 15789 4906
rect 15841 4910 15920 4926
rect 15952 4926 16124 4928
rect 15952 4910 16031 4926
rect 16038 4924 16068 4926
rect 15616 4888 15645 4898
rect 15659 4888 15688 4898
rect 15703 4888 15733 4902
rect 15776 4888 15819 4902
rect 15841 4898 16031 4910
rect 16096 4906 16102 4926
rect 15826 4888 15856 4898
rect 15857 4888 16015 4898
rect 16019 4888 16049 4898
rect 16053 4888 16083 4902
rect 16111 4888 16124 4926
rect 16196 4940 16225 4956
rect 16239 4940 16268 4956
rect 16283 4946 16313 4962
rect 16341 4940 16347 4988
rect 16350 4982 16369 4988
rect 16384 4982 16414 4990
rect 16350 4974 16414 4982
rect 16350 4958 16430 4974
rect 16446 4967 16508 4998
rect 16524 4967 16586 4998
rect 16655 4996 16704 5021
rect 16719 4996 16749 5012
rect 16618 4982 16648 4990
rect 16655 4988 16765 4996
rect 16618 4974 16663 4982
rect 16350 4956 16369 4958
rect 16384 4956 16430 4958
rect 16350 4940 16430 4956
rect 16457 4954 16492 4967
rect 16533 4964 16570 4967
rect 16533 4962 16575 4964
rect 16462 4951 16492 4954
rect 16471 4947 16478 4951
rect 16478 4946 16479 4947
rect 16437 4940 16447 4946
rect 16196 4932 16231 4940
rect 16196 4906 16197 4932
rect 16204 4906 16231 4932
rect 16139 4888 16169 4902
rect 16196 4898 16231 4906
rect 16233 4932 16274 4940
rect 16233 4906 16248 4932
rect 16255 4906 16274 4932
rect 16338 4928 16369 4940
rect 16384 4928 16487 4940
rect 16499 4930 16525 4956
rect 16540 4951 16570 4962
rect 16602 4958 16664 4974
rect 16602 4956 16648 4958
rect 16602 4940 16664 4956
rect 16676 4940 16682 4988
rect 16685 4980 16765 4988
rect 16685 4978 16704 4980
rect 16719 4978 16753 4980
rect 16685 4962 16765 4978
rect 16685 4940 16704 4962
rect 16719 4946 16749 4962
rect 16777 4956 16783 5030
rect 16786 4956 16805 5100
rect 16820 4956 16826 5100
rect 16835 5030 16848 5100
rect 16900 5096 16922 5100
rect 16893 5074 16922 5088
rect 16975 5074 16991 5088
rect 17029 5084 17035 5086
rect 17042 5084 17150 5100
rect 17157 5084 17163 5086
rect 17171 5084 17186 5100
rect 17252 5094 17271 5097
rect 16893 5072 16991 5074
rect 17018 5072 17186 5084
rect 17201 5074 17217 5088
rect 17252 5075 17274 5094
rect 17284 5088 17300 5089
rect 17283 5086 17300 5088
rect 17284 5081 17300 5086
rect 17274 5074 17280 5075
rect 17283 5074 17312 5081
rect 17201 5073 17312 5074
rect 17201 5072 17318 5073
rect 16877 5064 16928 5072
rect 16975 5064 17009 5072
rect 16877 5052 16902 5064
rect 16909 5052 16928 5064
rect 16982 5062 17009 5064
rect 17018 5062 17239 5072
rect 17274 5069 17280 5072
rect 16982 5058 17239 5062
rect 16877 5044 16928 5052
rect 16975 5044 17239 5058
rect 17283 5064 17318 5072
rect 16829 4996 16848 5030
rect 16893 5036 16922 5044
rect 16893 5030 16910 5036
rect 16893 5028 16927 5030
rect 16975 5028 16991 5044
rect 16992 5034 17200 5044
rect 17201 5034 17217 5044
rect 17265 5040 17280 5055
rect 17283 5052 17284 5064
rect 17291 5052 17318 5064
rect 17283 5044 17318 5052
rect 17283 5043 17312 5044
rect 17003 5030 17217 5034
rect 17018 5028 17217 5030
rect 17252 5030 17265 5040
rect 17283 5030 17300 5043
rect 17252 5028 17300 5030
rect 16894 5024 16927 5028
rect 16890 5022 16927 5024
rect 16890 5021 16957 5022
rect 16890 5016 16921 5021
rect 16927 5016 16957 5021
rect 16890 5012 16957 5016
rect 16863 5009 16957 5012
rect 16863 5002 16912 5009
rect 16863 4996 16893 5002
rect 16912 4997 16917 5002
rect 16829 4980 16909 4996
rect 16921 4988 16957 5009
rect 17018 5004 17207 5028
rect 17252 5027 17299 5028
rect 17265 5022 17299 5027
rect 17033 5001 17207 5004
rect 17026 4998 17207 5001
rect 17235 5021 17299 5022
rect 16829 4978 16848 4980
rect 16863 4978 16897 4980
rect 16829 4962 16909 4978
rect 16829 4956 16848 4962
rect 16545 4930 16648 4940
rect 16499 4928 16648 4930
rect 16669 4928 16704 4940
rect 16338 4926 16500 4928
rect 16350 4906 16369 4926
rect 16384 4924 16414 4926
rect 16233 4898 16274 4906
rect 16356 4902 16369 4906
rect 16421 4910 16500 4926
rect 16532 4926 16704 4928
rect 16532 4910 16611 4926
rect 16618 4924 16648 4926
rect 16196 4888 16225 4898
rect 16239 4888 16268 4898
rect 16283 4888 16313 4902
rect 16356 4888 16399 4902
rect 16421 4898 16611 4910
rect 16676 4906 16682 4926
rect 16406 4888 16436 4898
rect 16437 4888 16595 4898
rect 16599 4888 16629 4898
rect 16633 4888 16663 4902
rect 16691 4888 16704 4926
rect 16776 4940 16805 4956
rect 16819 4940 16848 4956
rect 16863 4946 16893 4962
rect 16921 4940 16927 4988
rect 16930 4982 16949 4988
rect 16964 4982 16994 4990
rect 16930 4974 16994 4982
rect 16930 4958 17010 4974
rect 17026 4967 17088 4998
rect 17104 4967 17166 4998
rect 17235 4996 17284 5021
rect 17299 4996 17329 5012
rect 17198 4982 17228 4990
rect 17235 4988 17345 4996
rect 17198 4974 17243 4982
rect 16930 4956 16949 4958
rect 16964 4956 17010 4958
rect 16930 4940 17010 4956
rect 17037 4954 17072 4967
rect 17113 4964 17150 4967
rect 17113 4962 17155 4964
rect 17042 4951 17072 4954
rect 17051 4947 17058 4951
rect 17058 4946 17059 4947
rect 17017 4940 17027 4946
rect 16776 4932 16811 4940
rect 16776 4906 16777 4932
rect 16784 4906 16811 4932
rect 16719 4888 16749 4902
rect 16776 4898 16811 4906
rect 16813 4932 16854 4940
rect 16813 4906 16828 4932
rect 16835 4906 16854 4932
rect 16918 4928 16949 4940
rect 16964 4928 17067 4940
rect 17079 4930 17105 4956
rect 17120 4951 17150 4962
rect 17182 4958 17244 4974
rect 17182 4956 17228 4958
rect 17182 4940 17244 4956
rect 17256 4940 17262 4988
rect 17265 4980 17345 4988
rect 17265 4978 17284 4980
rect 17299 4978 17333 4980
rect 17265 4962 17345 4978
rect 17265 4940 17284 4962
rect 17299 4946 17329 4962
rect 17357 4956 17363 5030
rect 17366 4956 17385 5100
rect 17400 4956 17406 5100
rect 17415 5030 17428 5100
rect 17480 5096 17502 5100
rect 17473 5074 17502 5088
rect 17555 5074 17571 5088
rect 17609 5084 17615 5086
rect 17622 5084 17730 5100
rect 17737 5084 17743 5086
rect 17751 5084 17766 5100
rect 17832 5094 17851 5097
rect 17473 5072 17571 5074
rect 17598 5072 17766 5084
rect 17781 5074 17797 5088
rect 17832 5075 17854 5094
rect 17864 5088 17880 5089
rect 17863 5086 17880 5088
rect 17864 5081 17880 5086
rect 17854 5074 17860 5075
rect 17863 5074 17892 5081
rect 17781 5073 17892 5074
rect 17781 5072 17898 5073
rect 17457 5064 17508 5072
rect 17555 5064 17589 5072
rect 17457 5052 17482 5064
rect 17489 5052 17508 5064
rect 17562 5062 17589 5064
rect 17598 5062 17819 5072
rect 17854 5069 17860 5072
rect 17562 5058 17819 5062
rect 17457 5044 17508 5052
rect 17555 5044 17819 5058
rect 17863 5064 17898 5072
rect 17409 4996 17428 5030
rect 17473 5036 17502 5044
rect 17473 5030 17490 5036
rect 17473 5028 17507 5030
rect 17555 5028 17571 5044
rect 17572 5034 17780 5044
rect 17781 5034 17797 5044
rect 17845 5040 17860 5055
rect 17863 5052 17864 5064
rect 17871 5052 17898 5064
rect 17863 5044 17898 5052
rect 17863 5043 17892 5044
rect 17583 5030 17797 5034
rect 17598 5028 17797 5030
rect 17832 5030 17845 5040
rect 17863 5030 17880 5043
rect 17832 5028 17880 5030
rect 17474 5024 17507 5028
rect 17470 5022 17507 5024
rect 17470 5021 17537 5022
rect 17470 5016 17501 5021
rect 17507 5016 17537 5021
rect 17470 5012 17537 5016
rect 17443 5009 17537 5012
rect 17443 5002 17492 5009
rect 17443 4996 17473 5002
rect 17492 4997 17497 5002
rect 17409 4980 17489 4996
rect 17501 4988 17537 5009
rect 17598 5004 17787 5028
rect 17832 5027 17879 5028
rect 17845 5022 17879 5027
rect 17613 5001 17787 5004
rect 17606 4998 17787 5001
rect 17815 5021 17879 5022
rect 17409 4978 17428 4980
rect 17443 4978 17477 4980
rect 17409 4962 17489 4978
rect 17409 4956 17428 4962
rect 17125 4930 17228 4940
rect 17079 4928 17228 4930
rect 17249 4928 17284 4940
rect 16918 4926 17080 4928
rect 16930 4906 16949 4926
rect 16964 4924 16994 4926
rect 16813 4898 16854 4906
rect 16936 4902 16949 4906
rect 17001 4910 17080 4926
rect 17112 4926 17284 4928
rect 17112 4910 17191 4926
rect 17198 4924 17228 4926
rect 16776 4888 16805 4898
rect 16819 4888 16848 4898
rect 16863 4888 16893 4902
rect 16936 4888 16979 4902
rect 17001 4898 17191 4910
rect 17256 4906 17262 4926
rect 16986 4888 17016 4898
rect 17017 4888 17175 4898
rect 17179 4888 17209 4898
rect 17213 4888 17243 4902
rect 17271 4888 17284 4926
rect 17356 4940 17385 4956
rect 17399 4940 17428 4956
rect 17443 4946 17473 4962
rect 17501 4940 17507 4988
rect 17510 4982 17529 4988
rect 17544 4982 17574 4990
rect 17510 4974 17574 4982
rect 17510 4958 17590 4974
rect 17606 4967 17668 4998
rect 17684 4967 17746 4998
rect 17815 4996 17864 5021
rect 17879 4996 17909 5012
rect 17778 4982 17808 4990
rect 17815 4988 17925 4996
rect 17778 4974 17823 4982
rect 17510 4956 17529 4958
rect 17544 4956 17590 4958
rect 17510 4940 17590 4956
rect 17617 4954 17652 4967
rect 17693 4964 17730 4967
rect 17693 4962 17735 4964
rect 17622 4951 17652 4954
rect 17631 4947 17638 4951
rect 17638 4946 17639 4947
rect 17597 4940 17607 4946
rect 17356 4932 17391 4940
rect 17356 4906 17357 4932
rect 17364 4906 17391 4932
rect 17299 4888 17329 4902
rect 17356 4898 17391 4906
rect 17393 4932 17434 4940
rect 17393 4906 17408 4932
rect 17415 4906 17434 4932
rect 17498 4928 17529 4940
rect 17544 4928 17647 4940
rect 17659 4930 17685 4956
rect 17700 4951 17730 4962
rect 17762 4958 17824 4974
rect 17762 4956 17808 4958
rect 17762 4940 17824 4956
rect 17836 4940 17842 4988
rect 17845 4980 17925 4988
rect 17845 4978 17864 4980
rect 17879 4978 17913 4980
rect 17845 4962 17925 4978
rect 17845 4940 17864 4962
rect 17879 4946 17909 4962
rect 17937 4956 17943 5030
rect 17946 4956 17965 5100
rect 17980 4956 17986 5100
rect 17995 5030 18008 5100
rect 18060 5096 18082 5100
rect 18053 5074 18082 5088
rect 18135 5074 18151 5088
rect 18189 5084 18195 5086
rect 18202 5084 18310 5100
rect 18317 5084 18323 5086
rect 18331 5084 18346 5100
rect 18412 5094 18431 5097
rect 18053 5072 18151 5074
rect 18178 5072 18346 5084
rect 18361 5074 18377 5088
rect 18412 5075 18434 5094
rect 18444 5088 18460 5089
rect 18443 5086 18460 5088
rect 18444 5081 18460 5086
rect 18434 5074 18440 5075
rect 18443 5074 18472 5081
rect 18361 5073 18472 5074
rect 18361 5072 18478 5073
rect 18037 5064 18088 5072
rect 18135 5064 18169 5072
rect 18037 5052 18062 5064
rect 18069 5052 18088 5064
rect 18142 5062 18169 5064
rect 18178 5062 18399 5072
rect 18434 5069 18440 5072
rect 18142 5058 18399 5062
rect 18037 5044 18088 5052
rect 18135 5044 18399 5058
rect 18443 5064 18478 5072
rect 17989 4996 18008 5030
rect 18053 5036 18082 5044
rect 18053 5030 18070 5036
rect 18053 5028 18087 5030
rect 18135 5028 18151 5044
rect 18152 5034 18360 5044
rect 18361 5034 18377 5044
rect 18425 5040 18440 5055
rect 18443 5052 18444 5064
rect 18451 5052 18478 5064
rect 18443 5044 18478 5052
rect 18443 5043 18472 5044
rect 18163 5030 18377 5034
rect 18178 5028 18377 5030
rect 18412 5030 18425 5040
rect 18443 5030 18460 5043
rect 18412 5028 18460 5030
rect 18054 5024 18087 5028
rect 18050 5022 18087 5024
rect 18050 5021 18117 5022
rect 18050 5016 18081 5021
rect 18087 5016 18117 5021
rect 18050 5012 18117 5016
rect 18023 5009 18117 5012
rect 18023 5002 18072 5009
rect 18023 4996 18053 5002
rect 18072 4997 18077 5002
rect 17989 4980 18069 4996
rect 18081 4988 18117 5009
rect 18178 5004 18367 5028
rect 18412 5027 18459 5028
rect 18425 5022 18459 5027
rect 18193 5001 18367 5004
rect 18186 4998 18367 5001
rect 18395 5021 18459 5022
rect 17989 4978 18008 4980
rect 18023 4978 18057 4980
rect 17989 4962 18069 4978
rect 17989 4956 18008 4962
rect 17705 4930 17808 4940
rect 17659 4928 17808 4930
rect 17829 4928 17864 4940
rect 17498 4926 17660 4928
rect 17510 4906 17529 4926
rect 17544 4924 17574 4926
rect 17393 4898 17434 4906
rect 17516 4902 17529 4906
rect 17581 4910 17660 4926
rect 17692 4926 17864 4928
rect 17692 4910 17771 4926
rect 17778 4924 17808 4926
rect 17356 4888 17385 4898
rect 17399 4888 17428 4898
rect 17443 4888 17473 4902
rect 17516 4888 17559 4902
rect 17581 4898 17771 4910
rect 17836 4906 17842 4926
rect 17566 4888 17596 4898
rect 17597 4888 17755 4898
rect 17759 4888 17789 4898
rect 17793 4888 17823 4902
rect 17851 4888 17864 4926
rect 17936 4940 17965 4956
rect 17979 4940 18008 4956
rect 18023 4946 18053 4962
rect 18081 4940 18087 4988
rect 18090 4982 18109 4988
rect 18124 4982 18154 4990
rect 18090 4974 18154 4982
rect 18090 4958 18170 4974
rect 18186 4967 18248 4998
rect 18264 4967 18326 4998
rect 18395 4996 18444 5021
rect 18459 4996 18489 5012
rect 18358 4982 18388 4990
rect 18395 4988 18505 4996
rect 18358 4974 18403 4982
rect 18090 4956 18109 4958
rect 18124 4956 18170 4958
rect 18090 4940 18170 4956
rect 18197 4954 18232 4967
rect 18273 4964 18310 4967
rect 18273 4962 18315 4964
rect 18202 4951 18232 4954
rect 18211 4947 18218 4951
rect 18218 4946 18219 4947
rect 18177 4940 18187 4946
rect 17936 4932 17971 4940
rect 17936 4906 17937 4932
rect 17944 4906 17971 4932
rect 17879 4888 17909 4902
rect 17936 4898 17971 4906
rect 17973 4932 18014 4940
rect 17973 4906 17988 4932
rect 17995 4906 18014 4932
rect 18078 4928 18109 4940
rect 18124 4928 18227 4940
rect 18239 4930 18265 4956
rect 18280 4951 18310 4962
rect 18342 4958 18404 4974
rect 18342 4956 18388 4958
rect 18342 4940 18404 4956
rect 18416 4940 18422 4988
rect 18425 4980 18505 4988
rect 18425 4978 18444 4980
rect 18459 4978 18493 4980
rect 18425 4962 18505 4978
rect 18425 4940 18444 4962
rect 18459 4946 18489 4962
rect 18517 4956 18523 5030
rect 18532 4956 18545 5100
rect 18285 4930 18388 4940
rect 18239 4928 18388 4930
rect 18409 4928 18444 4940
rect 18078 4926 18240 4928
rect 18090 4906 18109 4926
rect 18124 4924 18154 4926
rect 17973 4898 18014 4906
rect 18096 4902 18109 4906
rect 18161 4910 18240 4926
rect 18272 4926 18444 4928
rect 18272 4910 18351 4926
rect 18358 4924 18388 4926
rect 17936 4888 17965 4898
rect 17979 4888 18008 4898
rect 18023 4888 18053 4902
rect 18096 4888 18139 4902
rect 18161 4898 18351 4910
rect 18416 4906 18422 4926
rect 18146 4888 18176 4898
rect 18177 4888 18335 4898
rect 18339 4888 18369 4898
rect 18373 4888 18403 4902
rect 18431 4888 18444 4926
rect 18516 4940 18545 4956
rect 18516 4932 18551 4940
rect 18516 4906 18517 4932
rect 18524 4906 18551 4932
rect 18459 4888 18489 4902
rect 18516 4898 18551 4906
rect 18516 4888 18545 4898
rect -1 4882 18545 4888
rect 0 4874 18545 4882
rect 15 4844 28 4874
rect 43 4860 73 4874
rect 116 4860 159 4874
rect 166 4860 386 4874
rect 393 4860 423 4874
rect 83 4846 98 4858
rect 117 4846 130 4860
rect 198 4856 351 4860
rect 80 4844 102 4846
rect 180 4844 372 4856
rect 451 4844 464 4874
rect 479 4860 509 4874
rect 546 4844 565 4874
rect 580 4844 586 4874
rect 595 4844 608 4874
rect 623 4860 653 4874
rect 696 4860 739 4874
rect 746 4860 966 4874
rect 973 4860 1003 4874
rect 663 4846 678 4858
rect 697 4846 710 4860
rect 778 4856 931 4860
rect 660 4844 682 4846
rect 760 4844 952 4856
rect 1031 4844 1044 4874
rect 1059 4860 1089 4874
rect 1126 4844 1145 4874
rect 1160 4844 1166 4874
rect 1175 4844 1188 4874
rect 1203 4860 1233 4874
rect 1276 4860 1319 4874
rect 1326 4860 1546 4874
rect 1553 4860 1583 4874
rect 1243 4846 1258 4858
rect 1277 4846 1290 4860
rect 1358 4856 1511 4860
rect 1240 4844 1262 4846
rect 1340 4844 1532 4856
rect 1611 4844 1624 4874
rect 1639 4860 1669 4874
rect 1706 4844 1725 4874
rect 1740 4844 1746 4874
rect 1755 4844 1768 4874
rect 1783 4860 1813 4874
rect 1856 4860 1899 4874
rect 1906 4860 2126 4874
rect 2133 4860 2163 4874
rect 1823 4846 1838 4858
rect 1857 4846 1870 4860
rect 1938 4856 2091 4860
rect 1820 4844 1842 4846
rect 1920 4844 2112 4856
rect 2191 4844 2204 4874
rect 2219 4860 2249 4874
rect 2286 4844 2305 4874
rect 2320 4844 2326 4874
rect 2335 4844 2348 4874
rect 2363 4860 2393 4874
rect 2436 4860 2479 4874
rect 2486 4860 2706 4874
rect 2713 4860 2743 4874
rect 2403 4846 2418 4858
rect 2437 4846 2450 4860
rect 2518 4856 2671 4860
rect 2400 4844 2422 4846
rect 2500 4844 2692 4856
rect 2771 4844 2784 4874
rect 2799 4860 2829 4874
rect 2866 4844 2885 4874
rect 2900 4844 2906 4874
rect 2915 4844 2928 4874
rect 2943 4860 2973 4874
rect 3016 4860 3059 4874
rect 3066 4860 3286 4874
rect 3293 4860 3323 4874
rect 2983 4846 2998 4858
rect 3017 4846 3030 4860
rect 3098 4856 3251 4860
rect 2980 4844 3002 4846
rect 3080 4844 3272 4856
rect 3351 4844 3364 4874
rect 3379 4860 3409 4874
rect 3446 4844 3465 4874
rect 3480 4844 3486 4874
rect 3495 4844 3508 4874
rect 3523 4860 3553 4874
rect 3596 4860 3639 4874
rect 3646 4860 3866 4874
rect 3873 4860 3903 4874
rect 3563 4846 3578 4858
rect 3597 4846 3610 4860
rect 3678 4856 3831 4860
rect 3560 4844 3582 4846
rect 3660 4844 3852 4856
rect 3931 4844 3944 4874
rect 3959 4860 3989 4874
rect 4026 4844 4045 4874
rect 4060 4844 4066 4874
rect 4075 4844 4088 4874
rect 4103 4860 4133 4874
rect 4176 4860 4219 4874
rect 4226 4860 4446 4874
rect 4453 4860 4483 4874
rect 4143 4846 4158 4858
rect 4177 4846 4190 4860
rect 4258 4856 4411 4860
rect 4140 4844 4162 4846
rect 4240 4844 4432 4856
rect 4511 4844 4524 4874
rect 4539 4860 4569 4874
rect 4606 4844 4625 4874
rect 4640 4844 4646 4874
rect 4655 4844 4668 4874
rect 4683 4860 4713 4874
rect 4756 4860 4799 4874
rect 4806 4860 5026 4874
rect 5033 4860 5063 4874
rect 4723 4846 4738 4858
rect 4757 4846 4770 4860
rect 4838 4856 4991 4860
rect 4720 4844 4742 4846
rect 4820 4844 5012 4856
rect 5091 4844 5104 4874
rect 5119 4860 5149 4874
rect 5186 4844 5205 4874
rect 5220 4844 5226 4874
rect 5235 4844 5248 4874
rect 5263 4860 5293 4874
rect 5336 4860 5379 4874
rect 5386 4860 5606 4874
rect 5613 4860 5643 4874
rect 5303 4846 5318 4858
rect 5337 4846 5350 4860
rect 5418 4856 5571 4860
rect 5300 4844 5322 4846
rect 5400 4844 5592 4856
rect 5671 4844 5684 4874
rect 5699 4860 5729 4874
rect 5766 4844 5785 4874
rect 5800 4844 5806 4874
rect 5815 4844 5828 4874
rect 5843 4860 5873 4874
rect 5916 4860 5959 4874
rect 5966 4860 6186 4874
rect 6193 4860 6223 4874
rect 5883 4846 5898 4858
rect 5917 4846 5930 4860
rect 5998 4856 6151 4860
rect 5880 4844 5902 4846
rect 5980 4844 6172 4856
rect 6251 4844 6264 4874
rect 6279 4860 6309 4874
rect 6346 4844 6365 4874
rect 6380 4844 6386 4874
rect 6395 4844 6408 4874
rect 6423 4860 6453 4874
rect 6496 4860 6539 4874
rect 6546 4860 6766 4874
rect 6773 4860 6803 4874
rect 6463 4846 6478 4858
rect 6497 4846 6510 4860
rect 6578 4856 6731 4860
rect 6460 4844 6482 4846
rect 6560 4844 6752 4856
rect 6831 4844 6844 4874
rect 6859 4860 6889 4874
rect 6926 4844 6945 4874
rect 6960 4844 6966 4874
rect 6975 4844 6988 4874
rect 7003 4860 7033 4874
rect 7076 4860 7119 4874
rect 7126 4860 7346 4874
rect 7353 4860 7383 4874
rect 7043 4846 7058 4858
rect 7077 4846 7090 4860
rect 7158 4856 7311 4860
rect 7040 4844 7062 4846
rect 7140 4844 7332 4856
rect 7411 4844 7424 4874
rect 7439 4860 7469 4874
rect 7506 4844 7525 4874
rect 7540 4844 7546 4874
rect 7555 4844 7568 4874
rect 7583 4860 7613 4874
rect 7656 4860 7699 4874
rect 7706 4860 7926 4874
rect 7933 4860 7963 4874
rect 7623 4846 7638 4858
rect 7657 4846 7670 4860
rect 7738 4856 7891 4860
rect 7620 4844 7642 4846
rect 7720 4844 7912 4856
rect 7991 4844 8004 4874
rect 8019 4860 8049 4874
rect 8086 4844 8105 4874
rect 8120 4844 8126 4874
rect 8135 4844 8148 4874
rect 8163 4860 8193 4874
rect 8236 4860 8279 4874
rect 8286 4860 8506 4874
rect 8513 4860 8543 4874
rect 8203 4846 8218 4858
rect 8237 4846 8250 4860
rect 8318 4856 8471 4860
rect 8200 4844 8222 4846
rect 8300 4844 8492 4856
rect 8571 4844 8584 4874
rect 8599 4860 8629 4874
rect 8666 4844 8685 4874
rect 8700 4844 8706 4874
rect 8715 4844 8728 4874
rect 8743 4860 8773 4874
rect 8816 4860 8859 4874
rect 8866 4860 9086 4874
rect 9093 4860 9123 4874
rect 8783 4846 8798 4858
rect 8817 4846 8830 4860
rect 8898 4856 9051 4860
rect 8780 4844 8802 4846
rect 8880 4844 9072 4856
rect 9151 4844 9164 4874
rect 9179 4860 9209 4874
rect 9246 4844 9265 4874
rect 9280 4844 9286 4874
rect 9295 4844 9308 4874
rect 9323 4860 9353 4874
rect 9396 4860 9439 4874
rect 9446 4860 9666 4874
rect 9673 4860 9703 4874
rect 9363 4846 9378 4858
rect 9397 4846 9410 4860
rect 9478 4856 9631 4860
rect 9360 4844 9382 4846
rect 9460 4844 9652 4856
rect 9731 4844 9744 4874
rect 9759 4860 9789 4874
rect 9826 4844 9845 4874
rect 9860 4844 9866 4874
rect 9875 4844 9888 4874
rect 9903 4860 9933 4874
rect 9976 4860 10019 4874
rect 10026 4860 10246 4874
rect 10253 4860 10283 4874
rect 9943 4846 9958 4858
rect 9977 4846 9990 4860
rect 10058 4856 10211 4860
rect 9940 4844 9962 4846
rect 10040 4844 10232 4856
rect 10311 4844 10324 4874
rect 10339 4860 10369 4874
rect 10406 4844 10425 4874
rect 10440 4844 10446 4874
rect 10455 4844 10468 4874
rect 10483 4860 10513 4874
rect 10556 4860 10599 4874
rect 10606 4860 10826 4874
rect 10833 4860 10863 4874
rect 10523 4846 10538 4858
rect 10557 4846 10570 4860
rect 10638 4856 10791 4860
rect 10520 4844 10542 4846
rect 10620 4844 10812 4856
rect 10891 4844 10904 4874
rect 10919 4860 10949 4874
rect 10986 4844 11005 4874
rect 11020 4844 11026 4874
rect 11035 4844 11048 4874
rect 11063 4860 11093 4874
rect 11136 4860 11179 4874
rect 11186 4860 11406 4874
rect 11413 4860 11443 4874
rect 11103 4846 11118 4858
rect 11137 4846 11150 4860
rect 11218 4856 11371 4860
rect 11100 4844 11122 4846
rect 11200 4844 11392 4856
rect 11471 4844 11484 4874
rect 11499 4860 11529 4874
rect 11566 4844 11585 4874
rect 11600 4844 11606 4874
rect 11615 4844 11628 4874
rect 11643 4860 11673 4874
rect 11716 4860 11759 4874
rect 11766 4860 11986 4874
rect 11993 4860 12023 4874
rect 11683 4846 11698 4858
rect 11717 4846 11730 4860
rect 11798 4856 11951 4860
rect 11680 4844 11702 4846
rect 11780 4844 11972 4856
rect 12051 4844 12064 4874
rect 12079 4860 12109 4874
rect 12146 4844 12165 4874
rect 12180 4844 12186 4874
rect 12195 4844 12208 4874
rect 12223 4860 12253 4874
rect 12296 4860 12339 4874
rect 12346 4860 12566 4874
rect 12573 4860 12603 4874
rect 12263 4846 12278 4858
rect 12297 4846 12310 4860
rect 12378 4856 12531 4860
rect 12260 4844 12282 4846
rect 12360 4844 12552 4856
rect 12631 4844 12644 4874
rect 12659 4860 12689 4874
rect 12726 4844 12745 4874
rect 12760 4844 12766 4874
rect 12775 4844 12788 4874
rect 12803 4860 12833 4874
rect 12876 4860 12919 4874
rect 12926 4860 13146 4874
rect 13153 4860 13183 4874
rect 12843 4846 12858 4858
rect 12877 4846 12890 4860
rect 12958 4856 13111 4860
rect 12840 4844 12862 4846
rect 12940 4844 13132 4856
rect 13211 4844 13224 4874
rect 13239 4860 13269 4874
rect 13306 4844 13325 4874
rect 13340 4844 13346 4874
rect 13355 4844 13368 4874
rect 13383 4860 13413 4874
rect 13456 4860 13499 4874
rect 13506 4860 13726 4874
rect 13733 4860 13763 4874
rect 13423 4846 13438 4858
rect 13457 4846 13470 4860
rect 13538 4856 13691 4860
rect 13420 4844 13442 4846
rect 13520 4844 13712 4856
rect 13791 4844 13804 4874
rect 13819 4860 13849 4874
rect 13886 4844 13905 4874
rect 13920 4844 13926 4874
rect 13935 4844 13948 4874
rect 13963 4860 13993 4874
rect 14036 4860 14079 4874
rect 14086 4860 14306 4874
rect 14313 4860 14343 4874
rect 14003 4846 14018 4858
rect 14037 4846 14050 4860
rect 14118 4856 14271 4860
rect 14000 4844 14022 4846
rect 14100 4844 14292 4856
rect 14371 4844 14384 4874
rect 14399 4860 14429 4874
rect 14466 4844 14485 4874
rect 14500 4844 14506 4874
rect 14515 4844 14528 4874
rect 14543 4860 14573 4874
rect 14616 4860 14659 4874
rect 14666 4860 14886 4874
rect 14893 4860 14923 4874
rect 14583 4846 14598 4858
rect 14617 4846 14630 4860
rect 14698 4856 14851 4860
rect 14580 4844 14602 4846
rect 14680 4844 14872 4856
rect 14951 4844 14964 4874
rect 14979 4860 15009 4874
rect 15046 4844 15065 4874
rect 15080 4844 15086 4874
rect 15095 4844 15108 4874
rect 15123 4860 15153 4874
rect 15196 4860 15239 4874
rect 15246 4860 15466 4874
rect 15473 4860 15503 4874
rect 15163 4846 15178 4858
rect 15197 4846 15210 4860
rect 15278 4856 15431 4860
rect 15160 4844 15182 4846
rect 15260 4844 15452 4856
rect 15531 4844 15544 4874
rect 15559 4860 15589 4874
rect 15626 4844 15645 4874
rect 15660 4844 15666 4874
rect 15675 4844 15688 4874
rect 15703 4860 15733 4874
rect 15776 4860 15819 4874
rect 15826 4860 16046 4874
rect 16053 4860 16083 4874
rect 15743 4846 15758 4858
rect 15777 4846 15790 4860
rect 15858 4856 16011 4860
rect 15740 4844 15762 4846
rect 15840 4844 16032 4856
rect 16111 4844 16124 4874
rect 16139 4860 16169 4874
rect 16206 4844 16225 4874
rect 16240 4844 16246 4874
rect 16255 4844 16268 4874
rect 16283 4860 16313 4874
rect 16356 4860 16399 4874
rect 16406 4860 16626 4874
rect 16633 4860 16663 4874
rect 16323 4846 16338 4858
rect 16357 4846 16370 4860
rect 16438 4856 16591 4860
rect 16320 4844 16342 4846
rect 16420 4844 16612 4856
rect 16691 4844 16704 4874
rect 16719 4860 16749 4874
rect 16786 4844 16805 4874
rect 16820 4844 16826 4874
rect 16835 4844 16848 4874
rect 16863 4860 16893 4874
rect 16936 4860 16979 4874
rect 16986 4860 17206 4874
rect 17213 4860 17243 4874
rect 16903 4846 16918 4858
rect 16937 4846 16950 4860
rect 17018 4856 17171 4860
rect 16900 4844 16922 4846
rect 17000 4844 17192 4856
rect 17271 4844 17284 4874
rect 17299 4860 17329 4874
rect 17366 4844 17385 4874
rect 17400 4844 17406 4874
rect 17415 4844 17428 4874
rect 17443 4860 17473 4874
rect 17516 4860 17559 4874
rect 17566 4860 17786 4874
rect 17793 4860 17823 4874
rect 17483 4846 17498 4858
rect 17517 4846 17530 4860
rect 17598 4856 17751 4860
rect 17480 4844 17502 4846
rect 17580 4844 17772 4856
rect 17851 4844 17864 4874
rect 17879 4860 17909 4874
rect 17946 4844 17965 4874
rect 17980 4844 17986 4874
rect 17995 4844 18008 4874
rect 18023 4860 18053 4874
rect 18096 4860 18139 4874
rect 18146 4860 18366 4874
rect 18373 4860 18403 4874
rect 18063 4846 18078 4858
rect 18097 4846 18110 4860
rect 18178 4856 18331 4860
rect 18060 4844 18082 4846
rect 18160 4844 18352 4856
rect 18431 4844 18444 4874
rect 18459 4860 18489 4874
rect 18532 4844 18545 4874
rect 0 4830 18545 4844
rect 15 4760 28 4830
rect 80 4826 102 4830
rect 73 4804 102 4818
rect 155 4804 171 4818
rect 209 4814 215 4816
rect 222 4814 330 4830
rect 337 4814 343 4816
rect 351 4814 366 4830
rect 432 4824 451 4827
rect 73 4802 171 4804
rect 198 4802 366 4814
rect 381 4804 397 4818
rect 432 4805 454 4824
rect 464 4818 480 4819
rect 463 4816 480 4818
rect 464 4811 480 4816
rect 454 4804 460 4805
rect 463 4804 492 4811
rect 381 4803 492 4804
rect 381 4802 498 4803
rect 57 4794 108 4802
rect 155 4794 189 4802
rect 57 4782 82 4794
rect 89 4782 108 4794
rect 162 4792 189 4794
rect 198 4792 419 4802
rect 454 4799 460 4802
rect 162 4788 419 4792
rect 57 4774 108 4782
rect 155 4774 419 4788
rect 463 4794 498 4802
rect 9 4726 28 4760
rect 73 4766 102 4774
rect 73 4760 90 4766
rect 73 4758 107 4760
rect 155 4758 171 4774
rect 172 4764 380 4774
rect 381 4764 397 4774
rect 445 4770 460 4785
rect 463 4782 464 4794
rect 471 4782 498 4794
rect 463 4774 498 4782
rect 463 4773 492 4774
rect 183 4760 397 4764
rect 198 4758 397 4760
rect 432 4760 445 4770
rect 463 4760 480 4773
rect 432 4758 480 4760
rect 74 4754 107 4758
rect 70 4752 107 4754
rect 70 4751 137 4752
rect 70 4746 101 4751
rect 107 4746 137 4751
rect 70 4742 137 4746
rect 43 4739 137 4742
rect 43 4732 92 4739
rect 43 4726 73 4732
rect 92 4727 97 4732
rect 9 4710 89 4726
rect 101 4718 137 4739
rect 198 4734 387 4758
rect 432 4757 479 4758
rect 445 4752 479 4757
rect 213 4731 387 4734
rect 206 4728 387 4731
rect 415 4751 479 4752
rect 9 4708 28 4710
rect 43 4708 77 4710
rect 9 4692 89 4708
rect 9 4686 28 4692
rect -1 4670 28 4686
rect 43 4676 73 4692
rect 101 4670 107 4718
rect 110 4712 129 4718
rect 144 4712 174 4720
rect 110 4704 174 4712
rect 110 4688 190 4704
rect 206 4697 268 4728
rect 284 4697 346 4728
rect 415 4726 464 4751
rect 479 4726 509 4742
rect 378 4712 408 4720
rect 415 4718 525 4726
rect 378 4704 423 4712
rect 110 4686 129 4688
rect 144 4686 190 4688
rect 110 4670 190 4686
rect 217 4684 252 4697
rect 293 4694 330 4697
rect 293 4692 335 4694
rect 222 4681 252 4684
rect 231 4677 238 4681
rect 238 4676 239 4677
rect 197 4670 207 4676
rect -7 4662 34 4670
rect -7 4636 8 4662
rect 15 4636 34 4662
rect 98 4658 129 4670
rect 144 4658 247 4670
rect 259 4660 285 4686
rect 300 4681 330 4692
rect 362 4688 424 4704
rect 362 4686 408 4688
rect 362 4670 424 4686
rect 436 4670 442 4718
rect 445 4710 525 4718
rect 445 4708 464 4710
rect 479 4708 513 4710
rect 445 4692 525 4708
rect 445 4670 464 4692
rect 479 4676 509 4692
rect 537 4686 543 4760
rect 546 4686 565 4830
rect 580 4686 586 4830
rect 595 4760 608 4830
rect 660 4826 682 4830
rect 653 4804 682 4818
rect 735 4804 751 4818
rect 789 4814 795 4816
rect 802 4814 910 4830
rect 917 4814 923 4816
rect 931 4814 946 4830
rect 1012 4824 1031 4827
rect 653 4802 751 4804
rect 778 4802 946 4814
rect 961 4804 977 4818
rect 1012 4805 1034 4824
rect 1044 4818 1060 4819
rect 1043 4816 1060 4818
rect 1044 4811 1060 4816
rect 1034 4804 1040 4805
rect 1043 4804 1072 4811
rect 961 4803 1072 4804
rect 961 4802 1078 4803
rect 637 4794 688 4802
rect 735 4794 769 4802
rect 637 4782 662 4794
rect 669 4782 688 4794
rect 742 4792 769 4794
rect 778 4792 999 4802
rect 1034 4799 1040 4802
rect 742 4788 999 4792
rect 637 4774 688 4782
rect 735 4774 999 4788
rect 1043 4794 1078 4802
rect 589 4726 608 4760
rect 653 4766 682 4774
rect 653 4760 670 4766
rect 653 4758 687 4760
rect 735 4758 751 4774
rect 752 4764 960 4774
rect 961 4764 977 4774
rect 1025 4770 1040 4785
rect 1043 4782 1044 4794
rect 1051 4782 1078 4794
rect 1043 4774 1078 4782
rect 1043 4773 1072 4774
rect 763 4760 977 4764
rect 778 4758 977 4760
rect 1012 4760 1025 4770
rect 1043 4760 1060 4773
rect 1012 4758 1060 4760
rect 654 4754 687 4758
rect 650 4752 687 4754
rect 650 4751 717 4752
rect 650 4746 681 4751
rect 687 4746 717 4751
rect 650 4742 717 4746
rect 623 4739 717 4742
rect 623 4732 672 4739
rect 623 4726 653 4732
rect 672 4727 677 4732
rect 589 4710 669 4726
rect 681 4718 717 4739
rect 778 4734 967 4758
rect 1012 4757 1059 4758
rect 1025 4752 1059 4757
rect 793 4731 967 4734
rect 786 4728 967 4731
rect 995 4751 1059 4752
rect 589 4708 608 4710
rect 623 4708 657 4710
rect 589 4692 669 4708
rect 589 4686 608 4692
rect 305 4660 408 4670
rect 259 4658 408 4660
rect 429 4658 464 4670
rect 98 4656 260 4658
rect 110 4636 129 4656
rect 144 4654 174 4656
rect -7 4628 34 4636
rect 116 4632 129 4636
rect 181 4640 260 4656
rect 292 4656 464 4658
rect 292 4640 371 4656
rect 378 4654 408 4656
rect -1 4618 28 4628
rect 43 4618 73 4632
rect 116 4618 159 4632
rect 181 4628 371 4640
rect 436 4636 442 4656
rect 166 4618 196 4628
rect 197 4618 355 4628
rect 359 4618 389 4628
rect 393 4618 423 4632
rect 451 4618 464 4656
rect 536 4670 565 4686
rect 579 4670 608 4686
rect 623 4676 653 4692
rect 681 4670 687 4718
rect 690 4712 709 4718
rect 724 4712 754 4720
rect 690 4704 754 4712
rect 690 4688 770 4704
rect 786 4697 848 4728
rect 864 4697 926 4728
rect 995 4726 1044 4751
rect 1059 4726 1089 4742
rect 958 4712 988 4720
rect 995 4718 1105 4726
rect 958 4704 1003 4712
rect 690 4686 709 4688
rect 724 4686 770 4688
rect 690 4670 770 4686
rect 797 4684 832 4697
rect 873 4694 910 4697
rect 873 4692 915 4694
rect 802 4681 832 4684
rect 811 4677 818 4681
rect 818 4676 819 4677
rect 777 4670 787 4676
rect 536 4662 571 4670
rect 536 4636 537 4662
rect 544 4636 571 4662
rect 479 4618 509 4632
rect 536 4628 571 4636
rect 573 4662 614 4670
rect 573 4636 588 4662
rect 595 4636 614 4662
rect 678 4658 709 4670
rect 724 4658 827 4670
rect 839 4660 865 4686
rect 880 4681 910 4692
rect 942 4688 1004 4704
rect 942 4686 988 4688
rect 942 4670 1004 4686
rect 1016 4670 1022 4718
rect 1025 4710 1105 4718
rect 1025 4708 1044 4710
rect 1059 4708 1093 4710
rect 1025 4692 1105 4708
rect 1025 4670 1044 4692
rect 1059 4676 1089 4692
rect 1117 4686 1123 4760
rect 1126 4686 1145 4830
rect 1160 4686 1166 4830
rect 1175 4760 1188 4830
rect 1240 4826 1262 4830
rect 1233 4804 1262 4818
rect 1315 4804 1331 4818
rect 1369 4814 1375 4816
rect 1382 4814 1490 4830
rect 1497 4814 1503 4816
rect 1511 4814 1526 4830
rect 1592 4824 1611 4827
rect 1233 4802 1331 4804
rect 1358 4802 1526 4814
rect 1541 4804 1557 4818
rect 1592 4805 1614 4824
rect 1624 4818 1640 4819
rect 1623 4816 1640 4818
rect 1624 4811 1640 4816
rect 1614 4804 1620 4805
rect 1623 4804 1652 4811
rect 1541 4803 1652 4804
rect 1541 4802 1658 4803
rect 1217 4794 1268 4802
rect 1315 4794 1349 4802
rect 1217 4782 1242 4794
rect 1249 4782 1268 4794
rect 1322 4792 1349 4794
rect 1358 4792 1579 4802
rect 1614 4799 1620 4802
rect 1322 4788 1579 4792
rect 1217 4774 1268 4782
rect 1315 4774 1579 4788
rect 1623 4794 1658 4802
rect 1169 4726 1188 4760
rect 1233 4766 1262 4774
rect 1233 4760 1250 4766
rect 1233 4758 1267 4760
rect 1315 4758 1331 4774
rect 1332 4764 1540 4774
rect 1541 4764 1557 4774
rect 1605 4770 1620 4785
rect 1623 4782 1624 4794
rect 1631 4782 1658 4794
rect 1623 4774 1658 4782
rect 1623 4773 1652 4774
rect 1343 4760 1557 4764
rect 1358 4758 1557 4760
rect 1592 4760 1605 4770
rect 1623 4760 1640 4773
rect 1592 4758 1640 4760
rect 1234 4754 1267 4758
rect 1230 4752 1267 4754
rect 1230 4751 1297 4752
rect 1230 4746 1261 4751
rect 1267 4746 1297 4751
rect 1230 4742 1297 4746
rect 1203 4739 1297 4742
rect 1203 4732 1252 4739
rect 1203 4726 1233 4732
rect 1252 4727 1257 4732
rect 1169 4710 1249 4726
rect 1261 4718 1297 4739
rect 1358 4734 1547 4758
rect 1592 4757 1639 4758
rect 1605 4752 1639 4757
rect 1373 4731 1547 4734
rect 1366 4728 1547 4731
rect 1575 4751 1639 4752
rect 1169 4708 1188 4710
rect 1203 4708 1237 4710
rect 1169 4692 1249 4708
rect 1169 4686 1188 4692
rect 885 4660 988 4670
rect 839 4658 988 4660
rect 1009 4658 1044 4670
rect 678 4656 840 4658
rect 690 4636 709 4656
rect 724 4654 754 4656
rect 573 4628 614 4636
rect 696 4632 709 4636
rect 761 4640 840 4656
rect 872 4656 1044 4658
rect 872 4640 951 4656
rect 958 4654 988 4656
rect 536 4618 565 4628
rect 579 4618 608 4628
rect 623 4618 653 4632
rect 696 4618 739 4632
rect 761 4628 951 4640
rect 1016 4636 1022 4656
rect 746 4618 776 4628
rect 777 4618 935 4628
rect 939 4618 969 4628
rect 973 4618 1003 4632
rect 1031 4618 1044 4656
rect 1116 4670 1145 4686
rect 1159 4670 1188 4686
rect 1203 4676 1233 4692
rect 1261 4670 1267 4718
rect 1270 4712 1289 4718
rect 1304 4712 1334 4720
rect 1270 4704 1334 4712
rect 1270 4688 1350 4704
rect 1366 4697 1428 4728
rect 1444 4697 1506 4728
rect 1575 4726 1624 4751
rect 1639 4726 1669 4742
rect 1538 4712 1568 4720
rect 1575 4718 1685 4726
rect 1538 4704 1583 4712
rect 1270 4686 1289 4688
rect 1304 4686 1350 4688
rect 1270 4670 1350 4686
rect 1377 4684 1412 4697
rect 1453 4694 1490 4697
rect 1453 4692 1495 4694
rect 1382 4681 1412 4684
rect 1391 4677 1398 4681
rect 1398 4676 1399 4677
rect 1357 4670 1367 4676
rect 1116 4662 1151 4670
rect 1116 4636 1117 4662
rect 1124 4636 1151 4662
rect 1059 4618 1089 4632
rect 1116 4628 1151 4636
rect 1153 4662 1194 4670
rect 1153 4636 1168 4662
rect 1175 4636 1194 4662
rect 1258 4658 1289 4670
rect 1304 4658 1407 4670
rect 1419 4660 1445 4686
rect 1460 4681 1490 4692
rect 1522 4688 1584 4704
rect 1522 4686 1568 4688
rect 1522 4670 1584 4686
rect 1596 4670 1602 4718
rect 1605 4710 1685 4718
rect 1605 4708 1624 4710
rect 1639 4708 1673 4710
rect 1605 4692 1685 4708
rect 1605 4670 1624 4692
rect 1639 4676 1669 4692
rect 1697 4686 1703 4760
rect 1706 4686 1725 4830
rect 1740 4686 1746 4830
rect 1755 4760 1768 4830
rect 1820 4826 1842 4830
rect 1813 4804 1842 4818
rect 1895 4804 1911 4818
rect 1949 4814 1955 4816
rect 1962 4814 2070 4830
rect 2077 4814 2083 4816
rect 2091 4814 2106 4830
rect 2172 4824 2191 4827
rect 1813 4802 1911 4804
rect 1938 4802 2106 4814
rect 2121 4804 2137 4818
rect 2172 4805 2194 4824
rect 2204 4818 2220 4819
rect 2203 4816 2220 4818
rect 2204 4811 2220 4816
rect 2194 4804 2200 4805
rect 2203 4804 2232 4811
rect 2121 4803 2232 4804
rect 2121 4802 2238 4803
rect 1797 4794 1848 4802
rect 1895 4794 1929 4802
rect 1797 4782 1822 4794
rect 1829 4782 1848 4794
rect 1902 4792 1929 4794
rect 1938 4792 2159 4802
rect 2194 4799 2200 4802
rect 1902 4788 2159 4792
rect 1797 4774 1848 4782
rect 1895 4774 2159 4788
rect 2203 4794 2238 4802
rect 1749 4726 1768 4760
rect 1813 4766 1842 4774
rect 1813 4760 1830 4766
rect 1813 4758 1847 4760
rect 1895 4758 1911 4774
rect 1912 4764 2120 4774
rect 2121 4764 2137 4774
rect 2185 4770 2200 4785
rect 2203 4782 2204 4794
rect 2211 4782 2238 4794
rect 2203 4774 2238 4782
rect 2203 4773 2232 4774
rect 1923 4760 2137 4764
rect 1938 4758 2137 4760
rect 2172 4760 2185 4770
rect 2203 4760 2220 4773
rect 2172 4758 2220 4760
rect 1814 4754 1847 4758
rect 1810 4752 1847 4754
rect 1810 4751 1877 4752
rect 1810 4746 1841 4751
rect 1847 4746 1877 4751
rect 1810 4742 1877 4746
rect 1783 4739 1877 4742
rect 1783 4732 1832 4739
rect 1783 4726 1813 4732
rect 1832 4727 1837 4732
rect 1749 4710 1829 4726
rect 1841 4718 1877 4739
rect 1938 4734 2127 4758
rect 2172 4757 2219 4758
rect 2185 4752 2219 4757
rect 1953 4731 2127 4734
rect 1946 4728 2127 4731
rect 2155 4751 2219 4752
rect 1749 4708 1768 4710
rect 1783 4708 1817 4710
rect 1749 4692 1829 4708
rect 1749 4686 1768 4692
rect 1465 4660 1568 4670
rect 1419 4658 1568 4660
rect 1589 4658 1624 4670
rect 1258 4656 1420 4658
rect 1270 4636 1289 4656
rect 1304 4654 1334 4656
rect 1153 4628 1194 4636
rect 1276 4632 1289 4636
rect 1341 4640 1420 4656
rect 1452 4656 1624 4658
rect 1452 4640 1531 4656
rect 1538 4654 1568 4656
rect 1116 4618 1145 4628
rect 1159 4618 1188 4628
rect 1203 4618 1233 4632
rect 1276 4618 1319 4632
rect 1341 4628 1531 4640
rect 1596 4636 1602 4656
rect 1326 4618 1356 4628
rect 1357 4618 1515 4628
rect 1519 4618 1549 4628
rect 1553 4618 1583 4632
rect 1611 4618 1624 4656
rect 1696 4670 1725 4686
rect 1739 4670 1768 4686
rect 1783 4676 1813 4692
rect 1841 4670 1847 4718
rect 1850 4712 1869 4718
rect 1884 4712 1914 4720
rect 1850 4704 1914 4712
rect 1850 4688 1930 4704
rect 1946 4697 2008 4728
rect 2024 4697 2086 4728
rect 2155 4726 2204 4751
rect 2219 4726 2249 4742
rect 2118 4712 2148 4720
rect 2155 4718 2265 4726
rect 2118 4704 2163 4712
rect 1850 4686 1869 4688
rect 1884 4686 1930 4688
rect 1850 4670 1930 4686
rect 1957 4684 1992 4697
rect 2033 4694 2070 4697
rect 2033 4692 2075 4694
rect 1962 4681 1992 4684
rect 1971 4677 1978 4681
rect 1978 4676 1979 4677
rect 1937 4670 1947 4676
rect 1696 4662 1731 4670
rect 1696 4636 1697 4662
rect 1704 4636 1731 4662
rect 1639 4618 1669 4632
rect 1696 4628 1731 4636
rect 1733 4662 1774 4670
rect 1733 4636 1748 4662
rect 1755 4636 1774 4662
rect 1838 4658 1869 4670
rect 1884 4658 1987 4670
rect 1999 4660 2025 4686
rect 2040 4681 2070 4692
rect 2102 4688 2164 4704
rect 2102 4686 2148 4688
rect 2102 4670 2164 4686
rect 2176 4670 2182 4718
rect 2185 4710 2265 4718
rect 2185 4708 2204 4710
rect 2219 4708 2253 4710
rect 2185 4692 2265 4708
rect 2185 4670 2204 4692
rect 2219 4676 2249 4692
rect 2277 4686 2283 4760
rect 2286 4686 2305 4830
rect 2320 4686 2326 4830
rect 2335 4760 2348 4830
rect 2400 4826 2422 4830
rect 2393 4804 2422 4818
rect 2475 4804 2491 4818
rect 2529 4814 2535 4816
rect 2542 4814 2650 4830
rect 2657 4814 2663 4816
rect 2671 4814 2686 4830
rect 2752 4824 2771 4827
rect 2393 4802 2491 4804
rect 2518 4802 2686 4814
rect 2701 4804 2717 4818
rect 2752 4805 2774 4824
rect 2784 4818 2800 4819
rect 2783 4816 2800 4818
rect 2784 4811 2800 4816
rect 2774 4804 2780 4805
rect 2783 4804 2812 4811
rect 2701 4803 2812 4804
rect 2701 4802 2818 4803
rect 2377 4794 2428 4802
rect 2475 4794 2509 4802
rect 2377 4782 2402 4794
rect 2409 4782 2428 4794
rect 2482 4792 2509 4794
rect 2518 4792 2739 4802
rect 2774 4799 2780 4802
rect 2482 4788 2739 4792
rect 2377 4774 2428 4782
rect 2475 4774 2739 4788
rect 2783 4794 2818 4802
rect 2329 4726 2348 4760
rect 2393 4766 2422 4774
rect 2393 4760 2410 4766
rect 2393 4758 2427 4760
rect 2475 4758 2491 4774
rect 2492 4764 2700 4774
rect 2701 4764 2717 4774
rect 2765 4770 2780 4785
rect 2783 4782 2784 4794
rect 2791 4782 2818 4794
rect 2783 4774 2818 4782
rect 2783 4773 2812 4774
rect 2503 4760 2717 4764
rect 2518 4758 2717 4760
rect 2752 4760 2765 4770
rect 2783 4760 2800 4773
rect 2752 4758 2800 4760
rect 2394 4754 2427 4758
rect 2390 4752 2427 4754
rect 2390 4751 2457 4752
rect 2390 4746 2421 4751
rect 2427 4746 2457 4751
rect 2390 4742 2457 4746
rect 2363 4739 2457 4742
rect 2363 4732 2412 4739
rect 2363 4726 2393 4732
rect 2412 4727 2417 4732
rect 2329 4710 2409 4726
rect 2421 4718 2457 4739
rect 2518 4734 2707 4758
rect 2752 4757 2799 4758
rect 2765 4752 2799 4757
rect 2533 4731 2707 4734
rect 2526 4728 2707 4731
rect 2735 4751 2799 4752
rect 2329 4708 2348 4710
rect 2363 4708 2397 4710
rect 2329 4692 2409 4708
rect 2329 4686 2348 4692
rect 2045 4660 2148 4670
rect 1999 4658 2148 4660
rect 2169 4658 2204 4670
rect 1838 4656 2000 4658
rect 1850 4636 1869 4656
rect 1884 4654 1914 4656
rect 1733 4628 1774 4636
rect 1856 4632 1869 4636
rect 1921 4640 2000 4656
rect 2032 4656 2204 4658
rect 2032 4640 2111 4656
rect 2118 4654 2148 4656
rect 1696 4618 1725 4628
rect 1739 4618 1768 4628
rect 1783 4618 1813 4632
rect 1856 4618 1899 4632
rect 1921 4628 2111 4640
rect 2176 4636 2182 4656
rect 1906 4618 1936 4628
rect 1937 4618 2095 4628
rect 2099 4618 2129 4628
rect 2133 4618 2163 4632
rect 2191 4618 2204 4656
rect 2276 4670 2305 4686
rect 2319 4670 2348 4686
rect 2363 4676 2393 4692
rect 2421 4670 2427 4718
rect 2430 4712 2449 4718
rect 2464 4712 2494 4720
rect 2430 4704 2494 4712
rect 2430 4688 2510 4704
rect 2526 4697 2588 4728
rect 2604 4697 2666 4728
rect 2735 4726 2784 4751
rect 2799 4726 2829 4742
rect 2698 4712 2728 4720
rect 2735 4718 2845 4726
rect 2698 4704 2743 4712
rect 2430 4686 2449 4688
rect 2464 4686 2510 4688
rect 2430 4670 2510 4686
rect 2537 4684 2572 4697
rect 2613 4694 2650 4697
rect 2613 4692 2655 4694
rect 2542 4681 2572 4684
rect 2551 4677 2558 4681
rect 2558 4676 2559 4677
rect 2517 4670 2527 4676
rect 2276 4662 2311 4670
rect 2276 4636 2277 4662
rect 2284 4636 2311 4662
rect 2219 4618 2249 4632
rect 2276 4628 2311 4636
rect 2313 4662 2354 4670
rect 2313 4636 2328 4662
rect 2335 4636 2354 4662
rect 2418 4658 2449 4670
rect 2464 4658 2567 4670
rect 2579 4660 2605 4686
rect 2620 4681 2650 4692
rect 2682 4688 2744 4704
rect 2682 4686 2728 4688
rect 2682 4670 2744 4686
rect 2756 4670 2762 4718
rect 2765 4710 2845 4718
rect 2765 4708 2784 4710
rect 2799 4708 2833 4710
rect 2765 4692 2845 4708
rect 2765 4670 2784 4692
rect 2799 4676 2829 4692
rect 2857 4686 2863 4760
rect 2866 4686 2885 4830
rect 2900 4686 2906 4830
rect 2915 4760 2928 4830
rect 2980 4826 3002 4830
rect 2973 4804 3002 4818
rect 3055 4804 3071 4818
rect 3109 4814 3115 4816
rect 3122 4814 3230 4830
rect 3237 4814 3243 4816
rect 3251 4814 3266 4830
rect 3332 4824 3351 4827
rect 2973 4802 3071 4804
rect 3098 4802 3266 4814
rect 3281 4804 3297 4818
rect 3332 4805 3354 4824
rect 3364 4818 3380 4819
rect 3363 4816 3380 4818
rect 3364 4811 3380 4816
rect 3354 4804 3360 4805
rect 3363 4804 3392 4811
rect 3281 4803 3392 4804
rect 3281 4802 3398 4803
rect 2957 4794 3008 4802
rect 3055 4794 3089 4802
rect 2957 4782 2982 4794
rect 2989 4782 3008 4794
rect 3062 4792 3089 4794
rect 3098 4792 3319 4802
rect 3354 4799 3360 4802
rect 3062 4788 3319 4792
rect 2957 4774 3008 4782
rect 3055 4774 3319 4788
rect 3363 4794 3398 4802
rect 2909 4726 2928 4760
rect 2973 4766 3002 4774
rect 2973 4760 2990 4766
rect 2973 4758 3007 4760
rect 3055 4758 3071 4774
rect 3072 4764 3280 4774
rect 3281 4764 3297 4774
rect 3345 4770 3360 4785
rect 3363 4782 3364 4794
rect 3371 4782 3398 4794
rect 3363 4774 3398 4782
rect 3363 4773 3392 4774
rect 3083 4760 3297 4764
rect 3098 4758 3297 4760
rect 3332 4760 3345 4770
rect 3363 4760 3380 4773
rect 3332 4758 3380 4760
rect 2974 4754 3007 4758
rect 2970 4752 3007 4754
rect 2970 4751 3037 4752
rect 2970 4746 3001 4751
rect 3007 4746 3037 4751
rect 2970 4742 3037 4746
rect 2943 4739 3037 4742
rect 2943 4732 2992 4739
rect 2943 4726 2973 4732
rect 2992 4727 2997 4732
rect 2909 4710 2989 4726
rect 3001 4718 3037 4739
rect 3098 4734 3287 4758
rect 3332 4757 3379 4758
rect 3345 4752 3379 4757
rect 3113 4731 3287 4734
rect 3106 4728 3287 4731
rect 3315 4751 3379 4752
rect 2909 4708 2928 4710
rect 2943 4708 2977 4710
rect 2909 4692 2989 4708
rect 2909 4686 2928 4692
rect 2625 4660 2728 4670
rect 2579 4658 2728 4660
rect 2749 4658 2784 4670
rect 2418 4656 2580 4658
rect 2430 4636 2449 4656
rect 2464 4654 2494 4656
rect 2313 4628 2354 4636
rect 2436 4632 2449 4636
rect 2501 4640 2580 4656
rect 2612 4656 2784 4658
rect 2612 4640 2691 4656
rect 2698 4654 2728 4656
rect 2276 4618 2305 4628
rect 2319 4618 2348 4628
rect 2363 4618 2393 4632
rect 2436 4618 2479 4632
rect 2501 4628 2691 4640
rect 2756 4636 2762 4656
rect 2486 4618 2516 4628
rect 2517 4618 2675 4628
rect 2679 4618 2709 4628
rect 2713 4618 2743 4632
rect 2771 4618 2784 4656
rect 2856 4670 2885 4686
rect 2899 4670 2928 4686
rect 2943 4676 2973 4692
rect 3001 4670 3007 4718
rect 3010 4712 3029 4718
rect 3044 4712 3074 4720
rect 3010 4704 3074 4712
rect 3010 4688 3090 4704
rect 3106 4697 3168 4728
rect 3184 4697 3246 4728
rect 3315 4726 3364 4751
rect 3379 4726 3409 4742
rect 3278 4712 3308 4720
rect 3315 4718 3425 4726
rect 3278 4704 3323 4712
rect 3010 4686 3029 4688
rect 3044 4686 3090 4688
rect 3010 4670 3090 4686
rect 3117 4684 3152 4697
rect 3193 4694 3230 4697
rect 3193 4692 3235 4694
rect 3122 4681 3152 4684
rect 3131 4677 3138 4681
rect 3138 4676 3139 4677
rect 3097 4670 3107 4676
rect 2856 4662 2891 4670
rect 2856 4636 2857 4662
rect 2864 4636 2891 4662
rect 2799 4618 2829 4632
rect 2856 4628 2891 4636
rect 2893 4662 2934 4670
rect 2893 4636 2908 4662
rect 2915 4636 2934 4662
rect 2998 4658 3029 4670
rect 3044 4658 3147 4670
rect 3159 4660 3185 4686
rect 3200 4681 3230 4692
rect 3262 4688 3324 4704
rect 3262 4686 3308 4688
rect 3262 4670 3324 4686
rect 3336 4670 3342 4718
rect 3345 4710 3425 4718
rect 3345 4708 3364 4710
rect 3379 4708 3413 4710
rect 3345 4692 3425 4708
rect 3345 4670 3364 4692
rect 3379 4676 3409 4692
rect 3437 4686 3443 4760
rect 3446 4686 3465 4830
rect 3480 4686 3486 4830
rect 3495 4760 3508 4830
rect 3560 4826 3582 4830
rect 3553 4804 3582 4818
rect 3635 4804 3651 4818
rect 3689 4814 3695 4816
rect 3702 4814 3810 4830
rect 3817 4814 3823 4816
rect 3831 4814 3846 4830
rect 3912 4824 3931 4827
rect 3553 4802 3651 4804
rect 3678 4802 3846 4814
rect 3861 4804 3877 4818
rect 3912 4805 3934 4824
rect 3944 4818 3960 4819
rect 3943 4816 3960 4818
rect 3944 4811 3960 4816
rect 3934 4804 3940 4805
rect 3943 4804 3972 4811
rect 3861 4803 3972 4804
rect 3861 4802 3978 4803
rect 3537 4794 3588 4802
rect 3635 4794 3669 4802
rect 3537 4782 3562 4794
rect 3569 4782 3588 4794
rect 3642 4792 3669 4794
rect 3678 4792 3899 4802
rect 3934 4799 3940 4802
rect 3642 4788 3899 4792
rect 3537 4774 3588 4782
rect 3635 4774 3899 4788
rect 3943 4794 3978 4802
rect 3489 4726 3508 4760
rect 3553 4766 3582 4774
rect 3553 4760 3570 4766
rect 3553 4758 3587 4760
rect 3635 4758 3651 4774
rect 3652 4764 3860 4774
rect 3861 4764 3877 4774
rect 3925 4770 3940 4785
rect 3943 4782 3944 4794
rect 3951 4782 3978 4794
rect 3943 4774 3978 4782
rect 3943 4773 3972 4774
rect 3663 4760 3877 4764
rect 3678 4758 3877 4760
rect 3912 4760 3925 4770
rect 3943 4760 3960 4773
rect 3912 4758 3960 4760
rect 3554 4754 3587 4758
rect 3550 4752 3587 4754
rect 3550 4751 3617 4752
rect 3550 4746 3581 4751
rect 3587 4746 3617 4751
rect 3550 4742 3617 4746
rect 3523 4739 3617 4742
rect 3523 4732 3572 4739
rect 3523 4726 3553 4732
rect 3572 4727 3577 4732
rect 3489 4710 3569 4726
rect 3581 4718 3617 4739
rect 3678 4734 3867 4758
rect 3912 4757 3959 4758
rect 3925 4752 3959 4757
rect 3693 4731 3867 4734
rect 3686 4728 3867 4731
rect 3895 4751 3959 4752
rect 3489 4708 3508 4710
rect 3523 4708 3557 4710
rect 3489 4692 3569 4708
rect 3489 4686 3508 4692
rect 3205 4660 3308 4670
rect 3159 4658 3308 4660
rect 3329 4658 3364 4670
rect 2998 4656 3160 4658
rect 3010 4636 3029 4656
rect 3044 4654 3074 4656
rect 2893 4628 2934 4636
rect 3016 4632 3029 4636
rect 3081 4640 3160 4656
rect 3192 4656 3364 4658
rect 3192 4640 3271 4656
rect 3278 4654 3308 4656
rect 2856 4618 2885 4628
rect 2899 4618 2928 4628
rect 2943 4618 2973 4632
rect 3016 4618 3059 4632
rect 3081 4628 3271 4640
rect 3336 4636 3342 4656
rect 3066 4618 3096 4628
rect 3097 4618 3255 4628
rect 3259 4618 3289 4628
rect 3293 4618 3323 4632
rect 3351 4618 3364 4656
rect 3436 4670 3465 4686
rect 3479 4670 3508 4686
rect 3523 4676 3553 4692
rect 3581 4670 3587 4718
rect 3590 4712 3609 4718
rect 3624 4712 3654 4720
rect 3590 4704 3654 4712
rect 3590 4688 3670 4704
rect 3686 4697 3748 4728
rect 3764 4697 3826 4728
rect 3895 4726 3944 4751
rect 3959 4726 3989 4742
rect 3858 4712 3888 4720
rect 3895 4718 4005 4726
rect 3858 4704 3903 4712
rect 3590 4686 3609 4688
rect 3624 4686 3670 4688
rect 3590 4670 3670 4686
rect 3697 4684 3732 4697
rect 3773 4694 3810 4697
rect 3773 4692 3815 4694
rect 3702 4681 3732 4684
rect 3711 4677 3718 4681
rect 3718 4676 3719 4677
rect 3677 4670 3687 4676
rect 3436 4662 3471 4670
rect 3436 4636 3437 4662
rect 3444 4636 3471 4662
rect 3379 4618 3409 4632
rect 3436 4628 3471 4636
rect 3473 4662 3514 4670
rect 3473 4636 3488 4662
rect 3495 4636 3514 4662
rect 3578 4658 3609 4670
rect 3624 4658 3727 4670
rect 3739 4660 3765 4686
rect 3780 4681 3810 4692
rect 3842 4688 3904 4704
rect 3842 4686 3888 4688
rect 3842 4670 3904 4686
rect 3916 4670 3922 4718
rect 3925 4710 4005 4718
rect 3925 4708 3944 4710
rect 3959 4708 3993 4710
rect 3925 4692 4005 4708
rect 3925 4670 3944 4692
rect 3959 4676 3989 4692
rect 4017 4686 4023 4760
rect 4026 4686 4045 4830
rect 4060 4686 4066 4830
rect 4075 4760 4088 4830
rect 4140 4826 4162 4830
rect 4133 4804 4162 4818
rect 4215 4804 4231 4818
rect 4269 4814 4275 4816
rect 4282 4814 4390 4830
rect 4397 4814 4403 4816
rect 4411 4814 4426 4830
rect 4492 4824 4511 4827
rect 4133 4802 4231 4804
rect 4258 4802 4426 4814
rect 4441 4804 4457 4818
rect 4492 4805 4514 4824
rect 4524 4818 4540 4819
rect 4523 4816 4540 4818
rect 4524 4811 4540 4816
rect 4514 4804 4520 4805
rect 4523 4804 4552 4811
rect 4441 4803 4552 4804
rect 4441 4802 4558 4803
rect 4117 4794 4168 4802
rect 4215 4794 4249 4802
rect 4117 4782 4142 4794
rect 4149 4782 4168 4794
rect 4222 4792 4249 4794
rect 4258 4792 4479 4802
rect 4514 4799 4520 4802
rect 4222 4788 4479 4792
rect 4117 4774 4168 4782
rect 4215 4774 4479 4788
rect 4523 4794 4558 4802
rect 4069 4726 4088 4760
rect 4133 4766 4162 4774
rect 4133 4760 4150 4766
rect 4133 4758 4167 4760
rect 4215 4758 4231 4774
rect 4232 4764 4440 4774
rect 4441 4764 4457 4774
rect 4505 4770 4520 4785
rect 4523 4782 4524 4794
rect 4531 4782 4558 4794
rect 4523 4774 4558 4782
rect 4523 4773 4552 4774
rect 4243 4760 4457 4764
rect 4258 4758 4457 4760
rect 4492 4760 4505 4770
rect 4523 4760 4540 4773
rect 4492 4758 4540 4760
rect 4134 4754 4167 4758
rect 4130 4752 4167 4754
rect 4130 4751 4197 4752
rect 4130 4746 4161 4751
rect 4167 4746 4197 4751
rect 4130 4742 4197 4746
rect 4103 4739 4197 4742
rect 4103 4732 4152 4739
rect 4103 4726 4133 4732
rect 4152 4727 4157 4732
rect 4069 4710 4149 4726
rect 4161 4718 4197 4739
rect 4258 4734 4447 4758
rect 4492 4757 4539 4758
rect 4505 4752 4539 4757
rect 4273 4731 4447 4734
rect 4266 4728 4447 4731
rect 4475 4751 4539 4752
rect 4069 4708 4088 4710
rect 4103 4708 4137 4710
rect 4069 4692 4149 4708
rect 4069 4686 4088 4692
rect 3785 4660 3888 4670
rect 3739 4658 3888 4660
rect 3909 4658 3944 4670
rect 3578 4656 3740 4658
rect 3590 4636 3609 4656
rect 3624 4654 3654 4656
rect 3473 4628 3514 4636
rect 3596 4632 3609 4636
rect 3661 4640 3740 4656
rect 3772 4656 3944 4658
rect 3772 4640 3851 4656
rect 3858 4654 3888 4656
rect 3436 4618 3465 4628
rect 3479 4618 3508 4628
rect 3523 4618 3553 4632
rect 3596 4618 3639 4632
rect 3661 4628 3851 4640
rect 3916 4636 3922 4656
rect 3646 4618 3676 4628
rect 3677 4618 3835 4628
rect 3839 4618 3869 4628
rect 3873 4618 3903 4632
rect 3931 4618 3944 4656
rect 4016 4670 4045 4686
rect 4059 4670 4088 4686
rect 4103 4676 4133 4692
rect 4161 4670 4167 4718
rect 4170 4712 4189 4718
rect 4204 4712 4234 4720
rect 4170 4704 4234 4712
rect 4170 4688 4250 4704
rect 4266 4697 4328 4728
rect 4344 4697 4406 4728
rect 4475 4726 4524 4751
rect 4539 4726 4569 4742
rect 4438 4712 4468 4720
rect 4475 4718 4585 4726
rect 4438 4704 4483 4712
rect 4170 4686 4189 4688
rect 4204 4686 4250 4688
rect 4170 4670 4250 4686
rect 4277 4684 4312 4697
rect 4353 4694 4390 4697
rect 4353 4692 4395 4694
rect 4282 4681 4312 4684
rect 4291 4677 4298 4681
rect 4298 4676 4299 4677
rect 4257 4670 4267 4676
rect 4016 4662 4051 4670
rect 4016 4636 4017 4662
rect 4024 4636 4051 4662
rect 3959 4618 3989 4632
rect 4016 4628 4051 4636
rect 4053 4662 4094 4670
rect 4053 4636 4068 4662
rect 4075 4636 4094 4662
rect 4158 4658 4189 4670
rect 4204 4658 4307 4670
rect 4319 4660 4345 4686
rect 4360 4681 4390 4692
rect 4422 4688 4484 4704
rect 4422 4686 4468 4688
rect 4422 4670 4484 4686
rect 4496 4670 4502 4718
rect 4505 4710 4585 4718
rect 4505 4708 4524 4710
rect 4539 4708 4573 4710
rect 4505 4692 4585 4708
rect 4505 4670 4524 4692
rect 4539 4676 4569 4692
rect 4597 4686 4603 4760
rect 4606 4686 4625 4830
rect 4640 4686 4646 4830
rect 4655 4760 4668 4830
rect 4720 4826 4742 4830
rect 4713 4804 4742 4818
rect 4795 4804 4811 4818
rect 4849 4814 4855 4816
rect 4862 4814 4970 4830
rect 4977 4814 4983 4816
rect 4991 4814 5006 4830
rect 5072 4824 5091 4827
rect 4713 4802 4811 4804
rect 4838 4802 5006 4814
rect 5021 4804 5037 4818
rect 5072 4805 5094 4824
rect 5104 4818 5120 4819
rect 5103 4816 5120 4818
rect 5104 4811 5120 4816
rect 5094 4804 5100 4805
rect 5103 4804 5132 4811
rect 5021 4803 5132 4804
rect 5021 4802 5138 4803
rect 4697 4794 4748 4802
rect 4795 4794 4829 4802
rect 4697 4782 4722 4794
rect 4729 4782 4748 4794
rect 4802 4792 4829 4794
rect 4838 4792 5059 4802
rect 5094 4799 5100 4802
rect 4802 4788 5059 4792
rect 4697 4774 4748 4782
rect 4795 4774 5059 4788
rect 5103 4794 5138 4802
rect 4649 4726 4668 4760
rect 4713 4766 4742 4774
rect 4713 4760 4730 4766
rect 4713 4758 4747 4760
rect 4795 4758 4811 4774
rect 4812 4764 5020 4774
rect 5021 4764 5037 4774
rect 5085 4770 5100 4785
rect 5103 4782 5104 4794
rect 5111 4782 5138 4794
rect 5103 4774 5138 4782
rect 5103 4773 5132 4774
rect 4823 4760 5037 4764
rect 4838 4758 5037 4760
rect 5072 4760 5085 4770
rect 5103 4760 5120 4773
rect 5072 4758 5120 4760
rect 4714 4754 4747 4758
rect 4710 4752 4747 4754
rect 4710 4751 4777 4752
rect 4710 4746 4741 4751
rect 4747 4746 4777 4751
rect 4710 4742 4777 4746
rect 4683 4739 4777 4742
rect 4683 4732 4732 4739
rect 4683 4726 4713 4732
rect 4732 4727 4737 4732
rect 4649 4710 4729 4726
rect 4741 4718 4777 4739
rect 4838 4734 5027 4758
rect 5072 4757 5119 4758
rect 5085 4752 5119 4757
rect 4853 4731 5027 4734
rect 4846 4728 5027 4731
rect 5055 4751 5119 4752
rect 4649 4708 4668 4710
rect 4683 4708 4717 4710
rect 4649 4692 4729 4708
rect 4649 4686 4668 4692
rect 4365 4660 4468 4670
rect 4319 4658 4468 4660
rect 4489 4658 4524 4670
rect 4158 4656 4320 4658
rect 4170 4636 4189 4656
rect 4204 4654 4234 4656
rect 4053 4628 4094 4636
rect 4176 4632 4189 4636
rect 4241 4640 4320 4656
rect 4352 4656 4524 4658
rect 4352 4640 4431 4656
rect 4438 4654 4468 4656
rect 4016 4618 4045 4628
rect 4059 4618 4088 4628
rect 4103 4618 4133 4632
rect 4176 4618 4219 4632
rect 4241 4628 4431 4640
rect 4496 4636 4502 4656
rect 4226 4618 4256 4628
rect 4257 4618 4415 4628
rect 4419 4618 4449 4628
rect 4453 4618 4483 4632
rect 4511 4618 4524 4656
rect 4596 4670 4625 4686
rect 4639 4670 4668 4686
rect 4683 4676 4713 4692
rect 4741 4670 4747 4718
rect 4750 4712 4769 4718
rect 4784 4712 4814 4720
rect 4750 4704 4814 4712
rect 4750 4688 4830 4704
rect 4846 4697 4908 4728
rect 4924 4697 4986 4728
rect 5055 4726 5104 4751
rect 5119 4726 5149 4742
rect 5018 4712 5048 4720
rect 5055 4718 5165 4726
rect 5018 4704 5063 4712
rect 4750 4686 4769 4688
rect 4784 4686 4830 4688
rect 4750 4670 4830 4686
rect 4857 4684 4892 4697
rect 4933 4694 4970 4697
rect 4933 4692 4975 4694
rect 4862 4681 4892 4684
rect 4871 4677 4878 4681
rect 4878 4676 4879 4677
rect 4837 4670 4847 4676
rect 4596 4662 4631 4670
rect 4596 4636 4597 4662
rect 4604 4636 4631 4662
rect 4539 4618 4569 4632
rect 4596 4628 4631 4636
rect 4633 4662 4674 4670
rect 4633 4636 4648 4662
rect 4655 4636 4674 4662
rect 4738 4658 4769 4670
rect 4784 4658 4887 4670
rect 4899 4660 4925 4686
rect 4940 4681 4970 4692
rect 5002 4688 5064 4704
rect 5002 4686 5048 4688
rect 5002 4670 5064 4686
rect 5076 4670 5082 4718
rect 5085 4710 5165 4718
rect 5085 4708 5104 4710
rect 5119 4708 5153 4710
rect 5085 4692 5165 4708
rect 5085 4670 5104 4692
rect 5119 4676 5149 4692
rect 5177 4686 5183 4760
rect 5186 4686 5205 4830
rect 5220 4686 5226 4830
rect 5235 4760 5248 4830
rect 5300 4826 5322 4830
rect 5293 4804 5322 4818
rect 5375 4804 5391 4818
rect 5429 4814 5435 4816
rect 5442 4814 5550 4830
rect 5557 4814 5563 4816
rect 5571 4814 5586 4830
rect 5652 4824 5671 4827
rect 5293 4802 5391 4804
rect 5418 4802 5586 4814
rect 5601 4804 5617 4818
rect 5652 4805 5674 4824
rect 5684 4818 5700 4819
rect 5683 4816 5700 4818
rect 5684 4811 5700 4816
rect 5674 4804 5680 4805
rect 5683 4804 5712 4811
rect 5601 4803 5712 4804
rect 5601 4802 5718 4803
rect 5277 4794 5328 4802
rect 5375 4794 5409 4802
rect 5277 4782 5302 4794
rect 5309 4782 5328 4794
rect 5382 4792 5409 4794
rect 5418 4792 5639 4802
rect 5674 4799 5680 4802
rect 5382 4788 5639 4792
rect 5277 4774 5328 4782
rect 5375 4774 5639 4788
rect 5683 4794 5718 4802
rect 5229 4726 5248 4760
rect 5293 4766 5322 4774
rect 5293 4760 5310 4766
rect 5293 4758 5327 4760
rect 5375 4758 5391 4774
rect 5392 4764 5600 4774
rect 5601 4764 5617 4774
rect 5665 4770 5680 4785
rect 5683 4782 5684 4794
rect 5691 4782 5718 4794
rect 5683 4774 5718 4782
rect 5683 4773 5712 4774
rect 5403 4760 5617 4764
rect 5418 4758 5617 4760
rect 5652 4760 5665 4770
rect 5683 4760 5700 4773
rect 5652 4758 5700 4760
rect 5294 4754 5327 4758
rect 5290 4752 5327 4754
rect 5290 4751 5357 4752
rect 5290 4746 5321 4751
rect 5327 4746 5357 4751
rect 5290 4742 5357 4746
rect 5263 4739 5357 4742
rect 5263 4732 5312 4739
rect 5263 4726 5293 4732
rect 5312 4727 5317 4732
rect 5229 4710 5309 4726
rect 5321 4718 5357 4739
rect 5418 4734 5607 4758
rect 5652 4757 5699 4758
rect 5665 4752 5699 4757
rect 5433 4731 5607 4734
rect 5426 4728 5607 4731
rect 5635 4751 5699 4752
rect 5229 4708 5248 4710
rect 5263 4708 5297 4710
rect 5229 4692 5309 4708
rect 5229 4686 5248 4692
rect 4945 4660 5048 4670
rect 4899 4658 5048 4660
rect 5069 4658 5104 4670
rect 4738 4656 4900 4658
rect 4750 4636 4769 4656
rect 4784 4654 4814 4656
rect 4633 4628 4674 4636
rect 4756 4632 4769 4636
rect 4821 4640 4900 4656
rect 4932 4656 5104 4658
rect 4932 4640 5011 4656
rect 5018 4654 5048 4656
rect 4596 4618 4625 4628
rect 4639 4618 4668 4628
rect 4683 4618 4713 4632
rect 4756 4618 4799 4632
rect 4821 4628 5011 4640
rect 5076 4636 5082 4656
rect 4806 4618 4836 4628
rect 4837 4618 4995 4628
rect 4999 4618 5029 4628
rect 5033 4618 5063 4632
rect 5091 4618 5104 4656
rect 5176 4670 5205 4686
rect 5219 4670 5248 4686
rect 5263 4676 5293 4692
rect 5321 4670 5327 4718
rect 5330 4712 5349 4718
rect 5364 4712 5394 4720
rect 5330 4704 5394 4712
rect 5330 4688 5410 4704
rect 5426 4697 5488 4728
rect 5504 4697 5566 4728
rect 5635 4726 5684 4751
rect 5699 4726 5729 4742
rect 5598 4712 5628 4720
rect 5635 4718 5745 4726
rect 5598 4704 5643 4712
rect 5330 4686 5349 4688
rect 5364 4686 5410 4688
rect 5330 4670 5410 4686
rect 5437 4684 5472 4697
rect 5513 4694 5550 4697
rect 5513 4692 5555 4694
rect 5442 4681 5472 4684
rect 5451 4677 5458 4681
rect 5458 4676 5459 4677
rect 5417 4670 5427 4676
rect 5176 4662 5211 4670
rect 5176 4636 5177 4662
rect 5184 4636 5211 4662
rect 5119 4618 5149 4632
rect 5176 4628 5211 4636
rect 5213 4662 5254 4670
rect 5213 4636 5228 4662
rect 5235 4636 5254 4662
rect 5318 4658 5349 4670
rect 5364 4658 5467 4670
rect 5479 4660 5505 4686
rect 5520 4681 5550 4692
rect 5582 4688 5644 4704
rect 5582 4686 5628 4688
rect 5582 4670 5644 4686
rect 5656 4670 5662 4718
rect 5665 4710 5745 4718
rect 5665 4708 5684 4710
rect 5699 4708 5733 4710
rect 5665 4692 5745 4708
rect 5665 4670 5684 4692
rect 5699 4676 5729 4692
rect 5757 4686 5763 4760
rect 5766 4686 5785 4830
rect 5800 4686 5806 4830
rect 5815 4760 5828 4830
rect 5880 4826 5902 4830
rect 5873 4804 5902 4818
rect 5955 4804 5971 4818
rect 6009 4814 6015 4816
rect 6022 4814 6130 4830
rect 6137 4814 6143 4816
rect 6151 4814 6166 4830
rect 6232 4824 6251 4827
rect 5873 4802 5971 4804
rect 5998 4802 6166 4814
rect 6181 4804 6197 4818
rect 6232 4805 6254 4824
rect 6264 4818 6280 4819
rect 6263 4816 6280 4818
rect 6264 4811 6280 4816
rect 6254 4804 6260 4805
rect 6263 4804 6292 4811
rect 6181 4803 6292 4804
rect 6181 4802 6298 4803
rect 5857 4794 5908 4802
rect 5955 4794 5989 4802
rect 5857 4782 5882 4794
rect 5889 4782 5908 4794
rect 5962 4792 5989 4794
rect 5998 4792 6219 4802
rect 6254 4799 6260 4802
rect 5962 4788 6219 4792
rect 5857 4774 5908 4782
rect 5955 4774 6219 4788
rect 6263 4794 6298 4802
rect 5809 4726 5828 4760
rect 5873 4766 5902 4774
rect 5873 4760 5890 4766
rect 5873 4758 5907 4760
rect 5955 4758 5971 4774
rect 5972 4764 6180 4774
rect 6181 4764 6197 4774
rect 6245 4770 6260 4785
rect 6263 4782 6264 4794
rect 6271 4782 6298 4794
rect 6263 4774 6298 4782
rect 6263 4773 6292 4774
rect 5983 4760 6197 4764
rect 5998 4758 6197 4760
rect 6232 4760 6245 4770
rect 6263 4760 6280 4773
rect 6232 4758 6280 4760
rect 5874 4754 5907 4758
rect 5870 4752 5907 4754
rect 5870 4751 5937 4752
rect 5870 4746 5901 4751
rect 5907 4746 5937 4751
rect 5870 4742 5937 4746
rect 5843 4739 5937 4742
rect 5843 4732 5892 4739
rect 5843 4726 5873 4732
rect 5892 4727 5897 4732
rect 5809 4710 5889 4726
rect 5901 4718 5937 4739
rect 5998 4734 6187 4758
rect 6232 4757 6279 4758
rect 6245 4752 6279 4757
rect 6013 4731 6187 4734
rect 6006 4728 6187 4731
rect 6215 4751 6279 4752
rect 5809 4708 5828 4710
rect 5843 4708 5877 4710
rect 5809 4692 5889 4708
rect 5809 4686 5828 4692
rect 5525 4660 5628 4670
rect 5479 4658 5628 4660
rect 5649 4658 5684 4670
rect 5318 4656 5480 4658
rect 5330 4636 5349 4656
rect 5364 4654 5394 4656
rect 5213 4628 5254 4636
rect 5336 4632 5349 4636
rect 5401 4640 5480 4656
rect 5512 4656 5684 4658
rect 5512 4640 5591 4656
rect 5598 4654 5628 4656
rect 5176 4618 5205 4628
rect 5219 4618 5248 4628
rect 5263 4618 5293 4632
rect 5336 4618 5379 4632
rect 5401 4628 5591 4640
rect 5656 4636 5662 4656
rect 5386 4618 5416 4628
rect 5417 4618 5575 4628
rect 5579 4618 5609 4628
rect 5613 4618 5643 4632
rect 5671 4618 5684 4656
rect 5756 4670 5785 4686
rect 5799 4670 5828 4686
rect 5843 4676 5873 4692
rect 5901 4670 5907 4718
rect 5910 4712 5929 4718
rect 5944 4712 5974 4720
rect 5910 4704 5974 4712
rect 5910 4688 5990 4704
rect 6006 4697 6068 4728
rect 6084 4697 6146 4728
rect 6215 4726 6264 4751
rect 6279 4726 6309 4742
rect 6178 4712 6208 4720
rect 6215 4718 6325 4726
rect 6178 4704 6223 4712
rect 5910 4686 5929 4688
rect 5944 4686 5990 4688
rect 5910 4670 5990 4686
rect 6017 4684 6052 4697
rect 6093 4694 6130 4697
rect 6093 4692 6135 4694
rect 6022 4681 6052 4684
rect 6031 4677 6038 4681
rect 6038 4676 6039 4677
rect 5997 4670 6007 4676
rect 5756 4662 5791 4670
rect 5756 4636 5757 4662
rect 5764 4636 5791 4662
rect 5699 4618 5729 4632
rect 5756 4628 5791 4636
rect 5793 4662 5834 4670
rect 5793 4636 5808 4662
rect 5815 4636 5834 4662
rect 5898 4658 5929 4670
rect 5944 4658 6047 4670
rect 6059 4660 6085 4686
rect 6100 4681 6130 4692
rect 6162 4688 6224 4704
rect 6162 4686 6208 4688
rect 6162 4670 6224 4686
rect 6236 4670 6242 4718
rect 6245 4710 6325 4718
rect 6245 4708 6264 4710
rect 6279 4708 6313 4710
rect 6245 4692 6325 4708
rect 6245 4670 6264 4692
rect 6279 4676 6309 4692
rect 6337 4686 6343 4760
rect 6346 4686 6365 4830
rect 6380 4686 6386 4830
rect 6395 4760 6408 4830
rect 6460 4826 6482 4830
rect 6453 4804 6482 4818
rect 6535 4804 6551 4818
rect 6589 4814 6595 4816
rect 6602 4814 6710 4830
rect 6717 4814 6723 4816
rect 6731 4814 6746 4830
rect 6812 4824 6831 4827
rect 6453 4802 6551 4804
rect 6578 4802 6746 4814
rect 6761 4804 6777 4818
rect 6812 4805 6834 4824
rect 6844 4818 6860 4819
rect 6843 4816 6860 4818
rect 6844 4811 6860 4816
rect 6834 4804 6840 4805
rect 6843 4804 6872 4811
rect 6761 4803 6872 4804
rect 6761 4802 6878 4803
rect 6437 4794 6488 4802
rect 6535 4794 6569 4802
rect 6437 4782 6462 4794
rect 6469 4782 6488 4794
rect 6542 4792 6569 4794
rect 6578 4792 6799 4802
rect 6834 4799 6840 4802
rect 6542 4788 6799 4792
rect 6437 4774 6488 4782
rect 6535 4774 6799 4788
rect 6843 4794 6878 4802
rect 6389 4726 6408 4760
rect 6453 4766 6482 4774
rect 6453 4760 6470 4766
rect 6453 4758 6487 4760
rect 6535 4758 6551 4774
rect 6552 4764 6760 4774
rect 6761 4764 6777 4774
rect 6825 4770 6840 4785
rect 6843 4782 6844 4794
rect 6851 4782 6878 4794
rect 6843 4774 6878 4782
rect 6843 4773 6872 4774
rect 6563 4760 6777 4764
rect 6578 4758 6777 4760
rect 6812 4760 6825 4770
rect 6843 4760 6860 4773
rect 6812 4758 6860 4760
rect 6454 4754 6487 4758
rect 6450 4752 6487 4754
rect 6450 4751 6517 4752
rect 6450 4746 6481 4751
rect 6487 4746 6517 4751
rect 6450 4742 6517 4746
rect 6423 4739 6517 4742
rect 6423 4732 6472 4739
rect 6423 4726 6453 4732
rect 6472 4727 6477 4732
rect 6389 4710 6469 4726
rect 6481 4718 6517 4739
rect 6578 4734 6767 4758
rect 6812 4757 6859 4758
rect 6825 4752 6859 4757
rect 6593 4731 6767 4734
rect 6586 4728 6767 4731
rect 6795 4751 6859 4752
rect 6389 4708 6408 4710
rect 6423 4708 6457 4710
rect 6389 4692 6469 4708
rect 6389 4686 6408 4692
rect 6105 4660 6208 4670
rect 6059 4658 6208 4660
rect 6229 4658 6264 4670
rect 5898 4656 6060 4658
rect 5910 4636 5929 4656
rect 5944 4654 5974 4656
rect 5793 4628 5834 4636
rect 5916 4632 5929 4636
rect 5981 4640 6060 4656
rect 6092 4656 6264 4658
rect 6092 4640 6171 4656
rect 6178 4654 6208 4656
rect 5756 4618 5785 4628
rect 5799 4618 5828 4628
rect 5843 4618 5873 4632
rect 5916 4618 5959 4632
rect 5981 4628 6171 4640
rect 6236 4636 6242 4656
rect 5966 4618 5996 4628
rect 5997 4618 6155 4628
rect 6159 4618 6189 4628
rect 6193 4618 6223 4632
rect 6251 4618 6264 4656
rect 6336 4670 6365 4686
rect 6379 4670 6408 4686
rect 6423 4676 6453 4692
rect 6481 4670 6487 4718
rect 6490 4712 6509 4718
rect 6524 4712 6554 4720
rect 6490 4704 6554 4712
rect 6490 4688 6570 4704
rect 6586 4697 6648 4728
rect 6664 4697 6726 4728
rect 6795 4726 6844 4751
rect 6859 4726 6889 4742
rect 6758 4712 6788 4720
rect 6795 4718 6905 4726
rect 6758 4704 6803 4712
rect 6490 4686 6509 4688
rect 6524 4686 6570 4688
rect 6490 4670 6570 4686
rect 6597 4684 6632 4697
rect 6673 4694 6710 4697
rect 6673 4692 6715 4694
rect 6602 4681 6632 4684
rect 6611 4677 6618 4681
rect 6618 4676 6619 4677
rect 6577 4670 6587 4676
rect 6336 4662 6371 4670
rect 6336 4636 6337 4662
rect 6344 4636 6371 4662
rect 6279 4618 6309 4632
rect 6336 4628 6371 4636
rect 6373 4662 6414 4670
rect 6373 4636 6388 4662
rect 6395 4636 6414 4662
rect 6478 4658 6509 4670
rect 6524 4658 6627 4670
rect 6639 4660 6665 4686
rect 6680 4681 6710 4692
rect 6742 4688 6804 4704
rect 6742 4686 6788 4688
rect 6742 4670 6804 4686
rect 6816 4670 6822 4718
rect 6825 4710 6905 4718
rect 6825 4708 6844 4710
rect 6859 4708 6893 4710
rect 6825 4692 6905 4708
rect 6825 4670 6844 4692
rect 6859 4676 6889 4692
rect 6917 4686 6923 4760
rect 6926 4686 6945 4830
rect 6960 4686 6966 4830
rect 6975 4760 6988 4830
rect 7040 4826 7062 4830
rect 7033 4804 7062 4818
rect 7115 4804 7131 4818
rect 7169 4814 7175 4816
rect 7182 4814 7290 4830
rect 7297 4814 7303 4816
rect 7311 4814 7326 4830
rect 7392 4824 7411 4827
rect 7033 4802 7131 4804
rect 7158 4802 7326 4814
rect 7341 4804 7357 4818
rect 7392 4805 7414 4824
rect 7424 4818 7440 4819
rect 7423 4816 7440 4818
rect 7424 4811 7440 4816
rect 7414 4804 7420 4805
rect 7423 4804 7452 4811
rect 7341 4803 7452 4804
rect 7341 4802 7458 4803
rect 7017 4794 7068 4802
rect 7115 4794 7149 4802
rect 7017 4782 7042 4794
rect 7049 4782 7068 4794
rect 7122 4792 7149 4794
rect 7158 4792 7379 4802
rect 7414 4799 7420 4802
rect 7122 4788 7379 4792
rect 7017 4774 7068 4782
rect 7115 4774 7379 4788
rect 7423 4794 7458 4802
rect 6969 4726 6988 4760
rect 7033 4766 7062 4774
rect 7033 4760 7050 4766
rect 7033 4758 7067 4760
rect 7115 4758 7131 4774
rect 7132 4764 7340 4774
rect 7341 4764 7357 4774
rect 7405 4770 7420 4785
rect 7423 4782 7424 4794
rect 7431 4782 7458 4794
rect 7423 4774 7458 4782
rect 7423 4773 7452 4774
rect 7143 4760 7357 4764
rect 7158 4758 7357 4760
rect 7392 4760 7405 4770
rect 7423 4760 7440 4773
rect 7392 4758 7440 4760
rect 7034 4754 7067 4758
rect 7030 4752 7067 4754
rect 7030 4751 7097 4752
rect 7030 4746 7061 4751
rect 7067 4746 7097 4751
rect 7030 4742 7097 4746
rect 7003 4739 7097 4742
rect 7003 4732 7052 4739
rect 7003 4726 7033 4732
rect 7052 4727 7057 4732
rect 6969 4710 7049 4726
rect 7061 4718 7097 4739
rect 7158 4734 7347 4758
rect 7392 4757 7439 4758
rect 7405 4752 7439 4757
rect 7173 4731 7347 4734
rect 7166 4728 7347 4731
rect 7375 4751 7439 4752
rect 6969 4708 6988 4710
rect 7003 4708 7037 4710
rect 6969 4692 7049 4708
rect 6969 4686 6988 4692
rect 6685 4660 6788 4670
rect 6639 4658 6788 4660
rect 6809 4658 6844 4670
rect 6478 4656 6640 4658
rect 6490 4636 6509 4656
rect 6524 4654 6554 4656
rect 6373 4628 6414 4636
rect 6496 4632 6509 4636
rect 6561 4640 6640 4656
rect 6672 4656 6844 4658
rect 6672 4640 6751 4656
rect 6758 4654 6788 4656
rect 6336 4618 6365 4628
rect 6379 4618 6408 4628
rect 6423 4618 6453 4632
rect 6496 4618 6539 4632
rect 6561 4628 6751 4640
rect 6816 4636 6822 4656
rect 6546 4618 6576 4628
rect 6577 4618 6735 4628
rect 6739 4618 6769 4628
rect 6773 4618 6803 4632
rect 6831 4618 6844 4656
rect 6916 4670 6945 4686
rect 6959 4670 6988 4686
rect 7003 4676 7033 4692
rect 7061 4670 7067 4718
rect 7070 4712 7089 4718
rect 7104 4712 7134 4720
rect 7070 4704 7134 4712
rect 7070 4688 7150 4704
rect 7166 4697 7228 4728
rect 7244 4697 7306 4728
rect 7375 4726 7424 4751
rect 7439 4726 7469 4742
rect 7338 4712 7368 4720
rect 7375 4718 7485 4726
rect 7338 4704 7383 4712
rect 7070 4686 7089 4688
rect 7104 4686 7150 4688
rect 7070 4670 7150 4686
rect 7177 4684 7212 4697
rect 7253 4694 7290 4697
rect 7253 4692 7295 4694
rect 7182 4681 7212 4684
rect 7191 4677 7198 4681
rect 7198 4676 7199 4677
rect 7157 4670 7167 4676
rect 6916 4662 6951 4670
rect 6916 4636 6917 4662
rect 6924 4636 6951 4662
rect 6859 4618 6889 4632
rect 6916 4628 6951 4636
rect 6953 4662 6994 4670
rect 6953 4636 6968 4662
rect 6975 4636 6994 4662
rect 7058 4658 7089 4670
rect 7104 4658 7207 4670
rect 7219 4660 7245 4686
rect 7260 4681 7290 4692
rect 7322 4688 7384 4704
rect 7322 4686 7368 4688
rect 7322 4670 7384 4686
rect 7396 4670 7402 4718
rect 7405 4710 7485 4718
rect 7405 4708 7424 4710
rect 7439 4708 7473 4710
rect 7405 4692 7485 4708
rect 7405 4670 7424 4692
rect 7439 4676 7469 4692
rect 7497 4686 7503 4760
rect 7506 4686 7525 4830
rect 7540 4686 7546 4830
rect 7555 4760 7568 4830
rect 7620 4826 7642 4830
rect 7613 4804 7642 4818
rect 7695 4804 7711 4818
rect 7749 4814 7755 4816
rect 7762 4814 7870 4830
rect 7877 4814 7883 4816
rect 7891 4814 7906 4830
rect 7972 4824 7991 4827
rect 7613 4802 7711 4804
rect 7738 4802 7906 4814
rect 7921 4804 7937 4818
rect 7972 4805 7994 4824
rect 8004 4818 8020 4819
rect 8003 4816 8020 4818
rect 8004 4811 8020 4816
rect 7994 4804 8000 4805
rect 8003 4804 8032 4811
rect 7921 4803 8032 4804
rect 7921 4802 8038 4803
rect 7597 4794 7648 4802
rect 7695 4794 7729 4802
rect 7597 4782 7622 4794
rect 7629 4782 7648 4794
rect 7702 4792 7729 4794
rect 7738 4792 7959 4802
rect 7994 4799 8000 4802
rect 7702 4788 7959 4792
rect 7597 4774 7648 4782
rect 7695 4774 7959 4788
rect 8003 4794 8038 4802
rect 7549 4726 7568 4760
rect 7613 4766 7642 4774
rect 7613 4760 7630 4766
rect 7613 4758 7647 4760
rect 7695 4758 7711 4774
rect 7712 4764 7920 4774
rect 7921 4764 7937 4774
rect 7985 4770 8000 4785
rect 8003 4782 8004 4794
rect 8011 4782 8038 4794
rect 8003 4774 8038 4782
rect 8003 4773 8032 4774
rect 7723 4760 7937 4764
rect 7738 4758 7937 4760
rect 7972 4760 7985 4770
rect 8003 4760 8020 4773
rect 7972 4758 8020 4760
rect 7614 4754 7647 4758
rect 7610 4752 7647 4754
rect 7610 4751 7677 4752
rect 7610 4746 7641 4751
rect 7647 4746 7677 4751
rect 7610 4742 7677 4746
rect 7583 4739 7677 4742
rect 7583 4732 7632 4739
rect 7583 4726 7613 4732
rect 7632 4727 7637 4732
rect 7549 4710 7629 4726
rect 7641 4718 7677 4739
rect 7738 4734 7927 4758
rect 7972 4757 8019 4758
rect 7985 4752 8019 4757
rect 7753 4731 7927 4734
rect 7746 4728 7927 4731
rect 7955 4751 8019 4752
rect 7549 4708 7568 4710
rect 7583 4708 7617 4710
rect 7549 4692 7629 4708
rect 7549 4686 7568 4692
rect 7265 4660 7368 4670
rect 7219 4658 7368 4660
rect 7389 4658 7424 4670
rect 7058 4656 7220 4658
rect 7070 4636 7089 4656
rect 7104 4654 7134 4656
rect 6953 4628 6994 4636
rect 7076 4632 7089 4636
rect 7141 4640 7220 4656
rect 7252 4656 7424 4658
rect 7252 4640 7331 4656
rect 7338 4654 7368 4656
rect 6916 4618 6945 4628
rect 6959 4618 6988 4628
rect 7003 4618 7033 4632
rect 7076 4618 7119 4632
rect 7141 4628 7331 4640
rect 7396 4636 7402 4656
rect 7126 4618 7156 4628
rect 7157 4618 7315 4628
rect 7319 4618 7349 4628
rect 7353 4618 7383 4632
rect 7411 4618 7424 4656
rect 7496 4670 7525 4686
rect 7539 4670 7568 4686
rect 7583 4676 7613 4692
rect 7641 4670 7647 4718
rect 7650 4712 7669 4718
rect 7684 4712 7714 4720
rect 7650 4704 7714 4712
rect 7650 4688 7730 4704
rect 7746 4697 7808 4728
rect 7824 4697 7886 4728
rect 7955 4726 8004 4751
rect 8019 4726 8049 4742
rect 7918 4712 7948 4720
rect 7955 4718 8065 4726
rect 7918 4704 7963 4712
rect 7650 4686 7669 4688
rect 7684 4686 7730 4688
rect 7650 4670 7730 4686
rect 7757 4684 7792 4697
rect 7833 4694 7870 4697
rect 7833 4692 7875 4694
rect 7762 4681 7792 4684
rect 7771 4677 7778 4681
rect 7778 4676 7779 4677
rect 7737 4670 7747 4676
rect 7496 4662 7531 4670
rect 7496 4636 7497 4662
rect 7504 4636 7531 4662
rect 7439 4618 7469 4632
rect 7496 4628 7531 4636
rect 7533 4662 7574 4670
rect 7533 4636 7548 4662
rect 7555 4636 7574 4662
rect 7638 4658 7669 4670
rect 7684 4658 7787 4670
rect 7799 4660 7825 4686
rect 7840 4681 7870 4692
rect 7902 4688 7964 4704
rect 7902 4686 7948 4688
rect 7902 4670 7964 4686
rect 7976 4670 7982 4718
rect 7985 4710 8065 4718
rect 7985 4708 8004 4710
rect 8019 4708 8053 4710
rect 7985 4692 8065 4708
rect 7985 4670 8004 4692
rect 8019 4676 8049 4692
rect 8077 4686 8083 4760
rect 8086 4686 8105 4830
rect 8120 4686 8126 4830
rect 8135 4760 8148 4830
rect 8200 4826 8222 4830
rect 8193 4804 8222 4818
rect 8275 4804 8291 4818
rect 8329 4814 8335 4816
rect 8342 4814 8450 4830
rect 8457 4814 8463 4816
rect 8471 4814 8486 4830
rect 8552 4824 8571 4827
rect 8193 4802 8291 4804
rect 8318 4802 8486 4814
rect 8501 4804 8517 4818
rect 8552 4805 8574 4824
rect 8584 4818 8600 4819
rect 8583 4816 8600 4818
rect 8584 4811 8600 4816
rect 8574 4804 8580 4805
rect 8583 4804 8612 4811
rect 8501 4803 8612 4804
rect 8501 4802 8618 4803
rect 8177 4794 8228 4802
rect 8275 4794 8309 4802
rect 8177 4782 8202 4794
rect 8209 4782 8228 4794
rect 8282 4792 8309 4794
rect 8318 4792 8539 4802
rect 8574 4799 8580 4802
rect 8282 4788 8539 4792
rect 8177 4774 8228 4782
rect 8275 4774 8539 4788
rect 8583 4794 8618 4802
rect 8129 4726 8148 4760
rect 8193 4766 8222 4774
rect 8193 4760 8210 4766
rect 8193 4758 8227 4760
rect 8275 4758 8291 4774
rect 8292 4764 8500 4774
rect 8501 4764 8517 4774
rect 8565 4770 8580 4785
rect 8583 4782 8584 4794
rect 8591 4782 8618 4794
rect 8583 4774 8618 4782
rect 8583 4773 8612 4774
rect 8303 4760 8517 4764
rect 8318 4758 8517 4760
rect 8552 4760 8565 4770
rect 8583 4760 8600 4773
rect 8552 4758 8600 4760
rect 8194 4754 8227 4758
rect 8190 4752 8227 4754
rect 8190 4751 8257 4752
rect 8190 4746 8221 4751
rect 8227 4746 8257 4751
rect 8190 4742 8257 4746
rect 8163 4739 8257 4742
rect 8163 4732 8212 4739
rect 8163 4726 8193 4732
rect 8212 4727 8217 4732
rect 8129 4710 8209 4726
rect 8221 4718 8257 4739
rect 8318 4734 8507 4758
rect 8552 4757 8599 4758
rect 8565 4752 8599 4757
rect 8333 4731 8507 4734
rect 8326 4728 8507 4731
rect 8535 4751 8599 4752
rect 8129 4708 8148 4710
rect 8163 4708 8197 4710
rect 8129 4692 8209 4708
rect 8129 4686 8148 4692
rect 7845 4660 7948 4670
rect 7799 4658 7948 4660
rect 7969 4658 8004 4670
rect 7638 4656 7800 4658
rect 7650 4636 7669 4656
rect 7684 4654 7714 4656
rect 7533 4628 7574 4636
rect 7656 4632 7669 4636
rect 7721 4640 7800 4656
rect 7832 4656 8004 4658
rect 7832 4640 7911 4656
rect 7918 4654 7948 4656
rect 7496 4618 7525 4628
rect 7539 4618 7568 4628
rect 7583 4618 7613 4632
rect 7656 4618 7699 4632
rect 7721 4628 7911 4640
rect 7976 4636 7982 4656
rect 7706 4618 7736 4628
rect 7737 4618 7895 4628
rect 7899 4618 7929 4628
rect 7933 4618 7963 4632
rect 7991 4618 8004 4656
rect 8076 4670 8105 4686
rect 8119 4670 8148 4686
rect 8163 4676 8193 4692
rect 8221 4670 8227 4718
rect 8230 4712 8249 4718
rect 8264 4712 8294 4720
rect 8230 4704 8294 4712
rect 8230 4688 8310 4704
rect 8326 4697 8388 4728
rect 8404 4697 8466 4728
rect 8535 4726 8584 4751
rect 8599 4726 8629 4742
rect 8498 4712 8528 4720
rect 8535 4718 8645 4726
rect 8498 4704 8543 4712
rect 8230 4686 8249 4688
rect 8264 4686 8310 4688
rect 8230 4670 8310 4686
rect 8337 4684 8372 4697
rect 8413 4694 8450 4697
rect 8413 4692 8455 4694
rect 8342 4681 8372 4684
rect 8351 4677 8358 4681
rect 8358 4676 8359 4677
rect 8317 4670 8327 4676
rect 8076 4662 8111 4670
rect 8076 4636 8077 4662
rect 8084 4636 8111 4662
rect 8019 4618 8049 4632
rect 8076 4628 8111 4636
rect 8113 4662 8154 4670
rect 8113 4636 8128 4662
rect 8135 4636 8154 4662
rect 8218 4658 8249 4670
rect 8264 4658 8367 4670
rect 8379 4660 8405 4686
rect 8420 4681 8450 4692
rect 8482 4688 8544 4704
rect 8482 4686 8528 4688
rect 8482 4670 8544 4686
rect 8556 4670 8562 4718
rect 8565 4710 8645 4718
rect 8565 4708 8584 4710
rect 8599 4708 8633 4710
rect 8565 4692 8645 4708
rect 8565 4670 8584 4692
rect 8599 4676 8629 4692
rect 8657 4686 8663 4760
rect 8666 4686 8685 4830
rect 8700 4686 8706 4830
rect 8715 4760 8728 4830
rect 8780 4826 8802 4830
rect 8773 4804 8802 4818
rect 8855 4804 8871 4818
rect 8909 4814 8915 4816
rect 8922 4814 9030 4830
rect 9037 4814 9043 4816
rect 9051 4814 9066 4830
rect 9132 4824 9151 4827
rect 8773 4802 8871 4804
rect 8898 4802 9066 4814
rect 9081 4804 9097 4818
rect 9132 4805 9154 4824
rect 9164 4818 9180 4819
rect 9163 4816 9180 4818
rect 9164 4811 9180 4816
rect 9154 4804 9160 4805
rect 9163 4804 9192 4811
rect 9081 4803 9192 4804
rect 9081 4802 9198 4803
rect 8757 4794 8808 4802
rect 8855 4794 8889 4802
rect 8757 4782 8782 4794
rect 8789 4782 8808 4794
rect 8862 4792 8889 4794
rect 8898 4792 9119 4802
rect 9154 4799 9160 4802
rect 8862 4788 9119 4792
rect 8757 4774 8808 4782
rect 8855 4774 9119 4788
rect 9163 4794 9198 4802
rect 8709 4726 8728 4760
rect 8773 4766 8802 4774
rect 8773 4760 8790 4766
rect 8773 4758 8807 4760
rect 8855 4758 8871 4774
rect 8872 4764 9080 4774
rect 9081 4764 9097 4774
rect 9145 4770 9160 4785
rect 9163 4782 9164 4794
rect 9171 4782 9198 4794
rect 9163 4774 9198 4782
rect 9163 4773 9192 4774
rect 8883 4760 9097 4764
rect 8898 4758 9097 4760
rect 9132 4760 9145 4770
rect 9163 4760 9180 4773
rect 9132 4758 9180 4760
rect 8774 4754 8807 4758
rect 8770 4752 8807 4754
rect 8770 4751 8837 4752
rect 8770 4746 8801 4751
rect 8807 4746 8837 4751
rect 8770 4742 8837 4746
rect 8743 4739 8837 4742
rect 8743 4732 8792 4739
rect 8743 4726 8773 4732
rect 8792 4727 8797 4732
rect 8709 4710 8789 4726
rect 8801 4718 8837 4739
rect 8898 4734 9087 4758
rect 9132 4757 9179 4758
rect 9145 4752 9179 4757
rect 8913 4731 9087 4734
rect 8906 4728 9087 4731
rect 9115 4751 9179 4752
rect 8709 4708 8728 4710
rect 8743 4708 8777 4710
rect 8709 4692 8789 4708
rect 8709 4686 8728 4692
rect 8425 4660 8528 4670
rect 8379 4658 8528 4660
rect 8549 4658 8584 4670
rect 8218 4656 8380 4658
rect 8230 4636 8249 4656
rect 8264 4654 8294 4656
rect 8113 4628 8154 4636
rect 8236 4632 8249 4636
rect 8301 4640 8380 4656
rect 8412 4656 8584 4658
rect 8412 4640 8491 4656
rect 8498 4654 8528 4656
rect 8076 4618 8105 4628
rect 8119 4618 8148 4628
rect 8163 4618 8193 4632
rect 8236 4618 8279 4632
rect 8301 4628 8491 4640
rect 8556 4636 8562 4656
rect 8286 4618 8316 4628
rect 8317 4618 8475 4628
rect 8479 4618 8509 4628
rect 8513 4618 8543 4632
rect 8571 4618 8584 4656
rect 8656 4670 8685 4686
rect 8699 4670 8728 4686
rect 8743 4676 8773 4692
rect 8801 4670 8807 4718
rect 8810 4712 8829 4718
rect 8844 4712 8874 4720
rect 8810 4704 8874 4712
rect 8810 4688 8890 4704
rect 8906 4697 8968 4728
rect 8984 4697 9046 4728
rect 9115 4726 9164 4751
rect 9179 4726 9209 4742
rect 9078 4712 9108 4720
rect 9115 4718 9225 4726
rect 9078 4704 9123 4712
rect 8810 4686 8829 4688
rect 8844 4686 8890 4688
rect 8810 4670 8890 4686
rect 8917 4684 8952 4697
rect 8993 4694 9030 4697
rect 8993 4692 9035 4694
rect 8922 4681 8952 4684
rect 8931 4677 8938 4681
rect 8938 4676 8939 4677
rect 8897 4670 8907 4676
rect 8656 4662 8691 4670
rect 8656 4636 8657 4662
rect 8664 4636 8691 4662
rect 8599 4618 8629 4632
rect 8656 4628 8691 4636
rect 8693 4662 8734 4670
rect 8693 4636 8708 4662
rect 8715 4636 8734 4662
rect 8798 4658 8829 4670
rect 8844 4658 8947 4670
rect 8959 4660 8985 4686
rect 9000 4681 9030 4692
rect 9062 4688 9124 4704
rect 9062 4686 9108 4688
rect 9062 4670 9124 4686
rect 9136 4670 9142 4718
rect 9145 4710 9225 4718
rect 9145 4708 9164 4710
rect 9179 4708 9213 4710
rect 9145 4692 9225 4708
rect 9145 4670 9164 4692
rect 9179 4676 9209 4692
rect 9237 4686 9243 4760
rect 9246 4686 9265 4830
rect 9280 4686 9286 4830
rect 9295 4760 9308 4830
rect 9360 4826 9382 4830
rect 9353 4804 9382 4818
rect 9435 4804 9451 4818
rect 9489 4814 9495 4816
rect 9502 4814 9610 4830
rect 9617 4814 9623 4816
rect 9631 4814 9646 4830
rect 9712 4824 9731 4827
rect 9353 4802 9451 4804
rect 9478 4802 9646 4814
rect 9661 4804 9677 4818
rect 9712 4805 9734 4824
rect 9744 4818 9760 4819
rect 9743 4816 9760 4818
rect 9744 4811 9760 4816
rect 9734 4804 9740 4805
rect 9743 4804 9772 4811
rect 9661 4803 9772 4804
rect 9661 4802 9778 4803
rect 9337 4794 9388 4802
rect 9435 4794 9469 4802
rect 9337 4782 9362 4794
rect 9369 4782 9388 4794
rect 9442 4792 9469 4794
rect 9478 4792 9699 4802
rect 9734 4799 9740 4802
rect 9442 4788 9699 4792
rect 9337 4774 9388 4782
rect 9435 4774 9699 4788
rect 9743 4794 9778 4802
rect 9289 4726 9308 4760
rect 9353 4766 9382 4774
rect 9353 4760 9370 4766
rect 9353 4758 9387 4760
rect 9435 4758 9451 4774
rect 9452 4764 9660 4774
rect 9661 4764 9677 4774
rect 9725 4770 9740 4785
rect 9743 4782 9744 4794
rect 9751 4782 9778 4794
rect 9743 4774 9778 4782
rect 9743 4773 9772 4774
rect 9463 4760 9677 4764
rect 9478 4758 9677 4760
rect 9712 4760 9725 4770
rect 9743 4760 9760 4773
rect 9712 4758 9760 4760
rect 9354 4754 9387 4758
rect 9350 4752 9387 4754
rect 9350 4751 9417 4752
rect 9350 4746 9381 4751
rect 9387 4746 9417 4751
rect 9350 4742 9417 4746
rect 9323 4739 9417 4742
rect 9323 4732 9372 4739
rect 9323 4726 9353 4732
rect 9372 4727 9377 4732
rect 9289 4710 9369 4726
rect 9381 4718 9417 4739
rect 9478 4734 9667 4758
rect 9712 4757 9759 4758
rect 9725 4752 9759 4757
rect 9493 4731 9667 4734
rect 9486 4728 9667 4731
rect 9695 4751 9759 4752
rect 9289 4708 9308 4710
rect 9323 4708 9357 4710
rect 9289 4692 9369 4708
rect 9289 4686 9308 4692
rect 9005 4660 9108 4670
rect 8959 4658 9108 4660
rect 9129 4658 9164 4670
rect 8798 4656 8960 4658
rect 8810 4636 8829 4656
rect 8844 4654 8874 4656
rect 8693 4628 8734 4636
rect 8816 4632 8829 4636
rect 8881 4640 8960 4656
rect 8992 4656 9164 4658
rect 8992 4640 9071 4656
rect 9078 4654 9108 4656
rect 8656 4618 8685 4628
rect 8699 4618 8728 4628
rect 8743 4618 8773 4632
rect 8816 4618 8859 4632
rect 8881 4628 9071 4640
rect 9136 4636 9142 4656
rect 8866 4618 8896 4628
rect 8897 4618 9055 4628
rect 9059 4618 9089 4628
rect 9093 4618 9123 4632
rect 9151 4618 9164 4656
rect 9236 4670 9265 4686
rect 9279 4670 9308 4686
rect 9323 4676 9353 4692
rect 9381 4670 9387 4718
rect 9390 4712 9409 4718
rect 9424 4712 9454 4720
rect 9390 4704 9454 4712
rect 9390 4688 9470 4704
rect 9486 4697 9548 4728
rect 9564 4697 9626 4728
rect 9695 4726 9744 4751
rect 9759 4726 9789 4742
rect 9658 4712 9688 4720
rect 9695 4718 9805 4726
rect 9658 4704 9703 4712
rect 9390 4686 9409 4688
rect 9424 4686 9470 4688
rect 9390 4670 9470 4686
rect 9497 4684 9532 4697
rect 9573 4694 9610 4697
rect 9573 4692 9615 4694
rect 9502 4681 9532 4684
rect 9511 4677 9518 4681
rect 9518 4676 9519 4677
rect 9477 4670 9487 4676
rect 9236 4662 9271 4670
rect 9236 4636 9237 4662
rect 9244 4636 9271 4662
rect 9179 4618 9209 4632
rect 9236 4628 9271 4636
rect 9273 4662 9314 4670
rect 9273 4636 9288 4662
rect 9295 4636 9314 4662
rect 9378 4658 9409 4670
rect 9424 4658 9527 4670
rect 9539 4660 9565 4686
rect 9580 4681 9610 4692
rect 9642 4688 9704 4704
rect 9642 4686 9688 4688
rect 9642 4670 9704 4686
rect 9716 4670 9722 4718
rect 9725 4710 9805 4718
rect 9725 4708 9744 4710
rect 9759 4708 9793 4710
rect 9725 4692 9805 4708
rect 9725 4670 9744 4692
rect 9759 4676 9789 4692
rect 9817 4686 9823 4760
rect 9826 4686 9845 4830
rect 9860 4686 9866 4830
rect 9875 4760 9888 4830
rect 9940 4826 9962 4830
rect 9933 4804 9962 4818
rect 10015 4804 10031 4818
rect 10069 4814 10075 4816
rect 10082 4814 10190 4830
rect 10197 4814 10203 4816
rect 10211 4814 10226 4830
rect 10292 4824 10311 4827
rect 9933 4802 10031 4804
rect 10058 4802 10226 4814
rect 10241 4804 10257 4818
rect 10292 4805 10314 4824
rect 10324 4818 10340 4819
rect 10323 4816 10340 4818
rect 10324 4811 10340 4816
rect 10314 4804 10320 4805
rect 10323 4804 10352 4811
rect 10241 4803 10352 4804
rect 10241 4802 10358 4803
rect 9917 4794 9968 4802
rect 10015 4794 10049 4802
rect 9917 4782 9942 4794
rect 9949 4782 9968 4794
rect 10022 4792 10049 4794
rect 10058 4792 10279 4802
rect 10314 4799 10320 4802
rect 10022 4788 10279 4792
rect 9917 4774 9968 4782
rect 10015 4774 10279 4788
rect 10323 4794 10358 4802
rect 9869 4726 9888 4760
rect 9933 4766 9962 4774
rect 9933 4760 9950 4766
rect 9933 4758 9967 4760
rect 10015 4758 10031 4774
rect 10032 4764 10240 4774
rect 10241 4764 10257 4774
rect 10305 4770 10320 4785
rect 10323 4782 10324 4794
rect 10331 4782 10358 4794
rect 10323 4774 10358 4782
rect 10323 4773 10352 4774
rect 10043 4760 10257 4764
rect 10058 4758 10257 4760
rect 10292 4760 10305 4770
rect 10323 4760 10340 4773
rect 10292 4758 10340 4760
rect 9934 4754 9967 4758
rect 9930 4752 9967 4754
rect 9930 4751 9997 4752
rect 9930 4746 9961 4751
rect 9967 4746 9997 4751
rect 9930 4742 9997 4746
rect 9903 4739 9997 4742
rect 9903 4732 9952 4739
rect 9903 4726 9933 4732
rect 9952 4727 9957 4732
rect 9869 4710 9949 4726
rect 9961 4718 9997 4739
rect 10058 4734 10247 4758
rect 10292 4757 10339 4758
rect 10305 4752 10339 4757
rect 10073 4731 10247 4734
rect 10066 4728 10247 4731
rect 10275 4751 10339 4752
rect 9869 4708 9888 4710
rect 9903 4708 9937 4710
rect 9869 4692 9949 4708
rect 9869 4686 9888 4692
rect 9585 4660 9688 4670
rect 9539 4658 9688 4660
rect 9709 4658 9744 4670
rect 9378 4656 9540 4658
rect 9390 4636 9409 4656
rect 9424 4654 9454 4656
rect 9273 4628 9314 4636
rect 9396 4632 9409 4636
rect 9461 4640 9540 4656
rect 9572 4656 9744 4658
rect 9572 4640 9651 4656
rect 9658 4654 9688 4656
rect 9236 4618 9265 4628
rect 9279 4618 9308 4628
rect 9323 4618 9353 4632
rect 9396 4618 9439 4632
rect 9461 4628 9651 4640
rect 9716 4636 9722 4656
rect 9446 4618 9476 4628
rect 9477 4618 9635 4628
rect 9639 4618 9669 4628
rect 9673 4618 9703 4632
rect 9731 4618 9744 4656
rect 9816 4670 9845 4686
rect 9859 4670 9888 4686
rect 9903 4676 9933 4692
rect 9961 4670 9967 4718
rect 9970 4712 9989 4718
rect 10004 4712 10034 4720
rect 9970 4704 10034 4712
rect 9970 4688 10050 4704
rect 10066 4697 10128 4728
rect 10144 4697 10206 4728
rect 10275 4726 10324 4751
rect 10339 4726 10369 4742
rect 10238 4712 10268 4720
rect 10275 4718 10385 4726
rect 10238 4704 10283 4712
rect 9970 4686 9989 4688
rect 10004 4686 10050 4688
rect 9970 4670 10050 4686
rect 10077 4684 10112 4697
rect 10153 4694 10190 4697
rect 10153 4692 10195 4694
rect 10082 4681 10112 4684
rect 10091 4677 10098 4681
rect 10098 4676 10099 4677
rect 10057 4670 10067 4676
rect 9816 4662 9851 4670
rect 9816 4636 9817 4662
rect 9824 4636 9851 4662
rect 9759 4618 9789 4632
rect 9816 4628 9851 4636
rect 9853 4662 9894 4670
rect 9853 4636 9868 4662
rect 9875 4636 9894 4662
rect 9958 4658 9989 4670
rect 10004 4658 10107 4670
rect 10119 4660 10145 4686
rect 10160 4681 10190 4692
rect 10222 4688 10284 4704
rect 10222 4686 10268 4688
rect 10222 4670 10284 4686
rect 10296 4670 10302 4718
rect 10305 4710 10385 4718
rect 10305 4708 10324 4710
rect 10339 4708 10373 4710
rect 10305 4692 10385 4708
rect 10305 4670 10324 4692
rect 10339 4676 10369 4692
rect 10397 4686 10403 4760
rect 10406 4686 10425 4830
rect 10440 4686 10446 4830
rect 10455 4760 10468 4830
rect 10520 4826 10542 4830
rect 10513 4804 10542 4818
rect 10595 4804 10611 4818
rect 10649 4814 10655 4816
rect 10662 4814 10770 4830
rect 10777 4814 10783 4816
rect 10791 4814 10806 4830
rect 10872 4824 10891 4827
rect 10513 4802 10611 4804
rect 10638 4802 10806 4814
rect 10821 4804 10837 4818
rect 10872 4805 10894 4824
rect 10904 4818 10920 4819
rect 10903 4816 10920 4818
rect 10904 4811 10920 4816
rect 10894 4804 10900 4805
rect 10903 4804 10932 4811
rect 10821 4803 10932 4804
rect 10821 4802 10938 4803
rect 10497 4794 10548 4802
rect 10595 4794 10629 4802
rect 10497 4782 10522 4794
rect 10529 4782 10548 4794
rect 10602 4792 10629 4794
rect 10638 4792 10859 4802
rect 10894 4799 10900 4802
rect 10602 4788 10859 4792
rect 10497 4774 10548 4782
rect 10595 4774 10859 4788
rect 10903 4794 10938 4802
rect 10449 4726 10468 4760
rect 10513 4766 10542 4774
rect 10513 4760 10530 4766
rect 10513 4758 10547 4760
rect 10595 4758 10611 4774
rect 10612 4764 10820 4774
rect 10821 4764 10837 4774
rect 10885 4770 10900 4785
rect 10903 4782 10904 4794
rect 10911 4782 10938 4794
rect 10903 4774 10938 4782
rect 10903 4773 10932 4774
rect 10623 4760 10837 4764
rect 10638 4758 10837 4760
rect 10872 4760 10885 4770
rect 10903 4760 10920 4773
rect 10872 4758 10920 4760
rect 10514 4754 10547 4758
rect 10510 4752 10547 4754
rect 10510 4751 10577 4752
rect 10510 4746 10541 4751
rect 10547 4746 10577 4751
rect 10510 4742 10577 4746
rect 10483 4739 10577 4742
rect 10483 4732 10532 4739
rect 10483 4726 10513 4732
rect 10532 4727 10537 4732
rect 10449 4710 10529 4726
rect 10541 4718 10577 4739
rect 10638 4734 10827 4758
rect 10872 4757 10919 4758
rect 10885 4752 10919 4757
rect 10653 4731 10827 4734
rect 10646 4728 10827 4731
rect 10855 4751 10919 4752
rect 10449 4708 10468 4710
rect 10483 4708 10517 4710
rect 10449 4692 10529 4708
rect 10449 4686 10468 4692
rect 10165 4660 10268 4670
rect 10119 4658 10268 4660
rect 10289 4658 10324 4670
rect 9958 4656 10120 4658
rect 9970 4636 9989 4656
rect 10004 4654 10034 4656
rect 9853 4628 9894 4636
rect 9976 4632 9989 4636
rect 10041 4640 10120 4656
rect 10152 4656 10324 4658
rect 10152 4640 10231 4656
rect 10238 4654 10268 4656
rect 9816 4618 9845 4628
rect 9859 4618 9888 4628
rect 9903 4618 9933 4632
rect 9976 4618 10019 4632
rect 10041 4628 10231 4640
rect 10296 4636 10302 4656
rect 10026 4618 10056 4628
rect 10057 4618 10215 4628
rect 10219 4618 10249 4628
rect 10253 4618 10283 4632
rect 10311 4618 10324 4656
rect 10396 4670 10425 4686
rect 10439 4670 10468 4686
rect 10483 4676 10513 4692
rect 10541 4670 10547 4718
rect 10550 4712 10569 4718
rect 10584 4712 10614 4720
rect 10550 4704 10614 4712
rect 10550 4688 10630 4704
rect 10646 4697 10708 4728
rect 10724 4697 10786 4728
rect 10855 4726 10904 4751
rect 10919 4726 10949 4742
rect 10818 4712 10848 4720
rect 10855 4718 10965 4726
rect 10818 4704 10863 4712
rect 10550 4686 10569 4688
rect 10584 4686 10630 4688
rect 10550 4670 10630 4686
rect 10657 4684 10692 4697
rect 10733 4694 10770 4697
rect 10733 4692 10775 4694
rect 10662 4681 10692 4684
rect 10671 4677 10678 4681
rect 10678 4676 10679 4677
rect 10637 4670 10647 4676
rect 10396 4662 10431 4670
rect 10396 4636 10397 4662
rect 10404 4636 10431 4662
rect 10339 4618 10369 4632
rect 10396 4628 10431 4636
rect 10433 4662 10474 4670
rect 10433 4636 10448 4662
rect 10455 4636 10474 4662
rect 10538 4658 10569 4670
rect 10584 4658 10687 4670
rect 10699 4660 10725 4686
rect 10740 4681 10770 4692
rect 10802 4688 10864 4704
rect 10802 4686 10848 4688
rect 10802 4670 10864 4686
rect 10876 4670 10882 4718
rect 10885 4710 10965 4718
rect 10885 4708 10904 4710
rect 10919 4708 10953 4710
rect 10885 4692 10965 4708
rect 10885 4670 10904 4692
rect 10919 4676 10949 4692
rect 10977 4686 10983 4760
rect 10986 4686 11005 4830
rect 11020 4686 11026 4830
rect 11035 4760 11048 4830
rect 11100 4826 11122 4830
rect 11093 4804 11122 4818
rect 11175 4804 11191 4818
rect 11229 4814 11235 4816
rect 11242 4814 11350 4830
rect 11357 4814 11363 4816
rect 11371 4814 11386 4830
rect 11452 4824 11471 4827
rect 11093 4802 11191 4804
rect 11218 4802 11386 4814
rect 11401 4804 11417 4818
rect 11452 4805 11474 4824
rect 11484 4818 11500 4819
rect 11483 4816 11500 4818
rect 11484 4811 11500 4816
rect 11474 4804 11480 4805
rect 11483 4804 11512 4811
rect 11401 4803 11512 4804
rect 11401 4802 11518 4803
rect 11077 4794 11128 4802
rect 11175 4794 11209 4802
rect 11077 4782 11102 4794
rect 11109 4782 11128 4794
rect 11182 4792 11209 4794
rect 11218 4792 11439 4802
rect 11474 4799 11480 4802
rect 11182 4788 11439 4792
rect 11077 4774 11128 4782
rect 11175 4774 11439 4788
rect 11483 4794 11518 4802
rect 11029 4726 11048 4760
rect 11093 4766 11122 4774
rect 11093 4760 11110 4766
rect 11093 4758 11127 4760
rect 11175 4758 11191 4774
rect 11192 4764 11400 4774
rect 11401 4764 11417 4774
rect 11465 4770 11480 4785
rect 11483 4782 11484 4794
rect 11491 4782 11518 4794
rect 11483 4774 11518 4782
rect 11483 4773 11512 4774
rect 11203 4760 11417 4764
rect 11218 4758 11417 4760
rect 11452 4760 11465 4770
rect 11483 4760 11500 4773
rect 11452 4758 11500 4760
rect 11094 4754 11127 4758
rect 11090 4752 11127 4754
rect 11090 4751 11157 4752
rect 11090 4746 11121 4751
rect 11127 4746 11157 4751
rect 11090 4742 11157 4746
rect 11063 4739 11157 4742
rect 11063 4732 11112 4739
rect 11063 4726 11093 4732
rect 11112 4727 11117 4732
rect 11029 4710 11109 4726
rect 11121 4718 11157 4739
rect 11218 4734 11407 4758
rect 11452 4757 11499 4758
rect 11465 4752 11499 4757
rect 11233 4731 11407 4734
rect 11226 4728 11407 4731
rect 11435 4751 11499 4752
rect 11029 4708 11048 4710
rect 11063 4708 11097 4710
rect 11029 4692 11109 4708
rect 11029 4686 11048 4692
rect 10745 4660 10848 4670
rect 10699 4658 10848 4660
rect 10869 4658 10904 4670
rect 10538 4656 10700 4658
rect 10550 4636 10569 4656
rect 10584 4654 10614 4656
rect 10433 4628 10474 4636
rect 10556 4632 10569 4636
rect 10621 4640 10700 4656
rect 10732 4656 10904 4658
rect 10732 4640 10811 4656
rect 10818 4654 10848 4656
rect 10396 4618 10425 4628
rect 10439 4618 10468 4628
rect 10483 4618 10513 4632
rect 10556 4618 10599 4632
rect 10621 4628 10811 4640
rect 10876 4636 10882 4656
rect 10606 4618 10636 4628
rect 10637 4618 10795 4628
rect 10799 4618 10829 4628
rect 10833 4618 10863 4632
rect 10891 4618 10904 4656
rect 10976 4670 11005 4686
rect 11019 4670 11048 4686
rect 11063 4676 11093 4692
rect 11121 4670 11127 4718
rect 11130 4712 11149 4718
rect 11164 4712 11194 4720
rect 11130 4704 11194 4712
rect 11130 4688 11210 4704
rect 11226 4697 11288 4728
rect 11304 4697 11366 4728
rect 11435 4726 11484 4751
rect 11499 4726 11529 4742
rect 11398 4712 11428 4720
rect 11435 4718 11545 4726
rect 11398 4704 11443 4712
rect 11130 4686 11149 4688
rect 11164 4686 11210 4688
rect 11130 4670 11210 4686
rect 11237 4684 11272 4697
rect 11313 4694 11350 4697
rect 11313 4692 11355 4694
rect 11242 4681 11272 4684
rect 11251 4677 11258 4681
rect 11258 4676 11259 4677
rect 11217 4670 11227 4676
rect 10976 4662 11011 4670
rect 10976 4636 10977 4662
rect 10984 4636 11011 4662
rect 10919 4618 10949 4632
rect 10976 4628 11011 4636
rect 11013 4662 11054 4670
rect 11013 4636 11028 4662
rect 11035 4636 11054 4662
rect 11118 4658 11149 4670
rect 11164 4658 11267 4670
rect 11279 4660 11305 4686
rect 11320 4681 11350 4692
rect 11382 4688 11444 4704
rect 11382 4686 11428 4688
rect 11382 4670 11444 4686
rect 11456 4670 11462 4718
rect 11465 4710 11545 4718
rect 11465 4708 11484 4710
rect 11499 4708 11533 4710
rect 11465 4692 11545 4708
rect 11465 4670 11484 4692
rect 11499 4676 11529 4692
rect 11557 4686 11563 4760
rect 11566 4686 11585 4830
rect 11600 4686 11606 4830
rect 11615 4760 11628 4830
rect 11680 4826 11702 4830
rect 11673 4804 11702 4818
rect 11755 4804 11771 4818
rect 11809 4814 11815 4816
rect 11822 4814 11930 4830
rect 11937 4814 11943 4816
rect 11951 4814 11966 4830
rect 12032 4824 12051 4827
rect 11673 4802 11771 4804
rect 11798 4802 11966 4814
rect 11981 4804 11997 4818
rect 12032 4805 12054 4824
rect 12064 4818 12080 4819
rect 12063 4816 12080 4818
rect 12064 4811 12080 4816
rect 12054 4804 12060 4805
rect 12063 4804 12092 4811
rect 11981 4803 12092 4804
rect 11981 4802 12098 4803
rect 11657 4794 11708 4802
rect 11755 4794 11789 4802
rect 11657 4782 11682 4794
rect 11689 4782 11708 4794
rect 11762 4792 11789 4794
rect 11798 4792 12019 4802
rect 12054 4799 12060 4802
rect 11762 4788 12019 4792
rect 11657 4774 11708 4782
rect 11755 4774 12019 4788
rect 12063 4794 12098 4802
rect 11609 4726 11628 4760
rect 11673 4766 11702 4774
rect 11673 4760 11690 4766
rect 11673 4758 11707 4760
rect 11755 4758 11771 4774
rect 11772 4764 11980 4774
rect 11981 4764 11997 4774
rect 12045 4770 12060 4785
rect 12063 4782 12064 4794
rect 12071 4782 12098 4794
rect 12063 4774 12098 4782
rect 12063 4773 12092 4774
rect 11783 4760 11997 4764
rect 11798 4758 11997 4760
rect 12032 4760 12045 4770
rect 12063 4760 12080 4773
rect 12032 4758 12080 4760
rect 11674 4754 11707 4758
rect 11670 4752 11707 4754
rect 11670 4751 11737 4752
rect 11670 4746 11701 4751
rect 11707 4746 11737 4751
rect 11670 4742 11737 4746
rect 11643 4739 11737 4742
rect 11643 4732 11692 4739
rect 11643 4726 11673 4732
rect 11692 4727 11697 4732
rect 11609 4710 11689 4726
rect 11701 4718 11737 4739
rect 11798 4734 11987 4758
rect 12032 4757 12079 4758
rect 12045 4752 12079 4757
rect 11813 4731 11987 4734
rect 11806 4728 11987 4731
rect 12015 4751 12079 4752
rect 11609 4708 11628 4710
rect 11643 4708 11677 4710
rect 11609 4692 11689 4708
rect 11609 4686 11628 4692
rect 11325 4660 11428 4670
rect 11279 4658 11428 4660
rect 11449 4658 11484 4670
rect 11118 4656 11280 4658
rect 11130 4636 11149 4656
rect 11164 4654 11194 4656
rect 11013 4628 11054 4636
rect 11136 4632 11149 4636
rect 11201 4640 11280 4656
rect 11312 4656 11484 4658
rect 11312 4640 11391 4656
rect 11398 4654 11428 4656
rect 10976 4618 11005 4628
rect 11019 4618 11048 4628
rect 11063 4618 11093 4632
rect 11136 4618 11179 4632
rect 11201 4628 11391 4640
rect 11456 4636 11462 4656
rect 11186 4618 11216 4628
rect 11217 4618 11375 4628
rect 11379 4618 11409 4628
rect 11413 4618 11443 4632
rect 11471 4618 11484 4656
rect 11556 4670 11585 4686
rect 11599 4670 11628 4686
rect 11643 4676 11673 4692
rect 11701 4670 11707 4718
rect 11710 4712 11729 4718
rect 11744 4712 11774 4720
rect 11710 4704 11774 4712
rect 11710 4688 11790 4704
rect 11806 4697 11868 4728
rect 11884 4697 11946 4728
rect 12015 4726 12064 4751
rect 12079 4726 12109 4742
rect 11978 4712 12008 4720
rect 12015 4718 12125 4726
rect 11978 4704 12023 4712
rect 11710 4686 11729 4688
rect 11744 4686 11790 4688
rect 11710 4670 11790 4686
rect 11817 4684 11852 4697
rect 11893 4694 11930 4697
rect 11893 4692 11935 4694
rect 11822 4681 11852 4684
rect 11831 4677 11838 4681
rect 11838 4676 11839 4677
rect 11797 4670 11807 4676
rect 11556 4662 11591 4670
rect 11556 4636 11557 4662
rect 11564 4636 11591 4662
rect 11499 4618 11529 4632
rect 11556 4628 11591 4636
rect 11593 4662 11634 4670
rect 11593 4636 11608 4662
rect 11615 4636 11634 4662
rect 11698 4658 11729 4670
rect 11744 4658 11847 4670
rect 11859 4660 11885 4686
rect 11900 4681 11930 4692
rect 11962 4688 12024 4704
rect 11962 4686 12008 4688
rect 11962 4670 12024 4686
rect 12036 4670 12042 4718
rect 12045 4710 12125 4718
rect 12045 4708 12064 4710
rect 12079 4708 12113 4710
rect 12045 4692 12125 4708
rect 12045 4670 12064 4692
rect 12079 4676 12109 4692
rect 12137 4686 12143 4760
rect 12146 4686 12165 4830
rect 12180 4686 12186 4830
rect 12195 4760 12208 4830
rect 12260 4826 12282 4830
rect 12253 4804 12282 4818
rect 12335 4804 12351 4818
rect 12389 4814 12395 4816
rect 12402 4814 12510 4830
rect 12517 4814 12523 4816
rect 12531 4814 12546 4830
rect 12612 4824 12631 4827
rect 12253 4802 12351 4804
rect 12378 4802 12546 4814
rect 12561 4804 12577 4818
rect 12612 4805 12634 4824
rect 12644 4818 12660 4819
rect 12643 4816 12660 4818
rect 12644 4811 12660 4816
rect 12634 4804 12640 4805
rect 12643 4804 12672 4811
rect 12561 4803 12672 4804
rect 12561 4802 12678 4803
rect 12237 4794 12288 4802
rect 12335 4794 12369 4802
rect 12237 4782 12262 4794
rect 12269 4782 12288 4794
rect 12342 4792 12369 4794
rect 12378 4792 12599 4802
rect 12634 4799 12640 4802
rect 12342 4788 12599 4792
rect 12237 4774 12288 4782
rect 12335 4774 12599 4788
rect 12643 4794 12678 4802
rect 12189 4726 12208 4760
rect 12253 4766 12282 4774
rect 12253 4760 12270 4766
rect 12253 4758 12287 4760
rect 12335 4758 12351 4774
rect 12352 4764 12560 4774
rect 12561 4764 12577 4774
rect 12625 4770 12640 4785
rect 12643 4782 12644 4794
rect 12651 4782 12678 4794
rect 12643 4774 12678 4782
rect 12643 4773 12672 4774
rect 12363 4760 12577 4764
rect 12378 4758 12577 4760
rect 12612 4760 12625 4770
rect 12643 4760 12660 4773
rect 12612 4758 12660 4760
rect 12254 4754 12287 4758
rect 12250 4752 12287 4754
rect 12250 4751 12317 4752
rect 12250 4746 12281 4751
rect 12287 4746 12317 4751
rect 12250 4742 12317 4746
rect 12223 4739 12317 4742
rect 12223 4732 12272 4739
rect 12223 4726 12253 4732
rect 12272 4727 12277 4732
rect 12189 4710 12269 4726
rect 12281 4718 12317 4739
rect 12378 4734 12567 4758
rect 12612 4757 12659 4758
rect 12625 4752 12659 4757
rect 12393 4731 12567 4734
rect 12386 4728 12567 4731
rect 12595 4751 12659 4752
rect 12189 4708 12208 4710
rect 12223 4708 12257 4710
rect 12189 4692 12269 4708
rect 12189 4686 12208 4692
rect 11905 4660 12008 4670
rect 11859 4658 12008 4660
rect 12029 4658 12064 4670
rect 11698 4656 11860 4658
rect 11710 4636 11729 4656
rect 11744 4654 11774 4656
rect 11593 4628 11634 4636
rect 11716 4632 11729 4636
rect 11781 4640 11860 4656
rect 11892 4656 12064 4658
rect 11892 4640 11971 4656
rect 11978 4654 12008 4656
rect 11556 4618 11585 4628
rect 11599 4618 11628 4628
rect 11643 4618 11673 4632
rect 11716 4618 11759 4632
rect 11781 4628 11971 4640
rect 12036 4636 12042 4656
rect 11766 4618 11796 4628
rect 11797 4618 11955 4628
rect 11959 4618 11989 4628
rect 11993 4618 12023 4632
rect 12051 4618 12064 4656
rect 12136 4670 12165 4686
rect 12179 4670 12208 4686
rect 12223 4676 12253 4692
rect 12281 4670 12287 4718
rect 12290 4712 12309 4718
rect 12324 4712 12354 4720
rect 12290 4704 12354 4712
rect 12290 4688 12370 4704
rect 12386 4697 12448 4728
rect 12464 4697 12526 4728
rect 12595 4726 12644 4751
rect 12659 4726 12689 4742
rect 12558 4712 12588 4720
rect 12595 4718 12705 4726
rect 12558 4704 12603 4712
rect 12290 4686 12309 4688
rect 12324 4686 12370 4688
rect 12290 4670 12370 4686
rect 12397 4684 12432 4697
rect 12473 4694 12510 4697
rect 12473 4692 12515 4694
rect 12402 4681 12432 4684
rect 12411 4677 12418 4681
rect 12418 4676 12419 4677
rect 12377 4670 12387 4676
rect 12136 4662 12171 4670
rect 12136 4636 12137 4662
rect 12144 4636 12171 4662
rect 12079 4618 12109 4632
rect 12136 4628 12171 4636
rect 12173 4662 12214 4670
rect 12173 4636 12188 4662
rect 12195 4636 12214 4662
rect 12278 4658 12309 4670
rect 12324 4658 12427 4670
rect 12439 4660 12465 4686
rect 12480 4681 12510 4692
rect 12542 4688 12604 4704
rect 12542 4686 12588 4688
rect 12542 4670 12604 4686
rect 12616 4670 12622 4718
rect 12625 4710 12705 4718
rect 12625 4708 12644 4710
rect 12659 4708 12693 4710
rect 12625 4692 12705 4708
rect 12625 4670 12644 4692
rect 12659 4676 12689 4692
rect 12717 4686 12723 4760
rect 12726 4686 12745 4830
rect 12760 4686 12766 4830
rect 12775 4760 12788 4830
rect 12840 4826 12862 4830
rect 12833 4804 12862 4818
rect 12915 4804 12931 4818
rect 12969 4814 12975 4816
rect 12982 4814 13090 4830
rect 13097 4814 13103 4816
rect 13111 4814 13126 4830
rect 13192 4824 13211 4827
rect 12833 4802 12931 4804
rect 12958 4802 13126 4814
rect 13141 4804 13157 4818
rect 13192 4805 13214 4824
rect 13224 4818 13240 4819
rect 13223 4816 13240 4818
rect 13224 4811 13240 4816
rect 13214 4804 13220 4805
rect 13223 4804 13252 4811
rect 13141 4803 13252 4804
rect 13141 4802 13258 4803
rect 12817 4794 12868 4802
rect 12915 4794 12949 4802
rect 12817 4782 12842 4794
rect 12849 4782 12868 4794
rect 12922 4792 12949 4794
rect 12958 4792 13179 4802
rect 13214 4799 13220 4802
rect 12922 4788 13179 4792
rect 12817 4774 12868 4782
rect 12915 4774 13179 4788
rect 13223 4794 13258 4802
rect 12769 4726 12788 4760
rect 12833 4766 12862 4774
rect 12833 4760 12850 4766
rect 12833 4758 12867 4760
rect 12915 4758 12931 4774
rect 12932 4764 13140 4774
rect 13141 4764 13157 4774
rect 13205 4770 13220 4785
rect 13223 4782 13224 4794
rect 13231 4782 13258 4794
rect 13223 4774 13258 4782
rect 13223 4773 13252 4774
rect 12943 4760 13157 4764
rect 12958 4758 13157 4760
rect 13192 4760 13205 4770
rect 13223 4760 13240 4773
rect 13192 4758 13240 4760
rect 12834 4754 12867 4758
rect 12830 4752 12867 4754
rect 12830 4751 12897 4752
rect 12830 4746 12861 4751
rect 12867 4746 12897 4751
rect 12830 4742 12897 4746
rect 12803 4739 12897 4742
rect 12803 4732 12852 4739
rect 12803 4726 12833 4732
rect 12852 4727 12857 4732
rect 12769 4710 12849 4726
rect 12861 4718 12897 4739
rect 12958 4734 13147 4758
rect 13192 4757 13239 4758
rect 13205 4752 13239 4757
rect 12973 4731 13147 4734
rect 12966 4728 13147 4731
rect 13175 4751 13239 4752
rect 12769 4708 12788 4710
rect 12803 4708 12837 4710
rect 12769 4692 12849 4708
rect 12769 4686 12788 4692
rect 12485 4660 12588 4670
rect 12439 4658 12588 4660
rect 12609 4658 12644 4670
rect 12278 4656 12440 4658
rect 12290 4636 12309 4656
rect 12324 4654 12354 4656
rect 12173 4628 12214 4636
rect 12296 4632 12309 4636
rect 12361 4640 12440 4656
rect 12472 4656 12644 4658
rect 12472 4640 12551 4656
rect 12558 4654 12588 4656
rect 12136 4618 12165 4628
rect 12179 4618 12208 4628
rect 12223 4618 12253 4632
rect 12296 4618 12339 4632
rect 12361 4628 12551 4640
rect 12616 4636 12622 4656
rect 12346 4618 12376 4628
rect 12377 4618 12535 4628
rect 12539 4618 12569 4628
rect 12573 4618 12603 4632
rect 12631 4618 12644 4656
rect 12716 4670 12745 4686
rect 12759 4670 12788 4686
rect 12803 4676 12833 4692
rect 12861 4670 12867 4718
rect 12870 4712 12889 4718
rect 12904 4712 12934 4720
rect 12870 4704 12934 4712
rect 12870 4688 12950 4704
rect 12966 4697 13028 4728
rect 13044 4697 13106 4728
rect 13175 4726 13224 4751
rect 13239 4726 13269 4742
rect 13138 4712 13168 4720
rect 13175 4718 13285 4726
rect 13138 4704 13183 4712
rect 12870 4686 12889 4688
rect 12904 4686 12950 4688
rect 12870 4670 12950 4686
rect 12977 4684 13012 4697
rect 13053 4694 13090 4697
rect 13053 4692 13095 4694
rect 12982 4681 13012 4684
rect 12991 4677 12998 4681
rect 12998 4676 12999 4677
rect 12957 4670 12967 4676
rect 12716 4662 12751 4670
rect 12716 4636 12717 4662
rect 12724 4636 12751 4662
rect 12659 4618 12689 4632
rect 12716 4628 12751 4636
rect 12753 4662 12794 4670
rect 12753 4636 12768 4662
rect 12775 4636 12794 4662
rect 12858 4658 12889 4670
rect 12904 4658 13007 4670
rect 13019 4660 13045 4686
rect 13060 4681 13090 4692
rect 13122 4688 13184 4704
rect 13122 4686 13168 4688
rect 13122 4670 13184 4686
rect 13196 4670 13202 4718
rect 13205 4710 13285 4718
rect 13205 4708 13224 4710
rect 13239 4708 13273 4710
rect 13205 4692 13285 4708
rect 13205 4670 13224 4692
rect 13239 4676 13269 4692
rect 13297 4686 13303 4760
rect 13306 4686 13325 4830
rect 13340 4686 13346 4830
rect 13355 4760 13368 4830
rect 13420 4826 13442 4830
rect 13413 4804 13442 4818
rect 13495 4804 13511 4818
rect 13549 4814 13555 4816
rect 13562 4814 13670 4830
rect 13677 4814 13683 4816
rect 13691 4814 13706 4830
rect 13772 4824 13791 4827
rect 13413 4802 13511 4804
rect 13538 4802 13706 4814
rect 13721 4804 13737 4818
rect 13772 4805 13794 4824
rect 13804 4818 13820 4819
rect 13803 4816 13820 4818
rect 13804 4811 13820 4816
rect 13794 4804 13800 4805
rect 13803 4804 13832 4811
rect 13721 4803 13832 4804
rect 13721 4802 13838 4803
rect 13397 4794 13448 4802
rect 13495 4794 13529 4802
rect 13397 4782 13422 4794
rect 13429 4782 13448 4794
rect 13502 4792 13529 4794
rect 13538 4792 13759 4802
rect 13794 4799 13800 4802
rect 13502 4788 13759 4792
rect 13397 4774 13448 4782
rect 13495 4774 13759 4788
rect 13803 4794 13838 4802
rect 13349 4726 13368 4760
rect 13413 4766 13442 4774
rect 13413 4760 13430 4766
rect 13413 4758 13447 4760
rect 13495 4758 13511 4774
rect 13512 4764 13720 4774
rect 13721 4764 13737 4774
rect 13785 4770 13800 4785
rect 13803 4782 13804 4794
rect 13811 4782 13838 4794
rect 13803 4774 13838 4782
rect 13803 4773 13832 4774
rect 13523 4760 13737 4764
rect 13538 4758 13737 4760
rect 13772 4760 13785 4770
rect 13803 4760 13820 4773
rect 13772 4758 13820 4760
rect 13414 4754 13447 4758
rect 13410 4752 13447 4754
rect 13410 4751 13477 4752
rect 13410 4746 13441 4751
rect 13447 4746 13477 4751
rect 13410 4742 13477 4746
rect 13383 4739 13477 4742
rect 13383 4732 13432 4739
rect 13383 4726 13413 4732
rect 13432 4727 13437 4732
rect 13349 4710 13429 4726
rect 13441 4718 13477 4739
rect 13538 4734 13727 4758
rect 13772 4757 13819 4758
rect 13785 4752 13819 4757
rect 13553 4731 13727 4734
rect 13546 4728 13727 4731
rect 13755 4751 13819 4752
rect 13349 4708 13368 4710
rect 13383 4708 13417 4710
rect 13349 4692 13429 4708
rect 13349 4686 13368 4692
rect 13065 4660 13168 4670
rect 13019 4658 13168 4660
rect 13189 4658 13224 4670
rect 12858 4656 13020 4658
rect 12870 4636 12889 4656
rect 12904 4654 12934 4656
rect 12753 4628 12794 4636
rect 12876 4632 12889 4636
rect 12941 4640 13020 4656
rect 13052 4656 13224 4658
rect 13052 4640 13131 4656
rect 13138 4654 13168 4656
rect 12716 4618 12745 4628
rect 12759 4618 12788 4628
rect 12803 4618 12833 4632
rect 12876 4618 12919 4632
rect 12941 4628 13131 4640
rect 13196 4636 13202 4656
rect 12926 4618 12956 4628
rect 12957 4618 13115 4628
rect 13119 4618 13149 4628
rect 13153 4618 13183 4632
rect 13211 4618 13224 4656
rect 13296 4670 13325 4686
rect 13339 4670 13368 4686
rect 13383 4676 13413 4692
rect 13441 4670 13447 4718
rect 13450 4712 13469 4718
rect 13484 4712 13514 4720
rect 13450 4704 13514 4712
rect 13450 4688 13530 4704
rect 13546 4697 13608 4728
rect 13624 4697 13686 4728
rect 13755 4726 13804 4751
rect 13819 4726 13849 4742
rect 13718 4712 13748 4720
rect 13755 4718 13865 4726
rect 13718 4704 13763 4712
rect 13450 4686 13469 4688
rect 13484 4686 13530 4688
rect 13450 4670 13530 4686
rect 13557 4684 13592 4697
rect 13633 4694 13670 4697
rect 13633 4692 13675 4694
rect 13562 4681 13592 4684
rect 13571 4677 13578 4681
rect 13578 4676 13579 4677
rect 13537 4670 13547 4676
rect 13296 4662 13331 4670
rect 13296 4636 13297 4662
rect 13304 4636 13331 4662
rect 13239 4618 13269 4632
rect 13296 4628 13331 4636
rect 13333 4662 13374 4670
rect 13333 4636 13348 4662
rect 13355 4636 13374 4662
rect 13438 4658 13469 4670
rect 13484 4658 13587 4670
rect 13599 4660 13625 4686
rect 13640 4681 13670 4692
rect 13702 4688 13764 4704
rect 13702 4686 13748 4688
rect 13702 4670 13764 4686
rect 13776 4670 13782 4718
rect 13785 4710 13865 4718
rect 13785 4708 13804 4710
rect 13819 4708 13853 4710
rect 13785 4692 13865 4708
rect 13785 4670 13804 4692
rect 13819 4676 13849 4692
rect 13877 4686 13883 4760
rect 13886 4686 13905 4830
rect 13920 4686 13926 4830
rect 13935 4760 13948 4830
rect 14000 4826 14022 4830
rect 13993 4804 14022 4818
rect 14075 4804 14091 4818
rect 14129 4814 14135 4816
rect 14142 4814 14250 4830
rect 14257 4814 14263 4816
rect 14271 4814 14286 4830
rect 14352 4824 14371 4827
rect 13993 4802 14091 4804
rect 14118 4802 14286 4814
rect 14301 4804 14317 4818
rect 14352 4805 14374 4824
rect 14384 4818 14400 4819
rect 14383 4816 14400 4818
rect 14384 4811 14400 4816
rect 14374 4804 14380 4805
rect 14383 4804 14412 4811
rect 14301 4803 14412 4804
rect 14301 4802 14418 4803
rect 13977 4794 14028 4802
rect 14075 4794 14109 4802
rect 13977 4782 14002 4794
rect 14009 4782 14028 4794
rect 14082 4792 14109 4794
rect 14118 4792 14339 4802
rect 14374 4799 14380 4802
rect 14082 4788 14339 4792
rect 13977 4774 14028 4782
rect 14075 4774 14339 4788
rect 14383 4794 14418 4802
rect 13929 4726 13948 4760
rect 13993 4766 14022 4774
rect 13993 4760 14010 4766
rect 13993 4758 14027 4760
rect 14075 4758 14091 4774
rect 14092 4764 14300 4774
rect 14301 4764 14317 4774
rect 14365 4770 14380 4785
rect 14383 4782 14384 4794
rect 14391 4782 14418 4794
rect 14383 4774 14418 4782
rect 14383 4773 14412 4774
rect 14103 4760 14317 4764
rect 14118 4758 14317 4760
rect 14352 4760 14365 4770
rect 14383 4760 14400 4773
rect 14352 4758 14400 4760
rect 13994 4754 14027 4758
rect 13990 4752 14027 4754
rect 13990 4751 14057 4752
rect 13990 4746 14021 4751
rect 14027 4746 14057 4751
rect 13990 4742 14057 4746
rect 13963 4739 14057 4742
rect 13963 4732 14012 4739
rect 13963 4726 13993 4732
rect 14012 4727 14017 4732
rect 13929 4710 14009 4726
rect 14021 4718 14057 4739
rect 14118 4734 14307 4758
rect 14352 4757 14399 4758
rect 14365 4752 14399 4757
rect 14133 4731 14307 4734
rect 14126 4728 14307 4731
rect 14335 4751 14399 4752
rect 13929 4708 13948 4710
rect 13963 4708 13997 4710
rect 13929 4692 14009 4708
rect 13929 4686 13948 4692
rect 13645 4660 13748 4670
rect 13599 4658 13748 4660
rect 13769 4658 13804 4670
rect 13438 4656 13600 4658
rect 13450 4636 13469 4656
rect 13484 4654 13514 4656
rect 13333 4628 13374 4636
rect 13456 4632 13469 4636
rect 13521 4640 13600 4656
rect 13632 4656 13804 4658
rect 13632 4640 13711 4656
rect 13718 4654 13748 4656
rect 13296 4618 13325 4628
rect 13339 4618 13368 4628
rect 13383 4618 13413 4632
rect 13456 4618 13499 4632
rect 13521 4628 13711 4640
rect 13776 4636 13782 4656
rect 13506 4618 13536 4628
rect 13537 4618 13695 4628
rect 13699 4618 13729 4628
rect 13733 4618 13763 4632
rect 13791 4618 13804 4656
rect 13876 4670 13905 4686
rect 13919 4670 13948 4686
rect 13963 4676 13993 4692
rect 14021 4670 14027 4718
rect 14030 4712 14049 4718
rect 14064 4712 14094 4720
rect 14030 4704 14094 4712
rect 14030 4688 14110 4704
rect 14126 4697 14188 4728
rect 14204 4697 14266 4728
rect 14335 4726 14384 4751
rect 14399 4726 14429 4742
rect 14298 4712 14328 4720
rect 14335 4718 14445 4726
rect 14298 4704 14343 4712
rect 14030 4686 14049 4688
rect 14064 4686 14110 4688
rect 14030 4670 14110 4686
rect 14137 4684 14172 4697
rect 14213 4694 14250 4697
rect 14213 4692 14255 4694
rect 14142 4681 14172 4684
rect 14151 4677 14158 4681
rect 14158 4676 14159 4677
rect 14117 4670 14127 4676
rect 13876 4662 13911 4670
rect 13876 4636 13877 4662
rect 13884 4636 13911 4662
rect 13819 4618 13849 4632
rect 13876 4628 13911 4636
rect 13913 4662 13954 4670
rect 13913 4636 13928 4662
rect 13935 4636 13954 4662
rect 14018 4658 14049 4670
rect 14064 4658 14167 4670
rect 14179 4660 14205 4686
rect 14220 4681 14250 4692
rect 14282 4688 14344 4704
rect 14282 4686 14328 4688
rect 14282 4670 14344 4686
rect 14356 4670 14362 4718
rect 14365 4710 14445 4718
rect 14365 4708 14384 4710
rect 14399 4708 14433 4710
rect 14365 4692 14445 4708
rect 14365 4670 14384 4692
rect 14399 4676 14429 4692
rect 14457 4686 14463 4760
rect 14466 4686 14485 4830
rect 14500 4686 14506 4830
rect 14515 4760 14528 4830
rect 14580 4826 14602 4830
rect 14573 4804 14602 4818
rect 14655 4804 14671 4818
rect 14709 4814 14715 4816
rect 14722 4814 14830 4830
rect 14837 4814 14843 4816
rect 14851 4814 14866 4830
rect 14932 4824 14951 4827
rect 14573 4802 14671 4804
rect 14698 4802 14866 4814
rect 14881 4804 14897 4818
rect 14932 4805 14954 4824
rect 14964 4818 14980 4819
rect 14963 4816 14980 4818
rect 14964 4811 14980 4816
rect 14954 4804 14960 4805
rect 14963 4804 14992 4811
rect 14881 4803 14992 4804
rect 14881 4802 14998 4803
rect 14557 4794 14608 4802
rect 14655 4794 14689 4802
rect 14557 4782 14582 4794
rect 14589 4782 14608 4794
rect 14662 4792 14689 4794
rect 14698 4792 14919 4802
rect 14954 4799 14960 4802
rect 14662 4788 14919 4792
rect 14557 4774 14608 4782
rect 14655 4774 14919 4788
rect 14963 4794 14998 4802
rect 14509 4726 14528 4760
rect 14573 4766 14602 4774
rect 14573 4760 14590 4766
rect 14573 4758 14607 4760
rect 14655 4758 14671 4774
rect 14672 4764 14880 4774
rect 14881 4764 14897 4774
rect 14945 4770 14960 4785
rect 14963 4782 14964 4794
rect 14971 4782 14998 4794
rect 14963 4774 14998 4782
rect 14963 4773 14992 4774
rect 14683 4760 14897 4764
rect 14698 4758 14897 4760
rect 14932 4760 14945 4770
rect 14963 4760 14980 4773
rect 14932 4758 14980 4760
rect 14574 4754 14607 4758
rect 14570 4752 14607 4754
rect 14570 4751 14637 4752
rect 14570 4746 14601 4751
rect 14607 4746 14637 4751
rect 14570 4742 14637 4746
rect 14543 4739 14637 4742
rect 14543 4732 14592 4739
rect 14543 4726 14573 4732
rect 14592 4727 14597 4732
rect 14509 4710 14589 4726
rect 14601 4718 14637 4739
rect 14698 4734 14887 4758
rect 14932 4757 14979 4758
rect 14945 4752 14979 4757
rect 14713 4731 14887 4734
rect 14706 4728 14887 4731
rect 14915 4751 14979 4752
rect 14509 4708 14528 4710
rect 14543 4708 14577 4710
rect 14509 4692 14589 4708
rect 14509 4686 14528 4692
rect 14225 4660 14328 4670
rect 14179 4658 14328 4660
rect 14349 4658 14384 4670
rect 14018 4656 14180 4658
rect 14030 4636 14049 4656
rect 14064 4654 14094 4656
rect 13913 4628 13954 4636
rect 14036 4632 14049 4636
rect 14101 4640 14180 4656
rect 14212 4656 14384 4658
rect 14212 4640 14291 4656
rect 14298 4654 14328 4656
rect 13876 4618 13905 4628
rect 13919 4618 13948 4628
rect 13963 4618 13993 4632
rect 14036 4618 14079 4632
rect 14101 4628 14291 4640
rect 14356 4636 14362 4656
rect 14086 4618 14116 4628
rect 14117 4618 14275 4628
rect 14279 4618 14309 4628
rect 14313 4618 14343 4632
rect 14371 4618 14384 4656
rect 14456 4670 14485 4686
rect 14499 4670 14528 4686
rect 14543 4676 14573 4692
rect 14601 4670 14607 4718
rect 14610 4712 14629 4718
rect 14644 4712 14674 4720
rect 14610 4704 14674 4712
rect 14610 4688 14690 4704
rect 14706 4697 14768 4728
rect 14784 4697 14846 4728
rect 14915 4726 14964 4751
rect 14979 4726 15009 4742
rect 14878 4712 14908 4720
rect 14915 4718 15025 4726
rect 14878 4704 14923 4712
rect 14610 4686 14629 4688
rect 14644 4686 14690 4688
rect 14610 4670 14690 4686
rect 14717 4684 14752 4697
rect 14793 4694 14830 4697
rect 14793 4692 14835 4694
rect 14722 4681 14752 4684
rect 14731 4677 14738 4681
rect 14738 4676 14739 4677
rect 14697 4670 14707 4676
rect 14456 4662 14491 4670
rect 14456 4636 14457 4662
rect 14464 4636 14491 4662
rect 14399 4618 14429 4632
rect 14456 4628 14491 4636
rect 14493 4662 14534 4670
rect 14493 4636 14508 4662
rect 14515 4636 14534 4662
rect 14598 4658 14629 4670
rect 14644 4658 14747 4670
rect 14759 4660 14785 4686
rect 14800 4681 14830 4692
rect 14862 4688 14924 4704
rect 14862 4686 14908 4688
rect 14862 4670 14924 4686
rect 14936 4670 14942 4718
rect 14945 4710 15025 4718
rect 14945 4708 14964 4710
rect 14979 4708 15013 4710
rect 14945 4692 15025 4708
rect 14945 4670 14964 4692
rect 14979 4676 15009 4692
rect 15037 4686 15043 4760
rect 15046 4686 15065 4830
rect 15080 4686 15086 4830
rect 15095 4760 15108 4830
rect 15160 4826 15182 4830
rect 15153 4804 15182 4818
rect 15235 4804 15251 4818
rect 15289 4814 15295 4816
rect 15302 4814 15410 4830
rect 15417 4814 15423 4816
rect 15431 4814 15446 4830
rect 15512 4824 15531 4827
rect 15153 4802 15251 4804
rect 15278 4802 15446 4814
rect 15461 4804 15477 4818
rect 15512 4805 15534 4824
rect 15544 4818 15560 4819
rect 15543 4816 15560 4818
rect 15544 4811 15560 4816
rect 15534 4804 15540 4805
rect 15543 4804 15572 4811
rect 15461 4803 15572 4804
rect 15461 4802 15578 4803
rect 15137 4794 15188 4802
rect 15235 4794 15269 4802
rect 15137 4782 15162 4794
rect 15169 4782 15188 4794
rect 15242 4792 15269 4794
rect 15278 4792 15499 4802
rect 15534 4799 15540 4802
rect 15242 4788 15499 4792
rect 15137 4774 15188 4782
rect 15235 4774 15499 4788
rect 15543 4794 15578 4802
rect 15089 4726 15108 4760
rect 15153 4766 15182 4774
rect 15153 4760 15170 4766
rect 15153 4758 15187 4760
rect 15235 4758 15251 4774
rect 15252 4764 15460 4774
rect 15461 4764 15477 4774
rect 15525 4770 15540 4785
rect 15543 4782 15544 4794
rect 15551 4782 15578 4794
rect 15543 4774 15578 4782
rect 15543 4773 15572 4774
rect 15263 4760 15477 4764
rect 15278 4758 15477 4760
rect 15512 4760 15525 4770
rect 15543 4760 15560 4773
rect 15512 4758 15560 4760
rect 15154 4754 15187 4758
rect 15150 4752 15187 4754
rect 15150 4751 15217 4752
rect 15150 4746 15181 4751
rect 15187 4746 15217 4751
rect 15150 4742 15217 4746
rect 15123 4739 15217 4742
rect 15123 4732 15172 4739
rect 15123 4726 15153 4732
rect 15172 4727 15177 4732
rect 15089 4710 15169 4726
rect 15181 4718 15217 4739
rect 15278 4734 15467 4758
rect 15512 4757 15559 4758
rect 15525 4752 15559 4757
rect 15293 4731 15467 4734
rect 15286 4728 15467 4731
rect 15495 4751 15559 4752
rect 15089 4708 15108 4710
rect 15123 4708 15157 4710
rect 15089 4692 15169 4708
rect 15089 4686 15108 4692
rect 14805 4660 14908 4670
rect 14759 4658 14908 4660
rect 14929 4658 14964 4670
rect 14598 4656 14760 4658
rect 14610 4636 14629 4656
rect 14644 4654 14674 4656
rect 14493 4628 14534 4636
rect 14616 4632 14629 4636
rect 14681 4640 14760 4656
rect 14792 4656 14964 4658
rect 14792 4640 14871 4656
rect 14878 4654 14908 4656
rect 14456 4618 14485 4628
rect 14499 4618 14528 4628
rect 14543 4618 14573 4632
rect 14616 4618 14659 4632
rect 14681 4628 14871 4640
rect 14936 4636 14942 4656
rect 14666 4618 14696 4628
rect 14697 4618 14855 4628
rect 14859 4618 14889 4628
rect 14893 4618 14923 4632
rect 14951 4618 14964 4656
rect 15036 4670 15065 4686
rect 15079 4670 15108 4686
rect 15123 4676 15153 4692
rect 15181 4670 15187 4718
rect 15190 4712 15209 4718
rect 15224 4712 15254 4720
rect 15190 4704 15254 4712
rect 15190 4688 15270 4704
rect 15286 4697 15348 4728
rect 15364 4697 15426 4728
rect 15495 4726 15544 4751
rect 15559 4726 15589 4742
rect 15458 4712 15488 4720
rect 15495 4718 15605 4726
rect 15458 4704 15503 4712
rect 15190 4686 15209 4688
rect 15224 4686 15270 4688
rect 15190 4670 15270 4686
rect 15297 4684 15332 4697
rect 15373 4694 15410 4697
rect 15373 4692 15415 4694
rect 15302 4681 15332 4684
rect 15311 4677 15318 4681
rect 15318 4676 15319 4677
rect 15277 4670 15287 4676
rect 15036 4662 15071 4670
rect 15036 4636 15037 4662
rect 15044 4636 15071 4662
rect 14979 4618 15009 4632
rect 15036 4628 15071 4636
rect 15073 4662 15114 4670
rect 15073 4636 15088 4662
rect 15095 4636 15114 4662
rect 15178 4658 15209 4670
rect 15224 4658 15327 4670
rect 15339 4660 15365 4686
rect 15380 4681 15410 4692
rect 15442 4688 15504 4704
rect 15442 4686 15488 4688
rect 15442 4670 15504 4686
rect 15516 4670 15522 4718
rect 15525 4710 15605 4718
rect 15525 4708 15544 4710
rect 15559 4708 15593 4710
rect 15525 4692 15605 4708
rect 15525 4670 15544 4692
rect 15559 4676 15589 4692
rect 15617 4686 15623 4760
rect 15626 4686 15645 4830
rect 15660 4686 15666 4830
rect 15675 4760 15688 4830
rect 15740 4826 15762 4830
rect 15733 4804 15762 4818
rect 15815 4804 15831 4818
rect 15869 4814 15875 4816
rect 15882 4814 15990 4830
rect 15997 4814 16003 4816
rect 16011 4814 16026 4830
rect 16092 4824 16111 4827
rect 15733 4802 15831 4804
rect 15858 4802 16026 4814
rect 16041 4804 16057 4818
rect 16092 4805 16114 4824
rect 16124 4818 16140 4819
rect 16123 4816 16140 4818
rect 16124 4811 16140 4816
rect 16114 4804 16120 4805
rect 16123 4804 16152 4811
rect 16041 4803 16152 4804
rect 16041 4802 16158 4803
rect 15717 4794 15768 4802
rect 15815 4794 15849 4802
rect 15717 4782 15742 4794
rect 15749 4782 15768 4794
rect 15822 4792 15849 4794
rect 15858 4792 16079 4802
rect 16114 4799 16120 4802
rect 15822 4788 16079 4792
rect 15717 4774 15768 4782
rect 15815 4774 16079 4788
rect 16123 4794 16158 4802
rect 15669 4726 15688 4760
rect 15733 4766 15762 4774
rect 15733 4760 15750 4766
rect 15733 4758 15767 4760
rect 15815 4758 15831 4774
rect 15832 4764 16040 4774
rect 16041 4764 16057 4774
rect 16105 4770 16120 4785
rect 16123 4782 16124 4794
rect 16131 4782 16158 4794
rect 16123 4774 16158 4782
rect 16123 4773 16152 4774
rect 15843 4760 16057 4764
rect 15858 4758 16057 4760
rect 16092 4760 16105 4770
rect 16123 4760 16140 4773
rect 16092 4758 16140 4760
rect 15734 4754 15767 4758
rect 15730 4752 15767 4754
rect 15730 4751 15797 4752
rect 15730 4746 15761 4751
rect 15767 4746 15797 4751
rect 15730 4742 15797 4746
rect 15703 4739 15797 4742
rect 15703 4732 15752 4739
rect 15703 4726 15733 4732
rect 15752 4727 15757 4732
rect 15669 4710 15749 4726
rect 15761 4718 15797 4739
rect 15858 4734 16047 4758
rect 16092 4757 16139 4758
rect 16105 4752 16139 4757
rect 15873 4731 16047 4734
rect 15866 4728 16047 4731
rect 16075 4751 16139 4752
rect 15669 4708 15688 4710
rect 15703 4708 15737 4710
rect 15669 4692 15749 4708
rect 15669 4686 15688 4692
rect 15385 4660 15488 4670
rect 15339 4658 15488 4660
rect 15509 4658 15544 4670
rect 15178 4656 15340 4658
rect 15190 4636 15209 4656
rect 15224 4654 15254 4656
rect 15073 4628 15114 4636
rect 15196 4632 15209 4636
rect 15261 4640 15340 4656
rect 15372 4656 15544 4658
rect 15372 4640 15451 4656
rect 15458 4654 15488 4656
rect 15036 4618 15065 4628
rect 15079 4618 15108 4628
rect 15123 4618 15153 4632
rect 15196 4618 15239 4632
rect 15261 4628 15451 4640
rect 15516 4636 15522 4656
rect 15246 4618 15276 4628
rect 15277 4618 15435 4628
rect 15439 4618 15469 4628
rect 15473 4618 15503 4632
rect 15531 4618 15544 4656
rect 15616 4670 15645 4686
rect 15659 4670 15688 4686
rect 15703 4676 15733 4692
rect 15761 4670 15767 4718
rect 15770 4712 15789 4718
rect 15804 4712 15834 4720
rect 15770 4704 15834 4712
rect 15770 4688 15850 4704
rect 15866 4697 15928 4728
rect 15944 4697 16006 4728
rect 16075 4726 16124 4751
rect 16139 4726 16169 4742
rect 16038 4712 16068 4720
rect 16075 4718 16185 4726
rect 16038 4704 16083 4712
rect 15770 4686 15789 4688
rect 15804 4686 15850 4688
rect 15770 4670 15850 4686
rect 15877 4684 15912 4697
rect 15953 4694 15990 4697
rect 15953 4692 15995 4694
rect 15882 4681 15912 4684
rect 15891 4677 15898 4681
rect 15898 4676 15899 4677
rect 15857 4670 15867 4676
rect 15616 4662 15651 4670
rect 15616 4636 15617 4662
rect 15624 4636 15651 4662
rect 15559 4618 15589 4632
rect 15616 4628 15651 4636
rect 15653 4662 15694 4670
rect 15653 4636 15668 4662
rect 15675 4636 15694 4662
rect 15758 4658 15789 4670
rect 15804 4658 15907 4670
rect 15919 4660 15945 4686
rect 15960 4681 15990 4692
rect 16022 4688 16084 4704
rect 16022 4686 16068 4688
rect 16022 4670 16084 4686
rect 16096 4670 16102 4718
rect 16105 4710 16185 4718
rect 16105 4708 16124 4710
rect 16139 4708 16173 4710
rect 16105 4692 16185 4708
rect 16105 4670 16124 4692
rect 16139 4676 16169 4692
rect 16197 4686 16203 4760
rect 16206 4686 16225 4830
rect 16240 4686 16246 4830
rect 16255 4760 16268 4830
rect 16320 4826 16342 4830
rect 16313 4804 16342 4818
rect 16395 4804 16411 4818
rect 16449 4814 16455 4816
rect 16462 4814 16570 4830
rect 16577 4814 16583 4816
rect 16591 4814 16606 4830
rect 16672 4824 16691 4827
rect 16313 4802 16411 4804
rect 16438 4802 16606 4814
rect 16621 4804 16637 4818
rect 16672 4805 16694 4824
rect 16704 4818 16720 4819
rect 16703 4816 16720 4818
rect 16704 4811 16720 4816
rect 16694 4804 16700 4805
rect 16703 4804 16732 4811
rect 16621 4803 16732 4804
rect 16621 4802 16738 4803
rect 16297 4794 16348 4802
rect 16395 4794 16429 4802
rect 16297 4782 16322 4794
rect 16329 4782 16348 4794
rect 16402 4792 16429 4794
rect 16438 4792 16659 4802
rect 16694 4799 16700 4802
rect 16402 4788 16659 4792
rect 16297 4774 16348 4782
rect 16395 4774 16659 4788
rect 16703 4794 16738 4802
rect 16249 4726 16268 4760
rect 16313 4766 16342 4774
rect 16313 4760 16330 4766
rect 16313 4758 16347 4760
rect 16395 4758 16411 4774
rect 16412 4764 16620 4774
rect 16621 4764 16637 4774
rect 16685 4770 16700 4785
rect 16703 4782 16704 4794
rect 16711 4782 16738 4794
rect 16703 4774 16738 4782
rect 16703 4773 16732 4774
rect 16423 4760 16637 4764
rect 16438 4758 16637 4760
rect 16672 4760 16685 4770
rect 16703 4760 16720 4773
rect 16672 4758 16720 4760
rect 16314 4754 16347 4758
rect 16310 4752 16347 4754
rect 16310 4751 16377 4752
rect 16310 4746 16341 4751
rect 16347 4746 16377 4751
rect 16310 4742 16377 4746
rect 16283 4739 16377 4742
rect 16283 4732 16332 4739
rect 16283 4726 16313 4732
rect 16332 4727 16337 4732
rect 16249 4710 16329 4726
rect 16341 4718 16377 4739
rect 16438 4734 16627 4758
rect 16672 4757 16719 4758
rect 16685 4752 16719 4757
rect 16453 4731 16627 4734
rect 16446 4728 16627 4731
rect 16655 4751 16719 4752
rect 16249 4708 16268 4710
rect 16283 4708 16317 4710
rect 16249 4692 16329 4708
rect 16249 4686 16268 4692
rect 15965 4660 16068 4670
rect 15919 4658 16068 4660
rect 16089 4658 16124 4670
rect 15758 4656 15920 4658
rect 15770 4636 15789 4656
rect 15804 4654 15834 4656
rect 15653 4628 15694 4636
rect 15776 4632 15789 4636
rect 15841 4640 15920 4656
rect 15952 4656 16124 4658
rect 15952 4640 16031 4656
rect 16038 4654 16068 4656
rect 15616 4618 15645 4628
rect 15659 4618 15688 4628
rect 15703 4618 15733 4632
rect 15776 4618 15819 4632
rect 15841 4628 16031 4640
rect 16096 4636 16102 4656
rect 15826 4618 15856 4628
rect 15857 4618 16015 4628
rect 16019 4618 16049 4628
rect 16053 4618 16083 4632
rect 16111 4618 16124 4656
rect 16196 4670 16225 4686
rect 16239 4670 16268 4686
rect 16283 4676 16313 4692
rect 16341 4670 16347 4718
rect 16350 4712 16369 4718
rect 16384 4712 16414 4720
rect 16350 4704 16414 4712
rect 16350 4688 16430 4704
rect 16446 4697 16508 4728
rect 16524 4697 16586 4728
rect 16655 4726 16704 4751
rect 16719 4726 16749 4742
rect 16618 4712 16648 4720
rect 16655 4718 16765 4726
rect 16618 4704 16663 4712
rect 16350 4686 16369 4688
rect 16384 4686 16430 4688
rect 16350 4670 16430 4686
rect 16457 4684 16492 4697
rect 16533 4694 16570 4697
rect 16533 4692 16575 4694
rect 16462 4681 16492 4684
rect 16471 4677 16478 4681
rect 16478 4676 16479 4677
rect 16437 4670 16447 4676
rect 16196 4662 16231 4670
rect 16196 4636 16197 4662
rect 16204 4636 16231 4662
rect 16139 4618 16169 4632
rect 16196 4628 16231 4636
rect 16233 4662 16274 4670
rect 16233 4636 16248 4662
rect 16255 4636 16274 4662
rect 16338 4658 16369 4670
rect 16384 4658 16487 4670
rect 16499 4660 16525 4686
rect 16540 4681 16570 4692
rect 16602 4688 16664 4704
rect 16602 4686 16648 4688
rect 16602 4670 16664 4686
rect 16676 4670 16682 4718
rect 16685 4710 16765 4718
rect 16685 4708 16704 4710
rect 16719 4708 16753 4710
rect 16685 4692 16765 4708
rect 16685 4670 16704 4692
rect 16719 4676 16749 4692
rect 16777 4686 16783 4760
rect 16786 4686 16805 4830
rect 16820 4686 16826 4830
rect 16835 4760 16848 4830
rect 16900 4826 16922 4830
rect 16893 4804 16922 4818
rect 16975 4804 16991 4818
rect 17029 4814 17035 4816
rect 17042 4814 17150 4830
rect 17157 4814 17163 4816
rect 17171 4814 17186 4830
rect 17252 4824 17271 4827
rect 16893 4802 16991 4804
rect 17018 4802 17186 4814
rect 17201 4804 17217 4818
rect 17252 4805 17274 4824
rect 17284 4818 17300 4819
rect 17283 4816 17300 4818
rect 17284 4811 17300 4816
rect 17274 4804 17280 4805
rect 17283 4804 17312 4811
rect 17201 4803 17312 4804
rect 17201 4802 17318 4803
rect 16877 4794 16928 4802
rect 16975 4794 17009 4802
rect 16877 4782 16902 4794
rect 16909 4782 16928 4794
rect 16982 4792 17009 4794
rect 17018 4792 17239 4802
rect 17274 4799 17280 4802
rect 16982 4788 17239 4792
rect 16877 4774 16928 4782
rect 16975 4774 17239 4788
rect 17283 4794 17318 4802
rect 16829 4726 16848 4760
rect 16893 4766 16922 4774
rect 16893 4760 16910 4766
rect 16893 4758 16927 4760
rect 16975 4758 16991 4774
rect 16992 4764 17200 4774
rect 17201 4764 17217 4774
rect 17265 4770 17280 4785
rect 17283 4782 17284 4794
rect 17291 4782 17318 4794
rect 17283 4774 17318 4782
rect 17283 4773 17312 4774
rect 17003 4760 17217 4764
rect 17018 4758 17217 4760
rect 17252 4760 17265 4770
rect 17283 4760 17300 4773
rect 17252 4758 17300 4760
rect 16894 4754 16927 4758
rect 16890 4752 16927 4754
rect 16890 4751 16957 4752
rect 16890 4746 16921 4751
rect 16927 4746 16957 4751
rect 16890 4742 16957 4746
rect 16863 4739 16957 4742
rect 16863 4732 16912 4739
rect 16863 4726 16893 4732
rect 16912 4727 16917 4732
rect 16829 4710 16909 4726
rect 16921 4718 16957 4739
rect 17018 4734 17207 4758
rect 17252 4757 17299 4758
rect 17265 4752 17299 4757
rect 17033 4731 17207 4734
rect 17026 4728 17207 4731
rect 17235 4751 17299 4752
rect 16829 4708 16848 4710
rect 16863 4708 16897 4710
rect 16829 4692 16909 4708
rect 16829 4686 16848 4692
rect 16545 4660 16648 4670
rect 16499 4658 16648 4660
rect 16669 4658 16704 4670
rect 16338 4656 16500 4658
rect 16350 4636 16369 4656
rect 16384 4654 16414 4656
rect 16233 4628 16274 4636
rect 16356 4632 16369 4636
rect 16421 4640 16500 4656
rect 16532 4656 16704 4658
rect 16532 4640 16611 4656
rect 16618 4654 16648 4656
rect 16196 4618 16225 4628
rect 16239 4618 16268 4628
rect 16283 4618 16313 4632
rect 16356 4618 16399 4632
rect 16421 4628 16611 4640
rect 16676 4636 16682 4656
rect 16406 4618 16436 4628
rect 16437 4618 16595 4628
rect 16599 4618 16629 4628
rect 16633 4618 16663 4632
rect 16691 4618 16704 4656
rect 16776 4670 16805 4686
rect 16819 4670 16848 4686
rect 16863 4676 16893 4692
rect 16921 4670 16927 4718
rect 16930 4712 16949 4718
rect 16964 4712 16994 4720
rect 16930 4704 16994 4712
rect 16930 4688 17010 4704
rect 17026 4697 17088 4728
rect 17104 4697 17166 4728
rect 17235 4726 17284 4751
rect 17299 4726 17329 4742
rect 17198 4712 17228 4720
rect 17235 4718 17345 4726
rect 17198 4704 17243 4712
rect 16930 4686 16949 4688
rect 16964 4686 17010 4688
rect 16930 4670 17010 4686
rect 17037 4684 17072 4697
rect 17113 4694 17150 4697
rect 17113 4692 17155 4694
rect 17042 4681 17072 4684
rect 17051 4677 17058 4681
rect 17058 4676 17059 4677
rect 17017 4670 17027 4676
rect 16776 4662 16811 4670
rect 16776 4636 16777 4662
rect 16784 4636 16811 4662
rect 16719 4618 16749 4632
rect 16776 4628 16811 4636
rect 16813 4662 16854 4670
rect 16813 4636 16828 4662
rect 16835 4636 16854 4662
rect 16918 4658 16949 4670
rect 16964 4658 17067 4670
rect 17079 4660 17105 4686
rect 17120 4681 17150 4692
rect 17182 4688 17244 4704
rect 17182 4686 17228 4688
rect 17182 4670 17244 4686
rect 17256 4670 17262 4718
rect 17265 4710 17345 4718
rect 17265 4708 17284 4710
rect 17299 4708 17333 4710
rect 17265 4692 17345 4708
rect 17265 4670 17284 4692
rect 17299 4676 17329 4692
rect 17357 4686 17363 4760
rect 17366 4686 17385 4830
rect 17400 4686 17406 4830
rect 17415 4760 17428 4830
rect 17480 4826 17502 4830
rect 17473 4804 17502 4818
rect 17555 4804 17571 4818
rect 17609 4814 17615 4816
rect 17622 4814 17730 4830
rect 17737 4814 17743 4816
rect 17751 4814 17766 4830
rect 17832 4824 17851 4827
rect 17473 4802 17571 4804
rect 17598 4802 17766 4814
rect 17781 4804 17797 4818
rect 17832 4805 17854 4824
rect 17864 4818 17880 4819
rect 17863 4816 17880 4818
rect 17864 4811 17880 4816
rect 17854 4804 17860 4805
rect 17863 4804 17892 4811
rect 17781 4803 17892 4804
rect 17781 4802 17898 4803
rect 17457 4794 17508 4802
rect 17555 4794 17589 4802
rect 17457 4782 17482 4794
rect 17489 4782 17508 4794
rect 17562 4792 17589 4794
rect 17598 4792 17819 4802
rect 17854 4799 17860 4802
rect 17562 4788 17819 4792
rect 17457 4774 17508 4782
rect 17555 4774 17819 4788
rect 17863 4794 17898 4802
rect 17409 4726 17428 4760
rect 17473 4766 17502 4774
rect 17473 4760 17490 4766
rect 17473 4758 17507 4760
rect 17555 4758 17571 4774
rect 17572 4764 17780 4774
rect 17781 4764 17797 4774
rect 17845 4770 17860 4785
rect 17863 4782 17864 4794
rect 17871 4782 17898 4794
rect 17863 4774 17898 4782
rect 17863 4773 17892 4774
rect 17583 4760 17797 4764
rect 17598 4758 17797 4760
rect 17832 4760 17845 4770
rect 17863 4760 17880 4773
rect 17832 4758 17880 4760
rect 17474 4754 17507 4758
rect 17470 4752 17507 4754
rect 17470 4751 17537 4752
rect 17470 4746 17501 4751
rect 17507 4746 17537 4751
rect 17470 4742 17537 4746
rect 17443 4739 17537 4742
rect 17443 4732 17492 4739
rect 17443 4726 17473 4732
rect 17492 4727 17497 4732
rect 17409 4710 17489 4726
rect 17501 4718 17537 4739
rect 17598 4734 17787 4758
rect 17832 4757 17879 4758
rect 17845 4752 17879 4757
rect 17613 4731 17787 4734
rect 17606 4728 17787 4731
rect 17815 4751 17879 4752
rect 17409 4708 17428 4710
rect 17443 4708 17477 4710
rect 17409 4692 17489 4708
rect 17409 4686 17428 4692
rect 17125 4660 17228 4670
rect 17079 4658 17228 4660
rect 17249 4658 17284 4670
rect 16918 4656 17080 4658
rect 16930 4636 16949 4656
rect 16964 4654 16994 4656
rect 16813 4628 16854 4636
rect 16936 4632 16949 4636
rect 17001 4640 17080 4656
rect 17112 4656 17284 4658
rect 17112 4640 17191 4656
rect 17198 4654 17228 4656
rect 16776 4618 16805 4628
rect 16819 4618 16848 4628
rect 16863 4618 16893 4632
rect 16936 4618 16979 4632
rect 17001 4628 17191 4640
rect 17256 4636 17262 4656
rect 16986 4618 17016 4628
rect 17017 4618 17175 4628
rect 17179 4618 17209 4628
rect 17213 4618 17243 4632
rect 17271 4618 17284 4656
rect 17356 4670 17385 4686
rect 17399 4670 17428 4686
rect 17443 4676 17473 4692
rect 17501 4670 17507 4718
rect 17510 4712 17529 4718
rect 17544 4712 17574 4720
rect 17510 4704 17574 4712
rect 17510 4688 17590 4704
rect 17606 4697 17668 4728
rect 17684 4697 17746 4728
rect 17815 4726 17864 4751
rect 17879 4726 17909 4742
rect 17778 4712 17808 4720
rect 17815 4718 17925 4726
rect 17778 4704 17823 4712
rect 17510 4686 17529 4688
rect 17544 4686 17590 4688
rect 17510 4670 17590 4686
rect 17617 4684 17652 4697
rect 17693 4694 17730 4697
rect 17693 4692 17735 4694
rect 17622 4681 17652 4684
rect 17631 4677 17638 4681
rect 17638 4676 17639 4677
rect 17597 4670 17607 4676
rect 17356 4662 17391 4670
rect 17356 4636 17357 4662
rect 17364 4636 17391 4662
rect 17299 4618 17329 4632
rect 17356 4628 17391 4636
rect 17393 4662 17434 4670
rect 17393 4636 17408 4662
rect 17415 4636 17434 4662
rect 17498 4658 17529 4670
rect 17544 4658 17647 4670
rect 17659 4660 17685 4686
rect 17700 4681 17730 4692
rect 17762 4688 17824 4704
rect 17762 4686 17808 4688
rect 17762 4670 17824 4686
rect 17836 4670 17842 4718
rect 17845 4710 17925 4718
rect 17845 4708 17864 4710
rect 17879 4708 17913 4710
rect 17845 4692 17925 4708
rect 17845 4670 17864 4692
rect 17879 4676 17909 4692
rect 17937 4686 17943 4760
rect 17946 4686 17965 4830
rect 17980 4686 17986 4830
rect 17995 4760 18008 4830
rect 18060 4826 18082 4830
rect 18053 4804 18082 4818
rect 18135 4804 18151 4818
rect 18189 4814 18195 4816
rect 18202 4814 18310 4830
rect 18317 4814 18323 4816
rect 18331 4814 18346 4830
rect 18412 4824 18431 4827
rect 18053 4802 18151 4804
rect 18178 4802 18346 4814
rect 18361 4804 18377 4818
rect 18412 4805 18434 4824
rect 18444 4818 18460 4819
rect 18443 4816 18460 4818
rect 18444 4811 18460 4816
rect 18434 4804 18440 4805
rect 18443 4804 18472 4811
rect 18361 4803 18472 4804
rect 18361 4802 18478 4803
rect 18037 4794 18088 4802
rect 18135 4794 18169 4802
rect 18037 4782 18062 4794
rect 18069 4782 18088 4794
rect 18142 4792 18169 4794
rect 18178 4792 18399 4802
rect 18434 4799 18440 4802
rect 18142 4788 18399 4792
rect 18037 4774 18088 4782
rect 18135 4774 18399 4788
rect 18443 4794 18478 4802
rect 17989 4726 18008 4760
rect 18053 4766 18082 4774
rect 18053 4760 18070 4766
rect 18053 4758 18087 4760
rect 18135 4758 18151 4774
rect 18152 4764 18360 4774
rect 18361 4764 18377 4774
rect 18425 4770 18440 4785
rect 18443 4782 18444 4794
rect 18451 4782 18478 4794
rect 18443 4774 18478 4782
rect 18443 4773 18472 4774
rect 18163 4760 18377 4764
rect 18178 4758 18377 4760
rect 18412 4760 18425 4770
rect 18443 4760 18460 4773
rect 18412 4758 18460 4760
rect 18054 4754 18087 4758
rect 18050 4752 18087 4754
rect 18050 4751 18117 4752
rect 18050 4746 18081 4751
rect 18087 4746 18117 4751
rect 18050 4742 18117 4746
rect 18023 4739 18117 4742
rect 18023 4732 18072 4739
rect 18023 4726 18053 4732
rect 18072 4727 18077 4732
rect 17989 4710 18069 4726
rect 18081 4718 18117 4739
rect 18178 4734 18367 4758
rect 18412 4757 18459 4758
rect 18425 4752 18459 4757
rect 18193 4731 18367 4734
rect 18186 4728 18367 4731
rect 18395 4751 18459 4752
rect 17989 4708 18008 4710
rect 18023 4708 18057 4710
rect 17989 4692 18069 4708
rect 17989 4686 18008 4692
rect 17705 4660 17808 4670
rect 17659 4658 17808 4660
rect 17829 4658 17864 4670
rect 17498 4656 17660 4658
rect 17510 4636 17529 4656
rect 17544 4654 17574 4656
rect 17393 4628 17434 4636
rect 17516 4632 17529 4636
rect 17581 4640 17660 4656
rect 17692 4656 17864 4658
rect 17692 4640 17771 4656
rect 17778 4654 17808 4656
rect 17356 4618 17385 4628
rect 17399 4618 17428 4628
rect 17443 4618 17473 4632
rect 17516 4618 17559 4632
rect 17581 4628 17771 4640
rect 17836 4636 17842 4656
rect 17566 4618 17596 4628
rect 17597 4618 17755 4628
rect 17759 4618 17789 4628
rect 17793 4618 17823 4632
rect 17851 4618 17864 4656
rect 17936 4670 17965 4686
rect 17979 4670 18008 4686
rect 18023 4676 18053 4692
rect 18081 4670 18087 4718
rect 18090 4712 18109 4718
rect 18124 4712 18154 4720
rect 18090 4704 18154 4712
rect 18090 4688 18170 4704
rect 18186 4697 18248 4728
rect 18264 4697 18326 4728
rect 18395 4726 18444 4751
rect 18459 4726 18489 4742
rect 18358 4712 18388 4720
rect 18395 4718 18505 4726
rect 18358 4704 18403 4712
rect 18090 4686 18109 4688
rect 18124 4686 18170 4688
rect 18090 4670 18170 4686
rect 18197 4684 18232 4697
rect 18273 4694 18310 4697
rect 18273 4692 18315 4694
rect 18202 4681 18232 4684
rect 18211 4677 18218 4681
rect 18218 4676 18219 4677
rect 18177 4670 18187 4676
rect 17936 4662 17971 4670
rect 17936 4636 17937 4662
rect 17944 4636 17971 4662
rect 17879 4618 17909 4632
rect 17936 4628 17971 4636
rect 17973 4662 18014 4670
rect 17973 4636 17988 4662
rect 17995 4636 18014 4662
rect 18078 4658 18109 4670
rect 18124 4658 18227 4670
rect 18239 4660 18265 4686
rect 18280 4681 18310 4692
rect 18342 4688 18404 4704
rect 18342 4686 18388 4688
rect 18342 4670 18404 4686
rect 18416 4670 18422 4718
rect 18425 4710 18505 4718
rect 18425 4708 18444 4710
rect 18459 4708 18493 4710
rect 18425 4692 18505 4708
rect 18425 4670 18444 4692
rect 18459 4676 18489 4692
rect 18517 4686 18523 4760
rect 18532 4686 18545 4830
rect 18285 4660 18388 4670
rect 18239 4658 18388 4660
rect 18409 4658 18444 4670
rect 18078 4656 18240 4658
rect 18090 4636 18109 4656
rect 18124 4654 18154 4656
rect 17973 4628 18014 4636
rect 18096 4632 18109 4636
rect 18161 4640 18240 4656
rect 18272 4656 18444 4658
rect 18272 4640 18351 4656
rect 18358 4654 18388 4656
rect 17936 4618 17965 4628
rect 17979 4618 18008 4628
rect 18023 4618 18053 4632
rect 18096 4618 18139 4632
rect 18161 4628 18351 4640
rect 18416 4636 18422 4656
rect 18146 4618 18176 4628
rect 18177 4618 18335 4628
rect 18339 4618 18369 4628
rect 18373 4618 18403 4632
rect 18431 4618 18444 4656
rect 18516 4670 18545 4686
rect 18516 4662 18551 4670
rect 18516 4636 18517 4662
rect 18524 4636 18551 4662
rect 18459 4618 18489 4632
rect 18516 4628 18551 4636
rect 18516 4618 18545 4628
rect -1 4612 18545 4618
rect 0 4604 18545 4612
rect 15 4574 28 4604
rect 43 4590 73 4604
rect 116 4590 159 4604
rect 166 4590 386 4604
rect 393 4590 423 4604
rect 83 4576 98 4588
rect 117 4576 130 4590
rect 198 4586 351 4590
rect 80 4574 102 4576
rect 180 4574 372 4586
rect 451 4574 464 4604
rect 479 4590 509 4604
rect 546 4574 565 4604
rect 580 4574 586 4604
rect 595 4574 608 4604
rect 623 4590 653 4604
rect 696 4590 739 4604
rect 746 4590 966 4604
rect 973 4590 1003 4604
rect 663 4576 678 4588
rect 697 4576 710 4590
rect 778 4586 931 4590
rect 660 4574 682 4576
rect 760 4574 952 4586
rect 1031 4574 1044 4604
rect 1059 4590 1089 4604
rect 1126 4574 1145 4604
rect 1160 4574 1166 4604
rect 1175 4574 1188 4604
rect 1203 4590 1233 4604
rect 1276 4590 1319 4604
rect 1326 4590 1546 4604
rect 1553 4590 1583 4604
rect 1243 4576 1258 4588
rect 1277 4576 1290 4590
rect 1358 4586 1511 4590
rect 1240 4574 1262 4576
rect 1340 4574 1532 4586
rect 1611 4574 1624 4604
rect 1639 4590 1669 4604
rect 1706 4574 1725 4604
rect 1740 4574 1746 4604
rect 1755 4574 1768 4604
rect 1783 4590 1813 4604
rect 1856 4590 1899 4604
rect 1906 4590 2126 4604
rect 2133 4590 2163 4604
rect 1823 4576 1838 4588
rect 1857 4576 1870 4590
rect 1938 4586 2091 4590
rect 1820 4574 1842 4576
rect 1920 4574 2112 4586
rect 2191 4574 2204 4604
rect 2219 4590 2249 4604
rect 2286 4574 2305 4604
rect 2320 4574 2326 4604
rect 2335 4574 2348 4604
rect 2363 4590 2393 4604
rect 2436 4590 2479 4604
rect 2486 4590 2706 4604
rect 2713 4590 2743 4604
rect 2403 4576 2418 4588
rect 2437 4576 2450 4590
rect 2518 4586 2671 4590
rect 2400 4574 2422 4576
rect 2500 4574 2692 4586
rect 2771 4574 2784 4604
rect 2799 4590 2829 4604
rect 2866 4574 2885 4604
rect 2900 4574 2906 4604
rect 2915 4574 2928 4604
rect 2943 4590 2973 4604
rect 3016 4590 3059 4604
rect 3066 4590 3286 4604
rect 3293 4590 3323 4604
rect 2983 4576 2998 4588
rect 3017 4576 3030 4590
rect 3098 4586 3251 4590
rect 2980 4574 3002 4576
rect 3080 4574 3272 4586
rect 3351 4574 3364 4604
rect 3379 4590 3409 4604
rect 3446 4574 3465 4604
rect 3480 4574 3486 4604
rect 3495 4574 3508 4604
rect 3523 4590 3553 4604
rect 3596 4590 3639 4604
rect 3646 4590 3866 4604
rect 3873 4590 3903 4604
rect 3563 4576 3578 4588
rect 3597 4576 3610 4590
rect 3678 4586 3831 4590
rect 3560 4574 3582 4576
rect 3660 4574 3852 4586
rect 3931 4574 3944 4604
rect 3959 4590 3989 4604
rect 4026 4574 4045 4604
rect 4060 4574 4066 4604
rect 4075 4574 4088 4604
rect 4103 4590 4133 4604
rect 4176 4590 4219 4604
rect 4226 4590 4446 4604
rect 4453 4590 4483 4604
rect 4143 4576 4158 4588
rect 4177 4576 4190 4590
rect 4258 4586 4411 4590
rect 4140 4574 4162 4576
rect 4240 4574 4432 4586
rect 4511 4574 4524 4604
rect 4539 4590 4569 4604
rect 4606 4574 4625 4604
rect 4640 4574 4646 4604
rect 4655 4574 4668 4604
rect 4683 4590 4713 4604
rect 4756 4590 4799 4604
rect 4806 4590 5026 4604
rect 5033 4590 5063 4604
rect 4723 4576 4738 4588
rect 4757 4576 4770 4590
rect 4838 4586 4991 4590
rect 4720 4574 4742 4576
rect 4820 4574 5012 4586
rect 5091 4574 5104 4604
rect 5119 4590 5149 4604
rect 5186 4574 5205 4604
rect 5220 4574 5226 4604
rect 5235 4574 5248 4604
rect 5263 4590 5293 4604
rect 5336 4590 5379 4604
rect 5386 4590 5606 4604
rect 5613 4590 5643 4604
rect 5303 4576 5318 4588
rect 5337 4576 5350 4590
rect 5418 4586 5571 4590
rect 5300 4574 5322 4576
rect 5400 4574 5592 4586
rect 5671 4574 5684 4604
rect 5699 4590 5729 4604
rect 5766 4574 5785 4604
rect 5800 4574 5806 4604
rect 5815 4574 5828 4604
rect 5843 4590 5873 4604
rect 5916 4590 5959 4604
rect 5966 4590 6186 4604
rect 6193 4590 6223 4604
rect 5883 4576 5898 4588
rect 5917 4576 5930 4590
rect 5998 4586 6151 4590
rect 5880 4574 5902 4576
rect 5980 4574 6172 4586
rect 6251 4574 6264 4604
rect 6279 4590 6309 4604
rect 6346 4574 6365 4604
rect 6380 4574 6386 4604
rect 6395 4574 6408 4604
rect 6423 4590 6453 4604
rect 6496 4590 6539 4604
rect 6546 4590 6766 4604
rect 6773 4590 6803 4604
rect 6463 4576 6478 4588
rect 6497 4576 6510 4590
rect 6578 4586 6731 4590
rect 6460 4574 6482 4576
rect 6560 4574 6752 4586
rect 6831 4574 6844 4604
rect 6859 4590 6889 4604
rect 6926 4574 6945 4604
rect 6960 4574 6966 4604
rect 6975 4574 6988 4604
rect 7003 4590 7033 4604
rect 7076 4590 7119 4604
rect 7126 4590 7346 4604
rect 7353 4590 7383 4604
rect 7043 4576 7058 4588
rect 7077 4576 7090 4590
rect 7158 4586 7311 4590
rect 7040 4574 7062 4576
rect 7140 4574 7332 4586
rect 7411 4574 7424 4604
rect 7439 4590 7469 4604
rect 7506 4574 7525 4604
rect 7540 4574 7546 4604
rect 7555 4574 7568 4604
rect 7583 4590 7613 4604
rect 7656 4590 7699 4604
rect 7706 4590 7926 4604
rect 7933 4590 7963 4604
rect 7623 4576 7638 4588
rect 7657 4576 7670 4590
rect 7738 4586 7891 4590
rect 7620 4574 7642 4576
rect 7720 4574 7912 4586
rect 7991 4574 8004 4604
rect 8019 4590 8049 4604
rect 8086 4574 8105 4604
rect 8120 4574 8126 4604
rect 8135 4574 8148 4604
rect 8163 4590 8193 4604
rect 8236 4590 8279 4604
rect 8286 4590 8506 4604
rect 8513 4590 8543 4604
rect 8203 4576 8218 4588
rect 8237 4576 8250 4590
rect 8318 4586 8471 4590
rect 8200 4574 8222 4576
rect 8300 4574 8492 4586
rect 8571 4574 8584 4604
rect 8599 4590 8629 4604
rect 8666 4574 8685 4604
rect 8700 4574 8706 4604
rect 8715 4574 8728 4604
rect 8743 4590 8773 4604
rect 8816 4590 8859 4604
rect 8866 4590 9086 4604
rect 9093 4590 9123 4604
rect 8783 4576 8798 4588
rect 8817 4576 8830 4590
rect 8898 4586 9051 4590
rect 8780 4574 8802 4576
rect 8880 4574 9072 4586
rect 9151 4574 9164 4604
rect 9179 4590 9209 4604
rect 9246 4574 9265 4604
rect 9280 4574 9286 4604
rect 9295 4574 9308 4604
rect 9323 4590 9353 4604
rect 9396 4590 9439 4604
rect 9446 4590 9666 4604
rect 9673 4590 9703 4604
rect 9363 4576 9378 4588
rect 9397 4576 9410 4590
rect 9478 4586 9631 4590
rect 9360 4574 9382 4576
rect 9460 4574 9652 4586
rect 9731 4574 9744 4604
rect 9759 4590 9789 4604
rect 9826 4574 9845 4604
rect 9860 4574 9866 4604
rect 9875 4574 9888 4604
rect 9903 4590 9933 4604
rect 9976 4590 10019 4604
rect 10026 4590 10246 4604
rect 10253 4590 10283 4604
rect 9943 4576 9958 4588
rect 9977 4576 9990 4590
rect 10058 4586 10211 4590
rect 9940 4574 9962 4576
rect 10040 4574 10232 4586
rect 10311 4574 10324 4604
rect 10339 4590 10369 4604
rect 10406 4574 10425 4604
rect 10440 4574 10446 4604
rect 10455 4574 10468 4604
rect 10483 4590 10513 4604
rect 10556 4590 10599 4604
rect 10606 4590 10826 4604
rect 10833 4590 10863 4604
rect 10523 4576 10538 4588
rect 10557 4576 10570 4590
rect 10638 4586 10791 4590
rect 10520 4574 10542 4576
rect 10620 4574 10812 4586
rect 10891 4574 10904 4604
rect 10919 4590 10949 4604
rect 10986 4574 11005 4604
rect 11020 4574 11026 4604
rect 11035 4574 11048 4604
rect 11063 4590 11093 4604
rect 11136 4590 11179 4604
rect 11186 4590 11406 4604
rect 11413 4590 11443 4604
rect 11103 4576 11118 4588
rect 11137 4576 11150 4590
rect 11218 4586 11371 4590
rect 11100 4574 11122 4576
rect 11200 4574 11392 4586
rect 11471 4574 11484 4604
rect 11499 4590 11529 4604
rect 11566 4574 11585 4604
rect 11600 4574 11606 4604
rect 11615 4574 11628 4604
rect 11643 4590 11673 4604
rect 11716 4590 11759 4604
rect 11766 4590 11986 4604
rect 11993 4590 12023 4604
rect 11683 4576 11698 4588
rect 11717 4576 11730 4590
rect 11798 4586 11951 4590
rect 11680 4574 11702 4576
rect 11780 4574 11972 4586
rect 12051 4574 12064 4604
rect 12079 4590 12109 4604
rect 12146 4574 12165 4604
rect 12180 4574 12186 4604
rect 12195 4574 12208 4604
rect 12223 4590 12253 4604
rect 12296 4590 12339 4604
rect 12346 4590 12566 4604
rect 12573 4590 12603 4604
rect 12263 4576 12278 4588
rect 12297 4576 12310 4590
rect 12378 4586 12531 4590
rect 12260 4574 12282 4576
rect 12360 4574 12552 4586
rect 12631 4574 12644 4604
rect 12659 4590 12689 4604
rect 12726 4574 12745 4604
rect 12760 4574 12766 4604
rect 12775 4574 12788 4604
rect 12803 4590 12833 4604
rect 12876 4590 12919 4604
rect 12926 4590 13146 4604
rect 13153 4590 13183 4604
rect 12843 4576 12858 4588
rect 12877 4576 12890 4590
rect 12958 4586 13111 4590
rect 12840 4574 12862 4576
rect 12940 4574 13132 4586
rect 13211 4574 13224 4604
rect 13239 4590 13269 4604
rect 13306 4574 13325 4604
rect 13340 4574 13346 4604
rect 13355 4574 13368 4604
rect 13383 4590 13413 4604
rect 13456 4590 13499 4604
rect 13506 4590 13726 4604
rect 13733 4590 13763 4604
rect 13423 4576 13438 4588
rect 13457 4576 13470 4590
rect 13538 4586 13691 4590
rect 13420 4574 13442 4576
rect 13520 4574 13712 4586
rect 13791 4574 13804 4604
rect 13819 4590 13849 4604
rect 13886 4574 13905 4604
rect 13920 4574 13926 4604
rect 13935 4574 13948 4604
rect 13963 4590 13993 4604
rect 14036 4590 14079 4604
rect 14086 4590 14306 4604
rect 14313 4590 14343 4604
rect 14003 4576 14018 4588
rect 14037 4576 14050 4590
rect 14118 4586 14271 4590
rect 14000 4574 14022 4576
rect 14100 4574 14292 4586
rect 14371 4574 14384 4604
rect 14399 4590 14429 4604
rect 14466 4574 14485 4604
rect 14500 4574 14506 4604
rect 14515 4574 14528 4604
rect 14543 4590 14573 4604
rect 14616 4590 14659 4604
rect 14666 4590 14886 4604
rect 14893 4590 14923 4604
rect 14583 4576 14598 4588
rect 14617 4576 14630 4590
rect 14698 4586 14851 4590
rect 14580 4574 14602 4576
rect 14680 4574 14872 4586
rect 14951 4574 14964 4604
rect 14979 4590 15009 4604
rect 15046 4574 15065 4604
rect 15080 4574 15086 4604
rect 15095 4574 15108 4604
rect 15123 4590 15153 4604
rect 15196 4590 15239 4604
rect 15246 4590 15466 4604
rect 15473 4590 15503 4604
rect 15163 4576 15178 4588
rect 15197 4576 15210 4590
rect 15278 4586 15431 4590
rect 15160 4574 15182 4576
rect 15260 4574 15452 4586
rect 15531 4574 15544 4604
rect 15559 4590 15589 4604
rect 15626 4574 15645 4604
rect 15660 4574 15666 4604
rect 15675 4574 15688 4604
rect 15703 4590 15733 4604
rect 15776 4590 15819 4604
rect 15826 4590 16046 4604
rect 16053 4590 16083 4604
rect 15743 4576 15758 4588
rect 15777 4576 15790 4590
rect 15858 4586 16011 4590
rect 15740 4574 15762 4576
rect 15840 4574 16032 4586
rect 16111 4574 16124 4604
rect 16139 4590 16169 4604
rect 16206 4574 16225 4604
rect 16240 4574 16246 4604
rect 16255 4574 16268 4604
rect 16283 4590 16313 4604
rect 16356 4590 16399 4604
rect 16406 4590 16626 4604
rect 16633 4590 16663 4604
rect 16323 4576 16338 4588
rect 16357 4576 16370 4590
rect 16438 4586 16591 4590
rect 16320 4574 16342 4576
rect 16420 4574 16612 4586
rect 16691 4574 16704 4604
rect 16719 4590 16749 4604
rect 16786 4574 16805 4604
rect 16820 4574 16826 4604
rect 16835 4574 16848 4604
rect 16863 4590 16893 4604
rect 16936 4590 16979 4604
rect 16986 4590 17206 4604
rect 17213 4590 17243 4604
rect 16903 4576 16918 4588
rect 16937 4576 16950 4590
rect 17018 4586 17171 4590
rect 16900 4574 16922 4576
rect 17000 4574 17192 4586
rect 17271 4574 17284 4604
rect 17299 4590 17329 4604
rect 17366 4574 17385 4604
rect 17400 4574 17406 4604
rect 17415 4574 17428 4604
rect 17443 4590 17473 4604
rect 17516 4590 17559 4604
rect 17566 4590 17786 4604
rect 17793 4590 17823 4604
rect 17483 4576 17498 4588
rect 17517 4576 17530 4590
rect 17598 4586 17751 4590
rect 17480 4574 17502 4576
rect 17580 4574 17772 4586
rect 17851 4574 17864 4604
rect 17879 4590 17909 4604
rect 17946 4574 17965 4604
rect 17980 4574 17986 4604
rect 17995 4574 18008 4604
rect 18023 4590 18053 4604
rect 18096 4590 18139 4604
rect 18146 4590 18366 4604
rect 18373 4590 18403 4604
rect 18063 4576 18078 4588
rect 18097 4576 18110 4590
rect 18178 4586 18331 4590
rect 18060 4574 18082 4576
rect 18160 4574 18352 4586
rect 18431 4574 18444 4604
rect 18459 4590 18489 4604
rect 18532 4574 18545 4604
rect 0 4560 18545 4574
rect 15 4490 28 4560
rect 80 4556 102 4560
rect 73 4534 102 4548
rect 155 4534 171 4548
rect 209 4544 215 4546
rect 222 4544 330 4560
rect 337 4544 343 4546
rect 351 4544 366 4560
rect 432 4554 451 4557
rect 73 4532 171 4534
rect 198 4532 366 4544
rect 381 4534 397 4548
rect 432 4535 454 4554
rect 464 4548 480 4549
rect 463 4546 480 4548
rect 464 4541 480 4546
rect 454 4534 460 4535
rect 463 4534 492 4541
rect 381 4533 492 4534
rect 381 4532 498 4533
rect 57 4524 108 4532
rect 155 4524 189 4532
rect 57 4512 82 4524
rect 89 4512 108 4524
rect 162 4522 189 4524
rect 198 4522 419 4532
rect 454 4529 460 4532
rect 162 4518 419 4522
rect 57 4504 108 4512
rect 155 4504 419 4518
rect 463 4524 498 4532
rect 9 4456 28 4490
rect 73 4496 102 4504
rect 73 4490 90 4496
rect 73 4488 107 4490
rect 155 4488 171 4504
rect 172 4494 380 4504
rect 381 4494 397 4504
rect 445 4500 460 4515
rect 463 4512 464 4524
rect 471 4512 498 4524
rect 463 4504 498 4512
rect 463 4503 492 4504
rect 183 4490 397 4494
rect 198 4488 397 4490
rect 432 4490 445 4500
rect 463 4490 480 4503
rect 432 4488 480 4490
rect 74 4484 107 4488
rect 70 4482 107 4484
rect 70 4481 137 4482
rect 70 4476 101 4481
rect 107 4476 137 4481
rect 70 4472 137 4476
rect 43 4469 137 4472
rect 43 4462 92 4469
rect 43 4456 73 4462
rect 92 4457 97 4462
rect 9 4440 89 4456
rect 101 4448 137 4469
rect 198 4464 387 4488
rect 432 4487 479 4488
rect 445 4482 479 4487
rect 213 4461 387 4464
rect 206 4458 387 4461
rect 415 4481 479 4482
rect 9 4438 28 4440
rect 43 4438 77 4440
rect 9 4422 89 4438
rect 9 4416 28 4422
rect -1 4400 28 4416
rect 43 4406 73 4422
rect 101 4400 107 4448
rect 110 4442 129 4448
rect 144 4442 174 4450
rect 110 4434 174 4442
rect 110 4418 190 4434
rect 206 4427 268 4458
rect 284 4427 346 4458
rect 415 4456 464 4481
rect 479 4456 509 4472
rect 378 4442 408 4450
rect 415 4448 525 4456
rect 378 4434 423 4442
rect 110 4416 129 4418
rect 144 4416 190 4418
rect 110 4400 190 4416
rect 217 4414 252 4427
rect 293 4424 330 4427
rect 293 4422 335 4424
rect 222 4411 252 4414
rect 231 4407 238 4411
rect 238 4406 239 4407
rect 197 4400 207 4406
rect -7 4392 34 4400
rect -7 4366 8 4392
rect 15 4366 34 4392
rect 98 4388 129 4400
rect 144 4388 247 4400
rect 259 4390 285 4416
rect 300 4411 330 4422
rect 362 4418 424 4434
rect 362 4416 408 4418
rect 362 4400 424 4416
rect 436 4400 442 4448
rect 445 4440 525 4448
rect 445 4438 464 4440
rect 479 4438 513 4440
rect 445 4422 525 4438
rect 445 4400 464 4422
rect 479 4406 509 4422
rect 537 4416 543 4490
rect 546 4416 565 4560
rect 580 4416 586 4560
rect 595 4490 608 4560
rect 660 4556 682 4560
rect 653 4534 682 4548
rect 735 4534 751 4548
rect 789 4544 795 4546
rect 802 4544 910 4560
rect 917 4544 923 4546
rect 931 4544 946 4560
rect 1012 4554 1031 4557
rect 653 4532 751 4534
rect 778 4532 946 4544
rect 961 4534 977 4548
rect 1012 4535 1034 4554
rect 1044 4548 1060 4549
rect 1043 4546 1060 4548
rect 1044 4541 1060 4546
rect 1034 4534 1040 4535
rect 1043 4534 1072 4541
rect 961 4533 1072 4534
rect 961 4532 1078 4533
rect 637 4524 688 4532
rect 735 4524 769 4532
rect 637 4512 662 4524
rect 669 4512 688 4524
rect 742 4522 769 4524
rect 778 4522 999 4532
rect 1034 4529 1040 4532
rect 742 4518 999 4522
rect 637 4504 688 4512
rect 735 4504 999 4518
rect 1043 4524 1078 4532
rect 589 4456 608 4490
rect 653 4496 682 4504
rect 653 4490 670 4496
rect 653 4488 687 4490
rect 735 4488 751 4504
rect 752 4494 960 4504
rect 961 4494 977 4504
rect 1025 4500 1040 4515
rect 1043 4512 1044 4524
rect 1051 4512 1078 4524
rect 1043 4504 1078 4512
rect 1043 4503 1072 4504
rect 763 4490 977 4494
rect 778 4488 977 4490
rect 1012 4490 1025 4500
rect 1043 4490 1060 4503
rect 1012 4488 1060 4490
rect 654 4484 687 4488
rect 650 4482 687 4484
rect 650 4481 717 4482
rect 650 4476 681 4481
rect 687 4476 717 4481
rect 650 4472 717 4476
rect 623 4469 717 4472
rect 623 4462 672 4469
rect 623 4456 653 4462
rect 672 4457 677 4462
rect 589 4440 669 4456
rect 681 4448 717 4469
rect 778 4464 967 4488
rect 1012 4487 1059 4488
rect 1025 4482 1059 4487
rect 793 4461 967 4464
rect 786 4458 967 4461
rect 995 4481 1059 4482
rect 589 4438 608 4440
rect 623 4438 657 4440
rect 589 4422 669 4438
rect 589 4416 608 4422
rect 305 4390 408 4400
rect 259 4388 408 4390
rect 429 4388 464 4400
rect 98 4386 260 4388
rect 110 4366 129 4386
rect 144 4384 174 4386
rect -7 4358 34 4366
rect 116 4362 129 4366
rect 181 4370 260 4386
rect 292 4386 464 4388
rect 292 4370 371 4386
rect 378 4384 408 4386
rect -1 4348 28 4358
rect 43 4348 73 4362
rect 116 4348 159 4362
rect 181 4358 371 4370
rect 436 4366 442 4386
rect 166 4348 196 4358
rect 197 4348 355 4358
rect 359 4348 389 4358
rect 393 4348 423 4362
rect 451 4348 464 4386
rect 536 4400 565 4416
rect 579 4400 608 4416
rect 623 4406 653 4422
rect 681 4400 687 4448
rect 690 4442 709 4448
rect 724 4442 754 4450
rect 690 4434 754 4442
rect 690 4418 770 4434
rect 786 4427 848 4458
rect 864 4427 926 4458
rect 995 4456 1044 4481
rect 1059 4456 1089 4472
rect 958 4442 988 4450
rect 995 4448 1105 4456
rect 958 4434 1003 4442
rect 690 4416 709 4418
rect 724 4416 770 4418
rect 690 4400 770 4416
rect 797 4414 832 4427
rect 873 4424 910 4427
rect 873 4422 915 4424
rect 802 4411 832 4414
rect 811 4407 818 4411
rect 818 4406 819 4407
rect 777 4400 787 4406
rect 536 4392 571 4400
rect 536 4366 537 4392
rect 544 4366 571 4392
rect 479 4348 509 4362
rect 536 4358 571 4366
rect 573 4392 614 4400
rect 573 4366 588 4392
rect 595 4366 614 4392
rect 678 4388 709 4400
rect 724 4388 827 4400
rect 839 4390 865 4416
rect 880 4411 910 4422
rect 942 4418 1004 4434
rect 942 4416 988 4418
rect 942 4400 1004 4416
rect 1016 4400 1022 4448
rect 1025 4440 1105 4448
rect 1025 4438 1044 4440
rect 1059 4438 1093 4440
rect 1025 4422 1105 4438
rect 1025 4400 1044 4422
rect 1059 4406 1089 4422
rect 1117 4416 1123 4490
rect 1126 4416 1145 4560
rect 1160 4416 1166 4560
rect 1175 4490 1188 4560
rect 1240 4556 1262 4560
rect 1233 4534 1262 4548
rect 1315 4534 1331 4548
rect 1369 4544 1375 4546
rect 1382 4544 1490 4560
rect 1497 4544 1503 4546
rect 1511 4544 1526 4560
rect 1592 4554 1611 4557
rect 1233 4532 1331 4534
rect 1358 4532 1526 4544
rect 1541 4534 1557 4548
rect 1592 4535 1614 4554
rect 1624 4548 1640 4549
rect 1623 4546 1640 4548
rect 1624 4541 1640 4546
rect 1614 4534 1620 4535
rect 1623 4534 1652 4541
rect 1541 4533 1652 4534
rect 1541 4532 1658 4533
rect 1217 4524 1268 4532
rect 1315 4524 1349 4532
rect 1217 4512 1242 4524
rect 1249 4512 1268 4524
rect 1322 4522 1349 4524
rect 1358 4522 1579 4532
rect 1614 4529 1620 4532
rect 1322 4518 1579 4522
rect 1217 4504 1268 4512
rect 1315 4504 1579 4518
rect 1623 4524 1658 4532
rect 1169 4456 1188 4490
rect 1233 4496 1262 4504
rect 1233 4490 1250 4496
rect 1233 4488 1267 4490
rect 1315 4488 1331 4504
rect 1332 4494 1540 4504
rect 1541 4494 1557 4504
rect 1605 4500 1620 4515
rect 1623 4512 1624 4524
rect 1631 4512 1658 4524
rect 1623 4504 1658 4512
rect 1623 4503 1652 4504
rect 1343 4490 1557 4494
rect 1358 4488 1557 4490
rect 1592 4490 1605 4500
rect 1623 4490 1640 4503
rect 1592 4488 1640 4490
rect 1234 4484 1267 4488
rect 1230 4482 1267 4484
rect 1230 4481 1297 4482
rect 1230 4476 1261 4481
rect 1267 4476 1297 4481
rect 1230 4472 1297 4476
rect 1203 4469 1297 4472
rect 1203 4462 1252 4469
rect 1203 4456 1233 4462
rect 1252 4457 1257 4462
rect 1169 4440 1249 4456
rect 1261 4448 1297 4469
rect 1358 4464 1547 4488
rect 1592 4487 1639 4488
rect 1605 4482 1639 4487
rect 1373 4461 1547 4464
rect 1366 4458 1547 4461
rect 1575 4481 1639 4482
rect 1169 4438 1188 4440
rect 1203 4438 1237 4440
rect 1169 4422 1249 4438
rect 1169 4416 1188 4422
rect 885 4390 988 4400
rect 839 4388 988 4390
rect 1009 4388 1044 4400
rect 678 4386 840 4388
rect 690 4366 709 4386
rect 724 4384 754 4386
rect 573 4358 614 4366
rect 696 4362 709 4366
rect 761 4370 840 4386
rect 872 4386 1044 4388
rect 872 4370 951 4386
rect 958 4384 988 4386
rect 536 4348 565 4358
rect 579 4348 608 4358
rect 623 4348 653 4362
rect 696 4348 739 4362
rect 761 4358 951 4370
rect 1016 4366 1022 4386
rect 746 4348 776 4358
rect 777 4348 935 4358
rect 939 4348 969 4358
rect 973 4348 1003 4362
rect 1031 4348 1044 4386
rect 1116 4400 1145 4416
rect 1159 4400 1188 4416
rect 1203 4406 1233 4422
rect 1261 4400 1267 4448
rect 1270 4442 1289 4448
rect 1304 4442 1334 4450
rect 1270 4434 1334 4442
rect 1270 4418 1350 4434
rect 1366 4427 1428 4458
rect 1444 4427 1506 4458
rect 1575 4456 1624 4481
rect 1639 4456 1669 4472
rect 1538 4442 1568 4450
rect 1575 4448 1685 4456
rect 1538 4434 1583 4442
rect 1270 4416 1289 4418
rect 1304 4416 1350 4418
rect 1270 4400 1350 4416
rect 1377 4414 1412 4427
rect 1453 4424 1490 4427
rect 1453 4422 1495 4424
rect 1382 4411 1412 4414
rect 1391 4407 1398 4411
rect 1398 4406 1399 4407
rect 1357 4400 1367 4406
rect 1116 4392 1151 4400
rect 1116 4366 1117 4392
rect 1124 4366 1151 4392
rect 1059 4348 1089 4362
rect 1116 4358 1151 4366
rect 1153 4392 1194 4400
rect 1153 4366 1168 4392
rect 1175 4366 1194 4392
rect 1258 4388 1289 4400
rect 1304 4388 1407 4400
rect 1419 4390 1445 4416
rect 1460 4411 1490 4422
rect 1522 4418 1584 4434
rect 1522 4416 1568 4418
rect 1522 4400 1584 4416
rect 1596 4400 1602 4448
rect 1605 4440 1685 4448
rect 1605 4438 1624 4440
rect 1639 4438 1673 4440
rect 1605 4422 1685 4438
rect 1605 4400 1624 4422
rect 1639 4406 1669 4422
rect 1697 4416 1703 4490
rect 1706 4416 1725 4560
rect 1740 4416 1746 4560
rect 1755 4490 1768 4560
rect 1820 4556 1842 4560
rect 1813 4534 1842 4548
rect 1895 4534 1911 4548
rect 1949 4544 1955 4546
rect 1962 4544 2070 4560
rect 2077 4544 2083 4546
rect 2091 4544 2106 4560
rect 2172 4554 2191 4557
rect 1813 4532 1911 4534
rect 1938 4532 2106 4544
rect 2121 4534 2137 4548
rect 2172 4535 2194 4554
rect 2204 4548 2220 4549
rect 2203 4546 2220 4548
rect 2204 4541 2220 4546
rect 2194 4534 2200 4535
rect 2203 4534 2232 4541
rect 2121 4533 2232 4534
rect 2121 4532 2238 4533
rect 1797 4524 1848 4532
rect 1895 4524 1929 4532
rect 1797 4512 1822 4524
rect 1829 4512 1848 4524
rect 1902 4522 1929 4524
rect 1938 4522 2159 4532
rect 2194 4529 2200 4532
rect 1902 4518 2159 4522
rect 1797 4504 1848 4512
rect 1895 4504 2159 4518
rect 2203 4524 2238 4532
rect 1749 4456 1768 4490
rect 1813 4496 1842 4504
rect 1813 4490 1830 4496
rect 1813 4488 1847 4490
rect 1895 4488 1911 4504
rect 1912 4494 2120 4504
rect 2121 4494 2137 4504
rect 2185 4500 2200 4515
rect 2203 4512 2204 4524
rect 2211 4512 2238 4524
rect 2203 4504 2238 4512
rect 2203 4503 2232 4504
rect 1923 4490 2137 4494
rect 1938 4488 2137 4490
rect 2172 4490 2185 4500
rect 2203 4490 2220 4503
rect 2172 4488 2220 4490
rect 1814 4484 1847 4488
rect 1810 4482 1847 4484
rect 1810 4481 1877 4482
rect 1810 4476 1841 4481
rect 1847 4476 1877 4481
rect 1810 4472 1877 4476
rect 1783 4469 1877 4472
rect 1783 4462 1832 4469
rect 1783 4456 1813 4462
rect 1832 4457 1837 4462
rect 1749 4440 1829 4456
rect 1841 4448 1877 4469
rect 1938 4464 2127 4488
rect 2172 4487 2219 4488
rect 2185 4482 2219 4487
rect 1953 4461 2127 4464
rect 1946 4458 2127 4461
rect 2155 4481 2219 4482
rect 1749 4438 1768 4440
rect 1783 4438 1817 4440
rect 1749 4422 1829 4438
rect 1749 4416 1768 4422
rect 1465 4390 1568 4400
rect 1419 4388 1568 4390
rect 1589 4388 1624 4400
rect 1258 4386 1420 4388
rect 1270 4366 1289 4386
rect 1304 4384 1334 4386
rect 1153 4358 1194 4366
rect 1276 4362 1289 4366
rect 1341 4370 1420 4386
rect 1452 4386 1624 4388
rect 1452 4370 1531 4386
rect 1538 4384 1568 4386
rect 1116 4348 1145 4358
rect 1159 4348 1188 4358
rect 1203 4348 1233 4362
rect 1276 4348 1319 4362
rect 1341 4358 1531 4370
rect 1596 4366 1602 4386
rect 1326 4348 1356 4358
rect 1357 4348 1515 4358
rect 1519 4348 1549 4358
rect 1553 4348 1583 4362
rect 1611 4348 1624 4386
rect 1696 4400 1725 4416
rect 1739 4400 1768 4416
rect 1783 4406 1813 4422
rect 1841 4400 1847 4448
rect 1850 4442 1869 4448
rect 1884 4442 1914 4450
rect 1850 4434 1914 4442
rect 1850 4418 1930 4434
rect 1946 4427 2008 4458
rect 2024 4427 2086 4458
rect 2155 4456 2204 4481
rect 2219 4456 2249 4472
rect 2118 4442 2148 4450
rect 2155 4448 2265 4456
rect 2118 4434 2163 4442
rect 1850 4416 1869 4418
rect 1884 4416 1930 4418
rect 1850 4400 1930 4416
rect 1957 4414 1992 4427
rect 2033 4424 2070 4427
rect 2033 4422 2075 4424
rect 1962 4411 1992 4414
rect 1971 4407 1978 4411
rect 1978 4406 1979 4407
rect 1937 4400 1947 4406
rect 1696 4392 1731 4400
rect 1696 4366 1697 4392
rect 1704 4366 1731 4392
rect 1639 4348 1669 4362
rect 1696 4358 1731 4366
rect 1733 4392 1774 4400
rect 1733 4366 1748 4392
rect 1755 4366 1774 4392
rect 1838 4388 1869 4400
rect 1884 4388 1987 4400
rect 1999 4390 2025 4416
rect 2040 4411 2070 4422
rect 2102 4418 2164 4434
rect 2102 4416 2148 4418
rect 2102 4400 2164 4416
rect 2176 4400 2182 4448
rect 2185 4440 2265 4448
rect 2185 4438 2204 4440
rect 2219 4438 2253 4440
rect 2185 4422 2265 4438
rect 2185 4400 2204 4422
rect 2219 4406 2249 4422
rect 2277 4416 2283 4490
rect 2286 4416 2305 4560
rect 2320 4416 2326 4560
rect 2335 4490 2348 4560
rect 2400 4556 2422 4560
rect 2393 4534 2422 4548
rect 2475 4534 2491 4548
rect 2529 4544 2535 4546
rect 2542 4544 2650 4560
rect 2657 4544 2663 4546
rect 2671 4544 2686 4560
rect 2752 4554 2771 4557
rect 2393 4532 2491 4534
rect 2518 4532 2686 4544
rect 2701 4534 2717 4548
rect 2752 4535 2774 4554
rect 2784 4548 2800 4549
rect 2783 4546 2800 4548
rect 2784 4541 2800 4546
rect 2774 4534 2780 4535
rect 2783 4534 2812 4541
rect 2701 4533 2812 4534
rect 2701 4532 2818 4533
rect 2377 4524 2428 4532
rect 2475 4524 2509 4532
rect 2377 4512 2402 4524
rect 2409 4512 2428 4524
rect 2482 4522 2509 4524
rect 2518 4522 2739 4532
rect 2774 4529 2780 4532
rect 2482 4518 2739 4522
rect 2377 4504 2428 4512
rect 2475 4504 2739 4518
rect 2783 4524 2818 4532
rect 2329 4456 2348 4490
rect 2393 4496 2422 4504
rect 2393 4490 2410 4496
rect 2393 4488 2427 4490
rect 2475 4488 2491 4504
rect 2492 4494 2700 4504
rect 2701 4494 2717 4504
rect 2765 4500 2780 4515
rect 2783 4512 2784 4524
rect 2791 4512 2818 4524
rect 2783 4504 2818 4512
rect 2783 4503 2812 4504
rect 2503 4490 2717 4494
rect 2518 4488 2717 4490
rect 2752 4490 2765 4500
rect 2783 4490 2800 4503
rect 2752 4488 2800 4490
rect 2394 4484 2427 4488
rect 2390 4482 2427 4484
rect 2390 4481 2457 4482
rect 2390 4476 2421 4481
rect 2427 4476 2457 4481
rect 2390 4472 2457 4476
rect 2363 4469 2457 4472
rect 2363 4462 2412 4469
rect 2363 4456 2393 4462
rect 2412 4457 2417 4462
rect 2329 4440 2409 4456
rect 2421 4448 2457 4469
rect 2518 4464 2707 4488
rect 2752 4487 2799 4488
rect 2765 4482 2799 4487
rect 2533 4461 2707 4464
rect 2526 4458 2707 4461
rect 2735 4481 2799 4482
rect 2329 4438 2348 4440
rect 2363 4438 2397 4440
rect 2329 4422 2409 4438
rect 2329 4416 2348 4422
rect 2045 4390 2148 4400
rect 1999 4388 2148 4390
rect 2169 4388 2204 4400
rect 1838 4386 2000 4388
rect 1850 4366 1869 4386
rect 1884 4384 1914 4386
rect 1733 4358 1774 4366
rect 1856 4362 1869 4366
rect 1921 4370 2000 4386
rect 2032 4386 2204 4388
rect 2032 4370 2111 4386
rect 2118 4384 2148 4386
rect 1696 4348 1725 4358
rect 1739 4348 1768 4358
rect 1783 4348 1813 4362
rect 1856 4348 1899 4362
rect 1921 4358 2111 4370
rect 2176 4366 2182 4386
rect 1906 4348 1936 4358
rect 1937 4348 2095 4358
rect 2099 4348 2129 4358
rect 2133 4348 2163 4362
rect 2191 4348 2204 4386
rect 2276 4400 2305 4416
rect 2319 4400 2348 4416
rect 2363 4406 2393 4422
rect 2421 4400 2427 4448
rect 2430 4442 2449 4448
rect 2464 4442 2494 4450
rect 2430 4434 2494 4442
rect 2430 4418 2510 4434
rect 2526 4427 2588 4458
rect 2604 4427 2666 4458
rect 2735 4456 2784 4481
rect 2799 4456 2829 4472
rect 2698 4442 2728 4450
rect 2735 4448 2845 4456
rect 2698 4434 2743 4442
rect 2430 4416 2449 4418
rect 2464 4416 2510 4418
rect 2430 4400 2510 4416
rect 2537 4414 2572 4427
rect 2613 4424 2650 4427
rect 2613 4422 2655 4424
rect 2542 4411 2572 4414
rect 2551 4407 2558 4411
rect 2558 4406 2559 4407
rect 2517 4400 2527 4406
rect 2276 4392 2311 4400
rect 2276 4366 2277 4392
rect 2284 4366 2311 4392
rect 2219 4348 2249 4362
rect 2276 4358 2311 4366
rect 2313 4392 2354 4400
rect 2313 4366 2328 4392
rect 2335 4366 2354 4392
rect 2418 4388 2449 4400
rect 2464 4388 2567 4400
rect 2579 4390 2605 4416
rect 2620 4411 2650 4422
rect 2682 4418 2744 4434
rect 2682 4416 2728 4418
rect 2682 4400 2744 4416
rect 2756 4400 2762 4448
rect 2765 4440 2845 4448
rect 2765 4438 2784 4440
rect 2799 4438 2833 4440
rect 2765 4422 2845 4438
rect 2765 4400 2784 4422
rect 2799 4406 2829 4422
rect 2857 4416 2863 4490
rect 2866 4416 2885 4560
rect 2900 4416 2906 4560
rect 2915 4490 2928 4560
rect 2980 4556 3002 4560
rect 2973 4534 3002 4548
rect 3055 4534 3071 4548
rect 3109 4544 3115 4546
rect 3122 4544 3230 4560
rect 3237 4544 3243 4546
rect 3251 4544 3266 4560
rect 3332 4554 3351 4557
rect 2973 4532 3071 4534
rect 3098 4532 3266 4544
rect 3281 4534 3297 4548
rect 3332 4535 3354 4554
rect 3364 4548 3380 4549
rect 3363 4546 3380 4548
rect 3364 4541 3380 4546
rect 3354 4534 3360 4535
rect 3363 4534 3392 4541
rect 3281 4533 3392 4534
rect 3281 4532 3398 4533
rect 2957 4524 3008 4532
rect 3055 4524 3089 4532
rect 2957 4512 2982 4524
rect 2989 4512 3008 4524
rect 3062 4522 3089 4524
rect 3098 4522 3319 4532
rect 3354 4529 3360 4532
rect 3062 4518 3319 4522
rect 2957 4504 3008 4512
rect 3055 4504 3319 4518
rect 3363 4524 3398 4532
rect 2909 4456 2928 4490
rect 2973 4496 3002 4504
rect 2973 4490 2990 4496
rect 2973 4488 3007 4490
rect 3055 4488 3071 4504
rect 3072 4494 3280 4504
rect 3281 4494 3297 4504
rect 3345 4500 3360 4515
rect 3363 4512 3364 4524
rect 3371 4512 3398 4524
rect 3363 4504 3398 4512
rect 3363 4503 3392 4504
rect 3083 4490 3297 4494
rect 3098 4488 3297 4490
rect 3332 4490 3345 4500
rect 3363 4490 3380 4503
rect 3332 4488 3380 4490
rect 2974 4484 3007 4488
rect 2970 4482 3007 4484
rect 2970 4481 3037 4482
rect 2970 4476 3001 4481
rect 3007 4476 3037 4481
rect 2970 4472 3037 4476
rect 2943 4469 3037 4472
rect 2943 4462 2992 4469
rect 2943 4456 2973 4462
rect 2992 4457 2997 4462
rect 2909 4440 2989 4456
rect 3001 4448 3037 4469
rect 3098 4464 3287 4488
rect 3332 4487 3379 4488
rect 3345 4482 3379 4487
rect 3113 4461 3287 4464
rect 3106 4458 3287 4461
rect 3315 4481 3379 4482
rect 2909 4438 2928 4440
rect 2943 4438 2977 4440
rect 2909 4422 2989 4438
rect 2909 4416 2928 4422
rect 2625 4390 2728 4400
rect 2579 4388 2728 4390
rect 2749 4388 2784 4400
rect 2418 4386 2580 4388
rect 2430 4366 2449 4386
rect 2464 4384 2494 4386
rect 2313 4358 2354 4366
rect 2436 4362 2449 4366
rect 2501 4370 2580 4386
rect 2612 4386 2784 4388
rect 2612 4370 2691 4386
rect 2698 4384 2728 4386
rect 2276 4348 2305 4358
rect 2319 4348 2348 4358
rect 2363 4348 2393 4362
rect 2436 4348 2479 4362
rect 2501 4358 2691 4370
rect 2756 4366 2762 4386
rect 2486 4348 2516 4358
rect 2517 4348 2675 4358
rect 2679 4348 2709 4358
rect 2713 4348 2743 4362
rect 2771 4348 2784 4386
rect 2856 4400 2885 4416
rect 2899 4400 2928 4416
rect 2943 4406 2973 4422
rect 3001 4400 3007 4448
rect 3010 4442 3029 4448
rect 3044 4442 3074 4450
rect 3010 4434 3074 4442
rect 3010 4418 3090 4434
rect 3106 4427 3168 4458
rect 3184 4427 3246 4458
rect 3315 4456 3364 4481
rect 3379 4456 3409 4472
rect 3278 4442 3308 4450
rect 3315 4448 3425 4456
rect 3278 4434 3323 4442
rect 3010 4416 3029 4418
rect 3044 4416 3090 4418
rect 3010 4400 3090 4416
rect 3117 4414 3152 4427
rect 3193 4424 3230 4427
rect 3193 4422 3235 4424
rect 3122 4411 3152 4414
rect 3131 4407 3138 4411
rect 3138 4406 3139 4407
rect 3097 4400 3107 4406
rect 2856 4392 2891 4400
rect 2856 4366 2857 4392
rect 2864 4366 2891 4392
rect 2799 4348 2829 4362
rect 2856 4358 2891 4366
rect 2893 4392 2934 4400
rect 2893 4366 2908 4392
rect 2915 4366 2934 4392
rect 2998 4388 3029 4400
rect 3044 4388 3147 4400
rect 3159 4390 3185 4416
rect 3200 4411 3230 4422
rect 3262 4418 3324 4434
rect 3262 4416 3308 4418
rect 3262 4400 3324 4416
rect 3336 4400 3342 4448
rect 3345 4440 3425 4448
rect 3345 4438 3364 4440
rect 3379 4438 3413 4440
rect 3345 4422 3425 4438
rect 3345 4400 3364 4422
rect 3379 4406 3409 4422
rect 3437 4416 3443 4490
rect 3446 4416 3465 4560
rect 3480 4416 3486 4560
rect 3495 4490 3508 4560
rect 3560 4556 3582 4560
rect 3553 4534 3582 4548
rect 3635 4534 3651 4548
rect 3689 4544 3695 4546
rect 3702 4544 3810 4560
rect 3817 4544 3823 4546
rect 3831 4544 3846 4560
rect 3912 4554 3931 4557
rect 3553 4532 3651 4534
rect 3678 4532 3846 4544
rect 3861 4534 3877 4548
rect 3912 4535 3934 4554
rect 3944 4548 3960 4549
rect 3943 4546 3960 4548
rect 3944 4541 3960 4546
rect 3934 4534 3940 4535
rect 3943 4534 3972 4541
rect 3861 4533 3972 4534
rect 3861 4532 3978 4533
rect 3537 4524 3588 4532
rect 3635 4524 3669 4532
rect 3537 4512 3562 4524
rect 3569 4512 3588 4524
rect 3642 4522 3669 4524
rect 3678 4522 3899 4532
rect 3934 4529 3940 4532
rect 3642 4518 3899 4522
rect 3537 4504 3588 4512
rect 3635 4504 3899 4518
rect 3943 4524 3978 4532
rect 3489 4456 3508 4490
rect 3553 4496 3582 4504
rect 3553 4490 3570 4496
rect 3553 4488 3587 4490
rect 3635 4488 3651 4504
rect 3652 4494 3860 4504
rect 3861 4494 3877 4504
rect 3925 4500 3940 4515
rect 3943 4512 3944 4524
rect 3951 4512 3978 4524
rect 3943 4504 3978 4512
rect 3943 4503 3972 4504
rect 3663 4490 3877 4494
rect 3678 4488 3877 4490
rect 3912 4490 3925 4500
rect 3943 4490 3960 4503
rect 3912 4488 3960 4490
rect 3554 4484 3587 4488
rect 3550 4482 3587 4484
rect 3550 4481 3617 4482
rect 3550 4476 3581 4481
rect 3587 4476 3617 4481
rect 3550 4472 3617 4476
rect 3523 4469 3617 4472
rect 3523 4462 3572 4469
rect 3523 4456 3553 4462
rect 3572 4457 3577 4462
rect 3489 4440 3569 4456
rect 3581 4448 3617 4469
rect 3678 4464 3867 4488
rect 3912 4487 3959 4488
rect 3925 4482 3959 4487
rect 3693 4461 3867 4464
rect 3686 4458 3867 4461
rect 3895 4481 3959 4482
rect 3489 4438 3508 4440
rect 3523 4438 3557 4440
rect 3489 4422 3569 4438
rect 3489 4416 3508 4422
rect 3205 4390 3308 4400
rect 3159 4388 3308 4390
rect 3329 4388 3364 4400
rect 2998 4386 3160 4388
rect 3010 4366 3029 4386
rect 3044 4384 3074 4386
rect 2893 4358 2934 4366
rect 3016 4362 3029 4366
rect 3081 4370 3160 4386
rect 3192 4386 3364 4388
rect 3192 4370 3271 4386
rect 3278 4384 3308 4386
rect 2856 4348 2885 4358
rect 2899 4348 2928 4358
rect 2943 4348 2973 4362
rect 3016 4348 3059 4362
rect 3081 4358 3271 4370
rect 3336 4366 3342 4386
rect 3066 4348 3096 4358
rect 3097 4348 3255 4358
rect 3259 4348 3289 4358
rect 3293 4348 3323 4362
rect 3351 4348 3364 4386
rect 3436 4400 3465 4416
rect 3479 4400 3508 4416
rect 3523 4406 3553 4422
rect 3581 4400 3587 4448
rect 3590 4442 3609 4448
rect 3624 4442 3654 4450
rect 3590 4434 3654 4442
rect 3590 4418 3670 4434
rect 3686 4427 3748 4458
rect 3764 4427 3826 4458
rect 3895 4456 3944 4481
rect 3959 4456 3989 4472
rect 3858 4442 3888 4450
rect 3895 4448 4005 4456
rect 3858 4434 3903 4442
rect 3590 4416 3609 4418
rect 3624 4416 3670 4418
rect 3590 4400 3670 4416
rect 3697 4414 3732 4427
rect 3773 4424 3810 4427
rect 3773 4422 3815 4424
rect 3702 4411 3732 4414
rect 3711 4407 3718 4411
rect 3718 4406 3719 4407
rect 3677 4400 3687 4406
rect 3436 4392 3471 4400
rect 3436 4366 3437 4392
rect 3444 4366 3471 4392
rect 3379 4348 3409 4362
rect 3436 4358 3471 4366
rect 3473 4392 3514 4400
rect 3473 4366 3488 4392
rect 3495 4366 3514 4392
rect 3578 4388 3609 4400
rect 3624 4388 3727 4400
rect 3739 4390 3765 4416
rect 3780 4411 3810 4422
rect 3842 4418 3904 4434
rect 3842 4416 3888 4418
rect 3842 4400 3904 4416
rect 3916 4400 3922 4448
rect 3925 4440 4005 4448
rect 3925 4438 3944 4440
rect 3959 4438 3993 4440
rect 3925 4422 4005 4438
rect 3925 4400 3944 4422
rect 3959 4406 3989 4422
rect 4017 4416 4023 4490
rect 4026 4416 4045 4560
rect 4060 4416 4066 4560
rect 4075 4490 4088 4560
rect 4140 4556 4162 4560
rect 4133 4534 4162 4548
rect 4215 4534 4231 4548
rect 4269 4544 4275 4546
rect 4282 4544 4390 4560
rect 4397 4544 4403 4546
rect 4411 4544 4426 4560
rect 4492 4554 4511 4557
rect 4133 4532 4231 4534
rect 4258 4532 4426 4544
rect 4441 4534 4457 4548
rect 4492 4535 4514 4554
rect 4524 4548 4540 4549
rect 4523 4546 4540 4548
rect 4524 4541 4540 4546
rect 4514 4534 4520 4535
rect 4523 4534 4552 4541
rect 4441 4533 4552 4534
rect 4441 4532 4558 4533
rect 4117 4524 4168 4532
rect 4215 4524 4249 4532
rect 4117 4512 4142 4524
rect 4149 4512 4168 4524
rect 4222 4522 4249 4524
rect 4258 4522 4479 4532
rect 4514 4529 4520 4532
rect 4222 4518 4479 4522
rect 4117 4504 4168 4512
rect 4215 4504 4479 4518
rect 4523 4524 4558 4532
rect 4069 4456 4088 4490
rect 4133 4496 4162 4504
rect 4133 4490 4150 4496
rect 4133 4488 4167 4490
rect 4215 4488 4231 4504
rect 4232 4494 4440 4504
rect 4441 4494 4457 4504
rect 4505 4500 4520 4515
rect 4523 4512 4524 4524
rect 4531 4512 4558 4524
rect 4523 4504 4558 4512
rect 4523 4503 4552 4504
rect 4243 4490 4457 4494
rect 4258 4488 4457 4490
rect 4492 4490 4505 4500
rect 4523 4490 4540 4503
rect 4492 4488 4540 4490
rect 4134 4484 4167 4488
rect 4130 4482 4167 4484
rect 4130 4481 4197 4482
rect 4130 4476 4161 4481
rect 4167 4476 4197 4481
rect 4130 4472 4197 4476
rect 4103 4469 4197 4472
rect 4103 4462 4152 4469
rect 4103 4456 4133 4462
rect 4152 4457 4157 4462
rect 4069 4440 4149 4456
rect 4161 4448 4197 4469
rect 4258 4464 4447 4488
rect 4492 4487 4539 4488
rect 4505 4482 4539 4487
rect 4273 4461 4447 4464
rect 4266 4458 4447 4461
rect 4475 4481 4539 4482
rect 4069 4438 4088 4440
rect 4103 4438 4137 4440
rect 4069 4422 4149 4438
rect 4069 4416 4088 4422
rect 3785 4390 3888 4400
rect 3739 4388 3888 4390
rect 3909 4388 3944 4400
rect 3578 4386 3740 4388
rect 3590 4366 3609 4386
rect 3624 4384 3654 4386
rect 3473 4358 3514 4366
rect 3596 4362 3609 4366
rect 3661 4370 3740 4386
rect 3772 4386 3944 4388
rect 3772 4370 3851 4386
rect 3858 4384 3888 4386
rect 3436 4348 3465 4358
rect 3479 4348 3508 4358
rect 3523 4348 3553 4362
rect 3596 4348 3639 4362
rect 3661 4358 3851 4370
rect 3916 4366 3922 4386
rect 3646 4348 3676 4358
rect 3677 4348 3835 4358
rect 3839 4348 3869 4358
rect 3873 4348 3903 4362
rect 3931 4348 3944 4386
rect 4016 4400 4045 4416
rect 4059 4400 4088 4416
rect 4103 4406 4133 4422
rect 4161 4400 4167 4448
rect 4170 4442 4189 4448
rect 4204 4442 4234 4450
rect 4170 4434 4234 4442
rect 4170 4418 4250 4434
rect 4266 4427 4328 4458
rect 4344 4427 4406 4458
rect 4475 4456 4524 4481
rect 4539 4456 4569 4472
rect 4438 4442 4468 4450
rect 4475 4448 4585 4456
rect 4438 4434 4483 4442
rect 4170 4416 4189 4418
rect 4204 4416 4250 4418
rect 4170 4400 4250 4416
rect 4277 4414 4312 4427
rect 4353 4424 4390 4427
rect 4353 4422 4395 4424
rect 4282 4411 4312 4414
rect 4291 4407 4298 4411
rect 4298 4406 4299 4407
rect 4257 4400 4267 4406
rect 4016 4392 4051 4400
rect 4016 4366 4017 4392
rect 4024 4366 4051 4392
rect 3959 4348 3989 4362
rect 4016 4358 4051 4366
rect 4053 4392 4094 4400
rect 4053 4366 4068 4392
rect 4075 4366 4094 4392
rect 4158 4388 4189 4400
rect 4204 4388 4307 4400
rect 4319 4390 4345 4416
rect 4360 4411 4390 4422
rect 4422 4418 4484 4434
rect 4422 4416 4468 4418
rect 4422 4400 4484 4416
rect 4496 4400 4502 4448
rect 4505 4440 4585 4448
rect 4505 4438 4524 4440
rect 4539 4438 4573 4440
rect 4505 4422 4585 4438
rect 4505 4400 4524 4422
rect 4539 4406 4569 4422
rect 4597 4416 4603 4490
rect 4606 4416 4625 4560
rect 4640 4416 4646 4560
rect 4655 4490 4668 4560
rect 4720 4556 4742 4560
rect 4713 4534 4742 4548
rect 4795 4534 4811 4548
rect 4849 4544 4855 4546
rect 4862 4544 4970 4560
rect 4977 4544 4983 4546
rect 4991 4544 5006 4560
rect 5072 4554 5091 4557
rect 4713 4532 4811 4534
rect 4838 4532 5006 4544
rect 5021 4534 5037 4548
rect 5072 4535 5094 4554
rect 5104 4548 5120 4549
rect 5103 4546 5120 4548
rect 5104 4541 5120 4546
rect 5094 4534 5100 4535
rect 5103 4534 5132 4541
rect 5021 4533 5132 4534
rect 5021 4532 5138 4533
rect 4697 4524 4748 4532
rect 4795 4524 4829 4532
rect 4697 4512 4722 4524
rect 4729 4512 4748 4524
rect 4802 4522 4829 4524
rect 4838 4522 5059 4532
rect 5094 4529 5100 4532
rect 4802 4518 5059 4522
rect 4697 4504 4748 4512
rect 4795 4504 5059 4518
rect 5103 4524 5138 4532
rect 4649 4456 4668 4490
rect 4713 4496 4742 4504
rect 4713 4490 4730 4496
rect 4713 4488 4747 4490
rect 4795 4488 4811 4504
rect 4812 4494 5020 4504
rect 5021 4494 5037 4504
rect 5085 4500 5100 4515
rect 5103 4512 5104 4524
rect 5111 4512 5138 4524
rect 5103 4504 5138 4512
rect 5103 4503 5132 4504
rect 4823 4490 5037 4494
rect 4838 4488 5037 4490
rect 5072 4490 5085 4500
rect 5103 4490 5120 4503
rect 5072 4488 5120 4490
rect 4714 4484 4747 4488
rect 4710 4482 4747 4484
rect 4710 4481 4777 4482
rect 4710 4476 4741 4481
rect 4747 4476 4777 4481
rect 4710 4472 4777 4476
rect 4683 4469 4777 4472
rect 4683 4462 4732 4469
rect 4683 4456 4713 4462
rect 4732 4457 4737 4462
rect 4649 4440 4729 4456
rect 4741 4448 4777 4469
rect 4838 4464 5027 4488
rect 5072 4487 5119 4488
rect 5085 4482 5119 4487
rect 4853 4461 5027 4464
rect 4846 4458 5027 4461
rect 5055 4481 5119 4482
rect 4649 4438 4668 4440
rect 4683 4438 4717 4440
rect 4649 4422 4729 4438
rect 4649 4416 4668 4422
rect 4365 4390 4468 4400
rect 4319 4388 4468 4390
rect 4489 4388 4524 4400
rect 4158 4386 4320 4388
rect 4170 4366 4189 4386
rect 4204 4384 4234 4386
rect 4053 4358 4094 4366
rect 4176 4362 4189 4366
rect 4241 4370 4320 4386
rect 4352 4386 4524 4388
rect 4352 4370 4431 4386
rect 4438 4384 4468 4386
rect 4016 4348 4045 4358
rect 4059 4348 4088 4358
rect 4103 4348 4133 4362
rect 4176 4348 4219 4362
rect 4241 4358 4431 4370
rect 4496 4366 4502 4386
rect 4226 4348 4256 4358
rect 4257 4348 4415 4358
rect 4419 4348 4449 4358
rect 4453 4348 4483 4362
rect 4511 4348 4524 4386
rect 4596 4400 4625 4416
rect 4639 4400 4668 4416
rect 4683 4406 4713 4422
rect 4741 4400 4747 4448
rect 4750 4442 4769 4448
rect 4784 4442 4814 4450
rect 4750 4434 4814 4442
rect 4750 4418 4830 4434
rect 4846 4427 4908 4458
rect 4924 4427 4986 4458
rect 5055 4456 5104 4481
rect 5119 4456 5149 4472
rect 5018 4442 5048 4450
rect 5055 4448 5165 4456
rect 5018 4434 5063 4442
rect 4750 4416 4769 4418
rect 4784 4416 4830 4418
rect 4750 4400 4830 4416
rect 4857 4414 4892 4427
rect 4933 4424 4970 4427
rect 4933 4422 4975 4424
rect 4862 4411 4892 4414
rect 4871 4407 4878 4411
rect 4878 4406 4879 4407
rect 4837 4400 4847 4406
rect 4596 4392 4631 4400
rect 4596 4366 4597 4392
rect 4604 4366 4631 4392
rect 4539 4348 4569 4362
rect 4596 4358 4631 4366
rect 4633 4392 4674 4400
rect 4633 4366 4648 4392
rect 4655 4366 4674 4392
rect 4738 4388 4769 4400
rect 4784 4388 4887 4400
rect 4899 4390 4925 4416
rect 4940 4411 4970 4422
rect 5002 4418 5064 4434
rect 5002 4416 5048 4418
rect 5002 4400 5064 4416
rect 5076 4400 5082 4448
rect 5085 4440 5165 4448
rect 5085 4438 5104 4440
rect 5119 4438 5153 4440
rect 5085 4422 5165 4438
rect 5085 4400 5104 4422
rect 5119 4406 5149 4422
rect 5177 4416 5183 4490
rect 5186 4416 5205 4560
rect 5220 4416 5226 4560
rect 5235 4490 5248 4560
rect 5300 4556 5322 4560
rect 5293 4534 5322 4548
rect 5375 4534 5391 4548
rect 5429 4544 5435 4546
rect 5442 4544 5550 4560
rect 5557 4544 5563 4546
rect 5571 4544 5586 4560
rect 5652 4554 5671 4557
rect 5293 4532 5391 4534
rect 5418 4532 5586 4544
rect 5601 4534 5617 4548
rect 5652 4535 5674 4554
rect 5684 4548 5700 4549
rect 5683 4546 5700 4548
rect 5684 4541 5700 4546
rect 5674 4534 5680 4535
rect 5683 4534 5712 4541
rect 5601 4533 5712 4534
rect 5601 4532 5718 4533
rect 5277 4524 5328 4532
rect 5375 4524 5409 4532
rect 5277 4512 5302 4524
rect 5309 4512 5328 4524
rect 5382 4522 5409 4524
rect 5418 4522 5639 4532
rect 5674 4529 5680 4532
rect 5382 4518 5639 4522
rect 5277 4504 5328 4512
rect 5375 4504 5639 4518
rect 5683 4524 5718 4532
rect 5229 4456 5248 4490
rect 5293 4496 5322 4504
rect 5293 4490 5310 4496
rect 5293 4488 5327 4490
rect 5375 4488 5391 4504
rect 5392 4494 5600 4504
rect 5601 4494 5617 4504
rect 5665 4500 5680 4515
rect 5683 4512 5684 4524
rect 5691 4512 5718 4524
rect 5683 4504 5718 4512
rect 5683 4503 5712 4504
rect 5403 4490 5617 4494
rect 5418 4488 5617 4490
rect 5652 4490 5665 4500
rect 5683 4490 5700 4503
rect 5652 4488 5700 4490
rect 5294 4484 5327 4488
rect 5290 4482 5327 4484
rect 5290 4481 5357 4482
rect 5290 4476 5321 4481
rect 5327 4476 5357 4481
rect 5290 4472 5357 4476
rect 5263 4469 5357 4472
rect 5263 4462 5312 4469
rect 5263 4456 5293 4462
rect 5312 4457 5317 4462
rect 5229 4440 5309 4456
rect 5321 4448 5357 4469
rect 5418 4464 5607 4488
rect 5652 4487 5699 4488
rect 5665 4482 5699 4487
rect 5433 4461 5607 4464
rect 5426 4458 5607 4461
rect 5635 4481 5699 4482
rect 5229 4438 5248 4440
rect 5263 4438 5297 4440
rect 5229 4422 5309 4438
rect 5229 4416 5248 4422
rect 4945 4390 5048 4400
rect 4899 4388 5048 4390
rect 5069 4388 5104 4400
rect 4738 4386 4900 4388
rect 4750 4366 4769 4386
rect 4784 4384 4814 4386
rect 4633 4358 4674 4366
rect 4756 4362 4769 4366
rect 4821 4370 4900 4386
rect 4932 4386 5104 4388
rect 4932 4370 5011 4386
rect 5018 4384 5048 4386
rect 4596 4348 4625 4358
rect 4639 4348 4668 4358
rect 4683 4348 4713 4362
rect 4756 4348 4799 4362
rect 4821 4358 5011 4370
rect 5076 4366 5082 4386
rect 4806 4348 4836 4358
rect 4837 4348 4995 4358
rect 4999 4348 5029 4358
rect 5033 4348 5063 4362
rect 5091 4348 5104 4386
rect 5176 4400 5205 4416
rect 5219 4400 5248 4416
rect 5263 4406 5293 4422
rect 5321 4400 5327 4448
rect 5330 4442 5349 4448
rect 5364 4442 5394 4450
rect 5330 4434 5394 4442
rect 5330 4418 5410 4434
rect 5426 4427 5488 4458
rect 5504 4427 5566 4458
rect 5635 4456 5684 4481
rect 5699 4456 5729 4472
rect 5598 4442 5628 4450
rect 5635 4448 5745 4456
rect 5598 4434 5643 4442
rect 5330 4416 5349 4418
rect 5364 4416 5410 4418
rect 5330 4400 5410 4416
rect 5437 4414 5472 4427
rect 5513 4424 5550 4427
rect 5513 4422 5555 4424
rect 5442 4411 5472 4414
rect 5451 4407 5458 4411
rect 5458 4406 5459 4407
rect 5417 4400 5427 4406
rect 5176 4392 5211 4400
rect 5176 4366 5177 4392
rect 5184 4366 5211 4392
rect 5119 4348 5149 4362
rect 5176 4358 5211 4366
rect 5213 4392 5254 4400
rect 5213 4366 5228 4392
rect 5235 4366 5254 4392
rect 5318 4388 5349 4400
rect 5364 4388 5467 4400
rect 5479 4390 5505 4416
rect 5520 4411 5550 4422
rect 5582 4418 5644 4434
rect 5582 4416 5628 4418
rect 5582 4400 5644 4416
rect 5656 4400 5662 4448
rect 5665 4440 5745 4448
rect 5665 4438 5684 4440
rect 5699 4438 5733 4440
rect 5665 4422 5745 4438
rect 5665 4400 5684 4422
rect 5699 4406 5729 4422
rect 5757 4416 5763 4490
rect 5766 4416 5785 4560
rect 5800 4416 5806 4560
rect 5815 4490 5828 4560
rect 5880 4556 5902 4560
rect 5873 4534 5902 4548
rect 5955 4534 5971 4548
rect 6009 4544 6015 4546
rect 6022 4544 6130 4560
rect 6137 4544 6143 4546
rect 6151 4544 6166 4560
rect 6232 4554 6251 4557
rect 5873 4532 5971 4534
rect 5998 4532 6166 4544
rect 6181 4534 6197 4548
rect 6232 4535 6254 4554
rect 6264 4548 6280 4549
rect 6263 4546 6280 4548
rect 6264 4541 6280 4546
rect 6254 4534 6260 4535
rect 6263 4534 6292 4541
rect 6181 4533 6292 4534
rect 6181 4532 6298 4533
rect 5857 4524 5908 4532
rect 5955 4524 5989 4532
rect 5857 4512 5882 4524
rect 5889 4512 5908 4524
rect 5962 4522 5989 4524
rect 5998 4522 6219 4532
rect 6254 4529 6260 4532
rect 5962 4518 6219 4522
rect 5857 4504 5908 4512
rect 5955 4504 6219 4518
rect 6263 4524 6298 4532
rect 5809 4456 5828 4490
rect 5873 4496 5902 4504
rect 5873 4490 5890 4496
rect 5873 4488 5907 4490
rect 5955 4488 5971 4504
rect 5972 4494 6180 4504
rect 6181 4494 6197 4504
rect 6245 4500 6260 4515
rect 6263 4512 6264 4524
rect 6271 4512 6298 4524
rect 6263 4504 6298 4512
rect 6263 4503 6292 4504
rect 5983 4490 6197 4494
rect 5998 4488 6197 4490
rect 6232 4490 6245 4500
rect 6263 4490 6280 4503
rect 6232 4488 6280 4490
rect 5874 4484 5907 4488
rect 5870 4482 5907 4484
rect 5870 4481 5937 4482
rect 5870 4476 5901 4481
rect 5907 4476 5937 4481
rect 5870 4472 5937 4476
rect 5843 4469 5937 4472
rect 5843 4462 5892 4469
rect 5843 4456 5873 4462
rect 5892 4457 5897 4462
rect 5809 4440 5889 4456
rect 5901 4448 5937 4469
rect 5998 4464 6187 4488
rect 6232 4487 6279 4488
rect 6245 4482 6279 4487
rect 6013 4461 6187 4464
rect 6006 4458 6187 4461
rect 6215 4481 6279 4482
rect 5809 4438 5828 4440
rect 5843 4438 5877 4440
rect 5809 4422 5889 4438
rect 5809 4416 5828 4422
rect 5525 4390 5628 4400
rect 5479 4388 5628 4390
rect 5649 4388 5684 4400
rect 5318 4386 5480 4388
rect 5330 4366 5349 4386
rect 5364 4384 5394 4386
rect 5213 4358 5254 4366
rect 5336 4362 5349 4366
rect 5401 4370 5480 4386
rect 5512 4386 5684 4388
rect 5512 4370 5591 4386
rect 5598 4384 5628 4386
rect 5176 4348 5205 4358
rect 5219 4348 5248 4358
rect 5263 4348 5293 4362
rect 5336 4348 5379 4362
rect 5401 4358 5591 4370
rect 5656 4366 5662 4386
rect 5386 4348 5416 4358
rect 5417 4348 5575 4358
rect 5579 4348 5609 4358
rect 5613 4348 5643 4362
rect 5671 4348 5684 4386
rect 5756 4400 5785 4416
rect 5799 4400 5828 4416
rect 5843 4406 5873 4422
rect 5901 4400 5907 4448
rect 5910 4442 5929 4448
rect 5944 4442 5974 4450
rect 5910 4434 5974 4442
rect 5910 4418 5990 4434
rect 6006 4427 6068 4458
rect 6084 4427 6146 4458
rect 6215 4456 6264 4481
rect 6279 4456 6309 4472
rect 6178 4442 6208 4450
rect 6215 4448 6325 4456
rect 6178 4434 6223 4442
rect 5910 4416 5929 4418
rect 5944 4416 5990 4418
rect 5910 4400 5990 4416
rect 6017 4414 6052 4427
rect 6093 4424 6130 4427
rect 6093 4422 6135 4424
rect 6022 4411 6052 4414
rect 6031 4407 6038 4411
rect 6038 4406 6039 4407
rect 5997 4400 6007 4406
rect 5756 4392 5791 4400
rect 5756 4366 5757 4392
rect 5764 4366 5791 4392
rect 5699 4348 5729 4362
rect 5756 4358 5791 4366
rect 5793 4392 5834 4400
rect 5793 4366 5808 4392
rect 5815 4366 5834 4392
rect 5898 4388 5929 4400
rect 5944 4388 6047 4400
rect 6059 4390 6085 4416
rect 6100 4411 6130 4422
rect 6162 4418 6224 4434
rect 6162 4416 6208 4418
rect 6162 4400 6224 4416
rect 6236 4400 6242 4448
rect 6245 4440 6325 4448
rect 6245 4438 6264 4440
rect 6279 4438 6313 4440
rect 6245 4422 6325 4438
rect 6245 4400 6264 4422
rect 6279 4406 6309 4422
rect 6337 4416 6343 4490
rect 6346 4416 6365 4560
rect 6380 4416 6386 4560
rect 6395 4490 6408 4560
rect 6460 4556 6482 4560
rect 6453 4534 6482 4548
rect 6535 4534 6551 4548
rect 6589 4544 6595 4546
rect 6602 4544 6710 4560
rect 6717 4544 6723 4546
rect 6731 4544 6746 4560
rect 6812 4554 6831 4557
rect 6453 4532 6551 4534
rect 6578 4532 6746 4544
rect 6761 4534 6777 4548
rect 6812 4535 6834 4554
rect 6844 4548 6860 4549
rect 6843 4546 6860 4548
rect 6844 4541 6860 4546
rect 6834 4534 6840 4535
rect 6843 4534 6872 4541
rect 6761 4533 6872 4534
rect 6761 4532 6878 4533
rect 6437 4524 6488 4532
rect 6535 4524 6569 4532
rect 6437 4512 6462 4524
rect 6469 4512 6488 4524
rect 6542 4522 6569 4524
rect 6578 4522 6799 4532
rect 6834 4529 6840 4532
rect 6542 4518 6799 4522
rect 6437 4504 6488 4512
rect 6535 4504 6799 4518
rect 6843 4524 6878 4532
rect 6389 4456 6408 4490
rect 6453 4496 6482 4504
rect 6453 4490 6470 4496
rect 6453 4488 6487 4490
rect 6535 4488 6551 4504
rect 6552 4494 6760 4504
rect 6761 4494 6777 4504
rect 6825 4500 6840 4515
rect 6843 4512 6844 4524
rect 6851 4512 6878 4524
rect 6843 4504 6878 4512
rect 6843 4503 6872 4504
rect 6563 4490 6777 4494
rect 6578 4488 6777 4490
rect 6812 4490 6825 4500
rect 6843 4490 6860 4503
rect 6812 4488 6860 4490
rect 6454 4484 6487 4488
rect 6450 4482 6487 4484
rect 6450 4481 6517 4482
rect 6450 4476 6481 4481
rect 6487 4476 6517 4481
rect 6450 4472 6517 4476
rect 6423 4469 6517 4472
rect 6423 4462 6472 4469
rect 6423 4456 6453 4462
rect 6472 4457 6477 4462
rect 6389 4440 6469 4456
rect 6481 4448 6517 4469
rect 6578 4464 6767 4488
rect 6812 4487 6859 4488
rect 6825 4482 6859 4487
rect 6593 4461 6767 4464
rect 6586 4458 6767 4461
rect 6795 4481 6859 4482
rect 6389 4438 6408 4440
rect 6423 4438 6457 4440
rect 6389 4422 6469 4438
rect 6389 4416 6408 4422
rect 6105 4390 6208 4400
rect 6059 4388 6208 4390
rect 6229 4388 6264 4400
rect 5898 4386 6060 4388
rect 5910 4366 5929 4386
rect 5944 4384 5974 4386
rect 5793 4358 5834 4366
rect 5916 4362 5929 4366
rect 5981 4370 6060 4386
rect 6092 4386 6264 4388
rect 6092 4370 6171 4386
rect 6178 4384 6208 4386
rect 5756 4348 5785 4358
rect 5799 4348 5828 4358
rect 5843 4348 5873 4362
rect 5916 4348 5959 4362
rect 5981 4358 6171 4370
rect 6236 4366 6242 4386
rect 5966 4348 5996 4358
rect 5997 4348 6155 4358
rect 6159 4348 6189 4358
rect 6193 4348 6223 4362
rect 6251 4348 6264 4386
rect 6336 4400 6365 4416
rect 6379 4400 6408 4416
rect 6423 4406 6453 4422
rect 6481 4400 6487 4448
rect 6490 4442 6509 4448
rect 6524 4442 6554 4450
rect 6490 4434 6554 4442
rect 6490 4418 6570 4434
rect 6586 4427 6648 4458
rect 6664 4427 6726 4458
rect 6795 4456 6844 4481
rect 6859 4456 6889 4472
rect 6758 4442 6788 4450
rect 6795 4448 6905 4456
rect 6758 4434 6803 4442
rect 6490 4416 6509 4418
rect 6524 4416 6570 4418
rect 6490 4400 6570 4416
rect 6597 4414 6632 4427
rect 6673 4424 6710 4427
rect 6673 4422 6715 4424
rect 6602 4411 6632 4414
rect 6611 4407 6618 4411
rect 6618 4406 6619 4407
rect 6577 4400 6587 4406
rect 6336 4392 6371 4400
rect 6336 4366 6337 4392
rect 6344 4366 6371 4392
rect 6279 4348 6309 4362
rect 6336 4358 6371 4366
rect 6373 4392 6414 4400
rect 6373 4366 6388 4392
rect 6395 4366 6414 4392
rect 6478 4388 6509 4400
rect 6524 4388 6627 4400
rect 6639 4390 6665 4416
rect 6680 4411 6710 4422
rect 6742 4418 6804 4434
rect 6742 4416 6788 4418
rect 6742 4400 6804 4416
rect 6816 4400 6822 4448
rect 6825 4440 6905 4448
rect 6825 4438 6844 4440
rect 6859 4438 6893 4440
rect 6825 4422 6905 4438
rect 6825 4400 6844 4422
rect 6859 4406 6889 4422
rect 6917 4416 6923 4490
rect 6926 4416 6945 4560
rect 6960 4416 6966 4560
rect 6975 4490 6988 4560
rect 7040 4556 7062 4560
rect 7033 4534 7062 4548
rect 7115 4534 7131 4548
rect 7169 4544 7175 4546
rect 7182 4544 7290 4560
rect 7297 4544 7303 4546
rect 7311 4544 7326 4560
rect 7392 4554 7411 4557
rect 7033 4532 7131 4534
rect 7158 4532 7326 4544
rect 7341 4534 7357 4548
rect 7392 4535 7414 4554
rect 7424 4548 7440 4549
rect 7423 4546 7440 4548
rect 7424 4541 7440 4546
rect 7414 4534 7420 4535
rect 7423 4534 7452 4541
rect 7341 4533 7452 4534
rect 7341 4532 7458 4533
rect 7017 4524 7068 4532
rect 7115 4524 7149 4532
rect 7017 4512 7042 4524
rect 7049 4512 7068 4524
rect 7122 4522 7149 4524
rect 7158 4522 7379 4532
rect 7414 4529 7420 4532
rect 7122 4518 7379 4522
rect 7017 4504 7068 4512
rect 7115 4504 7379 4518
rect 7423 4524 7458 4532
rect 6969 4456 6988 4490
rect 7033 4496 7062 4504
rect 7033 4490 7050 4496
rect 7033 4488 7067 4490
rect 7115 4488 7131 4504
rect 7132 4494 7340 4504
rect 7341 4494 7357 4504
rect 7405 4500 7420 4515
rect 7423 4512 7424 4524
rect 7431 4512 7458 4524
rect 7423 4504 7458 4512
rect 7423 4503 7452 4504
rect 7143 4490 7357 4494
rect 7158 4488 7357 4490
rect 7392 4490 7405 4500
rect 7423 4490 7440 4503
rect 7392 4488 7440 4490
rect 7034 4484 7067 4488
rect 7030 4482 7067 4484
rect 7030 4481 7097 4482
rect 7030 4476 7061 4481
rect 7067 4476 7097 4481
rect 7030 4472 7097 4476
rect 7003 4469 7097 4472
rect 7003 4462 7052 4469
rect 7003 4456 7033 4462
rect 7052 4457 7057 4462
rect 6969 4440 7049 4456
rect 7061 4448 7097 4469
rect 7158 4464 7347 4488
rect 7392 4487 7439 4488
rect 7405 4482 7439 4487
rect 7173 4461 7347 4464
rect 7166 4458 7347 4461
rect 7375 4481 7439 4482
rect 6969 4438 6988 4440
rect 7003 4438 7037 4440
rect 6969 4422 7049 4438
rect 6969 4416 6988 4422
rect 6685 4390 6788 4400
rect 6639 4388 6788 4390
rect 6809 4388 6844 4400
rect 6478 4386 6640 4388
rect 6490 4366 6509 4386
rect 6524 4384 6554 4386
rect 6373 4358 6414 4366
rect 6496 4362 6509 4366
rect 6561 4370 6640 4386
rect 6672 4386 6844 4388
rect 6672 4370 6751 4386
rect 6758 4384 6788 4386
rect 6336 4348 6365 4358
rect 6379 4348 6408 4358
rect 6423 4348 6453 4362
rect 6496 4348 6539 4362
rect 6561 4358 6751 4370
rect 6816 4366 6822 4386
rect 6546 4348 6576 4358
rect 6577 4348 6735 4358
rect 6739 4348 6769 4358
rect 6773 4348 6803 4362
rect 6831 4348 6844 4386
rect 6916 4400 6945 4416
rect 6959 4400 6988 4416
rect 7003 4406 7033 4422
rect 7061 4400 7067 4448
rect 7070 4442 7089 4448
rect 7104 4442 7134 4450
rect 7070 4434 7134 4442
rect 7070 4418 7150 4434
rect 7166 4427 7228 4458
rect 7244 4427 7306 4458
rect 7375 4456 7424 4481
rect 7439 4456 7469 4472
rect 7338 4442 7368 4450
rect 7375 4448 7485 4456
rect 7338 4434 7383 4442
rect 7070 4416 7089 4418
rect 7104 4416 7150 4418
rect 7070 4400 7150 4416
rect 7177 4414 7212 4427
rect 7253 4424 7290 4427
rect 7253 4422 7295 4424
rect 7182 4411 7212 4414
rect 7191 4407 7198 4411
rect 7198 4406 7199 4407
rect 7157 4400 7167 4406
rect 6916 4392 6951 4400
rect 6916 4366 6917 4392
rect 6924 4366 6951 4392
rect 6859 4348 6889 4362
rect 6916 4358 6951 4366
rect 6953 4392 6994 4400
rect 6953 4366 6968 4392
rect 6975 4366 6994 4392
rect 7058 4388 7089 4400
rect 7104 4388 7207 4400
rect 7219 4390 7245 4416
rect 7260 4411 7290 4422
rect 7322 4418 7384 4434
rect 7322 4416 7368 4418
rect 7322 4400 7384 4416
rect 7396 4400 7402 4448
rect 7405 4440 7485 4448
rect 7405 4438 7424 4440
rect 7439 4438 7473 4440
rect 7405 4422 7485 4438
rect 7405 4400 7424 4422
rect 7439 4406 7469 4422
rect 7497 4416 7503 4490
rect 7506 4416 7525 4560
rect 7540 4416 7546 4560
rect 7555 4490 7568 4560
rect 7620 4556 7642 4560
rect 7613 4534 7642 4548
rect 7695 4534 7711 4548
rect 7749 4544 7755 4546
rect 7762 4544 7870 4560
rect 7877 4544 7883 4546
rect 7891 4544 7906 4560
rect 7972 4554 7991 4557
rect 7613 4532 7711 4534
rect 7738 4532 7906 4544
rect 7921 4534 7937 4548
rect 7972 4535 7994 4554
rect 8004 4548 8020 4549
rect 8003 4546 8020 4548
rect 8004 4541 8020 4546
rect 7994 4534 8000 4535
rect 8003 4534 8032 4541
rect 7921 4533 8032 4534
rect 7921 4532 8038 4533
rect 7597 4524 7648 4532
rect 7695 4524 7729 4532
rect 7597 4512 7622 4524
rect 7629 4512 7648 4524
rect 7702 4522 7729 4524
rect 7738 4522 7959 4532
rect 7994 4529 8000 4532
rect 7702 4518 7959 4522
rect 7597 4504 7648 4512
rect 7695 4504 7959 4518
rect 8003 4524 8038 4532
rect 7549 4456 7568 4490
rect 7613 4496 7642 4504
rect 7613 4490 7630 4496
rect 7613 4488 7647 4490
rect 7695 4488 7711 4504
rect 7712 4494 7920 4504
rect 7921 4494 7937 4504
rect 7985 4500 8000 4515
rect 8003 4512 8004 4524
rect 8011 4512 8038 4524
rect 8003 4504 8038 4512
rect 8003 4503 8032 4504
rect 7723 4490 7937 4494
rect 7738 4488 7937 4490
rect 7972 4490 7985 4500
rect 8003 4490 8020 4503
rect 7972 4488 8020 4490
rect 7614 4484 7647 4488
rect 7610 4482 7647 4484
rect 7610 4481 7677 4482
rect 7610 4476 7641 4481
rect 7647 4476 7677 4481
rect 7610 4472 7677 4476
rect 7583 4469 7677 4472
rect 7583 4462 7632 4469
rect 7583 4456 7613 4462
rect 7632 4457 7637 4462
rect 7549 4440 7629 4456
rect 7641 4448 7677 4469
rect 7738 4464 7927 4488
rect 7972 4487 8019 4488
rect 7985 4482 8019 4487
rect 7753 4461 7927 4464
rect 7746 4458 7927 4461
rect 7955 4481 8019 4482
rect 7549 4438 7568 4440
rect 7583 4438 7617 4440
rect 7549 4422 7629 4438
rect 7549 4416 7568 4422
rect 7265 4390 7368 4400
rect 7219 4388 7368 4390
rect 7389 4388 7424 4400
rect 7058 4386 7220 4388
rect 7070 4366 7089 4386
rect 7104 4384 7134 4386
rect 6953 4358 6994 4366
rect 7076 4362 7089 4366
rect 7141 4370 7220 4386
rect 7252 4386 7424 4388
rect 7252 4370 7331 4386
rect 7338 4384 7368 4386
rect 6916 4348 6945 4358
rect 6959 4348 6988 4358
rect 7003 4348 7033 4362
rect 7076 4348 7119 4362
rect 7141 4358 7331 4370
rect 7396 4366 7402 4386
rect 7126 4348 7156 4358
rect 7157 4348 7315 4358
rect 7319 4348 7349 4358
rect 7353 4348 7383 4362
rect 7411 4348 7424 4386
rect 7496 4400 7525 4416
rect 7539 4400 7568 4416
rect 7583 4406 7613 4422
rect 7641 4400 7647 4448
rect 7650 4442 7669 4448
rect 7684 4442 7714 4450
rect 7650 4434 7714 4442
rect 7650 4418 7730 4434
rect 7746 4427 7808 4458
rect 7824 4427 7886 4458
rect 7955 4456 8004 4481
rect 8019 4456 8049 4472
rect 7918 4442 7948 4450
rect 7955 4448 8065 4456
rect 7918 4434 7963 4442
rect 7650 4416 7669 4418
rect 7684 4416 7730 4418
rect 7650 4400 7730 4416
rect 7757 4414 7792 4427
rect 7833 4424 7870 4427
rect 7833 4422 7875 4424
rect 7762 4411 7792 4414
rect 7771 4407 7778 4411
rect 7778 4406 7779 4407
rect 7737 4400 7747 4406
rect 7496 4392 7531 4400
rect 7496 4366 7497 4392
rect 7504 4366 7531 4392
rect 7439 4348 7469 4362
rect 7496 4358 7531 4366
rect 7533 4392 7574 4400
rect 7533 4366 7548 4392
rect 7555 4366 7574 4392
rect 7638 4388 7669 4400
rect 7684 4388 7787 4400
rect 7799 4390 7825 4416
rect 7840 4411 7870 4422
rect 7902 4418 7964 4434
rect 7902 4416 7948 4418
rect 7902 4400 7964 4416
rect 7976 4400 7982 4448
rect 7985 4440 8065 4448
rect 7985 4438 8004 4440
rect 8019 4438 8053 4440
rect 7985 4422 8065 4438
rect 7985 4400 8004 4422
rect 8019 4406 8049 4422
rect 8077 4416 8083 4490
rect 8086 4416 8105 4560
rect 8120 4416 8126 4560
rect 8135 4490 8148 4560
rect 8200 4556 8222 4560
rect 8193 4534 8222 4548
rect 8275 4534 8291 4548
rect 8329 4544 8335 4546
rect 8342 4544 8450 4560
rect 8457 4544 8463 4546
rect 8471 4544 8486 4560
rect 8552 4554 8571 4557
rect 8193 4532 8291 4534
rect 8318 4532 8486 4544
rect 8501 4534 8517 4548
rect 8552 4535 8574 4554
rect 8584 4548 8600 4549
rect 8583 4546 8600 4548
rect 8584 4541 8600 4546
rect 8574 4534 8580 4535
rect 8583 4534 8612 4541
rect 8501 4533 8612 4534
rect 8501 4532 8618 4533
rect 8177 4524 8228 4532
rect 8275 4524 8309 4532
rect 8177 4512 8202 4524
rect 8209 4512 8228 4524
rect 8282 4522 8309 4524
rect 8318 4522 8539 4532
rect 8574 4529 8580 4532
rect 8282 4518 8539 4522
rect 8177 4504 8228 4512
rect 8275 4504 8539 4518
rect 8583 4524 8618 4532
rect 8129 4456 8148 4490
rect 8193 4496 8222 4504
rect 8193 4490 8210 4496
rect 8193 4488 8227 4490
rect 8275 4488 8291 4504
rect 8292 4494 8500 4504
rect 8501 4494 8517 4504
rect 8565 4500 8580 4515
rect 8583 4512 8584 4524
rect 8591 4512 8618 4524
rect 8583 4504 8618 4512
rect 8583 4503 8612 4504
rect 8303 4490 8517 4494
rect 8318 4488 8517 4490
rect 8552 4490 8565 4500
rect 8583 4490 8600 4503
rect 8552 4488 8600 4490
rect 8194 4484 8227 4488
rect 8190 4482 8227 4484
rect 8190 4481 8257 4482
rect 8190 4476 8221 4481
rect 8227 4476 8257 4481
rect 8190 4472 8257 4476
rect 8163 4469 8257 4472
rect 8163 4462 8212 4469
rect 8163 4456 8193 4462
rect 8212 4457 8217 4462
rect 8129 4440 8209 4456
rect 8221 4448 8257 4469
rect 8318 4464 8507 4488
rect 8552 4487 8599 4488
rect 8565 4482 8599 4487
rect 8333 4461 8507 4464
rect 8326 4458 8507 4461
rect 8535 4481 8599 4482
rect 8129 4438 8148 4440
rect 8163 4438 8197 4440
rect 8129 4422 8209 4438
rect 8129 4416 8148 4422
rect 7845 4390 7948 4400
rect 7799 4388 7948 4390
rect 7969 4388 8004 4400
rect 7638 4386 7800 4388
rect 7650 4366 7669 4386
rect 7684 4384 7714 4386
rect 7533 4358 7574 4366
rect 7656 4362 7669 4366
rect 7721 4370 7800 4386
rect 7832 4386 8004 4388
rect 7832 4370 7911 4386
rect 7918 4384 7948 4386
rect 7496 4348 7525 4358
rect 7539 4348 7568 4358
rect 7583 4348 7613 4362
rect 7656 4348 7699 4362
rect 7721 4358 7911 4370
rect 7976 4366 7982 4386
rect 7706 4348 7736 4358
rect 7737 4348 7895 4358
rect 7899 4348 7929 4358
rect 7933 4348 7963 4362
rect 7991 4348 8004 4386
rect 8076 4400 8105 4416
rect 8119 4400 8148 4416
rect 8163 4406 8193 4422
rect 8221 4400 8227 4448
rect 8230 4442 8249 4448
rect 8264 4442 8294 4450
rect 8230 4434 8294 4442
rect 8230 4418 8310 4434
rect 8326 4427 8388 4458
rect 8404 4427 8466 4458
rect 8535 4456 8584 4481
rect 8599 4456 8629 4472
rect 8498 4442 8528 4450
rect 8535 4448 8645 4456
rect 8498 4434 8543 4442
rect 8230 4416 8249 4418
rect 8264 4416 8310 4418
rect 8230 4400 8310 4416
rect 8337 4414 8372 4427
rect 8413 4424 8450 4427
rect 8413 4422 8455 4424
rect 8342 4411 8372 4414
rect 8351 4407 8358 4411
rect 8358 4406 8359 4407
rect 8317 4400 8327 4406
rect 8076 4392 8111 4400
rect 8076 4366 8077 4392
rect 8084 4366 8111 4392
rect 8019 4348 8049 4362
rect 8076 4358 8111 4366
rect 8113 4392 8154 4400
rect 8113 4366 8128 4392
rect 8135 4366 8154 4392
rect 8218 4388 8249 4400
rect 8264 4388 8367 4400
rect 8379 4390 8405 4416
rect 8420 4411 8450 4422
rect 8482 4418 8544 4434
rect 8482 4416 8528 4418
rect 8482 4400 8544 4416
rect 8556 4400 8562 4448
rect 8565 4440 8645 4448
rect 8565 4438 8584 4440
rect 8599 4438 8633 4440
rect 8565 4422 8645 4438
rect 8565 4400 8584 4422
rect 8599 4406 8629 4422
rect 8657 4416 8663 4490
rect 8666 4416 8685 4560
rect 8700 4416 8706 4560
rect 8715 4490 8728 4560
rect 8780 4556 8802 4560
rect 8773 4534 8802 4548
rect 8855 4534 8871 4548
rect 8909 4544 8915 4546
rect 8922 4544 9030 4560
rect 9037 4544 9043 4546
rect 9051 4544 9066 4560
rect 9132 4554 9151 4557
rect 8773 4532 8871 4534
rect 8898 4532 9066 4544
rect 9081 4534 9097 4548
rect 9132 4535 9154 4554
rect 9164 4548 9180 4549
rect 9163 4546 9180 4548
rect 9164 4541 9180 4546
rect 9154 4534 9160 4535
rect 9163 4534 9192 4541
rect 9081 4533 9192 4534
rect 9081 4532 9198 4533
rect 8757 4524 8808 4532
rect 8855 4524 8889 4532
rect 8757 4512 8782 4524
rect 8789 4512 8808 4524
rect 8862 4522 8889 4524
rect 8898 4522 9119 4532
rect 9154 4529 9160 4532
rect 8862 4518 9119 4522
rect 8757 4504 8808 4512
rect 8855 4504 9119 4518
rect 9163 4524 9198 4532
rect 8709 4456 8728 4490
rect 8773 4496 8802 4504
rect 8773 4490 8790 4496
rect 8773 4488 8807 4490
rect 8855 4488 8871 4504
rect 8872 4494 9080 4504
rect 9081 4494 9097 4504
rect 9145 4500 9160 4515
rect 9163 4512 9164 4524
rect 9171 4512 9198 4524
rect 9163 4504 9198 4512
rect 9163 4503 9192 4504
rect 8883 4490 9097 4494
rect 8898 4488 9097 4490
rect 9132 4490 9145 4500
rect 9163 4490 9180 4503
rect 9132 4488 9180 4490
rect 8774 4484 8807 4488
rect 8770 4482 8807 4484
rect 8770 4481 8837 4482
rect 8770 4476 8801 4481
rect 8807 4476 8837 4481
rect 8770 4472 8837 4476
rect 8743 4469 8837 4472
rect 8743 4462 8792 4469
rect 8743 4456 8773 4462
rect 8792 4457 8797 4462
rect 8709 4440 8789 4456
rect 8801 4448 8837 4469
rect 8898 4464 9087 4488
rect 9132 4487 9179 4488
rect 9145 4482 9179 4487
rect 8913 4461 9087 4464
rect 8906 4458 9087 4461
rect 9115 4481 9179 4482
rect 8709 4438 8728 4440
rect 8743 4438 8777 4440
rect 8709 4422 8789 4438
rect 8709 4416 8728 4422
rect 8425 4390 8528 4400
rect 8379 4388 8528 4390
rect 8549 4388 8584 4400
rect 8218 4386 8380 4388
rect 8230 4366 8249 4386
rect 8264 4384 8294 4386
rect 8113 4358 8154 4366
rect 8236 4362 8249 4366
rect 8301 4370 8380 4386
rect 8412 4386 8584 4388
rect 8412 4370 8491 4386
rect 8498 4384 8528 4386
rect 8076 4348 8105 4358
rect 8119 4348 8148 4358
rect 8163 4348 8193 4362
rect 8236 4348 8279 4362
rect 8301 4358 8491 4370
rect 8556 4366 8562 4386
rect 8286 4348 8316 4358
rect 8317 4348 8475 4358
rect 8479 4348 8509 4358
rect 8513 4348 8543 4362
rect 8571 4348 8584 4386
rect 8656 4400 8685 4416
rect 8699 4400 8728 4416
rect 8743 4406 8773 4422
rect 8801 4400 8807 4448
rect 8810 4442 8829 4448
rect 8844 4442 8874 4450
rect 8810 4434 8874 4442
rect 8810 4418 8890 4434
rect 8906 4427 8968 4458
rect 8984 4427 9046 4458
rect 9115 4456 9164 4481
rect 9179 4456 9209 4472
rect 9078 4442 9108 4450
rect 9115 4448 9225 4456
rect 9078 4434 9123 4442
rect 8810 4416 8829 4418
rect 8844 4416 8890 4418
rect 8810 4400 8890 4416
rect 8917 4414 8952 4427
rect 8993 4424 9030 4427
rect 8993 4422 9035 4424
rect 8922 4411 8952 4414
rect 8931 4407 8938 4411
rect 8938 4406 8939 4407
rect 8897 4400 8907 4406
rect 8656 4392 8691 4400
rect 8656 4366 8657 4392
rect 8664 4366 8691 4392
rect 8599 4348 8629 4362
rect 8656 4358 8691 4366
rect 8693 4392 8734 4400
rect 8693 4366 8708 4392
rect 8715 4366 8734 4392
rect 8798 4388 8829 4400
rect 8844 4388 8947 4400
rect 8959 4390 8985 4416
rect 9000 4411 9030 4422
rect 9062 4418 9124 4434
rect 9062 4416 9108 4418
rect 9062 4400 9124 4416
rect 9136 4400 9142 4448
rect 9145 4440 9225 4448
rect 9145 4438 9164 4440
rect 9179 4438 9213 4440
rect 9145 4422 9225 4438
rect 9145 4400 9164 4422
rect 9179 4406 9209 4422
rect 9237 4416 9243 4490
rect 9246 4416 9265 4560
rect 9280 4416 9286 4560
rect 9295 4490 9308 4560
rect 9360 4556 9382 4560
rect 9353 4534 9382 4548
rect 9435 4534 9451 4548
rect 9489 4544 9495 4546
rect 9502 4544 9610 4560
rect 9617 4544 9623 4546
rect 9631 4544 9646 4560
rect 9712 4554 9731 4557
rect 9353 4532 9451 4534
rect 9478 4532 9646 4544
rect 9661 4534 9677 4548
rect 9712 4535 9734 4554
rect 9744 4548 9760 4549
rect 9743 4546 9760 4548
rect 9744 4541 9760 4546
rect 9734 4534 9740 4535
rect 9743 4534 9772 4541
rect 9661 4533 9772 4534
rect 9661 4532 9778 4533
rect 9337 4524 9388 4532
rect 9435 4524 9469 4532
rect 9337 4512 9362 4524
rect 9369 4512 9388 4524
rect 9442 4522 9469 4524
rect 9478 4522 9699 4532
rect 9734 4529 9740 4532
rect 9442 4518 9699 4522
rect 9337 4504 9388 4512
rect 9435 4504 9699 4518
rect 9743 4524 9778 4532
rect 9289 4456 9308 4490
rect 9353 4496 9382 4504
rect 9353 4490 9370 4496
rect 9353 4488 9387 4490
rect 9435 4488 9451 4504
rect 9452 4494 9660 4504
rect 9661 4494 9677 4504
rect 9725 4500 9740 4515
rect 9743 4512 9744 4524
rect 9751 4512 9778 4524
rect 9743 4504 9778 4512
rect 9743 4503 9772 4504
rect 9463 4490 9677 4494
rect 9478 4488 9677 4490
rect 9712 4490 9725 4500
rect 9743 4490 9760 4503
rect 9712 4488 9760 4490
rect 9354 4484 9387 4488
rect 9350 4482 9387 4484
rect 9350 4481 9417 4482
rect 9350 4476 9381 4481
rect 9387 4476 9417 4481
rect 9350 4472 9417 4476
rect 9323 4469 9417 4472
rect 9323 4462 9372 4469
rect 9323 4456 9353 4462
rect 9372 4457 9377 4462
rect 9289 4440 9369 4456
rect 9381 4448 9417 4469
rect 9478 4464 9667 4488
rect 9712 4487 9759 4488
rect 9725 4482 9759 4487
rect 9493 4461 9667 4464
rect 9486 4458 9667 4461
rect 9695 4481 9759 4482
rect 9289 4438 9308 4440
rect 9323 4438 9357 4440
rect 9289 4422 9369 4438
rect 9289 4416 9308 4422
rect 9005 4390 9108 4400
rect 8959 4388 9108 4390
rect 9129 4388 9164 4400
rect 8798 4386 8960 4388
rect 8810 4366 8829 4386
rect 8844 4384 8874 4386
rect 8693 4358 8734 4366
rect 8816 4362 8829 4366
rect 8881 4370 8960 4386
rect 8992 4386 9164 4388
rect 8992 4370 9071 4386
rect 9078 4384 9108 4386
rect 8656 4348 8685 4358
rect 8699 4348 8728 4358
rect 8743 4348 8773 4362
rect 8816 4348 8859 4362
rect 8881 4358 9071 4370
rect 9136 4366 9142 4386
rect 8866 4348 8896 4358
rect 8897 4348 9055 4358
rect 9059 4348 9089 4358
rect 9093 4348 9123 4362
rect 9151 4348 9164 4386
rect 9236 4400 9265 4416
rect 9279 4400 9308 4416
rect 9323 4406 9353 4422
rect 9381 4400 9387 4448
rect 9390 4442 9409 4448
rect 9424 4442 9454 4450
rect 9390 4434 9454 4442
rect 9390 4418 9470 4434
rect 9486 4427 9548 4458
rect 9564 4427 9626 4458
rect 9695 4456 9744 4481
rect 9759 4456 9789 4472
rect 9658 4442 9688 4450
rect 9695 4448 9805 4456
rect 9658 4434 9703 4442
rect 9390 4416 9409 4418
rect 9424 4416 9470 4418
rect 9390 4400 9470 4416
rect 9497 4414 9532 4427
rect 9573 4424 9610 4427
rect 9573 4422 9615 4424
rect 9502 4411 9532 4414
rect 9511 4407 9518 4411
rect 9518 4406 9519 4407
rect 9477 4400 9487 4406
rect 9236 4392 9271 4400
rect 9236 4366 9237 4392
rect 9244 4366 9271 4392
rect 9179 4348 9209 4362
rect 9236 4358 9271 4366
rect 9273 4392 9314 4400
rect 9273 4366 9288 4392
rect 9295 4366 9314 4392
rect 9378 4388 9409 4400
rect 9424 4388 9527 4400
rect 9539 4390 9565 4416
rect 9580 4411 9610 4422
rect 9642 4418 9704 4434
rect 9642 4416 9688 4418
rect 9642 4400 9704 4416
rect 9716 4400 9722 4448
rect 9725 4440 9805 4448
rect 9725 4438 9744 4440
rect 9759 4438 9793 4440
rect 9725 4422 9805 4438
rect 9725 4400 9744 4422
rect 9759 4406 9789 4422
rect 9817 4416 9823 4490
rect 9826 4416 9845 4560
rect 9860 4416 9866 4560
rect 9875 4490 9888 4560
rect 9940 4556 9962 4560
rect 9933 4534 9962 4548
rect 10015 4534 10031 4548
rect 10069 4544 10075 4546
rect 10082 4544 10190 4560
rect 10197 4544 10203 4546
rect 10211 4544 10226 4560
rect 10292 4554 10311 4557
rect 9933 4532 10031 4534
rect 10058 4532 10226 4544
rect 10241 4534 10257 4548
rect 10292 4535 10314 4554
rect 10324 4548 10340 4549
rect 10323 4546 10340 4548
rect 10324 4541 10340 4546
rect 10314 4534 10320 4535
rect 10323 4534 10352 4541
rect 10241 4533 10352 4534
rect 10241 4532 10358 4533
rect 9917 4524 9968 4532
rect 10015 4524 10049 4532
rect 9917 4512 9942 4524
rect 9949 4512 9968 4524
rect 10022 4522 10049 4524
rect 10058 4522 10279 4532
rect 10314 4529 10320 4532
rect 10022 4518 10279 4522
rect 9917 4504 9968 4512
rect 10015 4504 10279 4518
rect 10323 4524 10358 4532
rect 9869 4456 9888 4490
rect 9933 4496 9962 4504
rect 9933 4490 9950 4496
rect 9933 4488 9967 4490
rect 10015 4488 10031 4504
rect 10032 4494 10240 4504
rect 10241 4494 10257 4504
rect 10305 4500 10320 4515
rect 10323 4512 10324 4524
rect 10331 4512 10358 4524
rect 10323 4504 10358 4512
rect 10323 4503 10352 4504
rect 10043 4490 10257 4494
rect 10058 4488 10257 4490
rect 10292 4490 10305 4500
rect 10323 4490 10340 4503
rect 10292 4488 10340 4490
rect 9934 4484 9967 4488
rect 9930 4482 9967 4484
rect 9930 4481 9997 4482
rect 9930 4476 9961 4481
rect 9967 4476 9997 4481
rect 9930 4472 9997 4476
rect 9903 4469 9997 4472
rect 9903 4462 9952 4469
rect 9903 4456 9933 4462
rect 9952 4457 9957 4462
rect 9869 4440 9949 4456
rect 9961 4448 9997 4469
rect 10058 4464 10247 4488
rect 10292 4487 10339 4488
rect 10305 4482 10339 4487
rect 10073 4461 10247 4464
rect 10066 4458 10247 4461
rect 10275 4481 10339 4482
rect 9869 4438 9888 4440
rect 9903 4438 9937 4440
rect 9869 4422 9949 4438
rect 9869 4416 9888 4422
rect 9585 4390 9688 4400
rect 9539 4388 9688 4390
rect 9709 4388 9744 4400
rect 9378 4386 9540 4388
rect 9390 4366 9409 4386
rect 9424 4384 9454 4386
rect 9273 4358 9314 4366
rect 9396 4362 9409 4366
rect 9461 4370 9540 4386
rect 9572 4386 9744 4388
rect 9572 4370 9651 4386
rect 9658 4384 9688 4386
rect 9236 4348 9265 4358
rect 9279 4348 9308 4358
rect 9323 4348 9353 4362
rect 9396 4348 9439 4362
rect 9461 4358 9651 4370
rect 9716 4366 9722 4386
rect 9446 4348 9476 4358
rect 9477 4348 9635 4358
rect 9639 4348 9669 4358
rect 9673 4348 9703 4362
rect 9731 4348 9744 4386
rect 9816 4400 9845 4416
rect 9859 4400 9888 4416
rect 9903 4406 9933 4422
rect 9961 4400 9967 4448
rect 9970 4442 9989 4448
rect 10004 4442 10034 4450
rect 9970 4434 10034 4442
rect 9970 4418 10050 4434
rect 10066 4427 10128 4458
rect 10144 4427 10206 4458
rect 10275 4456 10324 4481
rect 10339 4456 10369 4472
rect 10238 4442 10268 4450
rect 10275 4448 10385 4456
rect 10238 4434 10283 4442
rect 9970 4416 9989 4418
rect 10004 4416 10050 4418
rect 9970 4400 10050 4416
rect 10077 4414 10112 4427
rect 10153 4424 10190 4427
rect 10153 4422 10195 4424
rect 10082 4411 10112 4414
rect 10091 4407 10098 4411
rect 10098 4406 10099 4407
rect 10057 4400 10067 4406
rect 9816 4392 9851 4400
rect 9816 4366 9817 4392
rect 9824 4366 9851 4392
rect 9759 4348 9789 4362
rect 9816 4358 9851 4366
rect 9853 4392 9894 4400
rect 9853 4366 9868 4392
rect 9875 4366 9894 4392
rect 9958 4388 9989 4400
rect 10004 4388 10107 4400
rect 10119 4390 10145 4416
rect 10160 4411 10190 4422
rect 10222 4418 10284 4434
rect 10222 4416 10268 4418
rect 10222 4400 10284 4416
rect 10296 4400 10302 4448
rect 10305 4440 10385 4448
rect 10305 4438 10324 4440
rect 10339 4438 10373 4440
rect 10305 4422 10385 4438
rect 10305 4400 10324 4422
rect 10339 4406 10369 4422
rect 10397 4416 10403 4490
rect 10406 4416 10425 4560
rect 10440 4416 10446 4560
rect 10455 4490 10468 4560
rect 10520 4556 10542 4560
rect 10513 4534 10542 4548
rect 10595 4534 10611 4548
rect 10649 4544 10655 4546
rect 10662 4544 10770 4560
rect 10777 4544 10783 4546
rect 10791 4544 10806 4560
rect 10872 4554 10891 4557
rect 10513 4532 10611 4534
rect 10638 4532 10806 4544
rect 10821 4534 10837 4548
rect 10872 4535 10894 4554
rect 10904 4548 10920 4549
rect 10903 4546 10920 4548
rect 10904 4541 10920 4546
rect 10894 4534 10900 4535
rect 10903 4534 10932 4541
rect 10821 4533 10932 4534
rect 10821 4532 10938 4533
rect 10497 4524 10548 4532
rect 10595 4524 10629 4532
rect 10497 4512 10522 4524
rect 10529 4512 10548 4524
rect 10602 4522 10629 4524
rect 10638 4522 10859 4532
rect 10894 4529 10900 4532
rect 10602 4518 10859 4522
rect 10497 4504 10548 4512
rect 10595 4504 10859 4518
rect 10903 4524 10938 4532
rect 10449 4456 10468 4490
rect 10513 4496 10542 4504
rect 10513 4490 10530 4496
rect 10513 4488 10547 4490
rect 10595 4488 10611 4504
rect 10612 4494 10820 4504
rect 10821 4494 10837 4504
rect 10885 4500 10900 4515
rect 10903 4512 10904 4524
rect 10911 4512 10938 4524
rect 10903 4504 10938 4512
rect 10903 4503 10932 4504
rect 10623 4490 10837 4494
rect 10638 4488 10837 4490
rect 10872 4490 10885 4500
rect 10903 4490 10920 4503
rect 10872 4488 10920 4490
rect 10514 4484 10547 4488
rect 10510 4482 10547 4484
rect 10510 4481 10577 4482
rect 10510 4476 10541 4481
rect 10547 4476 10577 4481
rect 10510 4472 10577 4476
rect 10483 4469 10577 4472
rect 10483 4462 10532 4469
rect 10483 4456 10513 4462
rect 10532 4457 10537 4462
rect 10449 4440 10529 4456
rect 10541 4448 10577 4469
rect 10638 4464 10827 4488
rect 10872 4487 10919 4488
rect 10885 4482 10919 4487
rect 10653 4461 10827 4464
rect 10646 4458 10827 4461
rect 10855 4481 10919 4482
rect 10449 4438 10468 4440
rect 10483 4438 10517 4440
rect 10449 4422 10529 4438
rect 10449 4416 10468 4422
rect 10165 4390 10268 4400
rect 10119 4388 10268 4390
rect 10289 4388 10324 4400
rect 9958 4386 10120 4388
rect 9970 4366 9989 4386
rect 10004 4384 10034 4386
rect 9853 4358 9894 4366
rect 9976 4362 9989 4366
rect 10041 4370 10120 4386
rect 10152 4386 10324 4388
rect 10152 4370 10231 4386
rect 10238 4384 10268 4386
rect 9816 4348 9845 4358
rect 9859 4348 9888 4358
rect 9903 4348 9933 4362
rect 9976 4348 10019 4362
rect 10041 4358 10231 4370
rect 10296 4366 10302 4386
rect 10026 4348 10056 4358
rect 10057 4348 10215 4358
rect 10219 4348 10249 4358
rect 10253 4348 10283 4362
rect 10311 4348 10324 4386
rect 10396 4400 10425 4416
rect 10439 4400 10468 4416
rect 10483 4406 10513 4422
rect 10541 4400 10547 4448
rect 10550 4442 10569 4448
rect 10584 4442 10614 4450
rect 10550 4434 10614 4442
rect 10550 4418 10630 4434
rect 10646 4427 10708 4458
rect 10724 4427 10786 4458
rect 10855 4456 10904 4481
rect 10919 4456 10949 4472
rect 10818 4442 10848 4450
rect 10855 4448 10965 4456
rect 10818 4434 10863 4442
rect 10550 4416 10569 4418
rect 10584 4416 10630 4418
rect 10550 4400 10630 4416
rect 10657 4414 10692 4427
rect 10733 4424 10770 4427
rect 10733 4422 10775 4424
rect 10662 4411 10692 4414
rect 10671 4407 10678 4411
rect 10678 4406 10679 4407
rect 10637 4400 10647 4406
rect 10396 4392 10431 4400
rect 10396 4366 10397 4392
rect 10404 4366 10431 4392
rect 10339 4348 10369 4362
rect 10396 4358 10431 4366
rect 10433 4392 10474 4400
rect 10433 4366 10448 4392
rect 10455 4366 10474 4392
rect 10538 4388 10569 4400
rect 10584 4388 10687 4400
rect 10699 4390 10725 4416
rect 10740 4411 10770 4422
rect 10802 4418 10864 4434
rect 10802 4416 10848 4418
rect 10802 4400 10864 4416
rect 10876 4400 10882 4448
rect 10885 4440 10965 4448
rect 10885 4438 10904 4440
rect 10919 4438 10953 4440
rect 10885 4422 10965 4438
rect 10885 4400 10904 4422
rect 10919 4406 10949 4422
rect 10977 4416 10983 4490
rect 10986 4416 11005 4560
rect 11020 4416 11026 4560
rect 11035 4490 11048 4560
rect 11100 4556 11122 4560
rect 11093 4534 11122 4548
rect 11175 4534 11191 4548
rect 11229 4544 11235 4546
rect 11242 4544 11350 4560
rect 11357 4544 11363 4546
rect 11371 4544 11386 4560
rect 11452 4554 11471 4557
rect 11093 4532 11191 4534
rect 11218 4532 11386 4544
rect 11401 4534 11417 4548
rect 11452 4535 11474 4554
rect 11484 4548 11500 4549
rect 11483 4546 11500 4548
rect 11484 4541 11500 4546
rect 11474 4534 11480 4535
rect 11483 4534 11512 4541
rect 11401 4533 11512 4534
rect 11401 4532 11518 4533
rect 11077 4524 11128 4532
rect 11175 4524 11209 4532
rect 11077 4512 11102 4524
rect 11109 4512 11128 4524
rect 11182 4522 11209 4524
rect 11218 4522 11439 4532
rect 11474 4529 11480 4532
rect 11182 4518 11439 4522
rect 11077 4504 11128 4512
rect 11175 4504 11439 4518
rect 11483 4524 11518 4532
rect 11029 4456 11048 4490
rect 11093 4496 11122 4504
rect 11093 4490 11110 4496
rect 11093 4488 11127 4490
rect 11175 4488 11191 4504
rect 11192 4494 11400 4504
rect 11401 4494 11417 4504
rect 11465 4500 11480 4515
rect 11483 4512 11484 4524
rect 11491 4512 11518 4524
rect 11483 4504 11518 4512
rect 11483 4503 11512 4504
rect 11203 4490 11417 4494
rect 11218 4488 11417 4490
rect 11452 4490 11465 4500
rect 11483 4490 11500 4503
rect 11452 4488 11500 4490
rect 11094 4484 11127 4488
rect 11090 4482 11127 4484
rect 11090 4481 11157 4482
rect 11090 4476 11121 4481
rect 11127 4476 11157 4481
rect 11090 4472 11157 4476
rect 11063 4469 11157 4472
rect 11063 4462 11112 4469
rect 11063 4456 11093 4462
rect 11112 4457 11117 4462
rect 11029 4440 11109 4456
rect 11121 4448 11157 4469
rect 11218 4464 11407 4488
rect 11452 4487 11499 4488
rect 11465 4482 11499 4487
rect 11233 4461 11407 4464
rect 11226 4458 11407 4461
rect 11435 4481 11499 4482
rect 11029 4438 11048 4440
rect 11063 4438 11097 4440
rect 11029 4422 11109 4438
rect 11029 4416 11048 4422
rect 10745 4390 10848 4400
rect 10699 4388 10848 4390
rect 10869 4388 10904 4400
rect 10538 4386 10700 4388
rect 10550 4366 10569 4386
rect 10584 4384 10614 4386
rect 10433 4358 10474 4366
rect 10556 4362 10569 4366
rect 10621 4370 10700 4386
rect 10732 4386 10904 4388
rect 10732 4370 10811 4386
rect 10818 4384 10848 4386
rect 10396 4348 10425 4358
rect 10439 4348 10468 4358
rect 10483 4348 10513 4362
rect 10556 4348 10599 4362
rect 10621 4358 10811 4370
rect 10876 4366 10882 4386
rect 10606 4348 10636 4358
rect 10637 4348 10795 4358
rect 10799 4348 10829 4358
rect 10833 4348 10863 4362
rect 10891 4348 10904 4386
rect 10976 4400 11005 4416
rect 11019 4400 11048 4416
rect 11063 4406 11093 4422
rect 11121 4400 11127 4448
rect 11130 4442 11149 4448
rect 11164 4442 11194 4450
rect 11130 4434 11194 4442
rect 11130 4418 11210 4434
rect 11226 4427 11288 4458
rect 11304 4427 11366 4458
rect 11435 4456 11484 4481
rect 11499 4456 11529 4472
rect 11398 4442 11428 4450
rect 11435 4448 11545 4456
rect 11398 4434 11443 4442
rect 11130 4416 11149 4418
rect 11164 4416 11210 4418
rect 11130 4400 11210 4416
rect 11237 4414 11272 4427
rect 11313 4424 11350 4427
rect 11313 4422 11355 4424
rect 11242 4411 11272 4414
rect 11251 4407 11258 4411
rect 11258 4406 11259 4407
rect 11217 4400 11227 4406
rect 10976 4392 11011 4400
rect 10976 4366 10977 4392
rect 10984 4366 11011 4392
rect 10919 4348 10949 4362
rect 10976 4358 11011 4366
rect 11013 4392 11054 4400
rect 11013 4366 11028 4392
rect 11035 4366 11054 4392
rect 11118 4388 11149 4400
rect 11164 4388 11267 4400
rect 11279 4390 11305 4416
rect 11320 4411 11350 4422
rect 11382 4418 11444 4434
rect 11382 4416 11428 4418
rect 11382 4400 11444 4416
rect 11456 4400 11462 4448
rect 11465 4440 11545 4448
rect 11465 4438 11484 4440
rect 11499 4438 11533 4440
rect 11465 4422 11545 4438
rect 11465 4400 11484 4422
rect 11499 4406 11529 4422
rect 11557 4416 11563 4490
rect 11566 4416 11585 4560
rect 11600 4416 11606 4560
rect 11615 4490 11628 4560
rect 11680 4556 11702 4560
rect 11673 4534 11702 4548
rect 11755 4534 11771 4548
rect 11809 4544 11815 4546
rect 11822 4544 11930 4560
rect 11937 4544 11943 4546
rect 11951 4544 11966 4560
rect 12032 4554 12051 4557
rect 11673 4532 11771 4534
rect 11798 4532 11966 4544
rect 11981 4534 11997 4548
rect 12032 4535 12054 4554
rect 12064 4548 12080 4549
rect 12063 4546 12080 4548
rect 12064 4541 12080 4546
rect 12054 4534 12060 4535
rect 12063 4534 12092 4541
rect 11981 4533 12092 4534
rect 11981 4532 12098 4533
rect 11657 4524 11708 4532
rect 11755 4524 11789 4532
rect 11657 4512 11682 4524
rect 11689 4512 11708 4524
rect 11762 4522 11789 4524
rect 11798 4522 12019 4532
rect 12054 4529 12060 4532
rect 11762 4518 12019 4522
rect 11657 4504 11708 4512
rect 11755 4504 12019 4518
rect 12063 4524 12098 4532
rect 11609 4456 11628 4490
rect 11673 4496 11702 4504
rect 11673 4490 11690 4496
rect 11673 4488 11707 4490
rect 11755 4488 11771 4504
rect 11772 4494 11980 4504
rect 11981 4494 11997 4504
rect 12045 4500 12060 4515
rect 12063 4512 12064 4524
rect 12071 4512 12098 4524
rect 12063 4504 12098 4512
rect 12063 4503 12092 4504
rect 11783 4490 11997 4494
rect 11798 4488 11997 4490
rect 12032 4490 12045 4500
rect 12063 4490 12080 4503
rect 12032 4488 12080 4490
rect 11674 4484 11707 4488
rect 11670 4482 11707 4484
rect 11670 4481 11737 4482
rect 11670 4476 11701 4481
rect 11707 4476 11737 4481
rect 11670 4472 11737 4476
rect 11643 4469 11737 4472
rect 11643 4462 11692 4469
rect 11643 4456 11673 4462
rect 11692 4457 11697 4462
rect 11609 4440 11689 4456
rect 11701 4448 11737 4469
rect 11798 4464 11987 4488
rect 12032 4487 12079 4488
rect 12045 4482 12079 4487
rect 11813 4461 11987 4464
rect 11806 4458 11987 4461
rect 12015 4481 12079 4482
rect 11609 4438 11628 4440
rect 11643 4438 11677 4440
rect 11609 4422 11689 4438
rect 11609 4416 11628 4422
rect 11325 4390 11428 4400
rect 11279 4388 11428 4390
rect 11449 4388 11484 4400
rect 11118 4386 11280 4388
rect 11130 4366 11149 4386
rect 11164 4384 11194 4386
rect 11013 4358 11054 4366
rect 11136 4362 11149 4366
rect 11201 4370 11280 4386
rect 11312 4386 11484 4388
rect 11312 4370 11391 4386
rect 11398 4384 11428 4386
rect 10976 4348 11005 4358
rect 11019 4348 11048 4358
rect 11063 4348 11093 4362
rect 11136 4348 11179 4362
rect 11201 4358 11391 4370
rect 11456 4366 11462 4386
rect 11186 4348 11216 4358
rect 11217 4348 11375 4358
rect 11379 4348 11409 4358
rect 11413 4348 11443 4362
rect 11471 4348 11484 4386
rect 11556 4400 11585 4416
rect 11599 4400 11628 4416
rect 11643 4406 11673 4422
rect 11701 4400 11707 4448
rect 11710 4442 11729 4448
rect 11744 4442 11774 4450
rect 11710 4434 11774 4442
rect 11710 4418 11790 4434
rect 11806 4427 11868 4458
rect 11884 4427 11946 4458
rect 12015 4456 12064 4481
rect 12079 4456 12109 4472
rect 11978 4442 12008 4450
rect 12015 4448 12125 4456
rect 11978 4434 12023 4442
rect 11710 4416 11729 4418
rect 11744 4416 11790 4418
rect 11710 4400 11790 4416
rect 11817 4414 11852 4427
rect 11893 4424 11930 4427
rect 11893 4422 11935 4424
rect 11822 4411 11852 4414
rect 11831 4407 11838 4411
rect 11838 4406 11839 4407
rect 11797 4400 11807 4406
rect 11556 4392 11591 4400
rect 11556 4366 11557 4392
rect 11564 4366 11591 4392
rect 11499 4348 11529 4362
rect 11556 4358 11591 4366
rect 11593 4392 11634 4400
rect 11593 4366 11608 4392
rect 11615 4366 11634 4392
rect 11698 4388 11729 4400
rect 11744 4388 11847 4400
rect 11859 4390 11885 4416
rect 11900 4411 11930 4422
rect 11962 4418 12024 4434
rect 11962 4416 12008 4418
rect 11962 4400 12024 4416
rect 12036 4400 12042 4448
rect 12045 4440 12125 4448
rect 12045 4438 12064 4440
rect 12079 4438 12113 4440
rect 12045 4422 12125 4438
rect 12045 4400 12064 4422
rect 12079 4406 12109 4422
rect 12137 4416 12143 4490
rect 12146 4416 12165 4560
rect 12180 4416 12186 4560
rect 12195 4490 12208 4560
rect 12260 4556 12282 4560
rect 12253 4534 12282 4548
rect 12335 4534 12351 4548
rect 12389 4544 12395 4546
rect 12402 4544 12510 4560
rect 12517 4544 12523 4546
rect 12531 4544 12546 4560
rect 12612 4554 12631 4557
rect 12253 4532 12351 4534
rect 12378 4532 12546 4544
rect 12561 4534 12577 4548
rect 12612 4535 12634 4554
rect 12644 4548 12660 4549
rect 12643 4546 12660 4548
rect 12644 4541 12660 4546
rect 12634 4534 12640 4535
rect 12643 4534 12672 4541
rect 12561 4533 12672 4534
rect 12561 4532 12678 4533
rect 12237 4524 12288 4532
rect 12335 4524 12369 4532
rect 12237 4512 12262 4524
rect 12269 4512 12288 4524
rect 12342 4522 12369 4524
rect 12378 4522 12599 4532
rect 12634 4529 12640 4532
rect 12342 4518 12599 4522
rect 12237 4504 12288 4512
rect 12335 4504 12599 4518
rect 12643 4524 12678 4532
rect 12189 4456 12208 4490
rect 12253 4496 12282 4504
rect 12253 4490 12270 4496
rect 12253 4488 12287 4490
rect 12335 4488 12351 4504
rect 12352 4494 12560 4504
rect 12561 4494 12577 4504
rect 12625 4500 12640 4515
rect 12643 4512 12644 4524
rect 12651 4512 12678 4524
rect 12643 4504 12678 4512
rect 12643 4503 12672 4504
rect 12363 4490 12577 4494
rect 12378 4488 12577 4490
rect 12612 4490 12625 4500
rect 12643 4490 12660 4503
rect 12612 4488 12660 4490
rect 12254 4484 12287 4488
rect 12250 4482 12287 4484
rect 12250 4481 12317 4482
rect 12250 4476 12281 4481
rect 12287 4476 12317 4481
rect 12250 4472 12317 4476
rect 12223 4469 12317 4472
rect 12223 4462 12272 4469
rect 12223 4456 12253 4462
rect 12272 4457 12277 4462
rect 12189 4440 12269 4456
rect 12281 4448 12317 4469
rect 12378 4464 12567 4488
rect 12612 4487 12659 4488
rect 12625 4482 12659 4487
rect 12393 4461 12567 4464
rect 12386 4458 12567 4461
rect 12595 4481 12659 4482
rect 12189 4438 12208 4440
rect 12223 4438 12257 4440
rect 12189 4422 12269 4438
rect 12189 4416 12208 4422
rect 11905 4390 12008 4400
rect 11859 4388 12008 4390
rect 12029 4388 12064 4400
rect 11698 4386 11860 4388
rect 11710 4366 11729 4386
rect 11744 4384 11774 4386
rect 11593 4358 11634 4366
rect 11716 4362 11729 4366
rect 11781 4370 11860 4386
rect 11892 4386 12064 4388
rect 11892 4370 11971 4386
rect 11978 4384 12008 4386
rect 11556 4348 11585 4358
rect 11599 4348 11628 4358
rect 11643 4348 11673 4362
rect 11716 4348 11759 4362
rect 11781 4358 11971 4370
rect 12036 4366 12042 4386
rect 11766 4348 11796 4358
rect 11797 4348 11955 4358
rect 11959 4348 11989 4358
rect 11993 4348 12023 4362
rect 12051 4348 12064 4386
rect 12136 4400 12165 4416
rect 12179 4400 12208 4416
rect 12223 4406 12253 4422
rect 12281 4400 12287 4448
rect 12290 4442 12309 4448
rect 12324 4442 12354 4450
rect 12290 4434 12354 4442
rect 12290 4418 12370 4434
rect 12386 4427 12448 4458
rect 12464 4427 12526 4458
rect 12595 4456 12644 4481
rect 12659 4456 12689 4472
rect 12558 4442 12588 4450
rect 12595 4448 12705 4456
rect 12558 4434 12603 4442
rect 12290 4416 12309 4418
rect 12324 4416 12370 4418
rect 12290 4400 12370 4416
rect 12397 4414 12432 4427
rect 12473 4424 12510 4427
rect 12473 4422 12515 4424
rect 12402 4411 12432 4414
rect 12411 4407 12418 4411
rect 12418 4406 12419 4407
rect 12377 4400 12387 4406
rect 12136 4392 12171 4400
rect 12136 4366 12137 4392
rect 12144 4366 12171 4392
rect 12079 4348 12109 4362
rect 12136 4358 12171 4366
rect 12173 4392 12214 4400
rect 12173 4366 12188 4392
rect 12195 4366 12214 4392
rect 12278 4388 12309 4400
rect 12324 4388 12427 4400
rect 12439 4390 12465 4416
rect 12480 4411 12510 4422
rect 12542 4418 12604 4434
rect 12542 4416 12588 4418
rect 12542 4400 12604 4416
rect 12616 4400 12622 4448
rect 12625 4440 12705 4448
rect 12625 4438 12644 4440
rect 12659 4438 12693 4440
rect 12625 4422 12705 4438
rect 12625 4400 12644 4422
rect 12659 4406 12689 4422
rect 12717 4416 12723 4490
rect 12726 4416 12745 4560
rect 12760 4416 12766 4560
rect 12775 4490 12788 4560
rect 12840 4556 12862 4560
rect 12833 4534 12862 4548
rect 12915 4534 12931 4548
rect 12969 4544 12975 4546
rect 12982 4544 13090 4560
rect 13097 4544 13103 4546
rect 13111 4544 13126 4560
rect 13192 4554 13211 4557
rect 12833 4532 12931 4534
rect 12958 4532 13126 4544
rect 13141 4534 13157 4548
rect 13192 4535 13214 4554
rect 13224 4548 13240 4549
rect 13223 4546 13240 4548
rect 13224 4541 13240 4546
rect 13214 4534 13220 4535
rect 13223 4534 13252 4541
rect 13141 4533 13252 4534
rect 13141 4532 13258 4533
rect 12817 4524 12868 4532
rect 12915 4524 12949 4532
rect 12817 4512 12842 4524
rect 12849 4512 12868 4524
rect 12922 4522 12949 4524
rect 12958 4522 13179 4532
rect 13214 4529 13220 4532
rect 12922 4518 13179 4522
rect 12817 4504 12868 4512
rect 12915 4504 13179 4518
rect 13223 4524 13258 4532
rect 12769 4456 12788 4490
rect 12833 4496 12862 4504
rect 12833 4490 12850 4496
rect 12833 4488 12867 4490
rect 12915 4488 12931 4504
rect 12932 4494 13140 4504
rect 13141 4494 13157 4504
rect 13205 4500 13220 4515
rect 13223 4512 13224 4524
rect 13231 4512 13258 4524
rect 13223 4504 13258 4512
rect 13223 4503 13252 4504
rect 12943 4490 13157 4494
rect 12958 4488 13157 4490
rect 13192 4490 13205 4500
rect 13223 4490 13240 4503
rect 13192 4488 13240 4490
rect 12834 4484 12867 4488
rect 12830 4482 12867 4484
rect 12830 4481 12897 4482
rect 12830 4476 12861 4481
rect 12867 4476 12897 4481
rect 12830 4472 12897 4476
rect 12803 4469 12897 4472
rect 12803 4462 12852 4469
rect 12803 4456 12833 4462
rect 12852 4457 12857 4462
rect 12769 4440 12849 4456
rect 12861 4448 12897 4469
rect 12958 4464 13147 4488
rect 13192 4487 13239 4488
rect 13205 4482 13239 4487
rect 12973 4461 13147 4464
rect 12966 4458 13147 4461
rect 13175 4481 13239 4482
rect 12769 4438 12788 4440
rect 12803 4438 12837 4440
rect 12769 4422 12849 4438
rect 12769 4416 12788 4422
rect 12485 4390 12588 4400
rect 12439 4388 12588 4390
rect 12609 4388 12644 4400
rect 12278 4386 12440 4388
rect 12290 4366 12309 4386
rect 12324 4384 12354 4386
rect 12173 4358 12214 4366
rect 12296 4362 12309 4366
rect 12361 4370 12440 4386
rect 12472 4386 12644 4388
rect 12472 4370 12551 4386
rect 12558 4384 12588 4386
rect 12136 4348 12165 4358
rect 12179 4348 12208 4358
rect 12223 4348 12253 4362
rect 12296 4348 12339 4362
rect 12361 4358 12551 4370
rect 12616 4366 12622 4386
rect 12346 4348 12376 4358
rect 12377 4348 12535 4358
rect 12539 4348 12569 4358
rect 12573 4348 12603 4362
rect 12631 4348 12644 4386
rect 12716 4400 12745 4416
rect 12759 4400 12788 4416
rect 12803 4406 12833 4422
rect 12861 4400 12867 4448
rect 12870 4442 12889 4448
rect 12904 4442 12934 4450
rect 12870 4434 12934 4442
rect 12870 4418 12950 4434
rect 12966 4427 13028 4458
rect 13044 4427 13106 4458
rect 13175 4456 13224 4481
rect 13239 4456 13269 4472
rect 13138 4442 13168 4450
rect 13175 4448 13285 4456
rect 13138 4434 13183 4442
rect 12870 4416 12889 4418
rect 12904 4416 12950 4418
rect 12870 4400 12950 4416
rect 12977 4414 13012 4427
rect 13053 4424 13090 4427
rect 13053 4422 13095 4424
rect 12982 4411 13012 4414
rect 12991 4407 12998 4411
rect 12998 4406 12999 4407
rect 12957 4400 12967 4406
rect 12716 4392 12751 4400
rect 12716 4366 12717 4392
rect 12724 4366 12751 4392
rect 12659 4348 12689 4362
rect 12716 4358 12751 4366
rect 12753 4392 12794 4400
rect 12753 4366 12768 4392
rect 12775 4366 12794 4392
rect 12858 4388 12889 4400
rect 12904 4388 13007 4400
rect 13019 4390 13045 4416
rect 13060 4411 13090 4422
rect 13122 4418 13184 4434
rect 13122 4416 13168 4418
rect 13122 4400 13184 4416
rect 13196 4400 13202 4448
rect 13205 4440 13285 4448
rect 13205 4438 13224 4440
rect 13239 4438 13273 4440
rect 13205 4422 13285 4438
rect 13205 4400 13224 4422
rect 13239 4406 13269 4422
rect 13297 4416 13303 4490
rect 13306 4416 13325 4560
rect 13340 4416 13346 4560
rect 13355 4490 13368 4560
rect 13420 4556 13442 4560
rect 13413 4534 13442 4548
rect 13495 4534 13511 4548
rect 13549 4544 13555 4546
rect 13562 4544 13670 4560
rect 13677 4544 13683 4546
rect 13691 4544 13706 4560
rect 13772 4554 13791 4557
rect 13413 4532 13511 4534
rect 13538 4532 13706 4544
rect 13721 4534 13737 4548
rect 13772 4535 13794 4554
rect 13804 4548 13820 4549
rect 13803 4546 13820 4548
rect 13804 4541 13820 4546
rect 13794 4534 13800 4535
rect 13803 4534 13832 4541
rect 13721 4533 13832 4534
rect 13721 4532 13838 4533
rect 13397 4524 13448 4532
rect 13495 4524 13529 4532
rect 13397 4512 13422 4524
rect 13429 4512 13448 4524
rect 13502 4522 13529 4524
rect 13538 4522 13759 4532
rect 13794 4529 13800 4532
rect 13502 4518 13759 4522
rect 13397 4504 13448 4512
rect 13495 4504 13759 4518
rect 13803 4524 13838 4532
rect 13349 4456 13368 4490
rect 13413 4496 13442 4504
rect 13413 4490 13430 4496
rect 13413 4488 13447 4490
rect 13495 4488 13511 4504
rect 13512 4494 13720 4504
rect 13721 4494 13737 4504
rect 13785 4500 13800 4515
rect 13803 4512 13804 4524
rect 13811 4512 13838 4524
rect 13803 4504 13838 4512
rect 13803 4503 13832 4504
rect 13523 4490 13737 4494
rect 13538 4488 13737 4490
rect 13772 4490 13785 4500
rect 13803 4490 13820 4503
rect 13772 4488 13820 4490
rect 13414 4484 13447 4488
rect 13410 4482 13447 4484
rect 13410 4481 13477 4482
rect 13410 4476 13441 4481
rect 13447 4476 13477 4481
rect 13410 4472 13477 4476
rect 13383 4469 13477 4472
rect 13383 4462 13432 4469
rect 13383 4456 13413 4462
rect 13432 4457 13437 4462
rect 13349 4440 13429 4456
rect 13441 4448 13477 4469
rect 13538 4464 13727 4488
rect 13772 4487 13819 4488
rect 13785 4482 13819 4487
rect 13553 4461 13727 4464
rect 13546 4458 13727 4461
rect 13755 4481 13819 4482
rect 13349 4438 13368 4440
rect 13383 4438 13417 4440
rect 13349 4422 13429 4438
rect 13349 4416 13368 4422
rect 13065 4390 13168 4400
rect 13019 4388 13168 4390
rect 13189 4388 13224 4400
rect 12858 4386 13020 4388
rect 12870 4366 12889 4386
rect 12904 4384 12934 4386
rect 12753 4358 12794 4366
rect 12876 4362 12889 4366
rect 12941 4370 13020 4386
rect 13052 4386 13224 4388
rect 13052 4370 13131 4386
rect 13138 4384 13168 4386
rect 12716 4348 12745 4358
rect 12759 4348 12788 4358
rect 12803 4348 12833 4362
rect 12876 4348 12919 4362
rect 12941 4358 13131 4370
rect 13196 4366 13202 4386
rect 12926 4348 12956 4358
rect 12957 4348 13115 4358
rect 13119 4348 13149 4358
rect 13153 4348 13183 4362
rect 13211 4348 13224 4386
rect 13296 4400 13325 4416
rect 13339 4400 13368 4416
rect 13383 4406 13413 4422
rect 13441 4400 13447 4448
rect 13450 4442 13469 4448
rect 13484 4442 13514 4450
rect 13450 4434 13514 4442
rect 13450 4418 13530 4434
rect 13546 4427 13608 4458
rect 13624 4427 13686 4458
rect 13755 4456 13804 4481
rect 13819 4456 13849 4472
rect 13718 4442 13748 4450
rect 13755 4448 13865 4456
rect 13718 4434 13763 4442
rect 13450 4416 13469 4418
rect 13484 4416 13530 4418
rect 13450 4400 13530 4416
rect 13557 4414 13592 4427
rect 13633 4424 13670 4427
rect 13633 4422 13675 4424
rect 13562 4411 13592 4414
rect 13571 4407 13578 4411
rect 13578 4406 13579 4407
rect 13537 4400 13547 4406
rect 13296 4392 13331 4400
rect 13296 4366 13297 4392
rect 13304 4366 13331 4392
rect 13239 4348 13269 4362
rect 13296 4358 13331 4366
rect 13333 4392 13374 4400
rect 13333 4366 13348 4392
rect 13355 4366 13374 4392
rect 13438 4388 13469 4400
rect 13484 4388 13587 4400
rect 13599 4390 13625 4416
rect 13640 4411 13670 4422
rect 13702 4418 13764 4434
rect 13702 4416 13748 4418
rect 13702 4400 13764 4416
rect 13776 4400 13782 4448
rect 13785 4440 13865 4448
rect 13785 4438 13804 4440
rect 13819 4438 13853 4440
rect 13785 4422 13865 4438
rect 13785 4400 13804 4422
rect 13819 4406 13849 4422
rect 13877 4416 13883 4490
rect 13886 4416 13905 4560
rect 13920 4416 13926 4560
rect 13935 4490 13948 4560
rect 14000 4556 14022 4560
rect 13993 4534 14022 4548
rect 14075 4534 14091 4548
rect 14129 4544 14135 4546
rect 14142 4544 14250 4560
rect 14257 4544 14263 4546
rect 14271 4544 14286 4560
rect 14352 4554 14371 4557
rect 13993 4532 14091 4534
rect 14118 4532 14286 4544
rect 14301 4534 14317 4548
rect 14352 4535 14374 4554
rect 14384 4548 14400 4549
rect 14383 4546 14400 4548
rect 14384 4541 14400 4546
rect 14374 4534 14380 4535
rect 14383 4534 14412 4541
rect 14301 4533 14412 4534
rect 14301 4532 14418 4533
rect 13977 4524 14028 4532
rect 14075 4524 14109 4532
rect 13977 4512 14002 4524
rect 14009 4512 14028 4524
rect 14082 4522 14109 4524
rect 14118 4522 14339 4532
rect 14374 4529 14380 4532
rect 14082 4518 14339 4522
rect 13977 4504 14028 4512
rect 14075 4504 14339 4518
rect 14383 4524 14418 4532
rect 13929 4456 13948 4490
rect 13993 4496 14022 4504
rect 13993 4490 14010 4496
rect 13993 4488 14027 4490
rect 14075 4488 14091 4504
rect 14092 4494 14300 4504
rect 14301 4494 14317 4504
rect 14365 4500 14380 4515
rect 14383 4512 14384 4524
rect 14391 4512 14418 4524
rect 14383 4504 14418 4512
rect 14383 4503 14412 4504
rect 14103 4490 14317 4494
rect 14118 4488 14317 4490
rect 14352 4490 14365 4500
rect 14383 4490 14400 4503
rect 14352 4488 14400 4490
rect 13994 4484 14027 4488
rect 13990 4482 14027 4484
rect 13990 4481 14057 4482
rect 13990 4476 14021 4481
rect 14027 4476 14057 4481
rect 13990 4472 14057 4476
rect 13963 4469 14057 4472
rect 13963 4462 14012 4469
rect 13963 4456 13993 4462
rect 14012 4457 14017 4462
rect 13929 4440 14009 4456
rect 14021 4448 14057 4469
rect 14118 4464 14307 4488
rect 14352 4487 14399 4488
rect 14365 4482 14399 4487
rect 14133 4461 14307 4464
rect 14126 4458 14307 4461
rect 14335 4481 14399 4482
rect 13929 4438 13948 4440
rect 13963 4438 13997 4440
rect 13929 4422 14009 4438
rect 13929 4416 13948 4422
rect 13645 4390 13748 4400
rect 13599 4388 13748 4390
rect 13769 4388 13804 4400
rect 13438 4386 13600 4388
rect 13450 4366 13469 4386
rect 13484 4384 13514 4386
rect 13333 4358 13374 4366
rect 13456 4362 13469 4366
rect 13521 4370 13600 4386
rect 13632 4386 13804 4388
rect 13632 4370 13711 4386
rect 13718 4384 13748 4386
rect 13296 4348 13325 4358
rect 13339 4348 13368 4358
rect 13383 4348 13413 4362
rect 13456 4348 13499 4362
rect 13521 4358 13711 4370
rect 13776 4366 13782 4386
rect 13506 4348 13536 4358
rect 13537 4348 13695 4358
rect 13699 4348 13729 4358
rect 13733 4348 13763 4362
rect 13791 4348 13804 4386
rect 13876 4400 13905 4416
rect 13919 4400 13948 4416
rect 13963 4406 13993 4422
rect 14021 4400 14027 4448
rect 14030 4442 14049 4448
rect 14064 4442 14094 4450
rect 14030 4434 14094 4442
rect 14030 4418 14110 4434
rect 14126 4427 14188 4458
rect 14204 4427 14266 4458
rect 14335 4456 14384 4481
rect 14399 4456 14429 4472
rect 14298 4442 14328 4450
rect 14335 4448 14445 4456
rect 14298 4434 14343 4442
rect 14030 4416 14049 4418
rect 14064 4416 14110 4418
rect 14030 4400 14110 4416
rect 14137 4414 14172 4427
rect 14213 4424 14250 4427
rect 14213 4422 14255 4424
rect 14142 4411 14172 4414
rect 14151 4407 14158 4411
rect 14158 4406 14159 4407
rect 14117 4400 14127 4406
rect 13876 4392 13911 4400
rect 13876 4366 13877 4392
rect 13884 4366 13911 4392
rect 13819 4348 13849 4362
rect 13876 4358 13911 4366
rect 13913 4392 13954 4400
rect 13913 4366 13928 4392
rect 13935 4366 13954 4392
rect 14018 4388 14049 4400
rect 14064 4388 14167 4400
rect 14179 4390 14205 4416
rect 14220 4411 14250 4422
rect 14282 4418 14344 4434
rect 14282 4416 14328 4418
rect 14282 4400 14344 4416
rect 14356 4400 14362 4448
rect 14365 4440 14445 4448
rect 14365 4438 14384 4440
rect 14399 4438 14433 4440
rect 14365 4422 14445 4438
rect 14365 4400 14384 4422
rect 14399 4406 14429 4422
rect 14457 4416 14463 4490
rect 14466 4416 14485 4560
rect 14500 4416 14506 4560
rect 14515 4490 14528 4560
rect 14580 4556 14602 4560
rect 14573 4534 14602 4548
rect 14655 4534 14671 4548
rect 14709 4544 14715 4546
rect 14722 4544 14830 4560
rect 14837 4544 14843 4546
rect 14851 4544 14866 4560
rect 14932 4554 14951 4557
rect 14573 4532 14671 4534
rect 14698 4532 14866 4544
rect 14881 4534 14897 4548
rect 14932 4535 14954 4554
rect 14964 4548 14980 4549
rect 14963 4546 14980 4548
rect 14964 4541 14980 4546
rect 14954 4534 14960 4535
rect 14963 4534 14992 4541
rect 14881 4533 14992 4534
rect 14881 4532 14998 4533
rect 14557 4524 14608 4532
rect 14655 4524 14689 4532
rect 14557 4512 14582 4524
rect 14589 4512 14608 4524
rect 14662 4522 14689 4524
rect 14698 4522 14919 4532
rect 14954 4529 14960 4532
rect 14662 4518 14919 4522
rect 14557 4504 14608 4512
rect 14655 4504 14919 4518
rect 14963 4524 14998 4532
rect 14509 4456 14528 4490
rect 14573 4496 14602 4504
rect 14573 4490 14590 4496
rect 14573 4488 14607 4490
rect 14655 4488 14671 4504
rect 14672 4494 14880 4504
rect 14881 4494 14897 4504
rect 14945 4500 14960 4515
rect 14963 4512 14964 4524
rect 14971 4512 14998 4524
rect 14963 4504 14998 4512
rect 14963 4503 14992 4504
rect 14683 4490 14897 4494
rect 14698 4488 14897 4490
rect 14932 4490 14945 4500
rect 14963 4490 14980 4503
rect 14932 4488 14980 4490
rect 14574 4484 14607 4488
rect 14570 4482 14607 4484
rect 14570 4481 14637 4482
rect 14570 4476 14601 4481
rect 14607 4476 14637 4481
rect 14570 4472 14637 4476
rect 14543 4469 14637 4472
rect 14543 4462 14592 4469
rect 14543 4456 14573 4462
rect 14592 4457 14597 4462
rect 14509 4440 14589 4456
rect 14601 4448 14637 4469
rect 14698 4464 14887 4488
rect 14932 4487 14979 4488
rect 14945 4482 14979 4487
rect 14713 4461 14887 4464
rect 14706 4458 14887 4461
rect 14915 4481 14979 4482
rect 14509 4438 14528 4440
rect 14543 4438 14577 4440
rect 14509 4422 14589 4438
rect 14509 4416 14528 4422
rect 14225 4390 14328 4400
rect 14179 4388 14328 4390
rect 14349 4388 14384 4400
rect 14018 4386 14180 4388
rect 14030 4366 14049 4386
rect 14064 4384 14094 4386
rect 13913 4358 13954 4366
rect 14036 4362 14049 4366
rect 14101 4370 14180 4386
rect 14212 4386 14384 4388
rect 14212 4370 14291 4386
rect 14298 4384 14328 4386
rect 13876 4348 13905 4358
rect 13919 4348 13948 4358
rect 13963 4348 13993 4362
rect 14036 4348 14079 4362
rect 14101 4358 14291 4370
rect 14356 4366 14362 4386
rect 14086 4348 14116 4358
rect 14117 4348 14275 4358
rect 14279 4348 14309 4358
rect 14313 4348 14343 4362
rect 14371 4348 14384 4386
rect 14456 4400 14485 4416
rect 14499 4400 14528 4416
rect 14543 4406 14573 4422
rect 14601 4400 14607 4448
rect 14610 4442 14629 4448
rect 14644 4442 14674 4450
rect 14610 4434 14674 4442
rect 14610 4418 14690 4434
rect 14706 4427 14768 4458
rect 14784 4427 14846 4458
rect 14915 4456 14964 4481
rect 14979 4456 15009 4472
rect 14878 4442 14908 4450
rect 14915 4448 15025 4456
rect 14878 4434 14923 4442
rect 14610 4416 14629 4418
rect 14644 4416 14690 4418
rect 14610 4400 14690 4416
rect 14717 4414 14752 4427
rect 14793 4424 14830 4427
rect 14793 4422 14835 4424
rect 14722 4411 14752 4414
rect 14731 4407 14738 4411
rect 14738 4406 14739 4407
rect 14697 4400 14707 4406
rect 14456 4392 14491 4400
rect 14456 4366 14457 4392
rect 14464 4366 14491 4392
rect 14399 4348 14429 4362
rect 14456 4358 14491 4366
rect 14493 4392 14534 4400
rect 14493 4366 14508 4392
rect 14515 4366 14534 4392
rect 14598 4388 14629 4400
rect 14644 4388 14747 4400
rect 14759 4390 14785 4416
rect 14800 4411 14830 4422
rect 14862 4418 14924 4434
rect 14862 4416 14908 4418
rect 14862 4400 14924 4416
rect 14936 4400 14942 4448
rect 14945 4440 15025 4448
rect 14945 4438 14964 4440
rect 14979 4438 15013 4440
rect 14945 4422 15025 4438
rect 14945 4400 14964 4422
rect 14979 4406 15009 4422
rect 15037 4416 15043 4490
rect 15046 4416 15065 4560
rect 15080 4416 15086 4560
rect 15095 4490 15108 4560
rect 15160 4556 15182 4560
rect 15153 4534 15182 4548
rect 15235 4534 15251 4548
rect 15289 4544 15295 4546
rect 15302 4544 15410 4560
rect 15417 4544 15423 4546
rect 15431 4544 15446 4560
rect 15512 4554 15531 4557
rect 15153 4532 15251 4534
rect 15278 4532 15446 4544
rect 15461 4534 15477 4548
rect 15512 4535 15534 4554
rect 15544 4548 15560 4549
rect 15543 4546 15560 4548
rect 15544 4541 15560 4546
rect 15534 4534 15540 4535
rect 15543 4534 15572 4541
rect 15461 4533 15572 4534
rect 15461 4532 15578 4533
rect 15137 4524 15188 4532
rect 15235 4524 15269 4532
rect 15137 4512 15162 4524
rect 15169 4512 15188 4524
rect 15242 4522 15269 4524
rect 15278 4522 15499 4532
rect 15534 4529 15540 4532
rect 15242 4518 15499 4522
rect 15137 4504 15188 4512
rect 15235 4504 15499 4518
rect 15543 4524 15578 4532
rect 15089 4456 15108 4490
rect 15153 4496 15182 4504
rect 15153 4490 15170 4496
rect 15153 4488 15187 4490
rect 15235 4488 15251 4504
rect 15252 4494 15460 4504
rect 15461 4494 15477 4504
rect 15525 4500 15540 4515
rect 15543 4512 15544 4524
rect 15551 4512 15578 4524
rect 15543 4504 15578 4512
rect 15543 4503 15572 4504
rect 15263 4490 15477 4494
rect 15278 4488 15477 4490
rect 15512 4490 15525 4500
rect 15543 4490 15560 4503
rect 15512 4488 15560 4490
rect 15154 4484 15187 4488
rect 15150 4482 15187 4484
rect 15150 4481 15217 4482
rect 15150 4476 15181 4481
rect 15187 4476 15217 4481
rect 15150 4472 15217 4476
rect 15123 4469 15217 4472
rect 15123 4462 15172 4469
rect 15123 4456 15153 4462
rect 15172 4457 15177 4462
rect 15089 4440 15169 4456
rect 15181 4448 15217 4469
rect 15278 4464 15467 4488
rect 15512 4487 15559 4488
rect 15525 4482 15559 4487
rect 15293 4461 15467 4464
rect 15286 4458 15467 4461
rect 15495 4481 15559 4482
rect 15089 4438 15108 4440
rect 15123 4438 15157 4440
rect 15089 4422 15169 4438
rect 15089 4416 15108 4422
rect 14805 4390 14908 4400
rect 14759 4388 14908 4390
rect 14929 4388 14964 4400
rect 14598 4386 14760 4388
rect 14610 4366 14629 4386
rect 14644 4384 14674 4386
rect 14493 4358 14534 4366
rect 14616 4362 14629 4366
rect 14681 4370 14760 4386
rect 14792 4386 14964 4388
rect 14792 4370 14871 4386
rect 14878 4384 14908 4386
rect 14456 4348 14485 4358
rect 14499 4348 14528 4358
rect 14543 4348 14573 4362
rect 14616 4348 14659 4362
rect 14681 4358 14871 4370
rect 14936 4366 14942 4386
rect 14666 4348 14696 4358
rect 14697 4348 14855 4358
rect 14859 4348 14889 4358
rect 14893 4348 14923 4362
rect 14951 4348 14964 4386
rect 15036 4400 15065 4416
rect 15079 4400 15108 4416
rect 15123 4406 15153 4422
rect 15181 4400 15187 4448
rect 15190 4442 15209 4448
rect 15224 4442 15254 4450
rect 15190 4434 15254 4442
rect 15190 4418 15270 4434
rect 15286 4427 15348 4458
rect 15364 4427 15426 4458
rect 15495 4456 15544 4481
rect 15559 4456 15589 4472
rect 15458 4442 15488 4450
rect 15495 4448 15605 4456
rect 15458 4434 15503 4442
rect 15190 4416 15209 4418
rect 15224 4416 15270 4418
rect 15190 4400 15270 4416
rect 15297 4414 15332 4427
rect 15373 4424 15410 4427
rect 15373 4422 15415 4424
rect 15302 4411 15332 4414
rect 15311 4407 15318 4411
rect 15318 4406 15319 4407
rect 15277 4400 15287 4406
rect 15036 4392 15071 4400
rect 15036 4366 15037 4392
rect 15044 4366 15071 4392
rect 14979 4348 15009 4362
rect 15036 4358 15071 4366
rect 15073 4392 15114 4400
rect 15073 4366 15088 4392
rect 15095 4366 15114 4392
rect 15178 4388 15209 4400
rect 15224 4388 15327 4400
rect 15339 4390 15365 4416
rect 15380 4411 15410 4422
rect 15442 4418 15504 4434
rect 15442 4416 15488 4418
rect 15442 4400 15504 4416
rect 15516 4400 15522 4448
rect 15525 4440 15605 4448
rect 15525 4438 15544 4440
rect 15559 4438 15593 4440
rect 15525 4422 15605 4438
rect 15525 4400 15544 4422
rect 15559 4406 15589 4422
rect 15617 4416 15623 4490
rect 15626 4416 15645 4560
rect 15660 4416 15666 4560
rect 15675 4490 15688 4560
rect 15740 4556 15762 4560
rect 15733 4534 15762 4548
rect 15815 4534 15831 4548
rect 15869 4544 15875 4546
rect 15882 4544 15990 4560
rect 15997 4544 16003 4546
rect 16011 4544 16026 4560
rect 16092 4554 16111 4557
rect 15733 4532 15831 4534
rect 15858 4532 16026 4544
rect 16041 4534 16057 4548
rect 16092 4535 16114 4554
rect 16124 4548 16140 4549
rect 16123 4546 16140 4548
rect 16124 4541 16140 4546
rect 16114 4534 16120 4535
rect 16123 4534 16152 4541
rect 16041 4533 16152 4534
rect 16041 4532 16158 4533
rect 15717 4524 15768 4532
rect 15815 4524 15849 4532
rect 15717 4512 15742 4524
rect 15749 4512 15768 4524
rect 15822 4522 15849 4524
rect 15858 4522 16079 4532
rect 16114 4529 16120 4532
rect 15822 4518 16079 4522
rect 15717 4504 15768 4512
rect 15815 4504 16079 4518
rect 16123 4524 16158 4532
rect 15669 4456 15688 4490
rect 15733 4496 15762 4504
rect 15733 4490 15750 4496
rect 15733 4488 15767 4490
rect 15815 4488 15831 4504
rect 15832 4494 16040 4504
rect 16041 4494 16057 4504
rect 16105 4500 16120 4515
rect 16123 4512 16124 4524
rect 16131 4512 16158 4524
rect 16123 4504 16158 4512
rect 16123 4503 16152 4504
rect 15843 4490 16057 4494
rect 15858 4488 16057 4490
rect 16092 4490 16105 4500
rect 16123 4490 16140 4503
rect 16092 4488 16140 4490
rect 15734 4484 15767 4488
rect 15730 4482 15767 4484
rect 15730 4481 15797 4482
rect 15730 4476 15761 4481
rect 15767 4476 15797 4481
rect 15730 4472 15797 4476
rect 15703 4469 15797 4472
rect 15703 4462 15752 4469
rect 15703 4456 15733 4462
rect 15752 4457 15757 4462
rect 15669 4440 15749 4456
rect 15761 4448 15797 4469
rect 15858 4464 16047 4488
rect 16092 4487 16139 4488
rect 16105 4482 16139 4487
rect 15873 4461 16047 4464
rect 15866 4458 16047 4461
rect 16075 4481 16139 4482
rect 15669 4438 15688 4440
rect 15703 4438 15737 4440
rect 15669 4422 15749 4438
rect 15669 4416 15688 4422
rect 15385 4390 15488 4400
rect 15339 4388 15488 4390
rect 15509 4388 15544 4400
rect 15178 4386 15340 4388
rect 15190 4366 15209 4386
rect 15224 4384 15254 4386
rect 15073 4358 15114 4366
rect 15196 4362 15209 4366
rect 15261 4370 15340 4386
rect 15372 4386 15544 4388
rect 15372 4370 15451 4386
rect 15458 4384 15488 4386
rect 15036 4348 15065 4358
rect 15079 4348 15108 4358
rect 15123 4348 15153 4362
rect 15196 4348 15239 4362
rect 15261 4358 15451 4370
rect 15516 4366 15522 4386
rect 15246 4348 15276 4358
rect 15277 4348 15435 4358
rect 15439 4348 15469 4358
rect 15473 4348 15503 4362
rect 15531 4348 15544 4386
rect 15616 4400 15645 4416
rect 15659 4400 15688 4416
rect 15703 4406 15733 4422
rect 15761 4400 15767 4448
rect 15770 4442 15789 4448
rect 15804 4442 15834 4450
rect 15770 4434 15834 4442
rect 15770 4418 15850 4434
rect 15866 4427 15928 4458
rect 15944 4427 16006 4458
rect 16075 4456 16124 4481
rect 16139 4456 16169 4472
rect 16038 4442 16068 4450
rect 16075 4448 16185 4456
rect 16038 4434 16083 4442
rect 15770 4416 15789 4418
rect 15804 4416 15850 4418
rect 15770 4400 15850 4416
rect 15877 4414 15912 4427
rect 15953 4424 15990 4427
rect 15953 4422 15995 4424
rect 15882 4411 15912 4414
rect 15891 4407 15898 4411
rect 15898 4406 15899 4407
rect 15857 4400 15867 4406
rect 15616 4392 15651 4400
rect 15616 4366 15617 4392
rect 15624 4366 15651 4392
rect 15559 4348 15589 4362
rect 15616 4358 15651 4366
rect 15653 4392 15694 4400
rect 15653 4366 15668 4392
rect 15675 4366 15694 4392
rect 15758 4388 15789 4400
rect 15804 4388 15907 4400
rect 15919 4390 15945 4416
rect 15960 4411 15990 4422
rect 16022 4418 16084 4434
rect 16022 4416 16068 4418
rect 16022 4400 16084 4416
rect 16096 4400 16102 4448
rect 16105 4440 16185 4448
rect 16105 4438 16124 4440
rect 16139 4438 16173 4440
rect 16105 4422 16185 4438
rect 16105 4400 16124 4422
rect 16139 4406 16169 4422
rect 16197 4416 16203 4490
rect 16206 4416 16225 4560
rect 16240 4416 16246 4560
rect 16255 4490 16268 4560
rect 16320 4556 16342 4560
rect 16313 4534 16342 4548
rect 16395 4534 16411 4548
rect 16449 4544 16455 4546
rect 16462 4544 16570 4560
rect 16577 4544 16583 4546
rect 16591 4544 16606 4560
rect 16672 4554 16691 4557
rect 16313 4532 16411 4534
rect 16438 4532 16606 4544
rect 16621 4534 16637 4548
rect 16672 4535 16694 4554
rect 16704 4548 16720 4549
rect 16703 4546 16720 4548
rect 16704 4541 16720 4546
rect 16694 4534 16700 4535
rect 16703 4534 16732 4541
rect 16621 4533 16732 4534
rect 16621 4532 16738 4533
rect 16297 4524 16348 4532
rect 16395 4524 16429 4532
rect 16297 4512 16322 4524
rect 16329 4512 16348 4524
rect 16402 4522 16429 4524
rect 16438 4522 16659 4532
rect 16694 4529 16700 4532
rect 16402 4518 16659 4522
rect 16297 4504 16348 4512
rect 16395 4504 16659 4518
rect 16703 4524 16738 4532
rect 16249 4456 16268 4490
rect 16313 4496 16342 4504
rect 16313 4490 16330 4496
rect 16313 4488 16347 4490
rect 16395 4488 16411 4504
rect 16412 4494 16620 4504
rect 16621 4494 16637 4504
rect 16685 4500 16700 4515
rect 16703 4512 16704 4524
rect 16711 4512 16738 4524
rect 16703 4504 16738 4512
rect 16703 4503 16732 4504
rect 16423 4490 16637 4494
rect 16438 4488 16637 4490
rect 16672 4490 16685 4500
rect 16703 4490 16720 4503
rect 16672 4488 16720 4490
rect 16314 4484 16347 4488
rect 16310 4482 16347 4484
rect 16310 4481 16377 4482
rect 16310 4476 16341 4481
rect 16347 4476 16377 4481
rect 16310 4472 16377 4476
rect 16283 4469 16377 4472
rect 16283 4462 16332 4469
rect 16283 4456 16313 4462
rect 16332 4457 16337 4462
rect 16249 4440 16329 4456
rect 16341 4448 16377 4469
rect 16438 4464 16627 4488
rect 16672 4487 16719 4488
rect 16685 4482 16719 4487
rect 16453 4461 16627 4464
rect 16446 4458 16627 4461
rect 16655 4481 16719 4482
rect 16249 4438 16268 4440
rect 16283 4438 16317 4440
rect 16249 4422 16329 4438
rect 16249 4416 16268 4422
rect 15965 4390 16068 4400
rect 15919 4388 16068 4390
rect 16089 4388 16124 4400
rect 15758 4386 15920 4388
rect 15770 4366 15789 4386
rect 15804 4384 15834 4386
rect 15653 4358 15694 4366
rect 15776 4362 15789 4366
rect 15841 4370 15920 4386
rect 15952 4386 16124 4388
rect 15952 4370 16031 4386
rect 16038 4384 16068 4386
rect 15616 4348 15645 4358
rect 15659 4348 15688 4358
rect 15703 4348 15733 4362
rect 15776 4348 15819 4362
rect 15841 4358 16031 4370
rect 16096 4366 16102 4386
rect 15826 4348 15856 4358
rect 15857 4348 16015 4358
rect 16019 4348 16049 4358
rect 16053 4348 16083 4362
rect 16111 4348 16124 4386
rect 16196 4400 16225 4416
rect 16239 4400 16268 4416
rect 16283 4406 16313 4422
rect 16341 4400 16347 4448
rect 16350 4442 16369 4448
rect 16384 4442 16414 4450
rect 16350 4434 16414 4442
rect 16350 4418 16430 4434
rect 16446 4427 16508 4458
rect 16524 4427 16586 4458
rect 16655 4456 16704 4481
rect 16719 4456 16749 4472
rect 16618 4442 16648 4450
rect 16655 4448 16765 4456
rect 16618 4434 16663 4442
rect 16350 4416 16369 4418
rect 16384 4416 16430 4418
rect 16350 4400 16430 4416
rect 16457 4414 16492 4427
rect 16533 4424 16570 4427
rect 16533 4422 16575 4424
rect 16462 4411 16492 4414
rect 16471 4407 16478 4411
rect 16478 4406 16479 4407
rect 16437 4400 16447 4406
rect 16196 4392 16231 4400
rect 16196 4366 16197 4392
rect 16204 4366 16231 4392
rect 16139 4348 16169 4362
rect 16196 4358 16231 4366
rect 16233 4392 16274 4400
rect 16233 4366 16248 4392
rect 16255 4366 16274 4392
rect 16338 4388 16369 4400
rect 16384 4388 16487 4400
rect 16499 4390 16525 4416
rect 16540 4411 16570 4422
rect 16602 4418 16664 4434
rect 16602 4416 16648 4418
rect 16602 4400 16664 4416
rect 16676 4400 16682 4448
rect 16685 4440 16765 4448
rect 16685 4438 16704 4440
rect 16719 4438 16753 4440
rect 16685 4422 16765 4438
rect 16685 4400 16704 4422
rect 16719 4406 16749 4422
rect 16777 4416 16783 4490
rect 16786 4416 16805 4560
rect 16820 4416 16826 4560
rect 16835 4490 16848 4560
rect 16900 4556 16922 4560
rect 16893 4534 16922 4548
rect 16975 4534 16991 4548
rect 17029 4544 17035 4546
rect 17042 4544 17150 4560
rect 17157 4544 17163 4546
rect 17171 4544 17186 4560
rect 17252 4554 17271 4557
rect 16893 4532 16991 4534
rect 17018 4532 17186 4544
rect 17201 4534 17217 4548
rect 17252 4535 17274 4554
rect 17284 4548 17300 4549
rect 17283 4546 17300 4548
rect 17284 4541 17300 4546
rect 17274 4534 17280 4535
rect 17283 4534 17312 4541
rect 17201 4533 17312 4534
rect 17201 4532 17318 4533
rect 16877 4524 16928 4532
rect 16975 4524 17009 4532
rect 16877 4512 16902 4524
rect 16909 4512 16928 4524
rect 16982 4522 17009 4524
rect 17018 4522 17239 4532
rect 17274 4529 17280 4532
rect 16982 4518 17239 4522
rect 16877 4504 16928 4512
rect 16975 4504 17239 4518
rect 17283 4524 17318 4532
rect 16829 4456 16848 4490
rect 16893 4496 16922 4504
rect 16893 4490 16910 4496
rect 16893 4488 16927 4490
rect 16975 4488 16991 4504
rect 16992 4494 17200 4504
rect 17201 4494 17217 4504
rect 17265 4500 17280 4515
rect 17283 4512 17284 4524
rect 17291 4512 17318 4524
rect 17283 4504 17318 4512
rect 17283 4503 17312 4504
rect 17003 4490 17217 4494
rect 17018 4488 17217 4490
rect 17252 4490 17265 4500
rect 17283 4490 17300 4503
rect 17252 4488 17300 4490
rect 16894 4484 16927 4488
rect 16890 4482 16927 4484
rect 16890 4481 16957 4482
rect 16890 4476 16921 4481
rect 16927 4476 16957 4481
rect 16890 4472 16957 4476
rect 16863 4469 16957 4472
rect 16863 4462 16912 4469
rect 16863 4456 16893 4462
rect 16912 4457 16917 4462
rect 16829 4440 16909 4456
rect 16921 4448 16957 4469
rect 17018 4464 17207 4488
rect 17252 4487 17299 4488
rect 17265 4482 17299 4487
rect 17033 4461 17207 4464
rect 17026 4458 17207 4461
rect 17235 4481 17299 4482
rect 16829 4438 16848 4440
rect 16863 4438 16897 4440
rect 16829 4422 16909 4438
rect 16829 4416 16848 4422
rect 16545 4390 16648 4400
rect 16499 4388 16648 4390
rect 16669 4388 16704 4400
rect 16338 4386 16500 4388
rect 16350 4366 16369 4386
rect 16384 4384 16414 4386
rect 16233 4358 16274 4366
rect 16356 4362 16369 4366
rect 16421 4370 16500 4386
rect 16532 4386 16704 4388
rect 16532 4370 16611 4386
rect 16618 4384 16648 4386
rect 16196 4348 16225 4358
rect 16239 4348 16268 4358
rect 16283 4348 16313 4362
rect 16356 4348 16399 4362
rect 16421 4358 16611 4370
rect 16676 4366 16682 4386
rect 16406 4348 16436 4358
rect 16437 4348 16595 4358
rect 16599 4348 16629 4358
rect 16633 4348 16663 4362
rect 16691 4348 16704 4386
rect 16776 4400 16805 4416
rect 16819 4400 16848 4416
rect 16863 4406 16893 4422
rect 16921 4400 16927 4448
rect 16930 4442 16949 4448
rect 16964 4442 16994 4450
rect 16930 4434 16994 4442
rect 16930 4418 17010 4434
rect 17026 4427 17088 4458
rect 17104 4427 17166 4458
rect 17235 4456 17284 4481
rect 17299 4456 17329 4472
rect 17198 4442 17228 4450
rect 17235 4448 17345 4456
rect 17198 4434 17243 4442
rect 16930 4416 16949 4418
rect 16964 4416 17010 4418
rect 16930 4400 17010 4416
rect 17037 4414 17072 4427
rect 17113 4424 17150 4427
rect 17113 4422 17155 4424
rect 17042 4411 17072 4414
rect 17051 4407 17058 4411
rect 17058 4406 17059 4407
rect 17017 4400 17027 4406
rect 16776 4392 16811 4400
rect 16776 4366 16777 4392
rect 16784 4366 16811 4392
rect 16719 4348 16749 4362
rect 16776 4358 16811 4366
rect 16813 4392 16854 4400
rect 16813 4366 16828 4392
rect 16835 4366 16854 4392
rect 16918 4388 16949 4400
rect 16964 4388 17067 4400
rect 17079 4390 17105 4416
rect 17120 4411 17150 4422
rect 17182 4418 17244 4434
rect 17182 4416 17228 4418
rect 17182 4400 17244 4416
rect 17256 4400 17262 4448
rect 17265 4440 17345 4448
rect 17265 4438 17284 4440
rect 17299 4438 17333 4440
rect 17265 4422 17345 4438
rect 17265 4400 17284 4422
rect 17299 4406 17329 4422
rect 17357 4416 17363 4490
rect 17366 4416 17385 4560
rect 17400 4416 17406 4560
rect 17415 4490 17428 4560
rect 17480 4556 17502 4560
rect 17473 4534 17502 4548
rect 17555 4534 17571 4548
rect 17609 4544 17615 4546
rect 17622 4544 17730 4560
rect 17737 4544 17743 4546
rect 17751 4544 17766 4560
rect 17832 4554 17851 4557
rect 17473 4532 17571 4534
rect 17598 4532 17766 4544
rect 17781 4534 17797 4548
rect 17832 4535 17854 4554
rect 17864 4548 17880 4549
rect 17863 4546 17880 4548
rect 17864 4541 17880 4546
rect 17854 4534 17860 4535
rect 17863 4534 17892 4541
rect 17781 4533 17892 4534
rect 17781 4532 17898 4533
rect 17457 4524 17508 4532
rect 17555 4524 17589 4532
rect 17457 4512 17482 4524
rect 17489 4512 17508 4524
rect 17562 4522 17589 4524
rect 17598 4522 17819 4532
rect 17854 4529 17860 4532
rect 17562 4518 17819 4522
rect 17457 4504 17508 4512
rect 17555 4504 17819 4518
rect 17863 4524 17898 4532
rect 17409 4456 17428 4490
rect 17473 4496 17502 4504
rect 17473 4490 17490 4496
rect 17473 4488 17507 4490
rect 17555 4488 17571 4504
rect 17572 4494 17780 4504
rect 17781 4494 17797 4504
rect 17845 4500 17860 4515
rect 17863 4512 17864 4524
rect 17871 4512 17898 4524
rect 17863 4504 17898 4512
rect 17863 4503 17892 4504
rect 17583 4490 17797 4494
rect 17598 4488 17797 4490
rect 17832 4490 17845 4500
rect 17863 4490 17880 4503
rect 17832 4488 17880 4490
rect 17474 4484 17507 4488
rect 17470 4482 17507 4484
rect 17470 4481 17537 4482
rect 17470 4476 17501 4481
rect 17507 4476 17537 4481
rect 17470 4472 17537 4476
rect 17443 4469 17537 4472
rect 17443 4462 17492 4469
rect 17443 4456 17473 4462
rect 17492 4457 17497 4462
rect 17409 4440 17489 4456
rect 17501 4448 17537 4469
rect 17598 4464 17787 4488
rect 17832 4487 17879 4488
rect 17845 4482 17879 4487
rect 17613 4461 17787 4464
rect 17606 4458 17787 4461
rect 17815 4481 17879 4482
rect 17409 4438 17428 4440
rect 17443 4438 17477 4440
rect 17409 4422 17489 4438
rect 17409 4416 17428 4422
rect 17125 4390 17228 4400
rect 17079 4388 17228 4390
rect 17249 4388 17284 4400
rect 16918 4386 17080 4388
rect 16930 4366 16949 4386
rect 16964 4384 16994 4386
rect 16813 4358 16854 4366
rect 16936 4362 16949 4366
rect 17001 4370 17080 4386
rect 17112 4386 17284 4388
rect 17112 4370 17191 4386
rect 17198 4384 17228 4386
rect 16776 4348 16805 4358
rect 16819 4348 16848 4358
rect 16863 4348 16893 4362
rect 16936 4348 16979 4362
rect 17001 4358 17191 4370
rect 17256 4366 17262 4386
rect 16986 4348 17016 4358
rect 17017 4348 17175 4358
rect 17179 4348 17209 4358
rect 17213 4348 17243 4362
rect 17271 4348 17284 4386
rect 17356 4400 17385 4416
rect 17399 4400 17428 4416
rect 17443 4406 17473 4422
rect 17501 4400 17507 4448
rect 17510 4442 17529 4448
rect 17544 4442 17574 4450
rect 17510 4434 17574 4442
rect 17510 4418 17590 4434
rect 17606 4427 17668 4458
rect 17684 4427 17746 4458
rect 17815 4456 17864 4481
rect 17879 4456 17909 4472
rect 17778 4442 17808 4450
rect 17815 4448 17925 4456
rect 17778 4434 17823 4442
rect 17510 4416 17529 4418
rect 17544 4416 17590 4418
rect 17510 4400 17590 4416
rect 17617 4414 17652 4427
rect 17693 4424 17730 4427
rect 17693 4422 17735 4424
rect 17622 4411 17652 4414
rect 17631 4407 17638 4411
rect 17638 4406 17639 4407
rect 17597 4400 17607 4406
rect 17356 4392 17391 4400
rect 17356 4366 17357 4392
rect 17364 4366 17391 4392
rect 17299 4348 17329 4362
rect 17356 4358 17391 4366
rect 17393 4392 17434 4400
rect 17393 4366 17408 4392
rect 17415 4366 17434 4392
rect 17498 4388 17529 4400
rect 17544 4388 17647 4400
rect 17659 4390 17685 4416
rect 17700 4411 17730 4422
rect 17762 4418 17824 4434
rect 17762 4416 17808 4418
rect 17762 4400 17824 4416
rect 17836 4400 17842 4448
rect 17845 4440 17925 4448
rect 17845 4438 17864 4440
rect 17879 4438 17913 4440
rect 17845 4422 17925 4438
rect 17845 4400 17864 4422
rect 17879 4406 17909 4422
rect 17937 4416 17943 4490
rect 17946 4416 17965 4560
rect 17980 4416 17986 4560
rect 17995 4490 18008 4560
rect 18060 4556 18082 4560
rect 18053 4534 18082 4548
rect 18135 4534 18151 4548
rect 18189 4544 18195 4546
rect 18202 4544 18310 4560
rect 18317 4544 18323 4546
rect 18331 4544 18346 4560
rect 18412 4554 18431 4557
rect 18053 4532 18151 4534
rect 18178 4532 18346 4544
rect 18361 4534 18377 4548
rect 18412 4535 18434 4554
rect 18444 4548 18460 4549
rect 18443 4546 18460 4548
rect 18444 4541 18460 4546
rect 18434 4534 18440 4535
rect 18443 4534 18472 4541
rect 18361 4533 18472 4534
rect 18361 4532 18478 4533
rect 18037 4524 18088 4532
rect 18135 4524 18169 4532
rect 18037 4512 18062 4524
rect 18069 4512 18088 4524
rect 18142 4522 18169 4524
rect 18178 4522 18399 4532
rect 18434 4529 18440 4532
rect 18142 4518 18399 4522
rect 18037 4504 18088 4512
rect 18135 4504 18399 4518
rect 18443 4524 18478 4532
rect 17989 4456 18008 4490
rect 18053 4496 18082 4504
rect 18053 4490 18070 4496
rect 18053 4488 18087 4490
rect 18135 4488 18151 4504
rect 18152 4494 18360 4504
rect 18361 4494 18377 4504
rect 18425 4500 18440 4515
rect 18443 4512 18444 4524
rect 18451 4512 18478 4524
rect 18443 4504 18478 4512
rect 18443 4503 18472 4504
rect 18163 4490 18377 4494
rect 18178 4488 18377 4490
rect 18412 4490 18425 4500
rect 18443 4490 18460 4503
rect 18412 4488 18460 4490
rect 18054 4484 18087 4488
rect 18050 4482 18087 4484
rect 18050 4481 18117 4482
rect 18050 4476 18081 4481
rect 18087 4476 18117 4481
rect 18050 4472 18117 4476
rect 18023 4469 18117 4472
rect 18023 4462 18072 4469
rect 18023 4456 18053 4462
rect 18072 4457 18077 4462
rect 17989 4440 18069 4456
rect 18081 4448 18117 4469
rect 18178 4464 18367 4488
rect 18412 4487 18459 4488
rect 18425 4482 18459 4487
rect 18193 4461 18367 4464
rect 18186 4458 18367 4461
rect 18395 4481 18459 4482
rect 17989 4438 18008 4440
rect 18023 4438 18057 4440
rect 17989 4422 18069 4438
rect 17989 4416 18008 4422
rect 17705 4390 17808 4400
rect 17659 4388 17808 4390
rect 17829 4388 17864 4400
rect 17498 4386 17660 4388
rect 17510 4366 17529 4386
rect 17544 4384 17574 4386
rect 17393 4358 17434 4366
rect 17516 4362 17529 4366
rect 17581 4370 17660 4386
rect 17692 4386 17864 4388
rect 17692 4370 17771 4386
rect 17778 4384 17808 4386
rect 17356 4348 17385 4358
rect 17399 4348 17428 4358
rect 17443 4348 17473 4362
rect 17516 4348 17559 4362
rect 17581 4358 17771 4370
rect 17836 4366 17842 4386
rect 17566 4348 17596 4358
rect 17597 4348 17755 4358
rect 17759 4348 17789 4358
rect 17793 4348 17823 4362
rect 17851 4348 17864 4386
rect 17936 4400 17965 4416
rect 17979 4400 18008 4416
rect 18023 4406 18053 4422
rect 18081 4400 18087 4448
rect 18090 4442 18109 4448
rect 18124 4442 18154 4450
rect 18090 4434 18154 4442
rect 18090 4418 18170 4434
rect 18186 4427 18248 4458
rect 18264 4427 18326 4458
rect 18395 4456 18444 4481
rect 18459 4456 18489 4472
rect 18358 4442 18388 4450
rect 18395 4448 18505 4456
rect 18358 4434 18403 4442
rect 18090 4416 18109 4418
rect 18124 4416 18170 4418
rect 18090 4400 18170 4416
rect 18197 4414 18232 4427
rect 18273 4424 18310 4427
rect 18273 4422 18315 4424
rect 18202 4411 18232 4414
rect 18211 4407 18218 4411
rect 18218 4406 18219 4407
rect 18177 4400 18187 4406
rect 17936 4392 17971 4400
rect 17936 4366 17937 4392
rect 17944 4366 17971 4392
rect 17879 4348 17909 4362
rect 17936 4358 17971 4366
rect 17973 4392 18014 4400
rect 17973 4366 17988 4392
rect 17995 4366 18014 4392
rect 18078 4388 18109 4400
rect 18124 4388 18227 4400
rect 18239 4390 18265 4416
rect 18280 4411 18310 4422
rect 18342 4418 18404 4434
rect 18342 4416 18388 4418
rect 18342 4400 18404 4416
rect 18416 4400 18422 4448
rect 18425 4440 18505 4448
rect 18425 4438 18444 4440
rect 18459 4438 18493 4440
rect 18425 4422 18505 4438
rect 18425 4400 18444 4422
rect 18459 4406 18489 4422
rect 18517 4416 18523 4490
rect 18532 4416 18545 4560
rect 18285 4390 18388 4400
rect 18239 4388 18388 4390
rect 18409 4388 18444 4400
rect 18078 4386 18240 4388
rect 18090 4366 18109 4386
rect 18124 4384 18154 4386
rect 17973 4358 18014 4366
rect 18096 4362 18109 4366
rect 18161 4370 18240 4386
rect 18272 4386 18444 4388
rect 18272 4370 18351 4386
rect 18358 4384 18388 4386
rect 17936 4348 17965 4358
rect 17979 4348 18008 4358
rect 18023 4348 18053 4362
rect 18096 4348 18139 4362
rect 18161 4358 18351 4370
rect 18416 4366 18422 4386
rect 18146 4348 18176 4358
rect 18177 4348 18335 4358
rect 18339 4348 18369 4358
rect 18373 4348 18403 4362
rect 18431 4348 18444 4386
rect 18516 4400 18545 4416
rect 18516 4392 18551 4400
rect 18516 4366 18517 4392
rect 18524 4366 18551 4392
rect 18459 4348 18489 4362
rect 18516 4358 18551 4366
rect 18516 4348 18545 4358
rect -1 4342 18545 4348
rect 0 4334 18545 4342
rect 15 4304 28 4334
rect 43 4320 73 4334
rect 116 4320 159 4334
rect 166 4320 386 4334
rect 393 4320 423 4334
rect 83 4306 98 4318
rect 117 4306 130 4320
rect 198 4316 351 4320
rect 80 4304 102 4306
rect 180 4304 372 4316
rect 451 4304 464 4334
rect 479 4320 509 4334
rect 546 4304 565 4334
rect 580 4304 586 4334
rect 595 4304 608 4334
rect 623 4320 653 4334
rect 696 4320 739 4334
rect 746 4320 966 4334
rect 973 4320 1003 4334
rect 663 4306 678 4318
rect 697 4306 710 4320
rect 778 4316 931 4320
rect 660 4304 682 4306
rect 760 4304 952 4316
rect 1031 4304 1044 4334
rect 1059 4320 1089 4334
rect 1126 4304 1145 4334
rect 1160 4304 1166 4334
rect 1175 4304 1188 4334
rect 1203 4320 1233 4334
rect 1276 4320 1319 4334
rect 1326 4320 1546 4334
rect 1553 4320 1583 4334
rect 1243 4306 1258 4318
rect 1277 4306 1290 4320
rect 1358 4316 1511 4320
rect 1240 4304 1262 4306
rect 1340 4304 1532 4316
rect 1611 4304 1624 4334
rect 1639 4320 1669 4334
rect 1706 4304 1725 4334
rect 1740 4304 1746 4334
rect 1755 4304 1768 4334
rect 1783 4320 1813 4334
rect 1856 4320 1899 4334
rect 1906 4320 2126 4334
rect 2133 4320 2163 4334
rect 1823 4306 1838 4318
rect 1857 4306 1870 4320
rect 1938 4316 2091 4320
rect 1820 4304 1842 4306
rect 1920 4304 2112 4316
rect 2191 4304 2204 4334
rect 2219 4320 2249 4334
rect 2286 4304 2305 4334
rect 2320 4304 2326 4334
rect 2335 4304 2348 4334
rect 2363 4320 2393 4334
rect 2436 4320 2479 4334
rect 2486 4320 2706 4334
rect 2713 4320 2743 4334
rect 2403 4306 2418 4318
rect 2437 4306 2450 4320
rect 2518 4316 2671 4320
rect 2400 4304 2422 4306
rect 2500 4304 2692 4316
rect 2771 4304 2784 4334
rect 2799 4320 2829 4334
rect 2866 4304 2885 4334
rect 2900 4304 2906 4334
rect 2915 4304 2928 4334
rect 2943 4320 2973 4334
rect 3016 4320 3059 4334
rect 3066 4320 3286 4334
rect 3293 4320 3323 4334
rect 2983 4306 2998 4318
rect 3017 4306 3030 4320
rect 3098 4316 3251 4320
rect 2980 4304 3002 4306
rect 3080 4304 3272 4316
rect 3351 4304 3364 4334
rect 3379 4320 3409 4334
rect 3446 4304 3465 4334
rect 3480 4304 3486 4334
rect 3495 4304 3508 4334
rect 3523 4320 3553 4334
rect 3596 4320 3639 4334
rect 3646 4320 3866 4334
rect 3873 4320 3903 4334
rect 3563 4306 3578 4318
rect 3597 4306 3610 4320
rect 3678 4316 3831 4320
rect 3560 4304 3582 4306
rect 3660 4304 3852 4316
rect 3931 4304 3944 4334
rect 3959 4320 3989 4334
rect 4026 4304 4045 4334
rect 4060 4304 4066 4334
rect 4075 4304 4088 4334
rect 4103 4320 4133 4334
rect 4176 4320 4219 4334
rect 4226 4320 4446 4334
rect 4453 4320 4483 4334
rect 4143 4306 4158 4318
rect 4177 4306 4190 4320
rect 4258 4316 4411 4320
rect 4140 4304 4162 4306
rect 4240 4304 4432 4316
rect 4511 4304 4524 4334
rect 4539 4320 4569 4334
rect 4606 4304 4625 4334
rect 4640 4304 4646 4334
rect 4655 4304 4668 4334
rect 4683 4320 4713 4334
rect 4756 4320 4799 4334
rect 4806 4320 5026 4334
rect 5033 4320 5063 4334
rect 4723 4306 4738 4318
rect 4757 4306 4770 4320
rect 4838 4316 4991 4320
rect 4720 4304 4742 4306
rect 4820 4304 5012 4316
rect 5091 4304 5104 4334
rect 5119 4320 5149 4334
rect 5186 4304 5205 4334
rect 5220 4304 5226 4334
rect 5235 4304 5248 4334
rect 5263 4320 5293 4334
rect 5336 4320 5379 4334
rect 5386 4320 5606 4334
rect 5613 4320 5643 4334
rect 5303 4306 5318 4318
rect 5337 4306 5350 4320
rect 5418 4316 5571 4320
rect 5300 4304 5322 4306
rect 5400 4304 5592 4316
rect 5671 4304 5684 4334
rect 5699 4320 5729 4334
rect 5766 4304 5785 4334
rect 5800 4304 5806 4334
rect 5815 4304 5828 4334
rect 5843 4320 5873 4334
rect 5916 4320 5959 4334
rect 5966 4320 6186 4334
rect 6193 4320 6223 4334
rect 5883 4306 5898 4318
rect 5917 4306 5930 4320
rect 5998 4316 6151 4320
rect 5880 4304 5902 4306
rect 5980 4304 6172 4316
rect 6251 4304 6264 4334
rect 6279 4320 6309 4334
rect 6346 4304 6365 4334
rect 6380 4304 6386 4334
rect 6395 4304 6408 4334
rect 6423 4320 6453 4334
rect 6496 4320 6539 4334
rect 6546 4320 6766 4334
rect 6773 4320 6803 4334
rect 6463 4306 6478 4318
rect 6497 4306 6510 4320
rect 6578 4316 6731 4320
rect 6460 4304 6482 4306
rect 6560 4304 6752 4316
rect 6831 4304 6844 4334
rect 6859 4320 6889 4334
rect 6926 4304 6945 4334
rect 6960 4304 6966 4334
rect 6975 4304 6988 4334
rect 7003 4320 7033 4334
rect 7076 4320 7119 4334
rect 7126 4320 7346 4334
rect 7353 4320 7383 4334
rect 7043 4306 7058 4318
rect 7077 4306 7090 4320
rect 7158 4316 7311 4320
rect 7040 4304 7062 4306
rect 7140 4304 7332 4316
rect 7411 4304 7424 4334
rect 7439 4320 7469 4334
rect 7506 4304 7525 4334
rect 7540 4304 7546 4334
rect 7555 4304 7568 4334
rect 7583 4320 7613 4334
rect 7656 4320 7699 4334
rect 7706 4320 7926 4334
rect 7933 4320 7963 4334
rect 7623 4306 7638 4318
rect 7657 4306 7670 4320
rect 7738 4316 7891 4320
rect 7620 4304 7642 4306
rect 7720 4304 7912 4316
rect 7991 4304 8004 4334
rect 8019 4320 8049 4334
rect 8086 4304 8105 4334
rect 8120 4304 8126 4334
rect 8135 4304 8148 4334
rect 8163 4320 8193 4334
rect 8236 4320 8279 4334
rect 8286 4320 8506 4334
rect 8513 4320 8543 4334
rect 8203 4306 8218 4318
rect 8237 4306 8250 4320
rect 8318 4316 8471 4320
rect 8200 4304 8222 4306
rect 8300 4304 8492 4316
rect 8571 4304 8584 4334
rect 8599 4320 8629 4334
rect 8666 4304 8685 4334
rect 8700 4304 8706 4334
rect 8715 4304 8728 4334
rect 8743 4320 8773 4334
rect 8816 4320 8859 4334
rect 8866 4320 9086 4334
rect 9093 4320 9123 4334
rect 8783 4306 8798 4318
rect 8817 4306 8830 4320
rect 8898 4316 9051 4320
rect 8780 4304 8802 4306
rect 8880 4304 9072 4316
rect 9151 4304 9164 4334
rect 9179 4320 9209 4334
rect 9246 4304 9265 4334
rect 9280 4304 9286 4334
rect 9295 4304 9308 4334
rect 9323 4320 9353 4334
rect 9396 4320 9439 4334
rect 9446 4320 9666 4334
rect 9673 4320 9703 4334
rect 9363 4306 9378 4318
rect 9397 4306 9410 4320
rect 9478 4316 9631 4320
rect 9360 4304 9382 4306
rect 9460 4304 9652 4316
rect 9731 4304 9744 4334
rect 9759 4320 9789 4334
rect 9826 4304 9845 4334
rect 9860 4304 9866 4334
rect 9875 4304 9888 4334
rect 9903 4320 9933 4334
rect 9976 4320 10019 4334
rect 10026 4320 10246 4334
rect 10253 4320 10283 4334
rect 9943 4306 9958 4318
rect 9977 4306 9990 4320
rect 10058 4316 10211 4320
rect 9940 4304 9962 4306
rect 10040 4304 10232 4316
rect 10311 4304 10324 4334
rect 10339 4320 10369 4334
rect 10406 4304 10425 4334
rect 10440 4304 10446 4334
rect 10455 4304 10468 4334
rect 10483 4320 10513 4334
rect 10556 4320 10599 4334
rect 10606 4320 10826 4334
rect 10833 4320 10863 4334
rect 10523 4306 10538 4318
rect 10557 4306 10570 4320
rect 10638 4316 10791 4320
rect 10520 4304 10542 4306
rect 10620 4304 10812 4316
rect 10891 4304 10904 4334
rect 10919 4320 10949 4334
rect 10986 4304 11005 4334
rect 11020 4304 11026 4334
rect 11035 4304 11048 4334
rect 11063 4320 11093 4334
rect 11136 4320 11179 4334
rect 11186 4320 11406 4334
rect 11413 4320 11443 4334
rect 11103 4306 11118 4318
rect 11137 4306 11150 4320
rect 11218 4316 11371 4320
rect 11100 4304 11122 4306
rect 11200 4304 11392 4316
rect 11471 4304 11484 4334
rect 11499 4320 11529 4334
rect 11566 4304 11585 4334
rect 11600 4304 11606 4334
rect 11615 4304 11628 4334
rect 11643 4320 11673 4334
rect 11716 4320 11759 4334
rect 11766 4320 11986 4334
rect 11993 4320 12023 4334
rect 11683 4306 11698 4318
rect 11717 4306 11730 4320
rect 11798 4316 11951 4320
rect 11680 4304 11702 4306
rect 11780 4304 11972 4316
rect 12051 4304 12064 4334
rect 12079 4320 12109 4334
rect 12146 4304 12165 4334
rect 12180 4304 12186 4334
rect 12195 4304 12208 4334
rect 12223 4320 12253 4334
rect 12296 4320 12339 4334
rect 12346 4320 12566 4334
rect 12573 4320 12603 4334
rect 12263 4306 12278 4318
rect 12297 4306 12310 4320
rect 12378 4316 12531 4320
rect 12260 4304 12282 4306
rect 12360 4304 12552 4316
rect 12631 4304 12644 4334
rect 12659 4320 12689 4334
rect 12726 4304 12745 4334
rect 12760 4304 12766 4334
rect 12775 4304 12788 4334
rect 12803 4320 12833 4334
rect 12876 4320 12919 4334
rect 12926 4320 13146 4334
rect 13153 4320 13183 4334
rect 12843 4306 12858 4318
rect 12877 4306 12890 4320
rect 12958 4316 13111 4320
rect 12840 4304 12862 4306
rect 12940 4304 13132 4316
rect 13211 4304 13224 4334
rect 13239 4320 13269 4334
rect 13306 4304 13325 4334
rect 13340 4304 13346 4334
rect 13355 4304 13368 4334
rect 13383 4320 13413 4334
rect 13456 4320 13499 4334
rect 13506 4320 13726 4334
rect 13733 4320 13763 4334
rect 13423 4306 13438 4318
rect 13457 4306 13470 4320
rect 13538 4316 13691 4320
rect 13420 4304 13442 4306
rect 13520 4304 13712 4316
rect 13791 4304 13804 4334
rect 13819 4320 13849 4334
rect 13886 4304 13905 4334
rect 13920 4304 13926 4334
rect 13935 4304 13948 4334
rect 13963 4320 13993 4334
rect 14036 4320 14079 4334
rect 14086 4320 14306 4334
rect 14313 4320 14343 4334
rect 14003 4306 14018 4318
rect 14037 4306 14050 4320
rect 14118 4316 14271 4320
rect 14000 4304 14022 4306
rect 14100 4304 14292 4316
rect 14371 4304 14384 4334
rect 14399 4320 14429 4334
rect 14466 4304 14485 4334
rect 14500 4304 14506 4334
rect 14515 4304 14528 4334
rect 14543 4320 14573 4334
rect 14616 4320 14659 4334
rect 14666 4320 14886 4334
rect 14893 4320 14923 4334
rect 14583 4306 14598 4318
rect 14617 4306 14630 4320
rect 14698 4316 14851 4320
rect 14580 4304 14602 4306
rect 14680 4304 14872 4316
rect 14951 4304 14964 4334
rect 14979 4320 15009 4334
rect 15046 4304 15065 4334
rect 15080 4304 15086 4334
rect 15095 4304 15108 4334
rect 15123 4320 15153 4334
rect 15196 4320 15239 4334
rect 15246 4320 15466 4334
rect 15473 4320 15503 4334
rect 15163 4306 15178 4318
rect 15197 4306 15210 4320
rect 15278 4316 15431 4320
rect 15160 4304 15182 4306
rect 15260 4304 15452 4316
rect 15531 4304 15544 4334
rect 15559 4320 15589 4334
rect 15626 4304 15645 4334
rect 15660 4304 15666 4334
rect 15675 4304 15688 4334
rect 15703 4320 15733 4334
rect 15776 4320 15819 4334
rect 15826 4320 16046 4334
rect 16053 4320 16083 4334
rect 15743 4306 15758 4318
rect 15777 4306 15790 4320
rect 15858 4316 16011 4320
rect 15740 4304 15762 4306
rect 15840 4304 16032 4316
rect 16111 4304 16124 4334
rect 16139 4320 16169 4334
rect 16206 4304 16225 4334
rect 16240 4304 16246 4334
rect 16255 4304 16268 4334
rect 16283 4320 16313 4334
rect 16356 4320 16399 4334
rect 16406 4320 16626 4334
rect 16633 4320 16663 4334
rect 16323 4306 16338 4318
rect 16357 4306 16370 4320
rect 16438 4316 16591 4320
rect 16320 4304 16342 4306
rect 16420 4304 16612 4316
rect 16691 4304 16704 4334
rect 16719 4320 16749 4334
rect 16786 4304 16805 4334
rect 16820 4304 16826 4334
rect 16835 4304 16848 4334
rect 16863 4320 16893 4334
rect 16936 4320 16979 4334
rect 16986 4320 17206 4334
rect 17213 4320 17243 4334
rect 16903 4306 16918 4318
rect 16937 4306 16950 4320
rect 17018 4316 17171 4320
rect 16900 4304 16922 4306
rect 17000 4304 17192 4316
rect 17271 4304 17284 4334
rect 17299 4320 17329 4334
rect 17366 4304 17385 4334
rect 17400 4304 17406 4334
rect 17415 4304 17428 4334
rect 17443 4320 17473 4334
rect 17516 4320 17559 4334
rect 17566 4320 17786 4334
rect 17793 4320 17823 4334
rect 17483 4306 17498 4318
rect 17517 4306 17530 4320
rect 17598 4316 17751 4320
rect 17480 4304 17502 4306
rect 17580 4304 17772 4316
rect 17851 4304 17864 4334
rect 17879 4320 17909 4334
rect 17946 4304 17965 4334
rect 17980 4304 17986 4334
rect 17995 4304 18008 4334
rect 18023 4320 18053 4334
rect 18096 4320 18139 4334
rect 18146 4320 18366 4334
rect 18373 4320 18403 4334
rect 18063 4306 18078 4318
rect 18097 4306 18110 4320
rect 18178 4316 18331 4320
rect 18060 4304 18082 4306
rect 18160 4304 18352 4316
rect 18431 4304 18444 4334
rect 18459 4320 18489 4334
rect 18532 4304 18545 4334
rect 0 4290 18545 4304
rect 15 4220 28 4290
rect 80 4286 102 4290
rect 73 4264 102 4278
rect 155 4264 171 4278
rect 209 4274 215 4276
rect 222 4274 330 4290
rect 337 4274 343 4276
rect 351 4274 366 4290
rect 432 4284 451 4287
rect 73 4262 171 4264
rect 198 4262 366 4274
rect 381 4264 397 4278
rect 432 4265 454 4284
rect 464 4278 480 4279
rect 463 4276 480 4278
rect 464 4271 480 4276
rect 454 4264 460 4265
rect 463 4264 492 4271
rect 381 4263 492 4264
rect 381 4262 498 4263
rect 57 4254 108 4262
rect 155 4254 189 4262
rect 57 4242 82 4254
rect 89 4242 108 4254
rect 162 4252 189 4254
rect 198 4252 419 4262
rect 454 4259 460 4262
rect 162 4248 419 4252
rect 57 4234 108 4242
rect 155 4234 419 4248
rect 463 4254 498 4262
rect 9 4186 28 4220
rect 73 4226 102 4234
rect 73 4220 90 4226
rect 73 4218 107 4220
rect 155 4218 171 4234
rect 172 4224 380 4234
rect 381 4224 397 4234
rect 445 4230 460 4245
rect 463 4242 464 4254
rect 471 4242 498 4254
rect 463 4234 498 4242
rect 463 4233 492 4234
rect 183 4220 397 4224
rect 198 4218 397 4220
rect 432 4220 445 4230
rect 463 4220 480 4233
rect 432 4218 480 4220
rect 74 4214 107 4218
rect 70 4212 107 4214
rect 70 4211 137 4212
rect 70 4206 101 4211
rect 107 4206 137 4211
rect 70 4202 137 4206
rect 43 4199 137 4202
rect 43 4192 92 4199
rect 43 4186 73 4192
rect 92 4187 97 4192
rect 9 4170 89 4186
rect 101 4178 137 4199
rect 198 4194 387 4218
rect 432 4217 479 4218
rect 445 4212 479 4217
rect 213 4191 387 4194
rect 206 4188 387 4191
rect 415 4211 479 4212
rect 9 4168 28 4170
rect 43 4168 77 4170
rect 9 4152 89 4168
rect 9 4146 28 4152
rect -1 4130 28 4146
rect 43 4136 73 4152
rect 101 4130 107 4178
rect 110 4172 129 4178
rect 144 4172 174 4180
rect 110 4164 174 4172
rect 110 4148 190 4164
rect 206 4157 268 4188
rect 284 4157 346 4188
rect 415 4186 464 4211
rect 479 4186 509 4202
rect 378 4172 408 4180
rect 415 4178 525 4186
rect 378 4164 423 4172
rect 110 4146 129 4148
rect 144 4146 190 4148
rect 110 4130 190 4146
rect 217 4144 252 4157
rect 293 4154 330 4157
rect 293 4152 335 4154
rect 222 4141 252 4144
rect 231 4137 238 4141
rect 238 4136 239 4137
rect 197 4130 207 4136
rect -7 4122 34 4130
rect -7 4096 8 4122
rect 15 4096 34 4122
rect 98 4118 129 4130
rect 144 4118 247 4130
rect 259 4120 285 4146
rect 300 4141 330 4152
rect 362 4148 424 4164
rect 362 4146 408 4148
rect 362 4130 424 4146
rect 436 4130 442 4178
rect 445 4170 525 4178
rect 445 4168 464 4170
rect 479 4168 513 4170
rect 445 4152 525 4168
rect 445 4130 464 4152
rect 479 4136 509 4152
rect 537 4146 543 4220
rect 546 4146 565 4290
rect 580 4146 586 4290
rect 595 4220 608 4290
rect 660 4286 682 4290
rect 653 4264 682 4278
rect 735 4264 751 4278
rect 789 4274 795 4276
rect 802 4274 910 4290
rect 917 4274 923 4276
rect 931 4274 946 4290
rect 1012 4284 1031 4287
rect 653 4262 751 4264
rect 778 4262 946 4274
rect 961 4264 977 4278
rect 1012 4265 1034 4284
rect 1044 4278 1060 4279
rect 1043 4276 1060 4278
rect 1044 4271 1060 4276
rect 1034 4264 1040 4265
rect 1043 4264 1072 4271
rect 961 4263 1072 4264
rect 961 4262 1078 4263
rect 637 4254 688 4262
rect 735 4254 769 4262
rect 637 4242 662 4254
rect 669 4242 688 4254
rect 742 4252 769 4254
rect 778 4252 999 4262
rect 1034 4259 1040 4262
rect 742 4248 999 4252
rect 637 4234 688 4242
rect 735 4234 999 4248
rect 1043 4254 1078 4262
rect 589 4186 608 4220
rect 653 4226 682 4234
rect 653 4220 670 4226
rect 653 4218 687 4220
rect 735 4218 751 4234
rect 752 4224 960 4234
rect 961 4224 977 4234
rect 1025 4230 1040 4245
rect 1043 4242 1044 4254
rect 1051 4242 1078 4254
rect 1043 4234 1078 4242
rect 1043 4233 1072 4234
rect 763 4220 977 4224
rect 778 4218 977 4220
rect 1012 4220 1025 4230
rect 1043 4220 1060 4233
rect 1012 4218 1060 4220
rect 654 4214 687 4218
rect 650 4212 687 4214
rect 650 4211 717 4212
rect 650 4206 681 4211
rect 687 4206 717 4211
rect 650 4202 717 4206
rect 623 4199 717 4202
rect 623 4192 672 4199
rect 623 4186 653 4192
rect 672 4187 677 4192
rect 589 4170 669 4186
rect 681 4178 717 4199
rect 778 4194 967 4218
rect 1012 4217 1059 4218
rect 1025 4212 1059 4217
rect 793 4191 967 4194
rect 786 4188 967 4191
rect 995 4211 1059 4212
rect 589 4168 608 4170
rect 623 4168 657 4170
rect 589 4152 669 4168
rect 589 4146 608 4152
rect 305 4120 408 4130
rect 259 4118 408 4120
rect 429 4118 464 4130
rect 98 4116 260 4118
rect 110 4096 129 4116
rect 144 4114 174 4116
rect -7 4088 34 4096
rect 116 4092 129 4096
rect 181 4100 260 4116
rect 292 4116 464 4118
rect 292 4100 371 4116
rect 378 4114 408 4116
rect -1 4078 28 4088
rect 43 4078 73 4092
rect 116 4078 159 4092
rect 181 4088 371 4100
rect 436 4096 442 4116
rect 166 4078 196 4088
rect 197 4078 355 4088
rect 359 4078 389 4088
rect 393 4078 423 4092
rect 451 4078 464 4116
rect 536 4130 565 4146
rect 579 4130 608 4146
rect 623 4136 653 4152
rect 681 4130 687 4178
rect 690 4172 709 4178
rect 724 4172 754 4180
rect 690 4164 754 4172
rect 690 4148 770 4164
rect 786 4157 848 4188
rect 864 4157 926 4188
rect 995 4186 1044 4211
rect 1059 4186 1089 4202
rect 958 4172 988 4180
rect 995 4178 1105 4186
rect 958 4164 1003 4172
rect 690 4146 709 4148
rect 724 4146 770 4148
rect 690 4130 770 4146
rect 797 4144 832 4157
rect 873 4154 910 4157
rect 873 4152 915 4154
rect 802 4141 832 4144
rect 811 4137 818 4141
rect 818 4136 819 4137
rect 777 4130 787 4136
rect 536 4122 571 4130
rect 536 4096 537 4122
rect 544 4096 571 4122
rect 479 4078 509 4092
rect 536 4088 571 4096
rect 573 4122 614 4130
rect 573 4096 588 4122
rect 595 4096 614 4122
rect 678 4118 709 4130
rect 724 4118 827 4130
rect 839 4120 865 4146
rect 880 4141 910 4152
rect 942 4148 1004 4164
rect 942 4146 988 4148
rect 942 4130 1004 4146
rect 1016 4130 1022 4178
rect 1025 4170 1105 4178
rect 1025 4168 1044 4170
rect 1059 4168 1093 4170
rect 1025 4152 1105 4168
rect 1025 4130 1044 4152
rect 1059 4136 1089 4152
rect 1117 4146 1123 4220
rect 1126 4146 1145 4290
rect 1160 4146 1166 4290
rect 1175 4220 1188 4290
rect 1240 4286 1262 4290
rect 1233 4264 1262 4278
rect 1315 4264 1331 4278
rect 1369 4274 1375 4276
rect 1382 4274 1490 4290
rect 1497 4274 1503 4276
rect 1511 4274 1526 4290
rect 1592 4284 1611 4287
rect 1233 4262 1331 4264
rect 1358 4262 1526 4274
rect 1541 4264 1557 4278
rect 1592 4265 1614 4284
rect 1624 4278 1640 4279
rect 1623 4276 1640 4278
rect 1624 4271 1640 4276
rect 1614 4264 1620 4265
rect 1623 4264 1652 4271
rect 1541 4263 1652 4264
rect 1541 4262 1658 4263
rect 1217 4254 1268 4262
rect 1315 4254 1349 4262
rect 1217 4242 1242 4254
rect 1249 4242 1268 4254
rect 1322 4252 1349 4254
rect 1358 4252 1579 4262
rect 1614 4259 1620 4262
rect 1322 4248 1579 4252
rect 1217 4234 1268 4242
rect 1315 4234 1579 4248
rect 1623 4254 1658 4262
rect 1169 4186 1188 4220
rect 1233 4226 1262 4234
rect 1233 4220 1250 4226
rect 1233 4218 1267 4220
rect 1315 4218 1331 4234
rect 1332 4224 1540 4234
rect 1541 4224 1557 4234
rect 1605 4230 1620 4245
rect 1623 4242 1624 4254
rect 1631 4242 1658 4254
rect 1623 4234 1658 4242
rect 1623 4233 1652 4234
rect 1343 4220 1557 4224
rect 1358 4218 1557 4220
rect 1592 4220 1605 4230
rect 1623 4220 1640 4233
rect 1592 4218 1640 4220
rect 1234 4214 1267 4218
rect 1230 4212 1267 4214
rect 1230 4211 1297 4212
rect 1230 4206 1261 4211
rect 1267 4206 1297 4211
rect 1230 4202 1297 4206
rect 1203 4199 1297 4202
rect 1203 4192 1252 4199
rect 1203 4186 1233 4192
rect 1252 4187 1257 4192
rect 1169 4170 1249 4186
rect 1261 4178 1297 4199
rect 1358 4194 1547 4218
rect 1592 4217 1639 4218
rect 1605 4212 1639 4217
rect 1373 4191 1547 4194
rect 1366 4188 1547 4191
rect 1575 4211 1639 4212
rect 1169 4168 1188 4170
rect 1203 4168 1237 4170
rect 1169 4152 1249 4168
rect 1169 4146 1188 4152
rect 885 4120 988 4130
rect 839 4118 988 4120
rect 1009 4118 1044 4130
rect 678 4116 840 4118
rect 690 4096 709 4116
rect 724 4114 754 4116
rect 573 4088 614 4096
rect 696 4092 709 4096
rect 761 4100 840 4116
rect 872 4116 1044 4118
rect 872 4100 951 4116
rect 958 4114 988 4116
rect 536 4078 565 4088
rect 579 4078 608 4088
rect 623 4078 653 4092
rect 696 4078 739 4092
rect 761 4088 951 4100
rect 1016 4096 1022 4116
rect 746 4078 776 4088
rect 777 4078 935 4088
rect 939 4078 969 4088
rect 973 4078 1003 4092
rect 1031 4078 1044 4116
rect 1116 4130 1145 4146
rect 1159 4130 1188 4146
rect 1203 4136 1233 4152
rect 1261 4130 1267 4178
rect 1270 4172 1289 4178
rect 1304 4172 1334 4180
rect 1270 4164 1334 4172
rect 1270 4148 1350 4164
rect 1366 4157 1428 4188
rect 1444 4157 1506 4188
rect 1575 4186 1624 4211
rect 1639 4186 1669 4202
rect 1538 4172 1568 4180
rect 1575 4178 1685 4186
rect 1538 4164 1583 4172
rect 1270 4146 1289 4148
rect 1304 4146 1350 4148
rect 1270 4130 1350 4146
rect 1377 4144 1412 4157
rect 1453 4154 1490 4157
rect 1453 4152 1495 4154
rect 1382 4141 1412 4144
rect 1391 4137 1398 4141
rect 1398 4136 1399 4137
rect 1357 4130 1367 4136
rect 1116 4122 1151 4130
rect 1116 4096 1117 4122
rect 1124 4096 1151 4122
rect 1059 4078 1089 4092
rect 1116 4088 1151 4096
rect 1153 4122 1194 4130
rect 1153 4096 1168 4122
rect 1175 4096 1194 4122
rect 1258 4118 1289 4130
rect 1304 4118 1407 4130
rect 1419 4120 1445 4146
rect 1460 4141 1490 4152
rect 1522 4148 1584 4164
rect 1522 4146 1568 4148
rect 1522 4130 1584 4146
rect 1596 4130 1602 4178
rect 1605 4170 1685 4178
rect 1605 4168 1624 4170
rect 1639 4168 1673 4170
rect 1605 4152 1685 4168
rect 1605 4130 1624 4152
rect 1639 4136 1669 4152
rect 1697 4146 1703 4220
rect 1706 4146 1725 4290
rect 1740 4146 1746 4290
rect 1755 4220 1768 4290
rect 1820 4286 1842 4290
rect 1813 4264 1842 4278
rect 1895 4264 1911 4278
rect 1949 4274 1955 4276
rect 1962 4274 2070 4290
rect 2077 4274 2083 4276
rect 2091 4274 2106 4290
rect 2172 4284 2191 4287
rect 1813 4262 1911 4264
rect 1938 4262 2106 4274
rect 2121 4264 2137 4278
rect 2172 4265 2194 4284
rect 2204 4278 2220 4279
rect 2203 4276 2220 4278
rect 2204 4271 2220 4276
rect 2194 4264 2200 4265
rect 2203 4264 2232 4271
rect 2121 4263 2232 4264
rect 2121 4262 2238 4263
rect 1797 4254 1848 4262
rect 1895 4254 1929 4262
rect 1797 4242 1822 4254
rect 1829 4242 1848 4254
rect 1902 4252 1929 4254
rect 1938 4252 2159 4262
rect 2194 4259 2200 4262
rect 1902 4248 2159 4252
rect 1797 4234 1848 4242
rect 1895 4234 2159 4248
rect 2203 4254 2238 4262
rect 1749 4186 1768 4220
rect 1813 4226 1842 4234
rect 1813 4220 1830 4226
rect 1813 4218 1847 4220
rect 1895 4218 1911 4234
rect 1912 4224 2120 4234
rect 2121 4224 2137 4234
rect 2185 4230 2200 4245
rect 2203 4242 2204 4254
rect 2211 4242 2238 4254
rect 2203 4234 2238 4242
rect 2203 4233 2232 4234
rect 1923 4220 2137 4224
rect 1938 4218 2137 4220
rect 2172 4220 2185 4230
rect 2203 4220 2220 4233
rect 2172 4218 2220 4220
rect 1814 4214 1847 4218
rect 1810 4212 1847 4214
rect 1810 4211 1877 4212
rect 1810 4206 1841 4211
rect 1847 4206 1877 4211
rect 1810 4202 1877 4206
rect 1783 4199 1877 4202
rect 1783 4192 1832 4199
rect 1783 4186 1813 4192
rect 1832 4187 1837 4192
rect 1749 4170 1829 4186
rect 1841 4178 1877 4199
rect 1938 4194 2127 4218
rect 2172 4217 2219 4218
rect 2185 4212 2219 4217
rect 1953 4191 2127 4194
rect 1946 4188 2127 4191
rect 2155 4211 2219 4212
rect 1749 4168 1768 4170
rect 1783 4168 1817 4170
rect 1749 4152 1829 4168
rect 1749 4146 1768 4152
rect 1465 4120 1568 4130
rect 1419 4118 1568 4120
rect 1589 4118 1624 4130
rect 1258 4116 1420 4118
rect 1270 4096 1289 4116
rect 1304 4114 1334 4116
rect 1153 4088 1194 4096
rect 1276 4092 1289 4096
rect 1341 4100 1420 4116
rect 1452 4116 1624 4118
rect 1452 4100 1531 4116
rect 1538 4114 1568 4116
rect 1116 4078 1145 4088
rect 1159 4078 1188 4088
rect 1203 4078 1233 4092
rect 1276 4078 1319 4092
rect 1341 4088 1531 4100
rect 1596 4096 1602 4116
rect 1326 4078 1356 4088
rect 1357 4078 1515 4088
rect 1519 4078 1549 4088
rect 1553 4078 1583 4092
rect 1611 4078 1624 4116
rect 1696 4130 1725 4146
rect 1739 4130 1768 4146
rect 1783 4136 1813 4152
rect 1841 4130 1847 4178
rect 1850 4172 1869 4178
rect 1884 4172 1914 4180
rect 1850 4164 1914 4172
rect 1850 4148 1930 4164
rect 1946 4157 2008 4188
rect 2024 4157 2086 4188
rect 2155 4186 2204 4211
rect 2219 4186 2249 4202
rect 2118 4172 2148 4180
rect 2155 4178 2265 4186
rect 2118 4164 2163 4172
rect 1850 4146 1869 4148
rect 1884 4146 1930 4148
rect 1850 4130 1930 4146
rect 1957 4144 1992 4157
rect 2033 4154 2070 4157
rect 2033 4152 2075 4154
rect 1962 4141 1992 4144
rect 1971 4137 1978 4141
rect 1978 4136 1979 4137
rect 1937 4130 1947 4136
rect 1696 4122 1731 4130
rect 1696 4096 1697 4122
rect 1704 4096 1731 4122
rect 1639 4078 1669 4092
rect 1696 4088 1731 4096
rect 1733 4122 1774 4130
rect 1733 4096 1748 4122
rect 1755 4096 1774 4122
rect 1838 4118 1869 4130
rect 1884 4118 1987 4130
rect 1999 4120 2025 4146
rect 2040 4141 2070 4152
rect 2102 4148 2164 4164
rect 2102 4146 2148 4148
rect 2102 4130 2164 4146
rect 2176 4130 2182 4178
rect 2185 4170 2265 4178
rect 2185 4168 2204 4170
rect 2219 4168 2253 4170
rect 2185 4152 2265 4168
rect 2185 4130 2204 4152
rect 2219 4136 2249 4152
rect 2277 4146 2283 4220
rect 2286 4146 2305 4290
rect 2320 4146 2326 4290
rect 2335 4220 2348 4290
rect 2400 4286 2422 4290
rect 2393 4264 2422 4278
rect 2475 4264 2491 4278
rect 2529 4274 2535 4276
rect 2542 4274 2650 4290
rect 2657 4274 2663 4276
rect 2671 4274 2686 4290
rect 2752 4284 2771 4287
rect 2393 4262 2491 4264
rect 2518 4262 2686 4274
rect 2701 4264 2717 4278
rect 2752 4265 2774 4284
rect 2784 4278 2800 4279
rect 2783 4276 2800 4278
rect 2784 4271 2800 4276
rect 2774 4264 2780 4265
rect 2783 4264 2812 4271
rect 2701 4263 2812 4264
rect 2701 4262 2818 4263
rect 2377 4254 2428 4262
rect 2475 4254 2509 4262
rect 2377 4242 2402 4254
rect 2409 4242 2428 4254
rect 2482 4252 2509 4254
rect 2518 4252 2739 4262
rect 2774 4259 2780 4262
rect 2482 4248 2739 4252
rect 2377 4234 2428 4242
rect 2475 4234 2739 4248
rect 2783 4254 2818 4262
rect 2329 4186 2348 4220
rect 2393 4226 2422 4234
rect 2393 4220 2410 4226
rect 2393 4218 2427 4220
rect 2475 4218 2491 4234
rect 2492 4224 2700 4234
rect 2701 4224 2717 4234
rect 2765 4230 2780 4245
rect 2783 4242 2784 4254
rect 2791 4242 2818 4254
rect 2783 4234 2818 4242
rect 2783 4233 2812 4234
rect 2503 4220 2717 4224
rect 2518 4218 2717 4220
rect 2752 4220 2765 4230
rect 2783 4220 2800 4233
rect 2752 4218 2800 4220
rect 2394 4214 2427 4218
rect 2390 4212 2427 4214
rect 2390 4211 2457 4212
rect 2390 4206 2421 4211
rect 2427 4206 2457 4211
rect 2390 4202 2457 4206
rect 2363 4199 2457 4202
rect 2363 4192 2412 4199
rect 2363 4186 2393 4192
rect 2412 4187 2417 4192
rect 2329 4170 2409 4186
rect 2421 4178 2457 4199
rect 2518 4194 2707 4218
rect 2752 4217 2799 4218
rect 2765 4212 2799 4217
rect 2533 4191 2707 4194
rect 2526 4188 2707 4191
rect 2735 4211 2799 4212
rect 2329 4168 2348 4170
rect 2363 4168 2397 4170
rect 2329 4152 2409 4168
rect 2329 4146 2348 4152
rect 2045 4120 2148 4130
rect 1999 4118 2148 4120
rect 2169 4118 2204 4130
rect 1838 4116 2000 4118
rect 1850 4096 1869 4116
rect 1884 4114 1914 4116
rect 1733 4088 1774 4096
rect 1856 4092 1869 4096
rect 1921 4100 2000 4116
rect 2032 4116 2204 4118
rect 2032 4100 2111 4116
rect 2118 4114 2148 4116
rect 1696 4078 1725 4088
rect 1739 4078 1768 4088
rect 1783 4078 1813 4092
rect 1856 4078 1899 4092
rect 1921 4088 2111 4100
rect 2176 4096 2182 4116
rect 1906 4078 1936 4088
rect 1937 4078 2095 4088
rect 2099 4078 2129 4088
rect 2133 4078 2163 4092
rect 2191 4078 2204 4116
rect 2276 4130 2305 4146
rect 2319 4130 2348 4146
rect 2363 4136 2393 4152
rect 2421 4130 2427 4178
rect 2430 4172 2449 4178
rect 2464 4172 2494 4180
rect 2430 4164 2494 4172
rect 2430 4148 2510 4164
rect 2526 4157 2588 4188
rect 2604 4157 2666 4188
rect 2735 4186 2784 4211
rect 2799 4186 2829 4202
rect 2698 4172 2728 4180
rect 2735 4178 2845 4186
rect 2698 4164 2743 4172
rect 2430 4146 2449 4148
rect 2464 4146 2510 4148
rect 2430 4130 2510 4146
rect 2537 4144 2572 4157
rect 2613 4154 2650 4157
rect 2613 4152 2655 4154
rect 2542 4141 2572 4144
rect 2551 4137 2558 4141
rect 2558 4136 2559 4137
rect 2517 4130 2527 4136
rect 2276 4122 2311 4130
rect 2276 4096 2277 4122
rect 2284 4096 2311 4122
rect 2219 4078 2249 4092
rect 2276 4088 2311 4096
rect 2313 4122 2354 4130
rect 2313 4096 2328 4122
rect 2335 4096 2354 4122
rect 2418 4118 2449 4130
rect 2464 4118 2567 4130
rect 2579 4120 2605 4146
rect 2620 4141 2650 4152
rect 2682 4148 2744 4164
rect 2682 4146 2728 4148
rect 2682 4130 2744 4146
rect 2756 4130 2762 4178
rect 2765 4170 2845 4178
rect 2765 4168 2784 4170
rect 2799 4168 2833 4170
rect 2765 4152 2845 4168
rect 2765 4130 2784 4152
rect 2799 4136 2829 4152
rect 2857 4146 2863 4220
rect 2866 4146 2885 4290
rect 2900 4146 2906 4290
rect 2915 4220 2928 4290
rect 2980 4286 3002 4290
rect 2973 4264 3002 4278
rect 3055 4264 3071 4278
rect 3109 4274 3115 4276
rect 3122 4274 3230 4290
rect 3237 4274 3243 4276
rect 3251 4274 3266 4290
rect 3332 4284 3351 4287
rect 2973 4262 3071 4264
rect 3098 4262 3266 4274
rect 3281 4264 3297 4278
rect 3332 4265 3354 4284
rect 3364 4278 3380 4279
rect 3363 4276 3380 4278
rect 3364 4271 3380 4276
rect 3354 4264 3360 4265
rect 3363 4264 3392 4271
rect 3281 4263 3392 4264
rect 3281 4262 3398 4263
rect 2957 4254 3008 4262
rect 3055 4254 3089 4262
rect 2957 4242 2982 4254
rect 2989 4242 3008 4254
rect 3062 4252 3089 4254
rect 3098 4252 3319 4262
rect 3354 4259 3360 4262
rect 3062 4248 3319 4252
rect 2957 4234 3008 4242
rect 3055 4234 3319 4248
rect 3363 4254 3398 4262
rect 2909 4186 2928 4220
rect 2973 4226 3002 4234
rect 2973 4220 2990 4226
rect 2973 4218 3007 4220
rect 3055 4218 3071 4234
rect 3072 4224 3280 4234
rect 3281 4224 3297 4234
rect 3345 4230 3360 4245
rect 3363 4242 3364 4254
rect 3371 4242 3398 4254
rect 3363 4234 3398 4242
rect 3363 4233 3392 4234
rect 3083 4220 3297 4224
rect 3098 4218 3297 4220
rect 3332 4220 3345 4230
rect 3363 4220 3380 4233
rect 3332 4218 3380 4220
rect 2974 4214 3007 4218
rect 2970 4212 3007 4214
rect 2970 4211 3037 4212
rect 2970 4206 3001 4211
rect 3007 4206 3037 4211
rect 2970 4202 3037 4206
rect 2943 4199 3037 4202
rect 2943 4192 2992 4199
rect 2943 4186 2973 4192
rect 2992 4187 2997 4192
rect 2909 4170 2989 4186
rect 3001 4178 3037 4199
rect 3098 4194 3287 4218
rect 3332 4217 3379 4218
rect 3345 4212 3379 4217
rect 3113 4191 3287 4194
rect 3106 4188 3287 4191
rect 3315 4211 3379 4212
rect 2909 4168 2928 4170
rect 2943 4168 2977 4170
rect 2909 4152 2989 4168
rect 2909 4146 2928 4152
rect 2625 4120 2728 4130
rect 2579 4118 2728 4120
rect 2749 4118 2784 4130
rect 2418 4116 2580 4118
rect 2430 4096 2449 4116
rect 2464 4114 2494 4116
rect 2313 4088 2354 4096
rect 2436 4092 2449 4096
rect 2501 4100 2580 4116
rect 2612 4116 2784 4118
rect 2612 4100 2691 4116
rect 2698 4114 2728 4116
rect 2276 4078 2305 4088
rect 2319 4078 2348 4088
rect 2363 4078 2393 4092
rect 2436 4078 2479 4092
rect 2501 4088 2691 4100
rect 2756 4096 2762 4116
rect 2486 4078 2516 4088
rect 2517 4078 2675 4088
rect 2679 4078 2709 4088
rect 2713 4078 2743 4092
rect 2771 4078 2784 4116
rect 2856 4130 2885 4146
rect 2899 4130 2928 4146
rect 2943 4136 2973 4152
rect 3001 4130 3007 4178
rect 3010 4172 3029 4178
rect 3044 4172 3074 4180
rect 3010 4164 3074 4172
rect 3010 4148 3090 4164
rect 3106 4157 3168 4188
rect 3184 4157 3246 4188
rect 3315 4186 3364 4211
rect 3379 4186 3409 4202
rect 3278 4172 3308 4180
rect 3315 4178 3425 4186
rect 3278 4164 3323 4172
rect 3010 4146 3029 4148
rect 3044 4146 3090 4148
rect 3010 4130 3090 4146
rect 3117 4144 3152 4157
rect 3193 4154 3230 4157
rect 3193 4152 3235 4154
rect 3122 4141 3152 4144
rect 3131 4137 3138 4141
rect 3138 4136 3139 4137
rect 3097 4130 3107 4136
rect 2856 4122 2891 4130
rect 2856 4096 2857 4122
rect 2864 4096 2891 4122
rect 2799 4078 2829 4092
rect 2856 4088 2891 4096
rect 2893 4122 2934 4130
rect 2893 4096 2908 4122
rect 2915 4096 2934 4122
rect 2998 4118 3029 4130
rect 3044 4118 3147 4130
rect 3159 4120 3185 4146
rect 3200 4141 3230 4152
rect 3262 4148 3324 4164
rect 3262 4146 3308 4148
rect 3262 4130 3324 4146
rect 3336 4130 3342 4178
rect 3345 4170 3425 4178
rect 3345 4168 3364 4170
rect 3379 4168 3413 4170
rect 3345 4152 3425 4168
rect 3345 4130 3364 4152
rect 3379 4136 3409 4152
rect 3437 4146 3443 4220
rect 3446 4146 3465 4290
rect 3480 4146 3486 4290
rect 3495 4220 3508 4290
rect 3560 4286 3582 4290
rect 3553 4264 3582 4278
rect 3635 4264 3651 4278
rect 3689 4274 3695 4276
rect 3702 4274 3810 4290
rect 3817 4274 3823 4276
rect 3831 4274 3846 4290
rect 3912 4284 3931 4287
rect 3553 4262 3651 4264
rect 3678 4262 3846 4274
rect 3861 4264 3877 4278
rect 3912 4265 3934 4284
rect 3944 4278 3960 4279
rect 3943 4276 3960 4278
rect 3944 4271 3960 4276
rect 3934 4264 3940 4265
rect 3943 4264 3972 4271
rect 3861 4263 3972 4264
rect 3861 4262 3978 4263
rect 3537 4254 3588 4262
rect 3635 4254 3669 4262
rect 3537 4242 3562 4254
rect 3569 4242 3588 4254
rect 3642 4252 3669 4254
rect 3678 4252 3899 4262
rect 3934 4259 3940 4262
rect 3642 4248 3899 4252
rect 3537 4234 3588 4242
rect 3635 4234 3899 4248
rect 3943 4254 3978 4262
rect 3489 4186 3508 4220
rect 3553 4226 3582 4234
rect 3553 4220 3570 4226
rect 3553 4218 3587 4220
rect 3635 4218 3651 4234
rect 3652 4224 3860 4234
rect 3861 4224 3877 4234
rect 3925 4230 3940 4245
rect 3943 4242 3944 4254
rect 3951 4242 3978 4254
rect 3943 4234 3978 4242
rect 3943 4233 3972 4234
rect 3663 4220 3877 4224
rect 3678 4218 3877 4220
rect 3912 4220 3925 4230
rect 3943 4220 3960 4233
rect 3912 4218 3960 4220
rect 3554 4214 3587 4218
rect 3550 4212 3587 4214
rect 3550 4211 3617 4212
rect 3550 4206 3581 4211
rect 3587 4206 3617 4211
rect 3550 4202 3617 4206
rect 3523 4199 3617 4202
rect 3523 4192 3572 4199
rect 3523 4186 3553 4192
rect 3572 4187 3577 4192
rect 3489 4170 3569 4186
rect 3581 4178 3617 4199
rect 3678 4194 3867 4218
rect 3912 4217 3959 4218
rect 3925 4212 3959 4217
rect 3693 4191 3867 4194
rect 3686 4188 3867 4191
rect 3895 4211 3959 4212
rect 3489 4168 3508 4170
rect 3523 4168 3557 4170
rect 3489 4152 3569 4168
rect 3489 4146 3508 4152
rect 3205 4120 3308 4130
rect 3159 4118 3308 4120
rect 3329 4118 3364 4130
rect 2998 4116 3160 4118
rect 3010 4096 3029 4116
rect 3044 4114 3074 4116
rect 2893 4088 2934 4096
rect 3016 4092 3029 4096
rect 3081 4100 3160 4116
rect 3192 4116 3364 4118
rect 3192 4100 3271 4116
rect 3278 4114 3308 4116
rect 2856 4078 2885 4088
rect 2899 4078 2928 4088
rect 2943 4078 2973 4092
rect 3016 4078 3059 4092
rect 3081 4088 3271 4100
rect 3336 4096 3342 4116
rect 3066 4078 3096 4088
rect 3097 4078 3255 4088
rect 3259 4078 3289 4088
rect 3293 4078 3323 4092
rect 3351 4078 3364 4116
rect 3436 4130 3465 4146
rect 3479 4130 3508 4146
rect 3523 4136 3553 4152
rect 3581 4130 3587 4178
rect 3590 4172 3609 4178
rect 3624 4172 3654 4180
rect 3590 4164 3654 4172
rect 3590 4148 3670 4164
rect 3686 4157 3748 4188
rect 3764 4157 3826 4188
rect 3895 4186 3944 4211
rect 3959 4186 3989 4202
rect 3858 4172 3888 4180
rect 3895 4178 4005 4186
rect 3858 4164 3903 4172
rect 3590 4146 3609 4148
rect 3624 4146 3670 4148
rect 3590 4130 3670 4146
rect 3697 4144 3732 4157
rect 3773 4154 3810 4157
rect 3773 4152 3815 4154
rect 3702 4141 3732 4144
rect 3711 4137 3718 4141
rect 3718 4136 3719 4137
rect 3677 4130 3687 4136
rect 3436 4122 3471 4130
rect 3436 4096 3437 4122
rect 3444 4096 3471 4122
rect 3379 4078 3409 4092
rect 3436 4088 3471 4096
rect 3473 4122 3514 4130
rect 3473 4096 3488 4122
rect 3495 4096 3514 4122
rect 3578 4118 3609 4130
rect 3624 4118 3727 4130
rect 3739 4120 3765 4146
rect 3780 4141 3810 4152
rect 3842 4148 3904 4164
rect 3842 4146 3888 4148
rect 3842 4130 3904 4146
rect 3916 4130 3922 4178
rect 3925 4170 4005 4178
rect 3925 4168 3944 4170
rect 3959 4168 3993 4170
rect 3925 4152 4005 4168
rect 3925 4130 3944 4152
rect 3959 4136 3989 4152
rect 4017 4146 4023 4220
rect 4026 4146 4045 4290
rect 4060 4146 4066 4290
rect 4075 4220 4088 4290
rect 4140 4286 4162 4290
rect 4133 4264 4162 4278
rect 4215 4264 4231 4278
rect 4269 4274 4275 4276
rect 4282 4274 4390 4290
rect 4397 4274 4403 4276
rect 4411 4274 4426 4290
rect 4492 4284 4511 4287
rect 4133 4262 4231 4264
rect 4258 4262 4426 4274
rect 4441 4264 4457 4278
rect 4492 4265 4514 4284
rect 4524 4278 4540 4279
rect 4523 4276 4540 4278
rect 4524 4271 4540 4276
rect 4514 4264 4520 4265
rect 4523 4264 4552 4271
rect 4441 4263 4552 4264
rect 4441 4262 4558 4263
rect 4117 4254 4168 4262
rect 4215 4254 4249 4262
rect 4117 4242 4142 4254
rect 4149 4242 4168 4254
rect 4222 4252 4249 4254
rect 4258 4252 4479 4262
rect 4514 4259 4520 4262
rect 4222 4248 4479 4252
rect 4117 4234 4168 4242
rect 4215 4234 4479 4248
rect 4523 4254 4558 4262
rect 4069 4186 4088 4220
rect 4133 4226 4162 4234
rect 4133 4220 4150 4226
rect 4133 4218 4167 4220
rect 4215 4218 4231 4234
rect 4232 4224 4440 4234
rect 4441 4224 4457 4234
rect 4505 4230 4520 4245
rect 4523 4242 4524 4254
rect 4531 4242 4558 4254
rect 4523 4234 4558 4242
rect 4523 4233 4552 4234
rect 4243 4220 4457 4224
rect 4258 4218 4457 4220
rect 4492 4220 4505 4230
rect 4523 4220 4540 4233
rect 4492 4218 4540 4220
rect 4134 4214 4167 4218
rect 4130 4212 4167 4214
rect 4130 4211 4197 4212
rect 4130 4206 4161 4211
rect 4167 4206 4197 4211
rect 4130 4202 4197 4206
rect 4103 4199 4197 4202
rect 4103 4192 4152 4199
rect 4103 4186 4133 4192
rect 4152 4187 4157 4192
rect 4069 4170 4149 4186
rect 4161 4178 4197 4199
rect 4258 4194 4447 4218
rect 4492 4217 4539 4218
rect 4505 4212 4539 4217
rect 4273 4191 4447 4194
rect 4266 4188 4447 4191
rect 4475 4211 4539 4212
rect 4069 4168 4088 4170
rect 4103 4168 4137 4170
rect 4069 4152 4149 4168
rect 4069 4146 4088 4152
rect 3785 4120 3888 4130
rect 3739 4118 3888 4120
rect 3909 4118 3944 4130
rect 3578 4116 3740 4118
rect 3590 4096 3609 4116
rect 3624 4114 3654 4116
rect 3473 4088 3514 4096
rect 3596 4092 3609 4096
rect 3661 4100 3740 4116
rect 3772 4116 3944 4118
rect 3772 4100 3851 4116
rect 3858 4114 3888 4116
rect 3436 4078 3465 4088
rect 3479 4078 3508 4088
rect 3523 4078 3553 4092
rect 3596 4078 3639 4092
rect 3661 4088 3851 4100
rect 3916 4096 3922 4116
rect 3646 4078 3676 4088
rect 3677 4078 3835 4088
rect 3839 4078 3869 4088
rect 3873 4078 3903 4092
rect 3931 4078 3944 4116
rect 4016 4130 4045 4146
rect 4059 4130 4088 4146
rect 4103 4136 4133 4152
rect 4161 4130 4167 4178
rect 4170 4172 4189 4178
rect 4204 4172 4234 4180
rect 4170 4164 4234 4172
rect 4170 4148 4250 4164
rect 4266 4157 4328 4188
rect 4344 4157 4406 4188
rect 4475 4186 4524 4211
rect 4539 4186 4569 4202
rect 4438 4172 4468 4180
rect 4475 4178 4585 4186
rect 4438 4164 4483 4172
rect 4170 4146 4189 4148
rect 4204 4146 4250 4148
rect 4170 4130 4250 4146
rect 4277 4144 4312 4157
rect 4353 4154 4390 4157
rect 4353 4152 4395 4154
rect 4282 4141 4312 4144
rect 4291 4137 4298 4141
rect 4298 4136 4299 4137
rect 4257 4130 4267 4136
rect 4016 4122 4051 4130
rect 4016 4096 4017 4122
rect 4024 4096 4051 4122
rect 3959 4078 3989 4092
rect 4016 4088 4051 4096
rect 4053 4122 4094 4130
rect 4053 4096 4068 4122
rect 4075 4096 4094 4122
rect 4158 4118 4189 4130
rect 4204 4118 4307 4130
rect 4319 4120 4345 4146
rect 4360 4141 4390 4152
rect 4422 4148 4484 4164
rect 4422 4146 4468 4148
rect 4422 4130 4484 4146
rect 4496 4130 4502 4178
rect 4505 4170 4585 4178
rect 4505 4168 4524 4170
rect 4539 4168 4573 4170
rect 4505 4152 4585 4168
rect 4505 4130 4524 4152
rect 4539 4136 4569 4152
rect 4597 4146 4603 4220
rect 4606 4146 4625 4290
rect 4640 4146 4646 4290
rect 4655 4220 4668 4290
rect 4720 4286 4742 4290
rect 4713 4264 4742 4278
rect 4795 4264 4811 4278
rect 4849 4274 4855 4276
rect 4862 4274 4970 4290
rect 4977 4274 4983 4276
rect 4991 4274 5006 4290
rect 5072 4284 5091 4287
rect 4713 4262 4811 4264
rect 4838 4262 5006 4274
rect 5021 4264 5037 4278
rect 5072 4265 5094 4284
rect 5104 4278 5120 4279
rect 5103 4276 5120 4278
rect 5104 4271 5120 4276
rect 5094 4264 5100 4265
rect 5103 4264 5132 4271
rect 5021 4263 5132 4264
rect 5021 4262 5138 4263
rect 4697 4254 4748 4262
rect 4795 4254 4829 4262
rect 4697 4242 4722 4254
rect 4729 4242 4748 4254
rect 4802 4252 4829 4254
rect 4838 4252 5059 4262
rect 5094 4259 5100 4262
rect 4802 4248 5059 4252
rect 4697 4234 4748 4242
rect 4795 4234 5059 4248
rect 5103 4254 5138 4262
rect 4649 4186 4668 4220
rect 4713 4226 4742 4234
rect 4713 4220 4730 4226
rect 4713 4218 4747 4220
rect 4795 4218 4811 4234
rect 4812 4224 5020 4234
rect 5021 4224 5037 4234
rect 5085 4230 5100 4245
rect 5103 4242 5104 4254
rect 5111 4242 5138 4254
rect 5103 4234 5138 4242
rect 5103 4233 5132 4234
rect 4823 4220 5037 4224
rect 4838 4218 5037 4220
rect 5072 4220 5085 4230
rect 5103 4220 5120 4233
rect 5072 4218 5120 4220
rect 4714 4214 4747 4218
rect 4710 4212 4747 4214
rect 4710 4211 4777 4212
rect 4710 4206 4741 4211
rect 4747 4206 4777 4211
rect 4710 4202 4777 4206
rect 4683 4199 4777 4202
rect 4683 4192 4732 4199
rect 4683 4186 4713 4192
rect 4732 4187 4737 4192
rect 4649 4170 4729 4186
rect 4741 4178 4777 4199
rect 4838 4194 5027 4218
rect 5072 4217 5119 4218
rect 5085 4212 5119 4217
rect 4853 4191 5027 4194
rect 4846 4188 5027 4191
rect 5055 4211 5119 4212
rect 4649 4168 4668 4170
rect 4683 4168 4717 4170
rect 4649 4152 4729 4168
rect 4649 4146 4668 4152
rect 4365 4120 4468 4130
rect 4319 4118 4468 4120
rect 4489 4118 4524 4130
rect 4158 4116 4320 4118
rect 4170 4096 4189 4116
rect 4204 4114 4234 4116
rect 4053 4088 4094 4096
rect 4176 4092 4189 4096
rect 4241 4100 4320 4116
rect 4352 4116 4524 4118
rect 4352 4100 4431 4116
rect 4438 4114 4468 4116
rect 4016 4078 4045 4088
rect 4059 4078 4088 4088
rect 4103 4078 4133 4092
rect 4176 4078 4219 4092
rect 4241 4088 4431 4100
rect 4496 4096 4502 4116
rect 4226 4078 4256 4088
rect 4257 4078 4415 4088
rect 4419 4078 4449 4088
rect 4453 4078 4483 4092
rect 4511 4078 4524 4116
rect 4596 4130 4625 4146
rect 4639 4130 4668 4146
rect 4683 4136 4713 4152
rect 4741 4130 4747 4178
rect 4750 4172 4769 4178
rect 4784 4172 4814 4180
rect 4750 4164 4814 4172
rect 4750 4148 4830 4164
rect 4846 4157 4908 4188
rect 4924 4157 4986 4188
rect 5055 4186 5104 4211
rect 5119 4186 5149 4202
rect 5018 4172 5048 4180
rect 5055 4178 5165 4186
rect 5018 4164 5063 4172
rect 4750 4146 4769 4148
rect 4784 4146 4830 4148
rect 4750 4130 4830 4146
rect 4857 4144 4892 4157
rect 4933 4154 4970 4157
rect 4933 4152 4975 4154
rect 4862 4141 4892 4144
rect 4871 4137 4878 4141
rect 4878 4136 4879 4137
rect 4837 4130 4847 4136
rect 4596 4122 4631 4130
rect 4596 4096 4597 4122
rect 4604 4096 4631 4122
rect 4539 4078 4569 4092
rect 4596 4088 4631 4096
rect 4633 4122 4674 4130
rect 4633 4096 4648 4122
rect 4655 4096 4674 4122
rect 4738 4118 4769 4130
rect 4784 4118 4887 4130
rect 4899 4120 4925 4146
rect 4940 4141 4970 4152
rect 5002 4148 5064 4164
rect 5002 4146 5048 4148
rect 5002 4130 5064 4146
rect 5076 4130 5082 4178
rect 5085 4170 5165 4178
rect 5085 4168 5104 4170
rect 5119 4168 5153 4170
rect 5085 4152 5165 4168
rect 5085 4130 5104 4152
rect 5119 4136 5149 4152
rect 5177 4146 5183 4220
rect 5186 4146 5205 4290
rect 5220 4146 5226 4290
rect 5235 4220 5248 4290
rect 5300 4286 5322 4290
rect 5293 4264 5322 4278
rect 5375 4264 5391 4278
rect 5429 4274 5435 4276
rect 5442 4274 5550 4290
rect 5557 4274 5563 4276
rect 5571 4274 5586 4290
rect 5652 4284 5671 4287
rect 5293 4262 5391 4264
rect 5418 4262 5586 4274
rect 5601 4264 5617 4278
rect 5652 4265 5674 4284
rect 5684 4278 5700 4279
rect 5683 4276 5700 4278
rect 5684 4271 5700 4276
rect 5674 4264 5680 4265
rect 5683 4264 5712 4271
rect 5601 4263 5712 4264
rect 5601 4262 5718 4263
rect 5277 4254 5328 4262
rect 5375 4254 5409 4262
rect 5277 4242 5302 4254
rect 5309 4242 5328 4254
rect 5382 4252 5409 4254
rect 5418 4252 5639 4262
rect 5674 4259 5680 4262
rect 5382 4248 5639 4252
rect 5277 4234 5328 4242
rect 5375 4234 5639 4248
rect 5683 4254 5718 4262
rect 5229 4186 5248 4220
rect 5293 4226 5322 4234
rect 5293 4220 5310 4226
rect 5293 4218 5327 4220
rect 5375 4218 5391 4234
rect 5392 4224 5600 4234
rect 5601 4224 5617 4234
rect 5665 4230 5680 4245
rect 5683 4242 5684 4254
rect 5691 4242 5718 4254
rect 5683 4234 5718 4242
rect 5683 4233 5712 4234
rect 5403 4220 5617 4224
rect 5418 4218 5617 4220
rect 5652 4220 5665 4230
rect 5683 4220 5700 4233
rect 5652 4218 5700 4220
rect 5294 4214 5327 4218
rect 5290 4212 5327 4214
rect 5290 4211 5357 4212
rect 5290 4206 5321 4211
rect 5327 4206 5357 4211
rect 5290 4202 5357 4206
rect 5263 4199 5357 4202
rect 5263 4192 5312 4199
rect 5263 4186 5293 4192
rect 5312 4187 5317 4192
rect 5229 4170 5309 4186
rect 5321 4178 5357 4199
rect 5418 4194 5607 4218
rect 5652 4217 5699 4218
rect 5665 4212 5699 4217
rect 5433 4191 5607 4194
rect 5426 4188 5607 4191
rect 5635 4211 5699 4212
rect 5229 4168 5248 4170
rect 5263 4168 5297 4170
rect 5229 4152 5309 4168
rect 5229 4146 5248 4152
rect 4945 4120 5048 4130
rect 4899 4118 5048 4120
rect 5069 4118 5104 4130
rect 4738 4116 4900 4118
rect 4750 4096 4769 4116
rect 4784 4114 4814 4116
rect 4633 4088 4674 4096
rect 4756 4092 4769 4096
rect 4821 4100 4900 4116
rect 4932 4116 5104 4118
rect 4932 4100 5011 4116
rect 5018 4114 5048 4116
rect 4596 4078 4625 4088
rect 4639 4078 4668 4088
rect 4683 4078 4713 4092
rect 4756 4078 4799 4092
rect 4821 4088 5011 4100
rect 5076 4096 5082 4116
rect 4806 4078 4836 4088
rect 4837 4078 4995 4088
rect 4999 4078 5029 4088
rect 5033 4078 5063 4092
rect 5091 4078 5104 4116
rect 5176 4130 5205 4146
rect 5219 4130 5248 4146
rect 5263 4136 5293 4152
rect 5321 4130 5327 4178
rect 5330 4172 5349 4178
rect 5364 4172 5394 4180
rect 5330 4164 5394 4172
rect 5330 4148 5410 4164
rect 5426 4157 5488 4188
rect 5504 4157 5566 4188
rect 5635 4186 5684 4211
rect 5699 4186 5729 4202
rect 5598 4172 5628 4180
rect 5635 4178 5745 4186
rect 5598 4164 5643 4172
rect 5330 4146 5349 4148
rect 5364 4146 5410 4148
rect 5330 4130 5410 4146
rect 5437 4144 5472 4157
rect 5513 4154 5550 4157
rect 5513 4152 5555 4154
rect 5442 4141 5472 4144
rect 5451 4137 5458 4141
rect 5458 4136 5459 4137
rect 5417 4130 5427 4136
rect 5176 4122 5211 4130
rect 5176 4096 5177 4122
rect 5184 4096 5211 4122
rect 5119 4078 5149 4092
rect 5176 4088 5211 4096
rect 5213 4122 5254 4130
rect 5213 4096 5228 4122
rect 5235 4096 5254 4122
rect 5318 4118 5349 4130
rect 5364 4118 5467 4130
rect 5479 4120 5505 4146
rect 5520 4141 5550 4152
rect 5582 4148 5644 4164
rect 5582 4146 5628 4148
rect 5582 4130 5644 4146
rect 5656 4130 5662 4178
rect 5665 4170 5745 4178
rect 5665 4168 5684 4170
rect 5699 4168 5733 4170
rect 5665 4152 5745 4168
rect 5665 4130 5684 4152
rect 5699 4136 5729 4152
rect 5757 4146 5763 4220
rect 5766 4146 5785 4290
rect 5800 4146 5806 4290
rect 5815 4220 5828 4290
rect 5880 4286 5902 4290
rect 5873 4264 5902 4278
rect 5955 4264 5971 4278
rect 6009 4274 6015 4276
rect 6022 4274 6130 4290
rect 6137 4274 6143 4276
rect 6151 4274 6166 4290
rect 6232 4284 6251 4287
rect 5873 4262 5971 4264
rect 5998 4262 6166 4274
rect 6181 4264 6197 4278
rect 6232 4265 6254 4284
rect 6264 4278 6280 4279
rect 6263 4276 6280 4278
rect 6264 4271 6280 4276
rect 6254 4264 6260 4265
rect 6263 4264 6292 4271
rect 6181 4263 6292 4264
rect 6181 4262 6298 4263
rect 5857 4254 5908 4262
rect 5955 4254 5989 4262
rect 5857 4242 5882 4254
rect 5889 4242 5908 4254
rect 5962 4252 5989 4254
rect 5998 4252 6219 4262
rect 6254 4259 6260 4262
rect 5962 4248 6219 4252
rect 5857 4234 5908 4242
rect 5955 4234 6219 4248
rect 6263 4254 6298 4262
rect 5809 4186 5828 4220
rect 5873 4226 5902 4234
rect 5873 4220 5890 4226
rect 5873 4218 5907 4220
rect 5955 4218 5971 4234
rect 5972 4224 6180 4234
rect 6181 4224 6197 4234
rect 6245 4230 6260 4245
rect 6263 4242 6264 4254
rect 6271 4242 6298 4254
rect 6263 4234 6298 4242
rect 6263 4233 6292 4234
rect 5983 4220 6197 4224
rect 5998 4218 6197 4220
rect 6232 4220 6245 4230
rect 6263 4220 6280 4233
rect 6232 4218 6280 4220
rect 5874 4214 5907 4218
rect 5870 4212 5907 4214
rect 5870 4211 5937 4212
rect 5870 4206 5901 4211
rect 5907 4206 5937 4211
rect 5870 4202 5937 4206
rect 5843 4199 5937 4202
rect 5843 4192 5892 4199
rect 5843 4186 5873 4192
rect 5892 4187 5897 4192
rect 5809 4170 5889 4186
rect 5901 4178 5937 4199
rect 5998 4194 6187 4218
rect 6232 4217 6279 4218
rect 6245 4212 6279 4217
rect 6013 4191 6187 4194
rect 6006 4188 6187 4191
rect 6215 4211 6279 4212
rect 5809 4168 5828 4170
rect 5843 4168 5877 4170
rect 5809 4152 5889 4168
rect 5809 4146 5828 4152
rect 5525 4120 5628 4130
rect 5479 4118 5628 4120
rect 5649 4118 5684 4130
rect 5318 4116 5480 4118
rect 5330 4096 5349 4116
rect 5364 4114 5394 4116
rect 5213 4088 5254 4096
rect 5336 4092 5349 4096
rect 5401 4100 5480 4116
rect 5512 4116 5684 4118
rect 5512 4100 5591 4116
rect 5598 4114 5628 4116
rect 5176 4078 5205 4088
rect 5219 4078 5248 4088
rect 5263 4078 5293 4092
rect 5336 4078 5379 4092
rect 5401 4088 5591 4100
rect 5656 4096 5662 4116
rect 5386 4078 5416 4088
rect 5417 4078 5575 4088
rect 5579 4078 5609 4088
rect 5613 4078 5643 4092
rect 5671 4078 5684 4116
rect 5756 4130 5785 4146
rect 5799 4130 5828 4146
rect 5843 4136 5873 4152
rect 5901 4130 5907 4178
rect 5910 4172 5929 4178
rect 5944 4172 5974 4180
rect 5910 4164 5974 4172
rect 5910 4148 5990 4164
rect 6006 4157 6068 4188
rect 6084 4157 6146 4188
rect 6215 4186 6264 4211
rect 6279 4186 6309 4202
rect 6178 4172 6208 4180
rect 6215 4178 6325 4186
rect 6178 4164 6223 4172
rect 5910 4146 5929 4148
rect 5944 4146 5990 4148
rect 5910 4130 5990 4146
rect 6017 4144 6052 4157
rect 6093 4154 6130 4157
rect 6093 4152 6135 4154
rect 6022 4141 6052 4144
rect 6031 4137 6038 4141
rect 6038 4136 6039 4137
rect 5997 4130 6007 4136
rect 5756 4122 5791 4130
rect 5756 4096 5757 4122
rect 5764 4096 5791 4122
rect 5699 4078 5729 4092
rect 5756 4088 5791 4096
rect 5793 4122 5834 4130
rect 5793 4096 5808 4122
rect 5815 4096 5834 4122
rect 5898 4118 5929 4130
rect 5944 4118 6047 4130
rect 6059 4120 6085 4146
rect 6100 4141 6130 4152
rect 6162 4148 6224 4164
rect 6162 4146 6208 4148
rect 6162 4130 6224 4146
rect 6236 4130 6242 4178
rect 6245 4170 6325 4178
rect 6245 4168 6264 4170
rect 6279 4168 6313 4170
rect 6245 4152 6325 4168
rect 6245 4130 6264 4152
rect 6279 4136 6309 4152
rect 6337 4146 6343 4220
rect 6346 4146 6365 4290
rect 6380 4146 6386 4290
rect 6395 4220 6408 4290
rect 6460 4286 6482 4290
rect 6453 4264 6482 4278
rect 6535 4264 6551 4278
rect 6589 4274 6595 4276
rect 6602 4274 6710 4290
rect 6717 4274 6723 4276
rect 6731 4274 6746 4290
rect 6812 4284 6831 4287
rect 6453 4262 6551 4264
rect 6578 4262 6746 4274
rect 6761 4264 6777 4278
rect 6812 4265 6834 4284
rect 6844 4278 6860 4279
rect 6843 4276 6860 4278
rect 6844 4271 6860 4276
rect 6834 4264 6840 4265
rect 6843 4264 6872 4271
rect 6761 4263 6872 4264
rect 6761 4262 6878 4263
rect 6437 4254 6488 4262
rect 6535 4254 6569 4262
rect 6437 4242 6462 4254
rect 6469 4242 6488 4254
rect 6542 4252 6569 4254
rect 6578 4252 6799 4262
rect 6834 4259 6840 4262
rect 6542 4248 6799 4252
rect 6437 4234 6488 4242
rect 6535 4234 6799 4248
rect 6843 4254 6878 4262
rect 6389 4186 6408 4220
rect 6453 4226 6482 4234
rect 6453 4220 6470 4226
rect 6453 4218 6487 4220
rect 6535 4218 6551 4234
rect 6552 4224 6760 4234
rect 6761 4224 6777 4234
rect 6825 4230 6840 4245
rect 6843 4242 6844 4254
rect 6851 4242 6878 4254
rect 6843 4234 6878 4242
rect 6843 4233 6872 4234
rect 6563 4220 6777 4224
rect 6578 4218 6777 4220
rect 6812 4220 6825 4230
rect 6843 4220 6860 4233
rect 6812 4218 6860 4220
rect 6454 4214 6487 4218
rect 6450 4212 6487 4214
rect 6450 4211 6517 4212
rect 6450 4206 6481 4211
rect 6487 4206 6517 4211
rect 6450 4202 6517 4206
rect 6423 4199 6517 4202
rect 6423 4192 6472 4199
rect 6423 4186 6453 4192
rect 6472 4187 6477 4192
rect 6389 4170 6469 4186
rect 6481 4178 6517 4199
rect 6578 4194 6767 4218
rect 6812 4217 6859 4218
rect 6825 4212 6859 4217
rect 6593 4191 6767 4194
rect 6586 4188 6767 4191
rect 6795 4211 6859 4212
rect 6389 4168 6408 4170
rect 6423 4168 6457 4170
rect 6389 4152 6469 4168
rect 6389 4146 6408 4152
rect 6105 4120 6208 4130
rect 6059 4118 6208 4120
rect 6229 4118 6264 4130
rect 5898 4116 6060 4118
rect 5910 4096 5929 4116
rect 5944 4114 5974 4116
rect 5793 4088 5834 4096
rect 5916 4092 5929 4096
rect 5981 4100 6060 4116
rect 6092 4116 6264 4118
rect 6092 4100 6171 4116
rect 6178 4114 6208 4116
rect 5756 4078 5785 4088
rect 5799 4078 5828 4088
rect 5843 4078 5873 4092
rect 5916 4078 5959 4092
rect 5981 4088 6171 4100
rect 6236 4096 6242 4116
rect 5966 4078 5996 4088
rect 5997 4078 6155 4088
rect 6159 4078 6189 4088
rect 6193 4078 6223 4092
rect 6251 4078 6264 4116
rect 6336 4130 6365 4146
rect 6379 4130 6408 4146
rect 6423 4136 6453 4152
rect 6481 4130 6487 4178
rect 6490 4172 6509 4178
rect 6524 4172 6554 4180
rect 6490 4164 6554 4172
rect 6490 4148 6570 4164
rect 6586 4157 6648 4188
rect 6664 4157 6726 4188
rect 6795 4186 6844 4211
rect 6859 4186 6889 4202
rect 6758 4172 6788 4180
rect 6795 4178 6905 4186
rect 6758 4164 6803 4172
rect 6490 4146 6509 4148
rect 6524 4146 6570 4148
rect 6490 4130 6570 4146
rect 6597 4144 6632 4157
rect 6673 4154 6710 4157
rect 6673 4152 6715 4154
rect 6602 4141 6632 4144
rect 6611 4137 6618 4141
rect 6618 4136 6619 4137
rect 6577 4130 6587 4136
rect 6336 4122 6371 4130
rect 6336 4096 6337 4122
rect 6344 4096 6371 4122
rect 6279 4078 6309 4092
rect 6336 4088 6371 4096
rect 6373 4122 6414 4130
rect 6373 4096 6388 4122
rect 6395 4096 6414 4122
rect 6478 4118 6509 4130
rect 6524 4118 6627 4130
rect 6639 4120 6665 4146
rect 6680 4141 6710 4152
rect 6742 4148 6804 4164
rect 6742 4146 6788 4148
rect 6742 4130 6804 4146
rect 6816 4130 6822 4178
rect 6825 4170 6905 4178
rect 6825 4168 6844 4170
rect 6859 4168 6893 4170
rect 6825 4152 6905 4168
rect 6825 4130 6844 4152
rect 6859 4136 6889 4152
rect 6917 4146 6923 4220
rect 6926 4146 6945 4290
rect 6960 4146 6966 4290
rect 6975 4220 6988 4290
rect 7040 4286 7062 4290
rect 7033 4264 7062 4278
rect 7115 4264 7131 4278
rect 7169 4274 7175 4276
rect 7182 4274 7290 4290
rect 7297 4274 7303 4276
rect 7311 4274 7326 4290
rect 7392 4284 7411 4287
rect 7033 4262 7131 4264
rect 7158 4262 7326 4274
rect 7341 4264 7357 4278
rect 7392 4265 7414 4284
rect 7424 4278 7440 4279
rect 7423 4276 7440 4278
rect 7424 4271 7440 4276
rect 7414 4264 7420 4265
rect 7423 4264 7452 4271
rect 7341 4263 7452 4264
rect 7341 4262 7458 4263
rect 7017 4254 7068 4262
rect 7115 4254 7149 4262
rect 7017 4242 7042 4254
rect 7049 4242 7068 4254
rect 7122 4252 7149 4254
rect 7158 4252 7379 4262
rect 7414 4259 7420 4262
rect 7122 4248 7379 4252
rect 7017 4234 7068 4242
rect 7115 4234 7379 4248
rect 7423 4254 7458 4262
rect 6969 4186 6988 4220
rect 7033 4226 7062 4234
rect 7033 4220 7050 4226
rect 7033 4218 7067 4220
rect 7115 4218 7131 4234
rect 7132 4224 7340 4234
rect 7341 4224 7357 4234
rect 7405 4230 7420 4245
rect 7423 4242 7424 4254
rect 7431 4242 7458 4254
rect 7423 4234 7458 4242
rect 7423 4233 7452 4234
rect 7143 4220 7357 4224
rect 7158 4218 7357 4220
rect 7392 4220 7405 4230
rect 7423 4220 7440 4233
rect 7392 4218 7440 4220
rect 7034 4214 7067 4218
rect 7030 4212 7067 4214
rect 7030 4211 7097 4212
rect 7030 4206 7061 4211
rect 7067 4206 7097 4211
rect 7030 4202 7097 4206
rect 7003 4199 7097 4202
rect 7003 4192 7052 4199
rect 7003 4186 7033 4192
rect 7052 4187 7057 4192
rect 6969 4170 7049 4186
rect 7061 4178 7097 4199
rect 7158 4194 7347 4218
rect 7392 4217 7439 4218
rect 7405 4212 7439 4217
rect 7173 4191 7347 4194
rect 7166 4188 7347 4191
rect 7375 4211 7439 4212
rect 6969 4168 6988 4170
rect 7003 4168 7037 4170
rect 6969 4152 7049 4168
rect 6969 4146 6988 4152
rect 6685 4120 6788 4130
rect 6639 4118 6788 4120
rect 6809 4118 6844 4130
rect 6478 4116 6640 4118
rect 6490 4096 6509 4116
rect 6524 4114 6554 4116
rect 6373 4088 6414 4096
rect 6496 4092 6509 4096
rect 6561 4100 6640 4116
rect 6672 4116 6844 4118
rect 6672 4100 6751 4116
rect 6758 4114 6788 4116
rect 6336 4078 6365 4088
rect 6379 4078 6408 4088
rect 6423 4078 6453 4092
rect 6496 4078 6539 4092
rect 6561 4088 6751 4100
rect 6816 4096 6822 4116
rect 6546 4078 6576 4088
rect 6577 4078 6735 4088
rect 6739 4078 6769 4088
rect 6773 4078 6803 4092
rect 6831 4078 6844 4116
rect 6916 4130 6945 4146
rect 6959 4130 6988 4146
rect 7003 4136 7033 4152
rect 7061 4130 7067 4178
rect 7070 4172 7089 4178
rect 7104 4172 7134 4180
rect 7070 4164 7134 4172
rect 7070 4148 7150 4164
rect 7166 4157 7228 4188
rect 7244 4157 7306 4188
rect 7375 4186 7424 4211
rect 7439 4186 7469 4202
rect 7338 4172 7368 4180
rect 7375 4178 7485 4186
rect 7338 4164 7383 4172
rect 7070 4146 7089 4148
rect 7104 4146 7150 4148
rect 7070 4130 7150 4146
rect 7177 4144 7212 4157
rect 7253 4154 7290 4157
rect 7253 4152 7295 4154
rect 7182 4141 7212 4144
rect 7191 4137 7198 4141
rect 7198 4136 7199 4137
rect 7157 4130 7167 4136
rect 6916 4122 6951 4130
rect 6916 4096 6917 4122
rect 6924 4096 6951 4122
rect 6859 4078 6889 4092
rect 6916 4088 6951 4096
rect 6953 4122 6994 4130
rect 6953 4096 6968 4122
rect 6975 4096 6994 4122
rect 7058 4118 7089 4130
rect 7104 4118 7207 4130
rect 7219 4120 7245 4146
rect 7260 4141 7290 4152
rect 7322 4148 7384 4164
rect 7322 4146 7368 4148
rect 7322 4130 7384 4146
rect 7396 4130 7402 4178
rect 7405 4170 7485 4178
rect 7405 4168 7424 4170
rect 7439 4168 7473 4170
rect 7405 4152 7485 4168
rect 7405 4130 7424 4152
rect 7439 4136 7469 4152
rect 7497 4146 7503 4220
rect 7506 4146 7525 4290
rect 7540 4146 7546 4290
rect 7555 4220 7568 4290
rect 7620 4286 7642 4290
rect 7613 4264 7642 4278
rect 7695 4264 7711 4278
rect 7749 4274 7755 4276
rect 7762 4274 7870 4290
rect 7877 4274 7883 4276
rect 7891 4274 7906 4290
rect 7972 4284 7991 4287
rect 7613 4262 7711 4264
rect 7738 4262 7906 4274
rect 7921 4264 7937 4278
rect 7972 4265 7994 4284
rect 8004 4278 8020 4279
rect 8003 4276 8020 4278
rect 8004 4271 8020 4276
rect 7994 4264 8000 4265
rect 8003 4264 8032 4271
rect 7921 4263 8032 4264
rect 7921 4262 8038 4263
rect 7597 4254 7648 4262
rect 7695 4254 7729 4262
rect 7597 4242 7622 4254
rect 7629 4242 7648 4254
rect 7702 4252 7729 4254
rect 7738 4252 7959 4262
rect 7994 4259 8000 4262
rect 7702 4248 7959 4252
rect 7597 4234 7648 4242
rect 7695 4234 7959 4248
rect 8003 4254 8038 4262
rect 7549 4186 7568 4220
rect 7613 4226 7642 4234
rect 7613 4220 7630 4226
rect 7613 4218 7647 4220
rect 7695 4218 7711 4234
rect 7712 4224 7920 4234
rect 7921 4224 7937 4234
rect 7985 4230 8000 4245
rect 8003 4242 8004 4254
rect 8011 4242 8038 4254
rect 8003 4234 8038 4242
rect 8003 4233 8032 4234
rect 7723 4220 7937 4224
rect 7738 4218 7937 4220
rect 7972 4220 7985 4230
rect 8003 4220 8020 4233
rect 7972 4218 8020 4220
rect 7614 4214 7647 4218
rect 7610 4212 7647 4214
rect 7610 4211 7677 4212
rect 7610 4206 7641 4211
rect 7647 4206 7677 4211
rect 7610 4202 7677 4206
rect 7583 4199 7677 4202
rect 7583 4192 7632 4199
rect 7583 4186 7613 4192
rect 7632 4187 7637 4192
rect 7549 4170 7629 4186
rect 7641 4178 7677 4199
rect 7738 4194 7927 4218
rect 7972 4217 8019 4218
rect 7985 4212 8019 4217
rect 7753 4191 7927 4194
rect 7746 4188 7927 4191
rect 7955 4211 8019 4212
rect 7549 4168 7568 4170
rect 7583 4168 7617 4170
rect 7549 4152 7629 4168
rect 7549 4146 7568 4152
rect 7265 4120 7368 4130
rect 7219 4118 7368 4120
rect 7389 4118 7424 4130
rect 7058 4116 7220 4118
rect 7070 4096 7089 4116
rect 7104 4114 7134 4116
rect 6953 4088 6994 4096
rect 7076 4092 7089 4096
rect 7141 4100 7220 4116
rect 7252 4116 7424 4118
rect 7252 4100 7331 4116
rect 7338 4114 7368 4116
rect 6916 4078 6945 4088
rect 6959 4078 6988 4088
rect 7003 4078 7033 4092
rect 7076 4078 7119 4092
rect 7141 4088 7331 4100
rect 7396 4096 7402 4116
rect 7126 4078 7156 4088
rect 7157 4078 7315 4088
rect 7319 4078 7349 4088
rect 7353 4078 7383 4092
rect 7411 4078 7424 4116
rect 7496 4130 7525 4146
rect 7539 4130 7568 4146
rect 7583 4136 7613 4152
rect 7641 4130 7647 4178
rect 7650 4172 7669 4178
rect 7684 4172 7714 4180
rect 7650 4164 7714 4172
rect 7650 4148 7730 4164
rect 7746 4157 7808 4188
rect 7824 4157 7886 4188
rect 7955 4186 8004 4211
rect 8019 4186 8049 4202
rect 7918 4172 7948 4180
rect 7955 4178 8065 4186
rect 7918 4164 7963 4172
rect 7650 4146 7669 4148
rect 7684 4146 7730 4148
rect 7650 4130 7730 4146
rect 7757 4144 7792 4157
rect 7833 4154 7870 4157
rect 7833 4152 7875 4154
rect 7762 4141 7792 4144
rect 7771 4137 7778 4141
rect 7778 4136 7779 4137
rect 7737 4130 7747 4136
rect 7496 4122 7531 4130
rect 7496 4096 7497 4122
rect 7504 4096 7531 4122
rect 7439 4078 7469 4092
rect 7496 4088 7531 4096
rect 7533 4122 7574 4130
rect 7533 4096 7548 4122
rect 7555 4096 7574 4122
rect 7638 4118 7669 4130
rect 7684 4118 7787 4130
rect 7799 4120 7825 4146
rect 7840 4141 7870 4152
rect 7902 4148 7964 4164
rect 7902 4146 7948 4148
rect 7902 4130 7964 4146
rect 7976 4130 7982 4178
rect 7985 4170 8065 4178
rect 7985 4168 8004 4170
rect 8019 4168 8053 4170
rect 7985 4152 8065 4168
rect 7985 4130 8004 4152
rect 8019 4136 8049 4152
rect 8077 4146 8083 4220
rect 8086 4146 8105 4290
rect 8120 4146 8126 4290
rect 8135 4220 8148 4290
rect 8200 4286 8222 4290
rect 8193 4264 8222 4278
rect 8275 4264 8291 4278
rect 8329 4274 8335 4276
rect 8342 4274 8450 4290
rect 8457 4274 8463 4276
rect 8471 4274 8486 4290
rect 8552 4284 8571 4287
rect 8193 4262 8291 4264
rect 8318 4262 8486 4274
rect 8501 4264 8517 4278
rect 8552 4265 8574 4284
rect 8584 4278 8600 4279
rect 8583 4276 8600 4278
rect 8584 4271 8600 4276
rect 8574 4264 8580 4265
rect 8583 4264 8612 4271
rect 8501 4263 8612 4264
rect 8501 4262 8618 4263
rect 8177 4254 8228 4262
rect 8275 4254 8309 4262
rect 8177 4242 8202 4254
rect 8209 4242 8228 4254
rect 8282 4252 8309 4254
rect 8318 4252 8539 4262
rect 8574 4259 8580 4262
rect 8282 4248 8539 4252
rect 8177 4234 8228 4242
rect 8275 4234 8539 4248
rect 8583 4254 8618 4262
rect 8129 4186 8148 4220
rect 8193 4226 8222 4234
rect 8193 4220 8210 4226
rect 8193 4218 8227 4220
rect 8275 4218 8291 4234
rect 8292 4224 8500 4234
rect 8501 4224 8517 4234
rect 8565 4230 8580 4245
rect 8583 4242 8584 4254
rect 8591 4242 8618 4254
rect 8583 4234 8618 4242
rect 8583 4233 8612 4234
rect 8303 4220 8517 4224
rect 8318 4218 8517 4220
rect 8552 4220 8565 4230
rect 8583 4220 8600 4233
rect 8552 4218 8600 4220
rect 8194 4214 8227 4218
rect 8190 4212 8227 4214
rect 8190 4211 8257 4212
rect 8190 4206 8221 4211
rect 8227 4206 8257 4211
rect 8190 4202 8257 4206
rect 8163 4199 8257 4202
rect 8163 4192 8212 4199
rect 8163 4186 8193 4192
rect 8212 4187 8217 4192
rect 8129 4170 8209 4186
rect 8221 4178 8257 4199
rect 8318 4194 8507 4218
rect 8552 4217 8599 4218
rect 8565 4212 8599 4217
rect 8333 4191 8507 4194
rect 8326 4188 8507 4191
rect 8535 4211 8599 4212
rect 8129 4168 8148 4170
rect 8163 4168 8197 4170
rect 8129 4152 8209 4168
rect 8129 4146 8148 4152
rect 7845 4120 7948 4130
rect 7799 4118 7948 4120
rect 7969 4118 8004 4130
rect 7638 4116 7800 4118
rect 7650 4096 7669 4116
rect 7684 4114 7714 4116
rect 7533 4088 7574 4096
rect 7656 4092 7669 4096
rect 7721 4100 7800 4116
rect 7832 4116 8004 4118
rect 7832 4100 7911 4116
rect 7918 4114 7948 4116
rect 7496 4078 7525 4088
rect 7539 4078 7568 4088
rect 7583 4078 7613 4092
rect 7656 4078 7699 4092
rect 7721 4088 7911 4100
rect 7976 4096 7982 4116
rect 7706 4078 7736 4088
rect 7737 4078 7895 4088
rect 7899 4078 7929 4088
rect 7933 4078 7963 4092
rect 7991 4078 8004 4116
rect 8076 4130 8105 4146
rect 8119 4130 8148 4146
rect 8163 4136 8193 4152
rect 8221 4130 8227 4178
rect 8230 4172 8249 4178
rect 8264 4172 8294 4180
rect 8230 4164 8294 4172
rect 8230 4148 8310 4164
rect 8326 4157 8388 4188
rect 8404 4157 8466 4188
rect 8535 4186 8584 4211
rect 8599 4186 8629 4202
rect 8498 4172 8528 4180
rect 8535 4178 8645 4186
rect 8498 4164 8543 4172
rect 8230 4146 8249 4148
rect 8264 4146 8310 4148
rect 8230 4130 8310 4146
rect 8337 4144 8372 4157
rect 8413 4154 8450 4157
rect 8413 4152 8455 4154
rect 8342 4141 8372 4144
rect 8351 4137 8358 4141
rect 8358 4136 8359 4137
rect 8317 4130 8327 4136
rect 8076 4122 8111 4130
rect 8076 4096 8077 4122
rect 8084 4096 8111 4122
rect 8019 4078 8049 4092
rect 8076 4088 8111 4096
rect 8113 4122 8154 4130
rect 8113 4096 8128 4122
rect 8135 4096 8154 4122
rect 8218 4118 8249 4130
rect 8264 4118 8367 4130
rect 8379 4120 8405 4146
rect 8420 4141 8450 4152
rect 8482 4148 8544 4164
rect 8482 4146 8528 4148
rect 8482 4130 8544 4146
rect 8556 4130 8562 4178
rect 8565 4170 8645 4178
rect 8565 4168 8584 4170
rect 8599 4168 8633 4170
rect 8565 4152 8645 4168
rect 8565 4130 8584 4152
rect 8599 4136 8629 4152
rect 8657 4146 8663 4220
rect 8666 4146 8685 4290
rect 8700 4146 8706 4290
rect 8715 4220 8728 4290
rect 8780 4286 8802 4290
rect 8773 4264 8802 4278
rect 8855 4264 8871 4278
rect 8909 4274 8915 4276
rect 8922 4274 9030 4290
rect 9037 4274 9043 4276
rect 9051 4274 9066 4290
rect 9132 4284 9151 4287
rect 8773 4262 8871 4264
rect 8898 4262 9066 4274
rect 9081 4264 9097 4278
rect 9132 4265 9154 4284
rect 9164 4278 9180 4279
rect 9163 4276 9180 4278
rect 9164 4271 9180 4276
rect 9154 4264 9160 4265
rect 9163 4264 9192 4271
rect 9081 4263 9192 4264
rect 9081 4262 9198 4263
rect 8757 4254 8808 4262
rect 8855 4254 8889 4262
rect 8757 4242 8782 4254
rect 8789 4242 8808 4254
rect 8862 4252 8889 4254
rect 8898 4252 9119 4262
rect 9154 4259 9160 4262
rect 8862 4248 9119 4252
rect 8757 4234 8808 4242
rect 8855 4234 9119 4248
rect 9163 4254 9198 4262
rect 8709 4186 8728 4220
rect 8773 4226 8802 4234
rect 8773 4220 8790 4226
rect 8773 4218 8807 4220
rect 8855 4218 8871 4234
rect 8872 4224 9080 4234
rect 9081 4224 9097 4234
rect 9145 4230 9160 4245
rect 9163 4242 9164 4254
rect 9171 4242 9198 4254
rect 9163 4234 9198 4242
rect 9163 4233 9192 4234
rect 8883 4220 9097 4224
rect 8898 4218 9097 4220
rect 9132 4220 9145 4230
rect 9163 4220 9180 4233
rect 9132 4218 9180 4220
rect 8774 4214 8807 4218
rect 8770 4212 8807 4214
rect 8770 4211 8837 4212
rect 8770 4206 8801 4211
rect 8807 4206 8837 4211
rect 8770 4202 8837 4206
rect 8743 4199 8837 4202
rect 8743 4192 8792 4199
rect 8743 4186 8773 4192
rect 8792 4187 8797 4192
rect 8709 4170 8789 4186
rect 8801 4178 8837 4199
rect 8898 4194 9087 4218
rect 9132 4217 9179 4218
rect 9145 4212 9179 4217
rect 8913 4191 9087 4194
rect 8906 4188 9087 4191
rect 9115 4211 9179 4212
rect 8709 4168 8728 4170
rect 8743 4168 8777 4170
rect 8709 4152 8789 4168
rect 8709 4146 8728 4152
rect 8425 4120 8528 4130
rect 8379 4118 8528 4120
rect 8549 4118 8584 4130
rect 8218 4116 8380 4118
rect 8230 4096 8249 4116
rect 8264 4114 8294 4116
rect 8113 4088 8154 4096
rect 8236 4092 8249 4096
rect 8301 4100 8380 4116
rect 8412 4116 8584 4118
rect 8412 4100 8491 4116
rect 8498 4114 8528 4116
rect 8076 4078 8105 4088
rect 8119 4078 8148 4088
rect 8163 4078 8193 4092
rect 8236 4078 8279 4092
rect 8301 4088 8491 4100
rect 8556 4096 8562 4116
rect 8286 4078 8316 4088
rect 8317 4078 8475 4088
rect 8479 4078 8509 4088
rect 8513 4078 8543 4092
rect 8571 4078 8584 4116
rect 8656 4130 8685 4146
rect 8699 4130 8728 4146
rect 8743 4136 8773 4152
rect 8801 4130 8807 4178
rect 8810 4172 8829 4178
rect 8844 4172 8874 4180
rect 8810 4164 8874 4172
rect 8810 4148 8890 4164
rect 8906 4157 8968 4188
rect 8984 4157 9046 4188
rect 9115 4186 9164 4211
rect 9179 4186 9209 4202
rect 9078 4172 9108 4180
rect 9115 4178 9225 4186
rect 9078 4164 9123 4172
rect 8810 4146 8829 4148
rect 8844 4146 8890 4148
rect 8810 4130 8890 4146
rect 8917 4144 8952 4157
rect 8993 4154 9030 4157
rect 8993 4152 9035 4154
rect 8922 4141 8952 4144
rect 8931 4137 8938 4141
rect 8938 4136 8939 4137
rect 8897 4130 8907 4136
rect 8656 4122 8691 4130
rect 8656 4096 8657 4122
rect 8664 4096 8691 4122
rect 8599 4078 8629 4092
rect 8656 4088 8691 4096
rect 8693 4122 8734 4130
rect 8693 4096 8708 4122
rect 8715 4096 8734 4122
rect 8798 4118 8829 4130
rect 8844 4118 8947 4130
rect 8959 4120 8985 4146
rect 9000 4141 9030 4152
rect 9062 4148 9124 4164
rect 9062 4146 9108 4148
rect 9062 4130 9124 4146
rect 9136 4130 9142 4178
rect 9145 4170 9225 4178
rect 9145 4168 9164 4170
rect 9179 4168 9213 4170
rect 9145 4152 9225 4168
rect 9145 4130 9164 4152
rect 9179 4136 9209 4152
rect 9237 4146 9243 4220
rect 9246 4146 9265 4290
rect 9280 4146 9286 4290
rect 9295 4220 9308 4290
rect 9360 4286 9382 4290
rect 9353 4264 9382 4278
rect 9435 4264 9451 4278
rect 9489 4274 9495 4276
rect 9502 4274 9610 4290
rect 9617 4274 9623 4276
rect 9631 4274 9646 4290
rect 9712 4284 9731 4287
rect 9353 4262 9451 4264
rect 9478 4262 9646 4274
rect 9661 4264 9677 4278
rect 9712 4265 9734 4284
rect 9744 4278 9760 4279
rect 9743 4276 9760 4278
rect 9744 4271 9760 4276
rect 9734 4264 9740 4265
rect 9743 4264 9772 4271
rect 9661 4263 9772 4264
rect 9661 4262 9778 4263
rect 9337 4254 9388 4262
rect 9435 4254 9469 4262
rect 9337 4242 9362 4254
rect 9369 4242 9388 4254
rect 9442 4252 9469 4254
rect 9478 4252 9699 4262
rect 9734 4259 9740 4262
rect 9442 4248 9699 4252
rect 9337 4234 9388 4242
rect 9435 4234 9699 4248
rect 9743 4254 9778 4262
rect 9289 4186 9308 4220
rect 9353 4226 9382 4234
rect 9353 4220 9370 4226
rect 9353 4218 9387 4220
rect 9435 4218 9451 4234
rect 9452 4224 9660 4234
rect 9661 4224 9677 4234
rect 9725 4230 9740 4245
rect 9743 4242 9744 4254
rect 9751 4242 9778 4254
rect 9743 4234 9778 4242
rect 9743 4233 9772 4234
rect 9463 4220 9677 4224
rect 9478 4218 9677 4220
rect 9712 4220 9725 4230
rect 9743 4220 9760 4233
rect 9712 4218 9760 4220
rect 9354 4214 9387 4218
rect 9350 4212 9387 4214
rect 9350 4211 9417 4212
rect 9350 4206 9381 4211
rect 9387 4206 9417 4211
rect 9350 4202 9417 4206
rect 9323 4199 9417 4202
rect 9323 4192 9372 4199
rect 9323 4186 9353 4192
rect 9372 4187 9377 4192
rect 9289 4170 9369 4186
rect 9381 4178 9417 4199
rect 9478 4194 9667 4218
rect 9712 4217 9759 4218
rect 9725 4212 9759 4217
rect 9493 4191 9667 4194
rect 9486 4188 9667 4191
rect 9695 4211 9759 4212
rect 9289 4168 9308 4170
rect 9323 4168 9357 4170
rect 9289 4152 9369 4168
rect 9289 4146 9308 4152
rect 9005 4120 9108 4130
rect 8959 4118 9108 4120
rect 9129 4118 9164 4130
rect 8798 4116 8960 4118
rect 8810 4096 8829 4116
rect 8844 4114 8874 4116
rect 8693 4088 8734 4096
rect 8816 4092 8829 4096
rect 8881 4100 8960 4116
rect 8992 4116 9164 4118
rect 8992 4100 9071 4116
rect 9078 4114 9108 4116
rect 8656 4078 8685 4088
rect 8699 4078 8728 4088
rect 8743 4078 8773 4092
rect 8816 4078 8859 4092
rect 8881 4088 9071 4100
rect 9136 4096 9142 4116
rect 8866 4078 8896 4088
rect 8897 4078 9055 4088
rect 9059 4078 9089 4088
rect 9093 4078 9123 4092
rect 9151 4078 9164 4116
rect 9236 4130 9265 4146
rect 9279 4130 9308 4146
rect 9323 4136 9353 4152
rect 9381 4130 9387 4178
rect 9390 4172 9409 4178
rect 9424 4172 9454 4180
rect 9390 4164 9454 4172
rect 9390 4148 9470 4164
rect 9486 4157 9548 4188
rect 9564 4157 9626 4188
rect 9695 4186 9744 4211
rect 9759 4186 9789 4202
rect 9658 4172 9688 4180
rect 9695 4178 9805 4186
rect 9658 4164 9703 4172
rect 9390 4146 9409 4148
rect 9424 4146 9470 4148
rect 9390 4130 9470 4146
rect 9497 4144 9532 4157
rect 9573 4154 9610 4157
rect 9573 4152 9615 4154
rect 9502 4141 9532 4144
rect 9511 4137 9518 4141
rect 9518 4136 9519 4137
rect 9477 4130 9487 4136
rect 9236 4122 9271 4130
rect 9236 4096 9237 4122
rect 9244 4096 9271 4122
rect 9179 4078 9209 4092
rect 9236 4088 9271 4096
rect 9273 4122 9314 4130
rect 9273 4096 9288 4122
rect 9295 4096 9314 4122
rect 9378 4118 9409 4130
rect 9424 4118 9527 4130
rect 9539 4120 9565 4146
rect 9580 4141 9610 4152
rect 9642 4148 9704 4164
rect 9642 4146 9688 4148
rect 9642 4130 9704 4146
rect 9716 4130 9722 4178
rect 9725 4170 9805 4178
rect 9725 4168 9744 4170
rect 9759 4168 9793 4170
rect 9725 4152 9805 4168
rect 9725 4130 9744 4152
rect 9759 4136 9789 4152
rect 9817 4146 9823 4220
rect 9826 4146 9845 4290
rect 9860 4146 9866 4290
rect 9875 4220 9888 4290
rect 9940 4286 9962 4290
rect 9933 4264 9962 4278
rect 10015 4264 10031 4278
rect 10069 4274 10075 4276
rect 10082 4274 10190 4290
rect 10197 4274 10203 4276
rect 10211 4274 10226 4290
rect 10292 4284 10311 4287
rect 9933 4262 10031 4264
rect 10058 4262 10226 4274
rect 10241 4264 10257 4278
rect 10292 4265 10314 4284
rect 10324 4278 10340 4279
rect 10323 4276 10340 4278
rect 10324 4271 10340 4276
rect 10314 4264 10320 4265
rect 10323 4264 10352 4271
rect 10241 4263 10352 4264
rect 10241 4262 10358 4263
rect 9917 4254 9968 4262
rect 10015 4254 10049 4262
rect 9917 4242 9942 4254
rect 9949 4242 9968 4254
rect 10022 4252 10049 4254
rect 10058 4252 10279 4262
rect 10314 4259 10320 4262
rect 10022 4248 10279 4252
rect 9917 4234 9968 4242
rect 10015 4234 10279 4248
rect 10323 4254 10358 4262
rect 9869 4186 9888 4220
rect 9933 4226 9962 4234
rect 9933 4220 9950 4226
rect 9933 4218 9967 4220
rect 10015 4218 10031 4234
rect 10032 4224 10240 4234
rect 10241 4224 10257 4234
rect 10305 4230 10320 4245
rect 10323 4242 10324 4254
rect 10331 4242 10358 4254
rect 10323 4234 10358 4242
rect 10323 4233 10352 4234
rect 10043 4220 10257 4224
rect 10058 4218 10257 4220
rect 10292 4220 10305 4230
rect 10323 4220 10340 4233
rect 10292 4218 10340 4220
rect 9934 4214 9967 4218
rect 9930 4212 9967 4214
rect 9930 4211 9997 4212
rect 9930 4206 9961 4211
rect 9967 4206 9997 4211
rect 9930 4202 9997 4206
rect 9903 4199 9997 4202
rect 9903 4192 9952 4199
rect 9903 4186 9933 4192
rect 9952 4187 9957 4192
rect 9869 4170 9949 4186
rect 9961 4178 9997 4199
rect 10058 4194 10247 4218
rect 10292 4217 10339 4218
rect 10305 4212 10339 4217
rect 10073 4191 10247 4194
rect 10066 4188 10247 4191
rect 10275 4211 10339 4212
rect 9869 4168 9888 4170
rect 9903 4168 9937 4170
rect 9869 4152 9949 4168
rect 9869 4146 9888 4152
rect 9585 4120 9688 4130
rect 9539 4118 9688 4120
rect 9709 4118 9744 4130
rect 9378 4116 9540 4118
rect 9390 4096 9409 4116
rect 9424 4114 9454 4116
rect 9273 4088 9314 4096
rect 9396 4092 9409 4096
rect 9461 4100 9540 4116
rect 9572 4116 9744 4118
rect 9572 4100 9651 4116
rect 9658 4114 9688 4116
rect 9236 4078 9265 4088
rect 9279 4078 9308 4088
rect 9323 4078 9353 4092
rect 9396 4078 9439 4092
rect 9461 4088 9651 4100
rect 9716 4096 9722 4116
rect 9446 4078 9476 4088
rect 9477 4078 9635 4088
rect 9639 4078 9669 4088
rect 9673 4078 9703 4092
rect 9731 4078 9744 4116
rect 9816 4130 9845 4146
rect 9859 4130 9888 4146
rect 9903 4136 9933 4152
rect 9961 4130 9967 4178
rect 9970 4172 9989 4178
rect 10004 4172 10034 4180
rect 9970 4164 10034 4172
rect 9970 4148 10050 4164
rect 10066 4157 10128 4188
rect 10144 4157 10206 4188
rect 10275 4186 10324 4211
rect 10339 4186 10369 4202
rect 10238 4172 10268 4180
rect 10275 4178 10385 4186
rect 10238 4164 10283 4172
rect 9970 4146 9989 4148
rect 10004 4146 10050 4148
rect 9970 4130 10050 4146
rect 10077 4144 10112 4157
rect 10153 4154 10190 4157
rect 10153 4152 10195 4154
rect 10082 4141 10112 4144
rect 10091 4137 10098 4141
rect 10098 4136 10099 4137
rect 10057 4130 10067 4136
rect 9816 4122 9851 4130
rect 9816 4096 9817 4122
rect 9824 4096 9851 4122
rect 9759 4078 9789 4092
rect 9816 4088 9851 4096
rect 9853 4122 9894 4130
rect 9853 4096 9868 4122
rect 9875 4096 9894 4122
rect 9958 4118 9989 4130
rect 10004 4118 10107 4130
rect 10119 4120 10145 4146
rect 10160 4141 10190 4152
rect 10222 4148 10284 4164
rect 10222 4146 10268 4148
rect 10222 4130 10284 4146
rect 10296 4130 10302 4178
rect 10305 4170 10385 4178
rect 10305 4168 10324 4170
rect 10339 4168 10373 4170
rect 10305 4152 10385 4168
rect 10305 4130 10324 4152
rect 10339 4136 10369 4152
rect 10397 4146 10403 4220
rect 10406 4146 10425 4290
rect 10440 4146 10446 4290
rect 10455 4220 10468 4290
rect 10520 4286 10542 4290
rect 10513 4264 10542 4278
rect 10595 4264 10611 4278
rect 10649 4274 10655 4276
rect 10662 4274 10770 4290
rect 10777 4274 10783 4276
rect 10791 4274 10806 4290
rect 10872 4284 10891 4287
rect 10513 4262 10611 4264
rect 10638 4262 10806 4274
rect 10821 4264 10837 4278
rect 10872 4265 10894 4284
rect 10904 4278 10920 4279
rect 10903 4276 10920 4278
rect 10904 4271 10920 4276
rect 10894 4264 10900 4265
rect 10903 4264 10932 4271
rect 10821 4263 10932 4264
rect 10821 4262 10938 4263
rect 10497 4254 10548 4262
rect 10595 4254 10629 4262
rect 10497 4242 10522 4254
rect 10529 4242 10548 4254
rect 10602 4252 10629 4254
rect 10638 4252 10859 4262
rect 10894 4259 10900 4262
rect 10602 4248 10859 4252
rect 10497 4234 10548 4242
rect 10595 4234 10859 4248
rect 10903 4254 10938 4262
rect 10449 4186 10468 4220
rect 10513 4226 10542 4234
rect 10513 4220 10530 4226
rect 10513 4218 10547 4220
rect 10595 4218 10611 4234
rect 10612 4224 10820 4234
rect 10821 4224 10837 4234
rect 10885 4230 10900 4245
rect 10903 4242 10904 4254
rect 10911 4242 10938 4254
rect 10903 4234 10938 4242
rect 10903 4233 10932 4234
rect 10623 4220 10837 4224
rect 10638 4218 10837 4220
rect 10872 4220 10885 4230
rect 10903 4220 10920 4233
rect 10872 4218 10920 4220
rect 10514 4214 10547 4218
rect 10510 4212 10547 4214
rect 10510 4211 10577 4212
rect 10510 4206 10541 4211
rect 10547 4206 10577 4211
rect 10510 4202 10577 4206
rect 10483 4199 10577 4202
rect 10483 4192 10532 4199
rect 10483 4186 10513 4192
rect 10532 4187 10537 4192
rect 10449 4170 10529 4186
rect 10541 4178 10577 4199
rect 10638 4194 10827 4218
rect 10872 4217 10919 4218
rect 10885 4212 10919 4217
rect 10653 4191 10827 4194
rect 10646 4188 10827 4191
rect 10855 4211 10919 4212
rect 10449 4168 10468 4170
rect 10483 4168 10517 4170
rect 10449 4152 10529 4168
rect 10449 4146 10468 4152
rect 10165 4120 10268 4130
rect 10119 4118 10268 4120
rect 10289 4118 10324 4130
rect 9958 4116 10120 4118
rect 9970 4096 9989 4116
rect 10004 4114 10034 4116
rect 9853 4088 9894 4096
rect 9976 4092 9989 4096
rect 10041 4100 10120 4116
rect 10152 4116 10324 4118
rect 10152 4100 10231 4116
rect 10238 4114 10268 4116
rect 9816 4078 9845 4088
rect 9859 4078 9888 4088
rect 9903 4078 9933 4092
rect 9976 4078 10019 4092
rect 10041 4088 10231 4100
rect 10296 4096 10302 4116
rect 10026 4078 10056 4088
rect 10057 4078 10215 4088
rect 10219 4078 10249 4088
rect 10253 4078 10283 4092
rect 10311 4078 10324 4116
rect 10396 4130 10425 4146
rect 10439 4130 10468 4146
rect 10483 4136 10513 4152
rect 10541 4130 10547 4178
rect 10550 4172 10569 4178
rect 10584 4172 10614 4180
rect 10550 4164 10614 4172
rect 10550 4148 10630 4164
rect 10646 4157 10708 4188
rect 10724 4157 10786 4188
rect 10855 4186 10904 4211
rect 10919 4186 10949 4202
rect 10818 4172 10848 4180
rect 10855 4178 10965 4186
rect 10818 4164 10863 4172
rect 10550 4146 10569 4148
rect 10584 4146 10630 4148
rect 10550 4130 10630 4146
rect 10657 4144 10692 4157
rect 10733 4154 10770 4157
rect 10733 4152 10775 4154
rect 10662 4141 10692 4144
rect 10671 4137 10678 4141
rect 10678 4136 10679 4137
rect 10637 4130 10647 4136
rect 10396 4122 10431 4130
rect 10396 4096 10397 4122
rect 10404 4096 10431 4122
rect 10339 4078 10369 4092
rect 10396 4088 10431 4096
rect 10433 4122 10474 4130
rect 10433 4096 10448 4122
rect 10455 4096 10474 4122
rect 10538 4118 10569 4130
rect 10584 4118 10687 4130
rect 10699 4120 10725 4146
rect 10740 4141 10770 4152
rect 10802 4148 10864 4164
rect 10802 4146 10848 4148
rect 10802 4130 10864 4146
rect 10876 4130 10882 4178
rect 10885 4170 10965 4178
rect 10885 4168 10904 4170
rect 10919 4168 10953 4170
rect 10885 4152 10965 4168
rect 10885 4130 10904 4152
rect 10919 4136 10949 4152
rect 10977 4146 10983 4220
rect 10986 4146 11005 4290
rect 11020 4146 11026 4290
rect 11035 4220 11048 4290
rect 11100 4286 11122 4290
rect 11093 4264 11122 4278
rect 11175 4264 11191 4278
rect 11229 4274 11235 4276
rect 11242 4274 11350 4290
rect 11357 4274 11363 4276
rect 11371 4274 11386 4290
rect 11452 4284 11471 4287
rect 11093 4262 11191 4264
rect 11218 4262 11386 4274
rect 11401 4264 11417 4278
rect 11452 4265 11474 4284
rect 11484 4278 11500 4279
rect 11483 4276 11500 4278
rect 11484 4271 11500 4276
rect 11474 4264 11480 4265
rect 11483 4264 11512 4271
rect 11401 4263 11512 4264
rect 11401 4262 11518 4263
rect 11077 4254 11128 4262
rect 11175 4254 11209 4262
rect 11077 4242 11102 4254
rect 11109 4242 11128 4254
rect 11182 4252 11209 4254
rect 11218 4252 11439 4262
rect 11474 4259 11480 4262
rect 11182 4248 11439 4252
rect 11077 4234 11128 4242
rect 11175 4234 11439 4248
rect 11483 4254 11518 4262
rect 11029 4186 11048 4220
rect 11093 4226 11122 4234
rect 11093 4220 11110 4226
rect 11093 4218 11127 4220
rect 11175 4218 11191 4234
rect 11192 4224 11400 4234
rect 11401 4224 11417 4234
rect 11465 4230 11480 4245
rect 11483 4242 11484 4254
rect 11491 4242 11518 4254
rect 11483 4234 11518 4242
rect 11483 4233 11512 4234
rect 11203 4220 11417 4224
rect 11218 4218 11417 4220
rect 11452 4220 11465 4230
rect 11483 4220 11500 4233
rect 11452 4218 11500 4220
rect 11094 4214 11127 4218
rect 11090 4212 11127 4214
rect 11090 4211 11157 4212
rect 11090 4206 11121 4211
rect 11127 4206 11157 4211
rect 11090 4202 11157 4206
rect 11063 4199 11157 4202
rect 11063 4192 11112 4199
rect 11063 4186 11093 4192
rect 11112 4187 11117 4192
rect 11029 4170 11109 4186
rect 11121 4178 11157 4199
rect 11218 4194 11407 4218
rect 11452 4217 11499 4218
rect 11465 4212 11499 4217
rect 11233 4191 11407 4194
rect 11226 4188 11407 4191
rect 11435 4211 11499 4212
rect 11029 4168 11048 4170
rect 11063 4168 11097 4170
rect 11029 4152 11109 4168
rect 11029 4146 11048 4152
rect 10745 4120 10848 4130
rect 10699 4118 10848 4120
rect 10869 4118 10904 4130
rect 10538 4116 10700 4118
rect 10550 4096 10569 4116
rect 10584 4114 10614 4116
rect 10433 4088 10474 4096
rect 10556 4092 10569 4096
rect 10621 4100 10700 4116
rect 10732 4116 10904 4118
rect 10732 4100 10811 4116
rect 10818 4114 10848 4116
rect 10396 4078 10425 4088
rect 10439 4078 10468 4088
rect 10483 4078 10513 4092
rect 10556 4078 10599 4092
rect 10621 4088 10811 4100
rect 10876 4096 10882 4116
rect 10606 4078 10636 4088
rect 10637 4078 10795 4088
rect 10799 4078 10829 4088
rect 10833 4078 10863 4092
rect 10891 4078 10904 4116
rect 10976 4130 11005 4146
rect 11019 4130 11048 4146
rect 11063 4136 11093 4152
rect 11121 4130 11127 4178
rect 11130 4172 11149 4178
rect 11164 4172 11194 4180
rect 11130 4164 11194 4172
rect 11130 4148 11210 4164
rect 11226 4157 11288 4188
rect 11304 4157 11366 4188
rect 11435 4186 11484 4211
rect 11499 4186 11529 4202
rect 11398 4172 11428 4180
rect 11435 4178 11545 4186
rect 11398 4164 11443 4172
rect 11130 4146 11149 4148
rect 11164 4146 11210 4148
rect 11130 4130 11210 4146
rect 11237 4144 11272 4157
rect 11313 4154 11350 4157
rect 11313 4152 11355 4154
rect 11242 4141 11272 4144
rect 11251 4137 11258 4141
rect 11258 4136 11259 4137
rect 11217 4130 11227 4136
rect 10976 4122 11011 4130
rect 10976 4096 10977 4122
rect 10984 4096 11011 4122
rect 10919 4078 10949 4092
rect 10976 4088 11011 4096
rect 11013 4122 11054 4130
rect 11013 4096 11028 4122
rect 11035 4096 11054 4122
rect 11118 4118 11149 4130
rect 11164 4118 11267 4130
rect 11279 4120 11305 4146
rect 11320 4141 11350 4152
rect 11382 4148 11444 4164
rect 11382 4146 11428 4148
rect 11382 4130 11444 4146
rect 11456 4130 11462 4178
rect 11465 4170 11545 4178
rect 11465 4168 11484 4170
rect 11499 4168 11533 4170
rect 11465 4152 11545 4168
rect 11465 4130 11484 4152
rect 11499 4136 11529 4152
rect 11557 4146 11563 4220
rect 11566 4146 11585 4290
rect 11600 4146 11606 4290
rect 11615 4220 11628 4290
rect 11680 4286 11702 4290
rect 11673 4264 11702 4278
rect 11755 4264 11771 4278
rect 11809 4274 11815 4276
rect 11822 4274 11930 4290
rect 11937 4274 11943 4276
rect 11951 4274 11966 4290
rect 12032 4284 12051 4287
rect 11673 4262 11771 4264
rect 11798 4262 11966 4274
rect 11981 4264 11997 4278
rect 12032 4265 12054 4284
rect 12064 4278 12080 4279
rect 12063 4276 12080 4278
rect 12064 4271 12080 4276
rect 12054 4264 12060 4265
rect 12063 4264 12092 4271
rect 11981 4263 12092 4264
rect 11981 4262 12098 4263
rect 11657 4254 11708 4262
rect 11755 4254 11789 4262
rect 11657 4242 11682 4254
rect 11689 4242 11708 4254
rect 11762 4252 11789 4254
rect 11798 4252 12019 4262
rect 12054 4259 12060 4262
rect 11762 4248 12019 4252
rect 11657 4234 11708 4242
rect 11755 4234 12019 4248
rect 12063 4254 12098 4262
rect 11609 4186 11628 4220
rect 11673 4226 11702 4234
rect 11673 4220 11690 4226
rect 11673 4218 11707 4220
rect 11755 4218 11771 4234
rect 11772 4224 11980 4234
rect 11981 4224 11997 4234
rect 12045 4230 12060 4245
rect 12063 4242 12064 4254
rect 12071 4242 12098 4254
rect 12063 4234 12098 4242
rect 12063 4233 12092 4234
rect 11783 4220 11997 4224
rect 11798 4218 11997 4220
rect 12032 4220 12045 4230
rect 12063 4220 12080 4233
rect 12032 4218 12080 4220
rect 11674 4214 11707 4218
rect 11670 4212 11707 4214
rect 11670 4211 11737 4212
rect 11670 4206 11701 4211
rect 11707 4206 11737 4211
rect 11670 4202 11737 4206
rect 11643 4199 11737 4202
rect 11643 4192 11692 4199
rect 11643 4186 11673 4192
rect 11692 4187 11697 4192
rect 11609 4170 11689 4186
rect 11701 4178 11737 4199
rect 11798 4194 11987 4218
rect 12032 4217 12079 4218
rect 12045 4212 12079 4217
rect 11813 4191 11987 4194
rect 11806 4188 11987 4191
rect 12015 4211 12079 4212
rect 11609 4168 11628 4170
rect 11643 4168 11677 4170
rect 11609 4152 11689 4168
rect 11609 4146 11628 4152
rect 11325 4120 11428 4130
rect 11279 4118 11428 4120
rect 11449 4118 11484 4130
rect 11118 4116 11280 4118
rect 11130 4096 11149 4116
rect 11164 4114 11194 4116
rect 11013 4088 11054 4096
rect 11136 4092 11149 4096
rect 11201 4100 11280 4116
rect 11312 4116 11484 4118
rect 11312 4100 11391 4116
rect 11398 4114 11428 4116
rect 10976 4078 11005 4088
rect 11019 4078 11048 4088
rect 11063 4078 11093 4092
rect 11136 4078 11179 4092
rect 11201 4088 11391 4100
rect 11456 4096 11462 4116
rect 11186 4078 11216 4088
rect 11217 4078 11375 4088
rect 11379 4078 11409 4088
rect 11413 4078 11443 4092
rect 11471 4078 11484 4116
rect 11556 4130 11585 4146
rect 11599 4130 11628 4146
rect 11643 4136 11673 4152
rect 11701 4130 11707 4178
rect 11710 4172 11729 4178
rect 11744 4172 11774 4180
rect 11710 4164 11774 4172
rect 11710 4148 11790 4164
rect 11806 4157 11868 4188
rect 11884 4157 11946 4188
rect 12015 4186 12064 4211
rect 12079 4186 12109 4202
rect 11978 4172 12008 4180
rect 12015 4178 12125 4186
rect 11978 4164 12023 4172
rect 11710 4146 11729 4148
rect 11744 4146 11790 4148
rect 11710 4130 11790 4146
rect 11817 4144 11852 4157
rect 11893 4154 11930 4157
rect 11893 4152 11935 4154
rect 11822 4141 11852 4144
rect 11831 4137 11838 4141
rect 11838 4136 11839 4137
rect 11797 4130 11807 4136
rect 11556 4122 11591 4130
rect 11556 4096 11557 4122
rect 11564 4096 11591 4122
rect 11499 4078 11529 4092
rect 11556 4088 11591 4096
rect 11593 4122 11634 4130
rect 11593 4096 11608 4122
rect 11615 4096 11634 4122
rect 11698 4118 11729 4130
rect 11744 4118 11847 4130
rect 11859 4120 11885 4146
rect 11900 4141 11930 4152
rect 11962 4148 12024 4164
rect 11962 4146 12008 4148
rect 11962 4130 12024 4146
rect 12036 4130 12042 4178
rect 12045 4170 12125 4178
rect 12045 4168 12064 4170
rect 12079 4168 12113 4170
rect 12045 4152 12125 4168
rect 12045 4130 12064 4152
rect 12079 4136 12109 4152
rect 12137 4146 12143 4220
rect 12146 4146 12165 4290
rect 12180 4146 12186 4290
rect 12195 4220 12208 4290
rect 12260 4286 12282 4290
rect 12253 4264 12282 4278
rect 12335 4264 12351 4278
rect 12389 4274 12395 4276
rect 12402 4274 12510 4290
rect 12517 4274 12523 4276
rect 12531 4274 12546 4290
rect 12612 4284 12631 4287
rect 12253 4262 12351 4264
rect 12378 4262 12546 4274
rect 12561 4264 12577 4278
rect 12612 4265 12634 4284
rect 12644 4278 12660 4279
rect 12643 4276 12660 4278
rect 12644 4271 12660 4276
rect 12634 4264 12640 4265
rect 12643 4264 12672 4271
rect 12561 4263 12672 4264
rect 12561 4262 12678 4263
rect 12237 4254 12288 4262
rect 12335 4254 12369 4262
rect 12237 4242 12262 4254
rect 12269 4242 12288 4254
rect 12342 4252 12369 4254
rect 12378 4252 12599 4262
rect 12634 4259 12640 4262
rect 12342 4248 12599 4252
rect 12237 4234 12288 4242
rect 12335 4234 12599 4248
rect 12643 4254 12678 4262
rect 12189 4186 12208 4220
rect 12253 4226 12282 4234
rect 12253 4220 12270 4226
rect 12253 4218 12287 4220
rect 12335 4218 12351 4234
rect 12352 4224 12560 4234
rect 12561 4224 12577 4234
rect 12625 4230 12640 4245
rect 12643 4242 12644 4254
rect 12651 4242 12678 4254
rect 12643 4234 12678 4242
rect 12643 4233 12672 4234
rect 12363 4220 12577 4224
rect 12378 4218 12577 4220
rect 12612 4220 12625 4230
rect 12643 4220 12660 4233
rect 12612 4218 12660 4220
rect 12254 4214 12287 4218
rect 12250 4212 12287 4214
rect 12250 4211 12317 4212
rect 12250 4206 12281 4211
rect 12287 4206 12317 4211
rect 12250 4202 12317 4206
rect 12223 4199 12317 4202
rect 12223 4192 12272 4199
rect 12223 4186 12253 4192
rect 12272 4187 12277 4192
rect 12189 4170 12269 4186
rect 12281 4178 12317 4199
rect 12378 4194 12567 4218
rect 12612 4217 12659 4218
rect 12625 4212 12659 4217
rect 12393 4191 12567 4194
rect 12386 4188 12567 4191
rect 12595 4211 12659 4212
rect 12189 4168 12208 4170
rect 12223 4168 12257 4170
rect 12189 4152 12269 4168
rect 12189 4146 12208 4152
rect 11905 4120 12008 4130
rect 11859 4118 12008 4120
rect 12029 4118 12064 4130
rect 11698 4116 11860 4118
rect 11710 4096 11729 4116
rect 11744 4114 11774 4116
rect 11593 4088 11634 4096
rect 11716 4092 11729 4096
rect 11781 4100 11860 4116
rect 11892 4116 12064 4118
rect 11892 4100 11971 4116
rect 11978 4114 12008 4116
rect 11556 4078 11585 4088
rect 11599 4078 11628 4088
rect 11643 4078 11673 4092
rect 11716 4078 11759 4092
rect 11781 4088 11971 4100
rect 12036 4096 12042 4116
rect 11766 4078 11796 4088
rect 11797 4078 11955 4088
rect 11959 4078 11989 4088
rect 11993 4078 12023 4092
rect 12051 4078 12064 4116
rect 12136 4130 12165 4146
rect 12179 4130 12208 4146
rect 12223 4136 12253 4152
rect 12281 4130 12287 4178
rect 12290 4172 12309 4178
rect 12324 4172 12354 4180
rect 12290 4164 12354 4172
rect 12290 4148 12370 4164
rect 12386 4157 12448 4188
rect 12464 4157 12526 4188
rect 12595 4186 12644 4211
rect 12659 4186 12689 4202
rect 12558 4172 12588 4180
rect 12595 4178 12705 4186
rect 12558 4164 12603 4172
rect 12290 4146 12309 4148
rect 12324 4146 12370 4148
rect 12290 4130 12370 4146
rect 12397 4144 12432 4157
rect 12473 4154 12510 4157
rect 12473 4152 12515 4154
rect 12402 4141 12432 4144
rect 12411 4137 12418 4141
rect 12418 4136 12419 4137
rect 12377 4130 12387 4136
rect 12136 4122 12171 4130
rect 12136 4096 12137 4122
rect 12144 4096 12171 4122
rect 12079 4078 12109 4092
rect 12136 4088 12171 4096
rect 12173 4122 12214 4130
rect 12173 4096 12188 4122
rect 12195 4096 12214 4122
rect 12278 4118 12309 4130
rect 12324 4118 12427 4130
rect 12439 4120 12465 4146
rect 12480 4141 12510 4152
rect 12542 4148 12604 4164
rect 12542 4146 12588 4148
rect 12542 4130 12604 4146
rect 12616 4130 12622 4178
rect 12625 4170 12705 4178
rect 12625 4168 12644 4170
rect 12659 4168 12693 4170
rect 12625 4152 12705 4168
rect 12625 4130 12644 4152
rect 12659 4136 12689 4152
rect 12717 4146 12723 4220
rect 12726 4146 12745 4290
rect 12760 4146 12766 4290
rect 12775 4220 12788 4290
rect 12840 4286 12862 4290
rect 12833 4264 12862 4278
rect 12915 4264 12931 4278
rect 12969 4274 12975 4276
rect 12982 4274 13090 4290
rect 13097 4274 13103 4276
rect 13111 4274 13126 4290
rect 13192 4284 13211 4287
rect 12833 4262 12931 4264
rect 12958 4262 13126 4274
rect 13141 4264 13157 4278
rect 13192 4265 13214 4284
rect 13224 4278 13240 4279
rect 13223 4276 13240 4278
rect 13224 4271 13240 4276
rect 13214 4264 13220 4265
rect 13223 4264 13252 4271
rect 13141 4263 13252 4264
rect 13141 4262 13258 4263
rect 12817 4254 12868 4262
rect 12915 4254 12949 4262
rect 12817 4242 12842 4254
rect 12849 4242 12868 4254
rect 12922 4252 12949 4254
rect 12958 4252 13179 4262
rect 13214 4259 13220 4262
rect 12922 4248 13179 4252
rect 12817 4234 12868 4242
rect 12915 4234 13179 4248
rect 13223 4254 13258 4262
rect 12769 4186 12788 4220
rect 12833 4226 12862 4234
rect 12833 4220 12850 4226
rect 12833 4218 12867 4220
rect 12915 4218 12931 4234
rect 12932 4224 13140 4234
rect 13141 4224 13157 4234
rect 13205 4230 13220 4245
rect 13223 4242 13224 4254
rect 13231 4242 13258 4254
rect 13223 4234 13258 4242
rect 13223 4233 13252 4234
rect 12943 4220 13157 4224
rect 12958 4218 13157 4220
rect 13192 4220 13205 4230
rect 13223 4220 13240 4233
rect 13192 4218 13240 4220
rect 12834 4214 12867 4218
rect 12830 4212 12867 4214
rect 12830 4211 12897 4212
rect 12830 4206 12861 4211
rect 12867 4206 12897 4211
rect 12830 4202 12897 4206
rect 12803 4199 12897 4202
rect 12803 4192 12852 4199
rect 12803 4186 12833 4192
rect 12852 4187 12857 4192
rect 12769 4170 12849 4186
rect 12861 4178 12897 4199
rect 12958 4194 13147 4218
rect 13192 4217 13239 4218
rect 13205 4212 13239 4217
rect 12973 4191 13147 4194
rect 12966 4188 13147 4191
rect 13175 4211 13239 4212
rect 12769 4168 12788 4170
rect 12803 4168 12837 4170
rect 12769 4152 12849 4168
rect 12769 4146 12788 4152
rect 12485 4120 12588 4130
rect 12439 4118 12588 4120
rect 12609 4118 12644 4130
rect 12278 4116 12440 4118
rect 12290 4096 12309 4116
rect 12324 4114 12354 4116
rect 12173 4088 12214 4096
rect 12296 4092 12309 4096
rect 12361 4100 12440 4116
rect 12472 4116 12644 4118
rect 12472 4100 12551 4116
rect 12558 4114 12588 4116
rect 12136 4078 12165 4088
rect 12179 4078 12208 4088
rect 12223 4078 12253 4092
rect 12296 4078 12339 4092
rect 12361 4088 12551 4100
rect 12616 4096 12622 4116
rect 12346 4078 12376 4088
rect 12377 4078 12535 4088
rect 12539 4078 12569 4088
rect 12573 4078 12603 4092
rect 12631 4078 12644 4116
rect 12716 4130 12745 4146
rect 12759 4130 12788 4146
rect 12803 4136 12833 4152
rect 12861 4130 12867 4178
rect 12870 4172 12889 4178
rect 12904 4172 12934 4180
rect 12870 4164 12934 4172
rect 12870 4148 12950 4164
rect 12966 4157 13028 4188
rect 13044 4157 13106 4188
rect 13175 4186 13224 4211
rect 13239 4186 13269 4202
rect 13138 4172 13168 4180
rect 13175 4178 13285 4186
rect 13138 4164 13183 4172
rect 12870 4146 12889 4148
rect 12904 4146 12950 4148
rect 12870 4130 12950 4146
rect 12977 4144 13012 4157
rect 13053 4154 13090 4157
rect 13053 4152 13095 4154
rect 12982 4141 13012 4144
rect 12991 4137 12998 4141
rect 12998 4136 12999 4137
rect 12957 4130 12967 4136
rect 12716 4122 12751 4130
rect 12716 4096 12717 4122
rect 12724 4096 12751 4122
rect 12659 4078 12689 4092
rect 12716 4088 12751 4096
rect 12753 4122 12794 4130
rect 12753 4096 12768 4122
rect 12775 4096 12794 4122
rect 12858 4118 12889 4130
rect 12904 4118 13007 4130
rect 13019 4120 13045 4146
rect 13060 4141 13090 4152
rect 13122 4148 13184 4164
rect 13122 4146 13168 4148
rect 13122 4130 13184 4146
rect 13196 4130 13202 4178
rect 13205 4170 13285 4178
rect 13205 4168 13224 4170
rect 13239 4168 13273 4170
rect 13205 4152 13285 4168
rect 13205 4130 13224 4152
rect 13239 4136 13269 4152
rect 13297 4146 13303 4220
rect 13306 4146 13325 4290
rect 13340 4146 13346 4290
rect 13355 4220 13368 4290
rect 13420 4286 13442 4290
rect 13413 4264 13442 4278
rect 13495 4264 13511 4278
rect 13549 4274 13555 4276
rect 13562 4274 13670 4290
rect 13677 4274 13683 4276
rect 13691 4274 13706 4290
rect 13772 4284 13791 4287
rect 13413 4262 13511 4264
rect 13538 4262 13706 4274
rect 13721 4264 13737 4278
rect 13772 4265 13794 4284
rect 13804 4278 13820 4279
rect 13803 4276 13820 4278
rect 13804 4271 13820 4276
rect 13794 4264 13800 4265
rect 13803 4264 13832 4271
rect 13721 4263 13832 4264
rect 13721 4262 13838 4263
rect 13397 4254 13448 4262
rect 13495 4254 13529 4262
rect 13397 4242 13422 4254
rect 13429 4242 13448 4254
rect 13502 4252 13529 4254
rect 13538 4252 13759 4262
rect 13794 4259 13800 4262
rect 13502 4248 13759 4252
rect 13397 4234 13448 4242
rect 13495 4234 13759 4248
rect 13803 4254 13838 4262
rect 13349 4186 13368 4220
rect 13413 4226 13442 4234
rect 13413 4220 13430 4226
rect 13413 4218 13447 4220
rect 13495 4218 13511 4234
rect 13512 4224 13720 4234
rect 13721 4224 13737 4234
rect 13785 4230 13800 4245
rect 13803 4242 13804 4254
rect 13811 4242 13838 4254
rect 13803 4234 13838 4242
rect 13803 4233 13832 4234
rect 13523 4220 13737 4224
rect 13538 4218 13737 4220
rect 13772 4220 13785 4230
rect 13803 4220 13820 4233
rect 13772 4218 13820 4220
rect 13414 4214 13447 4218
rect 13410 4212 13447 4214
rect 13410 4211 13477 4212
rect 13410 4206 13441 4211
rect 13447 4206 13477 4211
rect 13410 4202 13477 4206
rect 13383 4199 13477 4202
rect 13383 4192 13432 4199
rect 13383 4186 13413 4192
rect 13432 4187 13437 4192
rect 13349 4170 13429 4186
rect 13441 4178 13477 4199
rect 13538 4194 13727 4218
rect 13772 4217 13819 4218
rect 13785 4212 13819 4217
rect 13553 4191 13727 4194
rect 13546 4188 13727 4191
rect 13755 4211 13819 4212
rect 13349 4168 13368 4170
rect 13383 4168 13417 4170
rect 13349 4152 13429 4168
rect 13349 4146 13368 4152
rect 13065 4120 13168 4130
rect 13019 4118 13168 4120
rect 13189 4118 13224 4130
rect 12858 4116 13020 4118
rect 12870 4096 12889 4116
rect 12904 4114 12934 4116
rect 12753 4088 12794 4096
rect 12876 4092 12889 4096
rect 12941 4100 13020 4116
rect 13052 4116 13224 4118
rect 13052 4100 13131 4116
rect 13138 4114 13168 4116
rect 12716 4078 12745 4088
rect 12759 4078 12788 4088
rect 12803 4078 12833 4092
rect 12876 4078 12919 4092
rect 12941 4088 13131 4100
rect 13196 4096 13202 4116
rect 12926 4078 12956 4088
rect 12957 4078 13115 4088
rect 13119 4078 13149 4088
rect 13153 4078 13183 4092
rect 13211 4078 13224 4116
rect 13296 4130 13325 4146
rect 13339 4130 13368 4146
rect 13383 4136 13413 4152
rect 13441 4130 13447 4178
rect 13450 4172 13469 4178
rect 13484 4172 13514 4180
rect 13450 4164 13514 4172
rect 13450 4148 13530 4164
rect 13546 4157 13608 4188
rect 13624 4157 13686 4188
rect 13755 4186 13804 4211
rect 13819 4186 13849 4202
rect 13718 4172 13748 4180
rect 13755 4178 13865 4186
rect 13718 4164 13763 4172
rect 13450 4146 13469 4148
rect 13484 4146 13530 4148
rect 13450 4130 13530 4146
rect 13557 4144 13592 4157
rect 13633 4154 13670 4157
rect 13633 4152 13675 4154
rect 13562 4141 13592 4144
rect 13571 4137 13578 4141
rect 13578 4136 13579 4137
rect 13537 4130 13547 4136
rect 13296 4122 13331 4130
rect 13296 4096 13297 4122
rect 13304 4096 13331 4122
rect 13239 4078 13269 4092
rect 13296 4088 13331 4096
rect 13333 4122 13374 4130
rect 13333 4096 13348 4122
rect 13355 4096 13374 4122
rect 13438 4118 13469 4130
rect 13484 4118 13587 4130
rect 13599 4120 13625 4146
rect 13640 4141 13670 4152
rect 13702 4148 13764 4164
rect 13702 4146 13748 4148
rect 13702 4130 13764 4146
rect 13776 4130 13782 4178
rect 13785 4170 13865 4178
rect 13785 4168 13804 4170
rect 13819 4168 13853 4170
rect 13785 4152 13865 4168
rect 13785 4130 13804 4152
rect 13819 4136 13849 4152
rect 13877 4146 13883 4220
rect 13886 4146 13905 4290
rect 13920 4146 13926 4290
rect 13935 4220 13948 4290
rect 14000 4286 14022 4290
rect 13993 4264 14022 4278
rect 14075 4264 14091 4278
rect 14129 4274 14135 4276
rect 14142 4274 14250 4290
rect 14257 4274 14263 4276
rect 14271 4274 14286 4290
rect 14352 4284 14371 4287
rect 13993 4262 14091 4264
rect 14118 4262 14286 4274
rect 14301 4264 14317 4278
rect 14352 4265 14374 4284
rect 14384 4278 14400 4279
rect 14383 4276 14400 4278
rect 14384 4271 14400 4276
rect 14374 4264 14380 4265
rect 14383 4264 14412 4271
rect 14301 4263 14412 4264
rect 14301 4262 14418 4263
rect 13977 4254 14028 4262
rect 14075 4254 14109 4262
rect 13977 4242 14002 4254
rect 14009 4242 14028 4254
rect 14082 4252 14109 4254
rect 14118 4252 14339 4262
rect 14374 4259 14380 4262
rect 14082 4248 14339 4252
rect 13977 4234 14028 4242
rect 14075 4234 14339 4248
rect 14383 4254 14418 4262
rect 13929 4186 13948 4220
rect 13993 4226 14022 4234
rect 13993 4220 14010 4226
rect 13993 4218 14027 4220
rect 14075 4218 14091 4234
rect 14092 4224 14300 4234
rect 14301 4224 14317 4234
rect 14365 4230 14380 4245
rect 14383 4242 14384 4254
rect 14391 4242 14418 4254
rect 14383 4234 14418 4242
rect 14383 4233 14412 4234
rect 14103 4220 14317 4224
rect 14118 4218 14317 4220
rect 14352 4220 14365 4230
rect 14383 4220 14400 4233
rect 14352 4218 14400 4220
rect 13994 4214 14027 4218
rect 13990 4212 14027 4214
rect 13990 4211 14057 4212
rect 13990 4206 14021 4211
rect 14027 4206 14057 4211
rect 13990 4202 14057 4206
rect 13963 4199 14057 4202
rect 13963 4192 14012 4199
rect 13963 4186 13993 4192
rect 14012 4187 14017 4192
rect 13929 4170 14009 4186
rect 14021 4178 14057 4199
rect 14118 4194 14307 4218
rect 14352 4217 14399 4218
rect 14365 4212 14399 4217
rect 14133 4191 14307 4194
rect 14126 4188 14307 4191
rect 14335 4211 14399 4212
rect 13929 4168 13948 4170
rect 13963 4168 13997 4170
rect 13929 4152 14009 4168
rect 13929 4146 13948 4152
rect 13645 4120 13748 4130
rect 13599 4118 13748 4120
rect 13769 4118 13804 4130
rect 13438 4116 13600 4118
rect 13450 4096 13469 4116
rect 13484 4114 13514 4116
rect 13333 4088 13374 4096
rect 13456 4092 13469 4096
rect 13521 4100 13600 4116
rect 13632 4116 13804 4118
rect 13632 4100 13711 4116
rect 13718 4114 13748 4116
rect 13296 4078 13325 4088
rect 13339 4078 13368 4088
rect 13383 4078 13413 4092
rect 13456 4078 13499 4092
rect 13521 4088 13711 4100
rect 13776 4096 13782 4116
rect 13506 4078 13536 4088
rect 13537 4078 13695 4088
rect 13699 4078 13729 4088
rect 13733 4078 13763 4092
rect 13791 4078 13804 4116
rect 13876 4130 13905 4146
rect 13919 4130 13948 4146
rect 13963 4136 13993 4152
rect 14021 4130 14027 4178
rect 14030 4172 14049 4178
rect 14064 4172 14094 4180
rect 14030 4164 14094 4172
rect 14030 4148 14110 4164
rect 14126 4157 14188 4188
rect 14204 4157 14266 4188
rect 14335 4186 14384 4211
rect 14399 4186 14429 4202
rect 14298 4172 14328 4180
rect 14335 4178 14445 4186
rect 14298 4164 14343 4172
rect 14030 4146 14049 4148
rect 14064 4146 14110 4148
rect 14030 4130 14110 4146
rect 14137 4144 14172 4157
rect 14213 4154 14250 4157
rect 14213 4152 14255 4154
rect 14142 4141 14172 4144
rect 14151 4137 14158 4141
rect 14158 4136 14159 4137
rect 14117 4130 14127 4136
rect 13876 4122 13911 4130
rect 13876 4096 13877 4122
rect 13884 4096 13911 4122
rect 13819 4078 13849 4092
rect 13876 4088 13911 4096
rect 13913 4122 13954 4130
rect 13913 4096 13928 4122
rect 13935 4096 13954 4122
rect 14018 4118 14049 4130
rect 14064 4118 14167 4130
rect 14179 4120 14205 4146
rect 14220 4141 14250 4152
rect 14282 4148 14344 4164
rect 14282 4146 14328 4148
rect 14282 4130 14344 4146
rect 14356 4130 14362 4178
rect 14365 4170 14445 4178
rect 14365 4168 14384 4170
rect 14399 4168 14433 4170
rect 14365 4152 14445 4168
rect 14365 4130 14384 4152
rect 14399 4136 14429 4152
rect 14457 4146 14463 4220
rect 14466 4146 14485 4290
rect 14500 4146 14506 4290
rect 14515 4220 14528 4290
rect 14580 4286 14602 4290
rect 14573 4264 14602 4278
rect 14655 4264 14671 4278
rect 14709 4274 14715 4276
rect 14722 4274 14830 4290
rect 14837 4274 14843 4276
rect 14851 4274 14866 4290
rect 14932 4284 14951 4287
rect 14573 4262 14671 4264
rect 14698 4262 14866 4274
rect 14881 4264 14897 4278
rect 14932 4265 14954 4284
rect 14964 4278 14980 4279
rect 14963 4276 14980 4278
rect 14964 4271 14980 4276
rect 14954 4264 14960 4265
rect 14963 4264 14992 4271
rect 14881 4263 14992 4264
rect 14881 4262 14998 4263
rect 14557 4254 14608 4262
rect 14655 4254 14689 4262
rect 14557 4242 14582 4254
rect 14589 4242 14608 4254
rect 14662 4252 14689 4254
rect 14698 4252 14919 4262
rect 14954 4259 14960 4262
rect 14662 4248 14919 4252
rect 14557 4234 14608 4242
rect 14655 4234 14919 4248
rect 14963 4254 14998 4262
rect 14509 4186 14528 4220
rect 14573 4226 14602 4234
rect 14573 4220 14590 4226
rect 14573 4218 14607 4220
rect 14655 4218 14671 4234
rect 14672 4224 14880 4234
rect 14881 4224 14897 4234
rect 14945 4230 14960 4245
rect 14963 4242 14964 4254
rect 14971 4242 14998 4254
rect 14963 4234 14998 4242
rect 14963 4233 14992 4234
rect 14683 4220 14897 4224
rect 14698 4218 14897 4220
rect 14932 4220 14945 4230
rect 14963 4220 14980 4233
rect 14932 4218 14980 4220
rect 14574 4214 14607 4218
rect 14570 4212 14607 4214
rect 14570 4211 14637 4212
rect 14570 4206 14601 4211
rect 14607 4206 14637 4211
rect 14570 4202 14637 4206
rect 14543 4199 14637 4202
rect 14543 4192 14592 4199
rect 14543 4186 14573 4192
rect 14592 4187 14597 4192
rect 14509 4170 14589 4186
rect 14601 4178 14637 4199
rect 14698 4194 14887 4218
rect 14932 4217 14979 4218
rect 14945 4212 14979 4217
rect 14713 4191 14887 4194
rect 14706 4188 14887 4191
rect 14915 4211 14979 4212
rect 14509 4168 14528 4170
rect 14543 4168 14577 4170
rect 14509 4152 14589 4168
rect 14509 4146 14528 4152
rect 14225 4120 14328 4130
rect 14179 4118 14328 4120
rect 14349 4118 14384 4130
rect 14018 4116 14180 4118
rect 14030 4096 14049 4116
rect 14064 4114 14094 4116
rect 13913 4088 13954 4096
rect 14036 4092 14049 4096
rect 14101 4100 14180 4116
rect 14212 4116 14384 4118
rect 14212 4100 14291 4116
rect 14298 4114 14328 4116
rect 13876 4078 13905 4088
rect 13919 4078 13948 4088
rect 13963 4078 13993 4092
rect 14036 4078 14079 4092
rect 14101 4088 14291 4100
rect 14356 4096 14362 4116
rect 14086 4078 14116 4088
rect 14117 4078 14275 4088
rect 14279 4078 14309 4088
rect 14313 4078 14343 4092
rect 14371 4078 14384 4116
rect 14456 4130 14485 4146
rect 14499 4130 14528 4146
rect 14543 4136 14573 4152
rect 14601 4130 14607 4178
rect 14610 4172 14629 4178
rect 14644 4172 14674 4180
rect 14610 4164 14674 4172
rect 14610 4148 14690 4164
rect 14706 4157 14768 4188
rect 14784 4157 14846 4188
rect 14915 4186 14964 4211
rect 14979 4186 15009 4202
rect 14878 4172 14908 4180
rect 14915 4178 15025 4186
rect 14878 4164 14923 4172
rect 14610 4146 14629 4148
rect 14644 4146 14690 4148
rect 14610 4130 14690 4146
rect 14717 4144 14752 4157
rect 14793 4154 14830 4157
rect 14793 4152 14835 4154
rect 14722 4141 14752 4144
rect 14731 4137 14738 4141
rect 14738 4136 14739 4137
rect 14697 4130 14707 4136
rect 14456 4122 14491 4130
rect 14456 4096 14457 4122
rect 14464 4096 14491 4122
rect 14399 4078 14429 4092
rect 14456 4088 14491 4096
rect 14493 4122 14534 4130
rect 14493 4096 14508 4122
rect 14515 4096 14534 4122
rect 14598 4118 14629 4130
rect 14644 4118 14747 4130
rect 14759 4120 14785 4146
rect 14800 4141 14830 4152
rect 14862 4148 14924 4164
rect 14862 4146 14908 4148
rect 14862 4130 14924 4146
rect 14936 4130 14942 4178
rect 14945 4170 15025 4178
rect 14945 4168 14964 4170
rect 14979 4168 15013 4170
rect 14945 4152 15025 4168
rect 14945 4130 14964 4152
rect 14979 4136 15009 4152
rect 15037 4146 15043 4220
rect 15046 4146 15065 4290
rect 15080 4146 15086 4290
rect 15095 4220 15108 4290
rect 15160 4286 15182 4290
rect 15153 4264 15182 4278
rect 15235 4264 15251 4278
rect 15289 4274 15295 4276
rect 15302 4274 15410 4290
rect 15417 4274 15423 4276
rect 15431 4274 15446 4290
rect 15512 4284 15531 4287
rect 15153 4262 15251 4264
rect 15278 4262 15446 4274
rect 15461 4264 15477 4278
rect 15512 4265 15534 4284
rect 15544 4278 15560 4279
rect 15543 4276 15560 4278
rect 15544 4271 15560 4276
rect 15534 4264 15540 4265
rect 15543 4264 15572 4271
rect 15461 4263 15572 4264
rect 15461 4262 15578 4263
rect 15137 4254 15188 4262
rect 15235 4254 15269 4262
rect 15137 4242 15162 4254
rect 15169 4242 15188 4254
rect 15242 4252 15269 4254
rect 15278 4252 15499 4262
rect 15534 4259 15540 4262
rect 15242 4248 15499 4252
rect 15137 4234 15188 4242
rect 15235 4234 15499 4248
rect 15543 4254 15578 4262
rect 15089 4186 15108 4220
rect 15153 4226 15182 4234
rect 15153 4220 15170 4226
rect 15153 4218 15187 4220
rect 15235 4218 15251 4234
rect 15252 4224 15460 4234
rect 15461 4224 15477 4234
rect 15525 4230 15540 4245
rect 15543 4242 15544 4254
rect 15551 4242 15578 4254
rect 15543 4234 15578 4242
rect 15543 4233 15572 4234
rect 15263 4220 15477 4224
rect 15278 4218 15477 4220
rect 15512 4220 15525 4230
rect 15543 4220 15560 4233
rect 15512 4218 15560 4220
rect 15154 4214 15187 4218
rect 15150 4212 15187 4214
rect 15150 4211 15217 4212
rect 15150 4206 15181 4211
rect 15187 4206 15217 4211
rect 15150 4202 15217 4206
rect 15123 4199 15217 4202
rect 15123 4192 15172 4199
rect 15123 4186 15153 4192
rect 15172 4187 15177 4192
rect 15089 4170 15169 4186
rect 15181 4178 15217 4199
rect 15278 4194 15467 4218
rect 15512 4217 15559 4218
rect 15525 4212 15559 4217
rect 15293 4191 15467 4194
rect 15286 4188 15467 4191
rect 15495 4211 15559 4212
rect 15089 4168 15108 4170
rect 15123 4168 15157 4170
rect 15089 4152 15169 4168
rect 15089 4146 15108 4152
rect 14805 4120 14908 4130
rect 14759 4118 14908 4120
rect 14929 4118 14964 4130
rect 14598 4116 14760 4118
rect 14610 4096 14629 4116
rect 14644 4114 14674 4116
rect 14493 4088 14534 4096
rect 14616 4092 14629 4096
rect 14681 4100 14760 4116
rect 14792 4116 14964 4118
rect 14792 4100 14871 4116
rect 14878 4114 14908 4116
rect 14456 4078 14485 4088
rect 14499 4078 14528 4088
rect 14543 4078 14573 4092
rect 14616 4078 14659 4092
rect 14681 4088 14871 4100
rect 14936 4096 14942 4116
rect 14666 4078 14696 4088
rect 14697 4078 14855 4088
rect 14859 4078 14889 4088
rect 14893 4078 14923 4092
rect 14951 4078 14964 4116
rect 15036 4130 15065 4146
rect 15079 4130 15108 4146
rect 15123 4136 15153 4152
rect 15181 4130 15187 4178
rect 15190 4172 15209 4178
rect 15224 4172 15254 4180
rect 15190 4164 15254 4172
rect 15190 4148 15270 4164
rect 15286 4157 15348 4188
rect 15364 4157 15426 4188
rect 15495 4186 15544 4211
rect 15559 4186 15589 4202
rect 15458 4172 15488 4180
rect 15495 4178 15605 4186
rect 15458 4164 15503 4172
rect 15190 4146 15209 4148
rect 15224 4146 15270 4148
rect 15190 4130 15270 4146
rect 15297 4144 15332 4157
rect 15373 4154 15410 4157
rect 15373 4152 15415 4154
rect 15302 4141 15332 4144
rect 15311 4137 15318 4141
rect 15318 4136 15319 4137
rect 15277 4130 15287 4136
rect 15036 4122 15071 4130
rect 15036 4096 15037 4122
rect 15044 4096 15071 4122
rect 14979 4078 15009 4092
rect 15036 4088 15071 4096
rect 15073 4122 15114 4130
rect 15073 4096 15088 4122
rect 15095 4096 15114 4122
rect 15178 4118 15209 4130
rect 15224 4118 15327 4130
rect 15339 4120 15365 4146
rect 15380 4141 15410 4152
rect 15442 4148 15504 4164
rect 15442 4146 15488 4148
rect 15442 4130 15504 4146
rect 15516 4130 15522 4178
rect 15525 4170 15605 4178
rect 15525 4168 15544 4170
rect 15559 4168 15593 4170
rect 15525 4152 15605 4168
rect 15525 4130 15544 4152
rect 15559 4136 15589 4152
rect 15617 4146 15623 4220
rect 15626 4146 15645 4290
rect 15660 4146 15666 4290
rect 15675 4220 15688 4290
rect 15740 4286 15762 4290
rect 15733 4264 15762 4278
rect 15815 4264 15831 4278
rect 15869 4274 15875 4276
rect 15882 4274 15990 4290
rect 15997 4274 16003 4276
rect 16011 4274 16026 4290
rect 16092 4284 16111 4287
rect 15733 4262 15831 4264
rect 15858 4262 16026 4274
rect 16041 4264 16057 4278
rect 16092 4265 16114 4284
rect 16124 4278 16140 4279
rect 16123 4276 16140 4278
rect 16124 4271 16140 4276
rect 16114 4264 16120 4265
rect 16123 4264 16152 4271
rect 16041 4263 16152 4264
rect 16041 4262 16158 4263
rect 15717 4254 15768 4262
rect 15815 4254 15849 4262
rect 15717 4242 15742 4254
rect 15749 4242 15768 4254
rect 15822 4252 15849 4254
rect 15858 4252 16079 4262
rect 16114 4259 16120 4262
rect 15822 4248 16079 4252
rect 15717 4234 15768 4242
rect 15815 4234 16079 4248
rect 16123 4254 16158 4262
rect 15669 4186 15688 4220
rect 15733 4226 15762 4234
rect 15733 4220 15750 4226
rect 15733 4218 15767 4220
rect 15815 4218 15831 4234
rect 15832 4224 16040 4234
rect 16041 4224 16057 4234
rect 16105 4230 16120 4245
rect 16123 4242 16124 4254
rect 16131 4242 16158 4254
rect 16123 4234 16158 4242
rect 16123 4233 16152 4234
rect 15843 4220 16057 4224
rect 15858 4218 16057 4220
rect 16092 4220 16105 4230
rect 16123 4220 16140 4233
rect 16092 4218 16140 4220
rect 15734 4214 15767 4218
rect 15730 4212 15767 4214
rect 15730 4211 15797 4212
rect 15730 4206 15761 4211
rect 15767 4206 15797 4211
rect 15730 4202 15797 4206
rect 15703 4199 15797 4202
rect 15703 4192 15752 4199
rect 15703 4186 15733 4192
rect 15752 4187 15757 4192
rect 15669 4170 15749 4186
rect 15761 4178 15797 4199
rect 15858 4194 16047 4218
rect 16092 4217 16139 4218
rect 16105 4212 16139 4217
rect 15873 4191 16047 4194
rect 15866 4188 16047 4191
rect 16075 4211 16139 4212
rect 15669 4168 15688 4170
rect 15703 4168 15737 4170
rect 15669 4152 15749 4168
rect 15669 4146 15688 4152
rect 15385 4120 15488 4130
rect 15339 4118 15488 4120
rect 15509 4118 15544 4130
rect 15178 4116 15340 4118
rect 15190 4096 15209 4116
rect 15224 4114 15254 4116
rect 15073 4088 15114 4096
rect 15196 4092 15209 4096
rect 15261 4100 15340 4116
rect 15372 4116 15544 4118
rect 15372 4100 15451 4116
rect 15458 4114 15488 4116
rect 15036 4078 15065 4088
rect 15079 4078 15108 4088
rect 15123 4078 15153 4092
rect 15196 4078 15239 4092
rect 15261 4088 15451 4100
rect 15516 4096 15522 4116
rect 15246 4078 15276 4088
rect 15277 4078 15435 4088
rect 15439 4078 15469 4088
rect 15473 4078 15503 4092
rect 15531 4078 15544 4116
rect 15616 4130 15645 4146
rect 15659 4130 15688 4146
rect 15703 4136 15733 4152
rect 15761 4130 15767 4178
rect 15770 4172 15789 4178
rect 15804 4172 15834 4180
rect 15770 4164 15834 4172
rect 15770 4148 15850 4164
rect 15866 4157 15928 4188
rect 15944 4157 16006 4188
rect 16075 4186 16124 4211
rect 16139 4186 16169 4202
rect 16038 4172 16068 4180
rect 16075 4178 16185 4186
rect 16038 4164 16083 4172
rect 15770 4146 15789 4148
rect 15804 4146 15850 4148
rect 15770 4130 15850 4146
rect 15877 4144 15912 4157
rect 15953 4154 15990 4157
rect 15953 4152 15995 4154
rect 15882 4141 15912 4144
rect 15891 4137 15898 4141
rect 15898 4136 15899 4137
rect 15857 4130 15867 4136
rect 15616 4122 15651 4130
rect 15616 4096 15617 4122
rect 15624 4096 15651 4122
rect 15559 4078 15589 4092
rect 15616 4088 15651 4096
rect 15653 4122 15694 4130
rect 15653 4096 15668 4122
rect 15675 4096 15694 4122
rect 15758 4118 15789 4130
rect 15804 4118 15907 4130
rect 15919 4120 15945 4146
rect 15960 4141 15990 4152
rect 16022 4148 16084 4164
rect 16022 4146 16068 4148
rect 16022 4130 16084 4146
rect 16096 4130 16102 4178
rect 16105 4170 16185 4178
rect 16105 4168 16124 4170
rect 16139 4168 16173 4170
rect 16105 4152 16185 4168
rect 16105 4130 16124 4152
rect 16139 4136 16169 4152
rect 16197 4146 16203 4220
rect 16206 4146 16225 4290
rect 16240 4146 16246 4290
rect 16255 4220 16268 4290
rect 16320 4286 16342 4290
rect 16313 4264 16342 4278
rect 16395 4264 16411 4278
rect 16449 4274 16455 4276
rect 16462 4274 16570 4290
rect 16577 4274 16583 4276
rect 16591 4274 16606 4290
rect 16672 4284 16691 4287
rect 16313 4262 16411 4264
rect 16438 4262 16606 4274
rect 16621 4264 16637 4278
rect 16672 4265 16694 4284
rect 16704 4278 16720 4279
rect 16703 4276 16720 4278
rect 16704 4271 16720 4276
rect 16694 4264 16700 4265
rect 16703 4264 16732 4271
rect 16621 4263 16732 4264
rect 16621 4262 16738 4263
rect 16297 4254 16348 4262
rect 16395 4254 16429 4262
rect 16297 4242 16322 4254
rect 16329 4242 16348 4254
rect 16402 4252 16429 4254
rect 16438 4252 16659 4262
rect 16694 4259 16700 4262
rect 16402 4248 16659 4252
rect 16297 4234 16348 4242
rect 16395 4234 16659 4248
rect 16703 4254 16738 4262
rect 16249 4186 16268 4220
rect 16313 4226 16342 4234
rect 16313 4220 16330 4226
rect 16313 4218 16347 4220
rect 16395 4218 16411 4234
rect 16412 4224 16620 4234
rect 16621 4224 16637 4234
rect 16685 4230 16700 4245
rect 16703 4242 16704 4254
rect 16711 4242 16738 4254
rect 16703 4234 16738 4242
rect 16703 4233 16732 4234
rect 16423 4220 16637 4224
rect 16438 4218 16637 4220
rect 16672 4220 16685 4230
rect 16703 4220 16720 4233
rect 16672 4218 16720 4220
rect 16314 4214 16347 4218
rect 16310 4212 16347 4214
rect 16310 4211 16377 4212
rect 16310 4206 16341 4211
rect 16347 4206 16377 4211
rect 16310 4202 16377 4206
rect 16283 4199 16377 4202
rect 16283 4192 16332 4199
rect 16283 4186 16313 4192
rect 16332 4187 16337 4192
rect 16249 4170 16329 4186
rect 16341 4178 16377 4199
rect 16438 4194 16627 4218
rect 16672 4217 16719 4218
rect 16685 4212 16719 4217
rect 16453 4191 16627 4194
rect 16446 4188 16627 4191
rect 16655 4211 16719 4212
rect 16249 4168 16268 4170
rect 16283 4168 16317 4170
rect 16249 4152 16329 4168
rect 16249 4146 16268 4152
rect 15965 4120 16068 4130
rect 15919 4118 16068 4120
rect 16089 4118 16124 4130
rect 15758 4116 15920 4118
rect 15770 4096 15789 4116
rect 15804 4114 15834 4116
rect 15653 4088 15694 4096
rect 15776 4092 15789 4096
rect 15841 4100 15920 4116
rect 15952 4116 16124 4118
rect 15952 4100 16031 4116
rect 16038 4114 16068 4116
rect 15616 4078 15645 4088
rect 15659 4078 15688 4088
rect 15703 4078 15733 4092
rect 15776 4078 15819 4092
rect 15841 4088 16031 4100
rect 16096 4096 16102 4116
rect 15826 4078 15856 4088
rect 15857 4078 16015 4088
rect 16019 4078 16049 4088
rect 16053 4078 16083 4092
rect 16111 4078 16124 4116
rect 16196 4130 16225 4146
rect 16239 4130 16268 4146
rect 16283 4136 16313 4152
rect 16341 4130 16347 4178
rect 16350 4172 16369 4178
rect 16384 4172 16414 4180
rect 16350 4164 16414 4172
rect 16350 4148 16430 4164
rect 16446 4157 16508 4188
rect 16524 4157 16586 4188
rect 16655 4186 16704 4211
rect 16719 4186 16749 4202
rect 16618 4172 16648 4180
rect 16655 4178 16765 4186
rect 16618 4164 16663 4172
rect 16350 4146 16369 4148
rect 16384 4146 16430 4148
rect 16350 4130 16430 4146
rect 16457 4144 16492 4157
rect 16533 4154 16570 4157
rect 16533 4152 16575 4154
rect 16462 4141 16492 4144
rect 16471 4137 16478 4141
rect 16478 4136 16479 4137
rect 16437 4130 16447 4136
rect 16196 4122 16231 4130
rect 16196 4096 16197 4122
rect 16204 4096 16231 4122
rect 16139 4078 16169 4092
rect 16196 4088 16231 4096
rect 16233 4122 16274 4130
rect 16233 4096 16248 4122
rect 16255 4096 16274 4122
rect 16338 4118 16369 4130
rect 16384 4118 16487 4130
rect 16499 4120 16525 4146
rect 16540 4141 16570 4152
rect 16602 4148 16664 4164
rect 16602 4146 16648 4148
rect 16602 4130 16664 4146
rect 16676 4130 16682 4178
rect 16685 4170 16765 4178
rect 16685 4168 16704 4170
rect 16719 4168 16753 4170
rect 16685 4152 16765 4168
rect 16685 4130 16704 4152
rect 16719 4136 16749 4152
rect 16777 4146 16783 4220
rect 16786 4146 16805 4290
rect 16820 4146 16826 4290
rect 16835 4220 16848 4290
rect 16900 4286 16922 4290
rect 16893 4264 16922 4278
rect 16975 4264 16991 4278
rect 17029 4274 17035 4276
rect 17042 4274 17150 4290
rect 17157 4274 17163 4276
rect 17171 4274 17186 4290
rect 17252 4284 17271 4287
rect 16893 4262 16991 4264
rect 17018 4262 17186 4274
rect 17201 4264 17217 4278
rect 17252 4265 17274 4284
rect 17284 4278 17300 4279
rect 17283 4276 17300 4278
rect 17284 4271 17300 4276
rect 17274 4264 17280 4265
rect 17283 4264 17312 4271
rect 17201 4263 17312 4264
rect 17201 4262 17318 4263
rect 16877 4254 16928 4262
rect 16975 4254 17009 4262
rect 16877 4242 16902 4254
rect 16909 4242 16928 4254
rect 16982 4252 17009 4254
rect 17018 4252 17239 4262
rect 17274 4259 17280 4262
rect 16982 4248 17239 4252
rect 16877 4234 16928 4242
rect 16975 4234 17239 4248
rect 17283 4254 17318 4262
rect 16829 4186 16848 4220
rect 16893 4226 16922 4234
rect 16893 4220 16910 4226
rect 16893 4218 16927 4220
rect 16975 4218 16991 4234
rect 16992 4224 17200 4234
rect 17201 4224 17217 4234
rect 17265 4230 17280 4245
rect 17283 4242 17284 4254
rect 17291 4242 17318 4254
rect 17283 4234 17318 4242
rect 17283 4233 17312 4234
rect 17003 4220 17217 4224
rect 17018 4218 17217 4220
rect 17252 4220 17265 4230
rect 17283 4220 17300 4233
rect 17252 4218 17300 4220
rect 16894 4214 16927 4218
rect 16890 4212 16927 4214
rect 16890 4211 16957 4212
rect 16890 4206 16921 4211
rect 16927 4206 16957 4211
rect 16890 4202 16957 4206
rect 16863 4199 16957 4202
rect 16863 4192 16912 4199
rect 16863 4186 16893 4192
rect 16912 4187 16917 4192
rect 16829 4170 16909 4186
rect 16921 4178 16957 4199
rect 17018 4194 17207 4218
rect 17252 4217 17299 4218
rect 17265 4212 17299 4217
rect 17033 4191 17207 4194
rect 17026 4188 17207 4191
rect 17235 4211 17299 4212
rect 16829 4168 16848 4170
rect 16863 4168 16897 4170
rect 16829 4152 16909 4168
rect 16829 4146 16848 4152
rect 16545 4120 16648 4130
rect 16499 4118 16648 4120
rect 16669 4118 16704 4130
rect 16338 4116 16500 4118
rect 16350 4096 16369 4116
rect 16384 4114 16414 4116
rect 16233 4088 16274 4096
rect 16356 4092 16369 4096
rect 16421 4100 16500 4116
rect 16532 4116 16704 4118
rect 16532 4100 16611 4116
rect 16618 4114 16648 4116
rect 16196 4078 16225 4088
rect 16239 4078 16268 4088
rect 16283 4078 16313 4092
rect 16356 4078 16399 4092
rect 16421 4088 16611 4100
rect 16676 4096 16682 4116
rect 16406 4078 16436 4088
rect 16437 4078 16595 4088
rect 16599 4078 16629 4088
rect 16633 4078 16663 4092
rect 16691 4078 16704 4116
rect 16776 4130 16805 4146
rect 16819 4130 16848 4146
rect 16863 4136 16893 4152
rect 16921 4130 16927 4178
rect 16930 4172 16949 4178
rect 16964 4172 16994 4180
rect 16930 4164 16994 4172
rect 16930 4148 17010 4164
rect 17026 4157 17088 4188
rect 17104 4157 17166 4188
rect 17235 4186 17284 4211
rect 17299 4186 17329 4202
rect 17198 4172 17228 4180
rect 17235 4178 17345 4186
rect 17198 4164 17243 4172
rect 16930 4146 16949 4148
rect 16964 4146 17010 4148
rect 16930 4130 17010 4146
rect 17037 4144 17072 4157
rect 17113 4154 17150 4157
rect 17113 4152 17155 4154
rect 17042 4141 17072 4144
rect 17051 4137 17058 4141
rect 17058 4136 17059 4137
rect 17017 4130 17027 4136
rect 16776 4122 16811 4130
rect 16776 4096 16777 4122
rect 16784 4096 16811 4122
rect 16719 4078 16749 4092
rect 16776 4088 16811 4096
rect 16813 4122 16854 4130
rect 16813 4096 16828 4122
rect 16835 4096 16854 4122
rect 16918 4118 16949 4130
rect 16964 4118 17067 4130
rect 17079 4120 17105 4146
rect 17120 4141 17150 4152
rect 17182 4148 17244 4164
rect 17182 4146 17228 4148
rect 17182 4130 17244 4146
rect 17256 4130 17262 4178
rect 17265 4170 17345 4178
rect 17265 4168 17284 4170
rect 17299 4168 17333 4170
rect 17265 4152 17345 4168
rect 17265 4130 17284 4152
rect 17299 4136 17329 4152
rect 17357 4146 17363 4220
rect 17366 4146 17385 4290
rect 17400 4146 17406 4290
rect 17415 4220 17428 4290
rect 17480 4286 17502 4290
rect 17473 4264 17502 4278
rect 17555 4264 17571 4278
rect 17609 4274 17615 4276
rect 17622 4274 17730 4290
rect 17737 4274 17743 4276
rect 17751 4274 17766 4290
rect 17832 4284 17851 4287
rect 17473 4262 17571 4264
rect 17598 4262 17766 4274
rect 17781 4264 17797 4278
rect 17832 4265 17854 4284
rect 17864 4278 17880 4279
rect 17863 4276 17880 4278
rect 17864 4271 17880 4276
rect 17854 4264 17860 4265
rect 17863 4264 17892 4271
rect 17781 4263 17892 4264
rect 17781 4262 17898 4263
rect 17457 4254 17508 4262
rect 17555 4254 17589 4262
rect 17457 4242 17482 4254
rect 17489 4242 17508 4254
rect 17562 4252 17589 4254
rect 17598 4252 17819 4262
rect 17854 4259 17860 4262
rect 17562 4248 17819 4252
rect 17457 4234 17508 4242
rect 17555 4234 17819 4248
rect 17863 4254 17898 4262
rect 17409 4186 17428 4220
rect 17473 4226 17502 4234
rect 17473 4220 17490 4226
rect 17473 4218 17507 4220
rect 17555 4218 17571 4234
rect 17572 4224 17780 4234
rect 17781 4224 17797 4234
rect 17845 4230 17860 4245
rect 17863 4242 17864 4254
rect 17871 4242 17898 4254
rect 17863 4234 17898 4242
rect 17863 4233 17892 4234
rect 17583 4220 17797 4224
rect 17598 4218 17797 4220
rect 17832 4220 17845 4230
rect 17863 4220 17880 4233
rect 17832 4218 17880 4220
rect 17474 4214 17507 4218
rect 17470 4212 17507 4214
rect 17470 4211 17537 4212
rect 17470 4206 17501 4211
rect 17507 4206 17537 4211
rect 17470 4202 17537 4206
rect 17443 4199 17537 4202
rect 17443 4192 17492 4199
rect 17443 4186 17473 4192
rect 17492 4187 17497 4192
rect 17409 4170 17489 4186
rect 17501 4178 17537 4199
rect 17598 4194 17787 4218
rect 17832 4217 17879 4218
rect 17845 4212 17879 4217
rect 17613 4191 17787 4194
rect 17606 4188 17787 4191
rect 17815 4211 17879 4212
rect 17409 4168 17428 4170
rect 17443 4168 17477 4170
rect 17409 4152 17489 4168
rect 17409 4146 17428 4152
rect 17125 4120 17228 4130
rect 17079 4118 17228 4120
rect 17249 4118 17284 4130
rect 16918 4116 17080 4118
rect 16930 4096 16949 4116
rect 16964 4114 16994 4116
rect 16813 4088 16854 4096
rect 16936 4092 16949 4096
rect 17001 4100 17080 4116
rect 17112 4116 17284 4118
rect 17112 4100 17191 4116
rect 17198 4114 17228 4116
rect 16776 4078 16805 4088
rect 16819 4078 16848 4088
rect 16863 4078 16893 4092
rect 16936 4078 16979 4092
rect 17001 4088 17191 4100
rect 17256 4096 17262 4116
rect 16986 4078 17016 4088
rect 17017 4078 17175 4088
rect 17179 4078 17209 4088
rect 17213 4078 17243 4092
rect 17271 4078 17284 4116
rect 17356 4130 17385 4146
rect 17399 4130 17428 4146
rect 17443 4136 17473 4152
rect 17501 4130 17507 4178
rect 17510 4172 17529 4178
rect 17544 4172 17574 4180
rect 17510 4164 17574 4172
rect 17510 4148 17590 4164
rect 17606 4157 17668 4188
rect 17684 4157 17746 4188
rect 17815 4186 17864 4211
rect 17879 4186 17909 4202
rect 17778 4172 17808 4180
rect 17815 4178 17925 4186
rect 17778 4164 17823 4172
rect 17510 4146 17529 4148
rect 17544 4146 17590 4148
rect 17510 4130 17590 4146
rect 17617 4144 17652 4157
rect 17693 4154 17730 4157
rect 17693 4152 17735 4154
rect 17622 4141 17652 4144
rect 17631 4137 17638 4141
rect 17638 4136 17639 4137
rect 17597 4130 17607 4136
rect 17356 4122 17391 4130
rect 17356 4096 17357 4122
rect 17364 4096 17391 4122
rect 17299 4078 17329 4092
rect 17356 4088 17391 4096
rect 17393 4122 17434 4130
rect 17393 4096 17408 4122
rect 17415 4096 17434 4122
rect 17498 4118 17529 4130
rect 17544 4118 17647 4130
rect 17659 4120 17685 4146
rect 17700 4141 17730 4152
rect 17762 4148 17824 4164
rect 17762 4146 17808 4148
rect 17762 4130 17824 4146
rect 17836 4130 17842 4178
rect 17845 4170 17925 4178
rect 17845 4168 17864 4170
rect 17879 4168 17913 4170
rect 17845 4152 17925 4168
rect 17845 4130 17864 4152
rect 17879 4136 17909 4152
rect 17937 4146 17943 4220
rect 17946 4146 17965 4290
rect 17980 4146 17986 4290
rect 17995 4220 18008 4290
rect 18060 4286 18082 4290
rect 18053 4264 18082 4278
rect 18135 4264 18151 4278
rect 18189 4274 18195 4276
rect 18202 4274 18310 4290
rect 18317 4274 18323 4276
rect 18331 4274 18346 4290
rect 18412 4284 18431 4287
rect 18053 4262 18151 4264
rect 18178 4262 18346 4274
rect 18361 4264 18377 4278
rect 18412 4265 18434 4284
rect 18444 4278 18460 4279
rect 18443 4276 18460 4278
rect 18444 4271 18460 4276
rect 18434 4264 18440 4265
rect 18443 4264 18472 4271
rect 18361 4263 18472 4264
rect 18361 4262 18478 4263
rect 18037 4254 18088 4262
rect 18135 4254 18169 4262
rect 18037 4242 18062 4254
rect 18069 4242 18088 4254
rect 18142 4252 18169 4254
rect 18178 4252 18399 4262
rect 18434 4259 18440 4262
rect 18142 4248 18399 4252
rect 18037 4234 18088 4242
rect 18135 4234 18399 4248
rect 18443 4254 18478 4262
rect 17989 4186 18008 4220
rect 18053 4226 18082 4234
rect 18053 4220 18070 4226
rect 18053 4218 18087 4220
rect 18135 4218 18151 4234
rect 18152 4224 18360 4234
rect 18361 4224 18377 4234
rect 18425 4230 18440 4245
rect 18443 4242 18444 4254
rect 18451 4242 18478 4254
rect 18443 4234 18478 4242
rect 18443 4233 18472 4234
rect 18163 4220 18377 4224
rect 18178 4218 18377 4220
rect 18412 4220 18425 4230
rect 18443 4220 18460 4233
rect 18412 4218 18460 4220
rect 18054 4214 18087 4218
rect 18050 4212 18087 4214
rect 18050 4211 18117 4212
rect 18050 4206 18081 4211
rect 18087 4206 18117 4211
rect 18050 4202 18117 4206
rect 18023 4199 18117 4202
rect 18023 4192 18072 4199
rect 18023 4186 18053 4192
rect 18072 4187 18077 4192
rect 17989 4170 18069 4186
rect 18081 4178 18117 4199
rect 18178 4194 18367 4218
rect 18412 4217 18459 4218
rect 18425 4212 18459 4217
rect 18193 4191 18367 4194
rect 18186 4188 18367 4191
rect 18395 4211 18459 4212
rect 17989 4168 18008 4170
rect 18023 4168 18057 4170
rect 17989 4152 18069 4168
rect 17989 4146 18008 4152
rect 17705 4120 17808 4130
rect 17659 4118 17808 4120
rect 17829 4118 17864 4130
rect 17498 4116 17660 4118
rect 17510 4096 17529 4116
rect 17544 4114 17574 4116
rect 17393 4088 17434 4096
rect 17516 4092 17529 4096
rect 17581 4100 17660 4116
rect 17692 4116 17864 4118
rect 17692 4100 17771 4116
rect 17778 4114 17808 4116
rect 17356 4078 17385 4088
rect 17399 4078 17428 4088
rect 17443 4078 17473 4092
rect 17516 4078 17559 4092
rect 17581 4088 17771 4100
rect 17836 4096 17842 4116
rect 17566 4078 17596 4088
rect 17597 4078 17755 4088
rect 17759 4078 17789 4088
rect 17793 4078 17823 4092
rect 17851 4078 17864 4116
rect 17936 4130 17965 4146
rect 17979 4130 18008 4146
rect 18023 4136 18053 4152
rect 18081 4130 18087 4178
rect 18090 4172 18109 4178
rect 18124 4172 18154 4180
rect 18090 4164 18154 4172
rect 18090 4148 18170 4164
rect 18186 4157 18248 4188
rect 18264 4157 18326 4188
rect 18395 4186 18444 4211
rect 18459 4186 18489 4202
rect 18358 4172 18388 4180
rect 18395 4178 18505 4186
rect 18358 4164 18403 4172
rect 18090 4146 18109 4148
rect 18124 4146 18170 4148
rect 18090 4130 18170 4146
rect 18197 4144 18232 4157
rect 18273 4154 18310 4157
rect 18273 4152 18315 4154
rect 18202 4141 18232 4144
rect 18211 4137 18218 4141
rect 18218 4136 18219 4137
rect 18177 4130 18187 4136
rect 17936 4122 17971 4130
rect 17936 4096 17937 4122
rect 17944 4096 17971 4122
rect 17879 4078 17909 4092
rect 17936 4088 17971 4096
rect 17973 4122 18014 4130
rect 17973 4096 17988 4122
rect 17995 4096 18014 4122
rect 18078 4118 18109 4130
rect 18124 4118 18227 4130
rect 18239 4120 18265 4146
rect 18280 4141 18310 4152
rect 18342 4148 18404 4164
rect 18342 4146 18388 4148
rect 18342 4130 18404 4146
rect 18416 4130 18422 4178
rect 18425 4170 18505 4178
rect 18425 4168 18444 4170
rect 18459 4168 18493 4170
rect 18425 4152 18505 4168
rect 18425 4130 18444 4152
rect 18459 4136 18489 4152
rect 18517 4146 18523 4220
rect 18532 4146 18545 4290
rect 18285 4120 18388 4130
rect 18239 4118 18388 4120
rect 18409 4118 18444 4130
rect 18078 4116 18240 4118
rect 18090 4096 18109 4116
rect 18124 4114 18154 4116
rect 17973 4088 18014 4096
rect 18096 4092 18109 4096
rect 18161 4100 18240 4116
rect 18272 4116 18444 4118
rect 18272 4100 18351 4116
rect 18358 4114 18388 4116
rect 17936 4078 17965 4088
rect 17979 4078 18008 4088
rect 18023 4078 18053 4092
rect 18096 4078 18139 4092
rect 18161 4088 18351 4100
rect 18416 4096 18422 4116
rect 18146 4078 18176 4088
rect 18177 4078 18335 4088
rect 18339 4078 18369 4088
rect 18373 4078 18403 4092
rect 18431 4078 18444 4116
rect 18516 4130 18545 4146
rect 18516 4122 18551 4130
rect 18516 4096 18517 4122
rect 18524 4096 18551 4122
rect 18459 4078 18489 4092
rect 18516 4088 18551 4096
rect 18516 4078 18545 4088
rect -1 4072 18545 4078
rect 0 4064 18545 4072
rect 15 4034 28 4064
rect 43 4050 73 4064
rect 116 4050 159 4064
rect 166 4050 386 4064
rect 393 4050 423 4064
rect 83 4036 98 4048
rect 117 4036 130 4050
rect 198 4046 351 4050
rect 80 4034 102 4036
rect 180 4034 372 4046
rect 451 4034 464 4064
rect 479 4050 509 4064
rect 546 4034 565 4064
rect 580 4034 586 4064
rect 595 4034 608 4064
rect 623 4050 653 4064
rect 696 4050 739 4064
rect 746 4050 966 4064
rect 973 4050 1003 4064
rect 663 4036 678 4048
rect 697 4036 710 4050
rect 778 4046 931 4050
rect 660 4034 682 4036
rect 760 4034 952 4046
rect 1031 4034 1044 4064
rect 1059 4050 1089 4064
rect 1126 4034 1145 4064
rect 1160 4034 1166 4064
rect 1175 4034 1188 4064
rect 1203 4050 1233 4064
rect 1276 4050 1319 4064
rect 1326 4050 1546 4064
rect 1553 4050 1583 4064
rect 1243 4036 1258 4048
rect 1277 4036 1290 4050
rect 1358 4046 1511 4050
rect 1240 4034 1262 4036
rect 1340 4034 1532 4046
rect 1611 4034 1624 4064
rect 1639 4050 1669 4064
rect 1706 4034 1725 4064
rect 1740 4034 1746 4064
rect 1755 4034 1768 4064
rect 1783 4050 1813 4064
rect 1856 4050 1899 4064
rect 1906 4050 2126 4064
rect 2133 4050 2163 4064
rect 1823 4036 1838 4048
rect 1857 4036 1870 4050
rect 1938 4046 2091 4050
rect 1820 4034 1842 4036
rect 1920 4034 2112 4046
rect 2191 4034 2204 4064
rect 2219 4050 2249 4064
rect 2286 4034 2305 4064
rect 2320 4034 2326 4064
rect 2335 4034 2348 4064
rect 2363 4050 2393 4064
rect 2436 4050 2479 4064
rect 2486 4050 2706 4064
rect 2713 4050 2743 4064
rect 2403 4036 2418 4048
rect 2437 4036 2450 4050
rect 2518 4046 2671 4050
rect 2400 4034 2422 4036
rect 2500 4034 2692 4046
rect 2771 4034 2784 4064
rect 2799 4050 2829 4064
rect 2866 4034 2885 4064
rect 2900 4034 2906 4064
rect 2915 4034 2928 4064
rect 2943 4050 2973 4064
rect 3016 4050 3059 4064
rect 3066 4050 3286 4064
rect 3293 4050 3323 4064
rect 2983 4036 2998 4048
rect 3017 4036 3030 4050
rect 3098 4046 3251 4050
rect 2980 4034 3002 4036
rect 3080 4034 3272 4046
rect 3351 4034 3364 4064
rect 3379 4050 3409 4064
rect 3446 4034 3465 4064
rect 3480 4034 3486 4064
rect 3495 4034 3508 4064
rect 3523 4050 3553 4064
rect 3596 4050 3639 4064
rect 3646 4050 3866 4064
rect 3873 4050 3903 4064
rect 3563 4036 3578 4048
rect 3597 4036 3610 4050
rect 3678 4046 3831 4050
rect 3560 4034 3582 4036
rect 3660 4034 3852 4046
rect 3931 4034 3944 4064
rect 3959 4050 3989 4064
rect 4026 4034 4045 4064
rect 4060 4034 4066 4064
rect 4075 4034 4088 4064
rect 4103 4050 4133 4064
rect 4176 4050 4219 4064
rect 4226 4050 4446 4064
rect 4453 4050 4483 4064
rect 4143 4036 4158 4048
rect 4177 4036 4190 4050
rect 4258 4046 4411 4050
rect 4140 4034 4162 4036
rect 4240 4034 4432 4046
rect 4511 4034 4524 4064
rect 4539 4050 4569 4064
rect 4606 4034 4625 4064
rect 4640 4034 4646 4064
rect 4655 4034 4668 4064
rect 4683 4050 4713 4064
rect 4756 4050 4799 4064
rect 4806 4050 5026 4064
rect 5033 4050 5063 4064
rect 4723 4036 4738 4048
rect 4757 4036 4770 4050
rect 4838 4046 4991 4050
rect 4720 4034 4742 4036
rect 4820 4034 5012 4046
rect 5091 4034 5104 4064
rect 5119 4050 5149 4064
rect 5186 4034 5205 4064
rect 5220 4034 5226 4064
rect 5235 4034 5248 4064
rect 5263 4050 5293 4064
rect 5336 4050 5379 4064
rect 5386 4050 5606 4064
rect 5613 4050 5643 4064
rect 5303 4036 5318 4048
rect 5337 4036 5350 4050
rect 5418 4046 5571 4050
rect 5300 4034 5322 4036
rect 5400 4034 5592 4046
rect 5671 4034 5684 4064
rect 5699 4050 5729 4064
rect 5766 4034 5785 4064
rect 5800 4034 5806 4064
rect 5815 4034 5828 4064
rect 5843 4050 5873 4064
rect 5916 4050 5959 4064
rect 5966 4050 6186 4064
rect 6193 4050 6223 4064
rect 5883 4036 5898 4048
rect 5917 4036 5930 4050
rect 5998 4046 6151 4050
rect 5880 4034 5902 4036
rect 5980 4034 6172 4046
rect 6251 4034 6264 4064
rect 6279 4050 6309 4064
rect 6346 4034 6365 4064
rect 6380 4034 6386 4064
rect 6395 4034 6408 4064
rect 6423 4050 6453 4064
rect 6496 4050 6539 4064
rect 6546 4050 6766 4064
rect 6773 4050 6803 4064
rect 6463 4036 6478 4048
rect 6497 4036 6510 4050
rect 6578 4046 6731 4050
rect 6460 4034 6482 4036
rect 6560 4034 6752 4046
rect 6831 4034 6844 4064
rect 6859 4050 6889 4064
rect 6926 4034 6945 4064
rect 6960 4034 6966 4064
rect 6975 4034 6988 4064
rect 7003 4050 7033 4064
rect 7076 4050 7119 4064
rect 7126 4050 7346 4064
rect 7353 4050 7383 4064
rect 7043 4036 7058 4048
rect 7077 4036 7090 4050
rect 7158 4046 7311 4050
rect 7040 4034 7062 4036
rect 7140 4034 7332 4046
rect 7411 4034 7424 4064
rect 7439 4050 7469 4064
rect 7506 4034 7525 4064
rect 7540 4034 7546 4064
rect 7555 4034 7568 4064
rect 7583 4050 7613 4064
rect 7656 4050 7699 4064
rect 7706 4050 7926 4064
rect 7933 4050 7963 4064
rect 7623 4036 7638 4048
rect 7657 4036 7670 4050
rect 7738 4046 7891 4050
rect 7620 4034 7642 4036
rect 7720 4034 7912 4046
rect 7991 4034 8004 4064
rect 8019 4050 8049 4064
rect 8086 4034 8105 4064
rect 8120 4034 8126 4064
rect 8135 4034 8148 4064
rect 8163 4050 8193 4064
rect 8236 4050 8279 4064
rect 8286 4050 8506 4064
rect 8513 4050 8543 4064
rect 8203 4036 8218 4048
rect 8237 4036 8250 4050
rect 8318 4046 8471 4050
rect 8200 4034 8222 4036
rect 8300 4034 8492 4046
rect 8571 4034 8584 4064
rect 8599 4050 8629 4064
rect 8666 4034 8685 4064
rect 8700 4034 8706 4064
rect 8715 4034 8728 4064
rect 8743 4050 8773 4064
rect 8816 4050 8859 4064
rect 8866 4050 9086 4064
rect 9093 4050 9123 4064
rect 8783 4036 8798 4048
rect 8817 4036 8830 4050
rect 8898 4046 9051 4050
rect 8780 4034 8802 4036
rect 8880 4034 9072 4046
rect 9151 4034 9164 4064
rect 9179 4050 9209 4064
rect 9246 4034 9265 4064
rect 9280 4034 9286 4064
rect 9295 4034 9308 4064
rect 9323 4050 9353 4064
rect 9396 4050 9439 4064
rect 9446 4050 9666 4064
rect 9673 4050 9703 4064
rect 9363 4036 9378 4048
rect 9397 4036 9410 4050
rect 9478 4046 9631 4050
rect 9360 4034 9382 4036
rect 9460 4034 9652 4046
rect 9731 4034 9744 4064
rect 9759 4050 9789 4064
rect 9826 4034 9845 4064
rect 9860 4034 9866 4064
rect 9875 4034 9888 4064
rect 9903 4050 9933 4064
rect 9976 4050 10019 4064
rect 10026 4050 10246 4064
rect 10253 4050 10283 4064
rect 9943 4036 9958 4048
rect 9977 4036 9990 4050
rect 10058 4046 10211 4050
rect 9940 4034 9962 4036
rect 10040 4034 10232 4046
rect 10311 4034 10324 4064
rect 10339 4050 10369 4064
rect 10406 4034 10425 4064
rect 10440 4034 10446 4064
rect 10455 4034 10468 4064
rect 10483 4050 10513 4064
rect 10556 4050 10599 4064
rect 10606 4050 10826 4064
rect 10833 4050 10863 4064
rect 10523 4036 10538 4048
rect 10557 4036 10570 4050
rect 10638 4046 10791 4050
rect 10520 4034 10542 4036
rect 10620 4034 10812 4046
rect 10891 4034 10904 4064
rect 10919 4050 10949 4064
rect 10986 4034 11005 4064
rect 11020 4034 11026 4064
rect 11035 4034 11048 4064
rect 11063 4050 11093 4064
rect 11136 4050 11179 4064
rect 11186 4050 11406 4064
rect 11413 4050 11443 4064
rect 11103 4036 11118 4048
rect 11137 4036 11150 4050
rect 11218 4046 11371 4050
rect 11100 4034 11122 4036
rect 11200 4034 11392 4046
rect 11471 4034 11484 4064
rect 11499 4050 11529 4064
rect 11566 4034 11585 4064
rect 11600 4034 11606 4064
rect 11615 4034 11628 4064
rect 11643 4050 11673 4064
rect 11716 4050 11759 4064
rect 11766 4050 11986 4064
rect 11993 4050 12023 4064
rect 11683 4036 11698 4048
rect 11717 4036 11730 4050
rect 11798 4046 11951 4050
rect 11680 4034 11702 4036
rect 11780 4034 11972 4046
rect 12051 4034 12064 4064
rect 12079 4050 12109 4064
rect 12146 4034 12165 4064
rect 12180 4034 12186 4064
rect 12195 4034 12208 4064
rect 12223 4050 12253 4064
rect 12296 4050 12339 4064
rect 12346 4050 12566 4064
rect 12573 4050 12603 4064
rect 12263 4036 12278 4048
rect 12297 4036 12310 4050
rect 12378 4046 12531 4050
rect 12260 4034 12282 4036
rect 12360 4034 12552 4046
rect 12631 4034 12644 4064
rect 12659 4050 12689 4064
rect 12726 4034 12745 4064
rect 12760 4034 12766 4064
rect 12775 4034 12788 4064
rect 12803 4050 12833 4064
rect 12876 4050 12919 4064
rect 12926 4050 13146 4064
rect 13153 4050 13183 4064
rect 12843 4036 12858 4048
rect 12877 4036 12890 4050
rect 12958 4046 13111 4050
rect 12840 4034 12862 4036
rect 12940 4034 13132 4046
rect 13211 4034 13224 4064
rect 13239 4050 13269 4064
rect 13306 4034 13325 4064
rect 13340 4034 13346 4064
rect 13355 4034 13368 4064
rect 13383 4050 13413 4064
rect 13456 4050 13499 4064
rect 13506 4050 13726 4064
rect 13733 4050 13763 4064
rect 13423 4036 13438 4048
rect 13457 4036 13470 4050
rect 13538 4046 13691 4050
rect 13420 4034 13442 4036
rect 13520 4034 13712 4046
rect 13791 4034 13804 4064
rect 13819 4050 13849 4064
rect 13886 4034 13905 4064
rect 13920 4034 13926 4064
rect 13935 4034 13948 4064
rect 13963 4050 13993 4064
rect 14036 4050 14079 4064
rect 14086 4050 14306 4064
rect 14313 4050 14343 4064
rect 14003 4036 14018 4048
rect 14037 4036 14050 4050
rect 14118 4046 14271 4050
rect 14000 4034 14022 4036
rect 14100 4034 14292 4046
rect 14371 4034 14384 4064
rect 14399 4050 14429 4064
rect 14466 4034 14485 4064
rect 14500 4034 14506 4064
rect 14515 4034 14528 4064
rect 14543 4050 14573 4064
rect 14616 4050 14659 4064
rect 14666 4050 14886 4064
rect 14893 4050 14923 4064
rect 14583 4036 14598 4048
rect 14617 4036 14630 4050
rect 14698 4046 14851 4050
rect 14580 4034 14602 4036
rect 14680 4034 14872 4046
rect 14951 4034 14964 4064
rect 14979 4050 15009 4064
rect 15046 4034 15065 4064
rect 15080 4034 15086 4064
rect 15095 4034 15108 4064
rect 15123 4050 15153 4064
rect 15196 4050 15239 4064
rect 15246 4050 15466 4064
rect 15473 4050 15503 4064
rect 15163 4036 15178 4048
rect 15197 4036 15210 4050
rect 15278 4046 15431 4050
rect 15160 4034 15182 4036
rect 15260 4034 15452 4046
rect 15531 4034 15544 4064
rect 15559 4050 15589 4064
rect 15626 4034 15645 4064
rect 15660 4034 15666 4064
rect 15675 4034 15688 4064
rect 15703 4050 15733 4064
rect 15776 4050 15819 4064
rect 15826 4050 16046 4064
rect 16053 4050 16083 4064
rect 15743 4036 15758 4048
rect 15777 4036 15790 4050
rect 15858 4046 16011 4050
rect 15740 4034 15762 4036
rect 15840 4034 16032 4046
rect 16111 4034 16124 4064
rect 16139 4050 16169 4064
rect 16206 4034 16225 4064
rect 16240 4034 16246 4064
rect 16255 4034 16268 4064
rect 16283 4050 16313 4064
rect 16356 4050 16399 4064
rect 16406 4050 16626 4064
rect 16633 4050 16663 4064
rect 16323 4036 16338 4048
rect 16357 4036 16370 4050
rect 16438 4046 16591 4050
rect 16320 4034 16342 4036
rect 16420 4034 16612 4046
rect 16691 4034 16704 4064
rect 16719 4050 16749 4064
rect 16786 4034 16805 4064
rect 16820 4034 16826 4064
rect 16835 4034 16848 4064
rect 16863 4050 16893 4064
rect 16936 4050 16979 4064
rect 16986 4050 17206 4064
rect 17213 4050 17243 4064
rect 16903 4036 16918 4048
rect 16937 4036 16950 4050
rect 17018 4046 17171 4050
rect 16900 4034 16922 4036
rect 17000 4034 17192 4046
rect 17271 4034 17284 4064
rect 17299 4050 17329 4064
rect 17366 4034 17385 4064
rect 17400 4034 17406 4064
rect 17415 4034 17428 4064
rect 17443 4050 17473 4064
rect 17516 4050 17559 4064
rect 17566 4050 17786 4064
rect 17793 4050 17823 4064
rect 17483 4036 17498 4048
rect 17517 4036 17530 4050
rect 17598 4046 17751 4050
rect 17480 4034 17502 4036
rect 17580 4034 17772 4046
rect 17851 4034 17864 4064
rect 17879 4050 17909 4064
rect 17946 4034 17965 4064
rect 17980 4034 17986 4064
rect 17995 4034 18008 4064
rect 18023 4050 18053 4064
rect 18096 4050 18139 4064
rect 18146 4050 18366 4064
rect 18373 4050 18403 4064
rect 18063 4036 18078 4048
rect 18097 4036 18110 4050
rect 18178 4046 18331 4050
rect 18060 4034 18082 4036
rect 18160 4034 18352 4046
rect 18431 4034 18444 4064
rect 18459 4050 18489 4064
rect 18532 4034 18545 4064
rect 0 4020 18545 4034
rect 15 3950 28 4020
rect 80 4016 102 4020
rect 73 3994 102 4008
rect 155 3994 171 4008
rect 209 4004 215 4006
rect 222 4004 330 4020
rect 337 4004 343 4006
rect 351 4004 366 4020
rect 432 4014 451 4017
rect 73 3992 171 3994
rect 198 3992 366 4004
rect 381 3994 397 4008
rect 432 3995 454 4014
rect 464 4008 480 4009
rect 463 4006 480 4008
rect 464 4001 480 4006
rect 454 3994 460 3995
rect 463 3994 492 4001
rect 381 3993 492 3994
rect 381 3992 498 3993
rect 57 3984 108 3992
rect 155 3984 189 3992
rect 57 3972 82 3984
rect 89 3972 108 3984
rect 162 3982 189 3984
rect 198 3982 419 3992
rect 454 3989 460 3992
rect 162 3978 419 3982
rect 57 3964 108 3972
rect 155 3964 419 3978
rect 463 3984 498 3992
rect 9 3916 28 3950
rect 73 3956 102 3964
rect 73 3950 90 3956
rect 73 3948 107 3950
rect 155 3948 171 3964
rect 172 3954 380 3964
rect 381 3954 397 3964
rect 445 3960 460 3975
rect 463 3972 464 3984
rect 471 3972 498 3984
rect 463 3964 498 3972
rect 463 3963 492 3964
rect 183 3950 397 3954
rect 198 3948 397 3950
rect 432 3950 445 3960
rect 463 3950 480 3963
rect 432 3948 480 3950
rect 74 3944 107 3948
rect 70 3942 107 3944
rect 70 3941 137 3942
rect 70 3936 101 3941
rect 107 3936 137 3941
rect 70 3932 137 3936
rect 43 3929 137 3932
rect 43 3922 92 3929
rect 43 3916 73 3922
rect 92 3917 97 3922
rect 9 3900 89 3916
rect 101 3908 137 3929
rect 198 3924 387 3948
rect 432 3947 479 3948
rect 445 3942 479 3947
rect 213 3921 387 3924
rect 206 3918 387 3921
rect 415 3941 479 3942
rect 9 3898 28 3900
rect 43 3898 77 3900
rect 9 3882 89 3898
rect 9 3876 28 3882
rect -1 3860 28 3876
rect 43 3866 73 3882
rect 101 3860 107 3908
rect 110 3902 129 3908
rect 144 3902 174 3910
rect 110 3894 174 3902
rect 110 3878 190 3894
rect 206 3887 268 3918
rect 284 3887 346 3918
rect 415 3916 464 3941
rect 479 3916 509 3932
rect 378 3902 408 3910
rect 415 3908 525 3916
rect 378 3894 423 3902
rect 110 3876 129 3878
rect 144 3876 190 3878
rect 110 3860 190 3876
rect 217 3874 252 3887
rect 293 3884 330 3887
rect 293 3882 335 3884
rect 222 3871 252 3874
rect 231 3867 238 3871
rect 238 3866 239 3867
rect 197 3860 207 3866
rect -7 3852 34 3860
rect -7 3826 8 3852
rect 15 3826 34 3852
rect 98 3848 129 3860
rect 144 3848 247 3860
rect 259 3850 285 3876
rect 300 3871 330 3882
rect 362 3878 424 3894
rect 362 3876 408 3878
rect 362 3860 424 3876
rect 436 3860 442 3908
rect 445 3900 525 3908
rect 445 3898 464 3900
rect 479 3898 513 3900
rect 445 3882 525 3898
rect 445 3860 464 3882
rect 479 3866 509 3882
rect 537 3876 543 3950
rect 546 3876 565 4020
rect 580 3876 586 4020
rect 595 3950 608 4020
rect 660 4016 682 4020
rect 653 3994 682 4008
rect 735 3994 751 4008
rect 789 4004 795 4006
rect 802 4004 910 4020
rect 917 4004 923 4006
rect 931 4004 946 4020
rect 1012 4014 1031 4017
rect 653 3992 751 3994
rect 778 3992 946 4004
rect 961 3994 977 4008
rect 1012 3995 1034 4014
rect 1044 4008 1060 4009
rect 1043 4006 1060 4008
rect 1044 4001 1060 4006
rect 1034 3994 1040 3995
rect 1043 3994 1072 4001
rect 961 3993 1072 3994
rect 961 3992 1078 3993
rect 637 3984 688 3992
rect 735 3984 769 3992
rect 637 3972 662 3984
rect 669 3972 688 3984
rect 742 3982 769 3984
rect 778 3982 999 3992
rect 1034 3989 1040 3992
rect 742 3978 999 3982
rect 637 3964 688 3972
rect 735 3964 999 3978
rect 1043 3984 1078 3992
rect 589 3916 608 3950
rect 653 3956 682 3964
rect 653 3950 670 3956
rect 653 3948 687 3950
rect 735 3948 751 3964
rect 752 3954 960 3964
rect 961 3954 977 3964
rect 1025 3960 1040 3975
rect 1043 3972 1044 3984
rect 1051 3972 1078 3984
rect 1043 3964 1078 3972
rect 1043 3963 1072 3964
rect 763 3950 977 3954
rect 778 3948 977 3950
rect 1012 3950 1025 3960
rect 1043 3950 1060 3963
rect 1012 3948 1060 3950
rect 654 3944 687 3948
rect 650 3942 687 3944
rect 650 3941 717 3942
rect 650 3936 681 3941
rect 687 3936 717 3941
rect 650 3932 717 3936
rect 623 3929 717 3932
rect 623 3922 672 3929
rect 623 3916 653 3922
rect 672 3917 677 3922
rect 589 3900 669 3916
rect 681 3908 717 3929
rect 778 3924 967 3948
rect 1012 3947 1059 3948
rect 1025 3942 1059 3947
rect 793 3921 967 3924
rect 786 3918 967 3921
rect 995 3941 1059 3942
rect 589 3898 608 3900
rect 623 3898 657 3900
rect 589 3882 669 3898
rect 589 3876 608 3882
rect 305 3850 408 3860
rect 259 3848 408 3850
rect 429 3848 464 3860
rect 98 3846 260 3848
rect 110 3826 129 3846
rect 144 3844 174 3846
rect -7 3818 34 3826
rect 116 3822 129 3826
rect 181 3830 260 3846
rect 292 3846 464 3848
rect 292 3830 371 3846
rect 378 3844 408 3846
rect -1 3808 28 3818
rect 43 3808 73 3822
rect 116 3808 159 3822
rect 181 3818 371 3830
rect 436 3826 442 3846
rect 166 3808 196 3818
rect 197 3808 355 3818
rect 359 3808 389 3818
rect 393 3808 423 3822
rect 451 3808 464 3846
rect 536 3860 565 3876
rect 579 3860 608 3876
rect 623 3866 653 3882
rect 681 3860 687 3908
rect 690 3902 709 3908
rect 724 3902 754 3910
rect 690 3894 754 3902
rect 690 3878 770 3894
rect 786 3887 848 3918
rect 864 3887 926 3918
rect 995 3916 1044 3941
rect 1059 3916 1089 3932
rect 958 3902 988 3910
rect 995 3908 1105 3916
rect 958 3894 1003 3902
rect 690 3876 709 3878
rect 724 3876 770 3878
rect 690 3860 770 3876
rect 797 3874 832 3887
rect 873 3884 910 3887
rect 873 3882 915 3884
rect 802 3871 832 3874
rect 811 3867 818 3871
rect 818 3866 819 3867
rect 777 3860 787 3866
rect 536 3852 571 3860
rect 536 3826 537 3852
rect 544 3826 571 3852
rect 479 3808 509 3822
rect 536 3818 571 3826
rect 573 3852 614 3860
rect 573 3826 588 3852
rect 595 3826 614 3852
rect 678 3848 709 3860
rect 724 3848 827 3860
rect 839 3850 865 3876
rect 880 3871 910 3882
rect 942 3878 1004 3894
rect 942 3876 988 3878
rect 942 3860 1004 3876
rect 1016 3860 1022 3908
rect 1025 3900 1105 3908
rect 1025 3898 1044 3900
rect 1059 3898 1093 3900
rect 1025 3882 1105 3898
rect 1025 3860 1044 3882
rect 1059 3866 1089 3882
rect 1117 3876 1123 3950
rect 1126 3876 1145 4020
rect 1160 3876 1166 4020
rect 1175 3950 1188 4020
rect 1240 4016 1262 4020
rect 1233 3994 1262 4008
rect 1315 3994 1331 4008
rect 1369 4004 1375 4006
rect 1382 4004 1490 4020
rect 1497 4004 1503 4006
rect 1511 4004 1526 4020
rect 1592 4014 1611 4017
rect 1233 3992 1331 3994
rect 1358 3992 1526 4004
rect 1541 3994 1557 4008
rect 1592 3995 1614 4014
rect 1624 4008 1640 4009
rect 1623 4006 1640 4008
rect 1624 4001 1640 4006
rect 1614 3994 1620 3995
rect 1623 3994 1652 4001
rect 1541 3993 1652 3994
rect 1541 3992 1658 3993
rect 1217 3984 1268 3992
rect 1315 3984 1349 3992
rect 1217 3972 1242 3984
rect 1249 3972 1268 3984
rect 1322 3982 1349 3984
rect 1358 3982 1579 3992
rect 1614 3989 1620 3992
rect 1322 3978 1579 3982
rect 1217 3964 1268 3972
rect 1315 3964 1579 3978
rect 1623 3984 1658 3992
rect 1169 3916 1188 3950
rect 1233 3956 1262 3964
rect 1233 3950 1250 3956
rect 1233 3948 1267 3950
rect 1315 3948 1331 3964
rect 1332 3954 1540 3964
rect 1541 3954 1557 3964
rect 1605 3960 1620 3975
rect 1623 3972 1624 3984
rect 1631 3972 1658 3984
rect 1623 3964 1658 3972
rect 1623 3963 1652 3964
rect 1343 3950 1557 3954
rect 1358 3948 1557 3950
rect 1592 3950 1605 3960
rect 1623 3950 1640 3963
rect 1592 3948 1640 3950
rect 1234 3944 1267 3948
rect 1230 3942 1267 3944
rect 1230 3941 1297 3942
rect 1230 3936 1261 3941
rect 1267 3936 1297 3941
rect 1230 3932 1297 3936
rect 1203 3929 1297 3932
rect 1203 3922 1252 3929
rect 1203 3916 1233 3922
rect 1252 3917 1257 3922
rect 1169 3900 1249 3916
rect 1261 3908 1297 3929
rect 1358 3924 1547 3948
rect 1592 3947 1639 3948
rect 1605 3942 1639 3947
rect 1373 3921 1547 3924
rect 1366 3918 1547 3921
rect 1575 3941 1639 3942
rect 1169 3898 1188 3900
rect 1203 3898 1237 3900
rect 1169 3882 1249 3898
rect 1169 3876 1188 3882
rect 885 3850 988 3860
rect 839 3848 988 3850
rect 1009 3848 1044 3860
rect 678 3846 840 3848
rect 690 3826 709 3846
rect 724 3844 754 3846
rect 573 3818 614 3826
rect 696 3822 709 3826
rect 761 3830 840 3846
rect 872 3846 1044 3848
rect 872 3830 951 3846
rect 958 3844 988 3846
rect 536 3808 565 3818
rect 579 3808 608 3818
rect 623 3808 653 3822
rect 696 3808 739 3822
rect 761 3818 951 3830
rect 1016 3826 1022 3846
rect 746 3808 776 3818
rect 777 3808 935 3818
rect 939 3808 969 3818
rect 973 3808 1003 3822
rect 1031 3808 1044 3846
rect 1116 3860 1145 3876
rect 1159 3860 1188 3876
rect 1203 3866 1233 3882
rect 1261 3860 1267 3908
rect 1270 3902 1289 3908
rect 1304 3902 1334 3910
rect 1270 3894 1334 3902
rect 1270 3878 1350 3894
rect 1366 3887 1428 3918
rect 1444 3887 1506 3918
rect 1575 3916 1624 3941
rect 1639 3916 1669 3932
rect 1538 3902 1568 3910
rect 1575 3908 1685 3916
rect 1538 3894 1583 3902
rect 1270 3876 1289 3878
rect 1304 3876 1350 3878
rect 1270 3860 1350 3876
rect 1377 3874 1412 3887
rect 1453 3884 1490 3887
rect 1453 3882 1495 3884
rect 1382 3871 1412 3874
rect 1391 3867 1398 3871
rect 1398 3866 1399 3867
rect 1357 3860 1367 3866
rect 1116 3852 1151 3860
rect 1116 3826 1117 3852
rect 1124 3826 1151 3852
rect 1059 3808 1089 3822
rect 1116 3818 1151 3826
rect 1153 3852 1194 3860
rect 1153 3826 1168 3852
rect 1175 3826 1194 3852
rect 1258 3848 1289 3860
rect 1304 3848 1407 3860
rect 1419 3850 1445 3876
rect 1460 3871 1490 3882
rect 1522 3878 1584 3894
rect 1522 3876 1568 3878
rect 1522 3860 1584 3876
rect 1596 3860 1602 3908
rect 1605 3900 1685 3908
rect 1605 3898 1624 3900
rect 1639 3898 1673 3900
rect 1605 3882 1685 3898
rect 1605 3860 1624 3882
rect 1639 3866 1669 3882
rect 1697 3876 1703 3950
rect 1706 3876 1725 4020
rect 1740 3876 1746 4020
rect 1755 3950 1768 4020
rect 1820 4016 1842 4020
rect 1813 3994 1842 4008
rect 1895 3994 1911 4008
rect 1949 4004 1955 4006
rect 1962 4004 2070 4020
rect 2077 4004 2083 4006
rect 2091 4004 2106 4020
rect 2172 4014 2191 4017
rect 1813 3992 1911 3994
rect 1938 3992 2106 4004
rect 2121 3994 2137 4008
rect 2172 3995 2194 4014
rect 2204 4008 2220 4009
rect 2203 4006 2220 4008
rect 2204 4001 2220 4006
rect 2194 3994 2200 3995
rect 2203 3994 2232 4001
rect 2121 3993 2232 3994
rect 2121 3992 2238 3993
rect 1797 3984 1848 3992
rect 1895 3984 1929 3992
rect 1797 3972 1822 3984
rect 1829 3972 1848 3984
rect 1902 3982 1929 3984
rect 1938 3982 2159 3992
rect 2194 3989 2200 3992
rect 1902 3978 2159 3982
rect 1797 3964 1848 3972
rect 1895 3964 2159 3978
rect 2203 3984 2238 3992
rect 1749 3916 1768 3950
rect 1813 3956 1842 3964
rect 1813 3950 1830 3956
rect 1813 3948 1847 3950
rect 1895 3948 1911 3964
rect 1912 3954 2120 3964
rect 2121 3954 2137 3964
rect 2185 3960 2200 3975
rect 2203 3972 2204 3984
rect 2211 3972 2238 3984
rect 2203 3964 2238 3972
rect 2203 3963 2232 3964
rect 1923 3950 2137 3954
rect 1938 3948 2137 3950
rect 2172 3950 2185 3960
rect 2203 3950 2220 3963
rect 2172 3948 2220 3950
rect 1814 3944 1847 3948
rect 1810 3942 1847 3944
rect 1810 3941 1877 3942
rect 1810 3936 1841 3941
rect 1847 3936 1877 3941
rect 1810 3932 1877 3936
rect 1783 3929 1877 3932
rect 1783 3922 1832 3929
rect 1783 3916 1813 3922
rect 1832 3917 1837 3922
rect 1749 3900 1829 3916
rect 1841 3908 1877 3929
rect 1938 3924 2127 3948
rect 2172 3947 2219 3948
rect 2185 3942 2219 3947
rect 1953 3921 2127 3924
rect 1946 3918 2127 3921
rect 2155 3941 2219 3942
rect 1749 3898 1768 3900
rect 1783 3898 1817 3900
rect 1749 3882 1829 3898
rect 1749 3876 1768 3882
rect 1465 3850 1568 3860
rect 1419 3848 1568 3850
rect 1589 3848 1624 3860
rect 1258 3846 1420 3848
rect 1270 3826 1289 3846
rect 1304 3844 1334 3846
rect 1153 3818 1194 3826
rect 1276 3822 1289 3826
rect 1341 3830 1420 3846
rect 1452 3846 1624 3848
rect 1452 3830 1531 3846
rect 1538 3844 1568 3846
rect 1116 3808 1145 3818
rect 1159 3808 1188 3818
rect 1203 3808 1233 3822
rect 1276 3808 1319 3822
rect 1341 3818 1531 3830
rect 1596 3826 1602 3846
rect 1326 3808 1356 3818
rect 1357 3808 1515 3818
rect 1519 3808 1549 3818
rect 1553 3808 1583 3822
rect 1611 3808 1624 3846
rect 1696 3860 1725 3876
rect 1739 3860 1768 3876
rect 1783 3866 1813 3882
rect 1841 3860 1847 3908
rect 1850 3902 1869 3908
rect 1884 3902 1914 3910
rect 1850 3894 1914 3902
rect 1850 3878 1930 3894
rect 1946 3887 2008 3918
rect 2024 3887 2086 3918
rect 2155 3916 2204 3941
rect 2219 3916 2249 3932
rect 2118 3902 2148 3910
rect 2155 3908 2265 3916
rect 2118 3894 2163 3902
rect 1850 3876 1869 3878
rect 1884 3876 1930 3878
rect 1850 3860 1930 3876
rect 1957 3874 1992 3887
rect 2033 3884 2070 3887
rect 2033 3882 2075 3884
rect 1962 3871 1992 3874
rect 1971 3867 1978 3871
rect 1978 3866 1979 3867
rect 1937 3860 1947 3866
rect 1696 3852 1731 3860
rect 1696 3826 1697 3852
rect 1704 3826 1731 3852
rect 1639 3808 1669 3822
rect 1696 3818 1731 3826
rect 1733 3852 1774 3860
rect 1733 3826 1748 3852
rect 1755 3826 1774 3852
rect 1838 3848 1869 3860
rect 1884 3848 1987 3860
rect 1999 3850 2025 3876
rect 2040 3871 2070 3882
rect 2102 3878 2164 3894
rect 2102 3876 2148 3878
rect 2102 3860 2164 3876
rect 2176 3860 2182 3908
rect 2185 3900 2265 3908
rect 2185 3898 2204 3900
rect 2219 3898 2253 3900
rect 2185 3882 2265 3898
rect 2185 3860 2204 3882
rect 2219 3866 2249 3882
rect 2277 3876 2283 3950
rect 2286 3876 2305 4020
rect 2320 3876 2326 4020
rect 2335 3950 2348 4020
rect 2400 4016 2422 4020
rect 2393 3994 2422 4008
rect 2475 3994 2491 4008
rect 2529 4004 2535 4006
rect 2542 4004 2650 4020
rect 2657 4004 2663 4006
rect 2671 4004 2686 4020
rect 2752 4014 2771 4017
rect 2393 3992 2491 3994
rect 2518 3992 2686 4004
rect 2701 3994 2717 4008
rect 2752 3995 2774 4014
rect 2784 4008 2800 4009
rect 2783 4006 2800 4008
rect 2784 4001 2800 4006
rect 2774 3994 2780 3995
rect 2783 3994 2812 4001
rect 2701 3993 2812 3994
rect 2701 3992 2818 3993
rect 2377 3984 2428 3992
rect 2475 3984 2509 3992
rect 2377 3972 2402 3984
rect 2409 3972 2428 3984
rect 2482 3982 2509 3984
rect 2518 3982 2739 3992
rect 2774 3989 2780 3992
rect 2482 3978 2739 3982
rect 2377 3964 2428 3972
rect 2475 3964 2739 3978
rect 2783 3984 2818 3992
rect 2329 3916 2348 3950
rect 2393 3956 2422 3964
rect 2393 3950 2410 3956
rect 2393 3948 2427 3950
rect 2475 3948 2491 3964
rect 2492 3954 2700 3964
rect 2701 3954 2717 3964
rect 2765 3960 2780 3975
rect 2783 3972 2784 3984
rect 2791 3972 2818 3984
rect 2783 3964 2818 3972
rect 2783 3963 2812 3964
rect 2503 3950 2717 3954
rect 2518 3948 2717 3950
rect 2752 3950 2765 3960
rect 2783 3950 2800 3963
rect 2752 3948 2800 3950
rect 2394 3944 2427 3948
rect 2390 3942 2427 3944
rect 2390 3941 2457 3942
rect 2390 3936 2421 3941
rect 2427 3936 2457 3941
rect 2390 3932 2457 3936
rect 2363 3929 2457 3932
rect 2363 3922 2412 3929
rect 2363 3916 2393 3922
rect 2412 3917 2417 3922
rect 2329 3900 2409 3916
rect 2421 3908 2457 3929
rect 2518 3924 2707 3948
rect 2752 3947 2799 3948
rect 2765 3942 2799 3947
rect 2533 3921 2707 3924
rect 2526 3918 2707 3921
rect 2735 3941 2799 3942
rect 2329 3898 2348 3900
rect 2363 3898 2397 3900
rect 2329 3882 2409 3898
rect 2329 3876 2348 3882
rect 2045 3850 2148 3860
rect 1999 3848 2148 3850
rect 2169 3848 2204 3860
rect 1838 3846 2000 3848
rect 1850 3826 1869 3846
rect 1884 3844 1914 3846
rect 1733 3818 1774 3826
rect 1856 3822 1869 3826
rect 1921 3830 2000 3846
rect 2032 3846 2204 3848
rect 2032 3830 2111 3846
rect 2118 3844 2148 3846
rect 1696 3808 1725 3818
rect 1739 3808 1768 3818
rect 1783 3808 1813 3822
rect 1856 3808 1899 3822
rect 1921 3818 2111 3830
rect 2176 3826 2182 3846
rect 1906 3808 1936 3818
rect 1937 3808 2095 3818
rect 2099 3808 2129 3818
rect 2133 3808 2163 3822
rect 2191 3808 2204 3846
rect 2276 3860 2305 3876
rect 2319 3860 2348 3876
rect 2363 3866 2393 3882
rect 2421 3860 2427 3908
rect 2430 3902 2449 3908
rect 2464 3902 2494 3910
rect 2430 3894 2494 3902
rect 2430 3878 2510 3894
rect 2526 3887 2588 3918
rect 2604 3887 2666 3918
rect 2735 3916 2784 3941
rect 2799 3916 2829 3932
rect 2698 3902 2728 3910
rect 2735 3908 2845 3916
rect 2698 3894 2743 3902
rect 2430 3876 2449 3878
rect 2464 3876 2510 3878
rect 2430 3860 2510 3876
rect 2537 3874 2572 3887
rect 2613 3884 2650 3887
rect 2613 3882 2655 3884
rect 2542 3871 2572 3874
rect 2551 3867 2558 3871
rect 2558 3866 2559 3867
rect 2517 3860 2527 3866
rect 2276 3852 2311 3860
rect 2276 3826 2277 3852
rect 2284 3826 2311 3852
rect 2219 3808 2249 3822
rect 2276 3818 2311 3826
rect 2313 3852 2354 3860
rect 2313 3826 2328 3852
rect 2335 3826 2354 3852
rect 2418 3848 2449 3860
rect 2464 3848 2567 3860
rect 2579 3850 2605 3876
rect 2620 3871 2650 3882
rect 2682 3878 2744 3894
rect 2682 3876 2728 3878
rect 2682 3860 2744 3876
rect 2756 3860 2762 3908
rect 2765 3900 2845 3908
rect 2765 3898 2784 3900
rect 2799 3898 2833 3900
rect 2765 3882 2845 3898
rect 2765 3860 2784 3882
rect 2799 3866 2829 3882
rect 2857 3876 2863 3950
rect 2866 3876 2885 4020
rect 2900 3876 2906 4020
rect 2915 3950 2928 4020
rect 2980 4016 3002 4020
rect 2973 3994 3002 4008
rect 3055 3994 3071 4008
rect 3109 4004 3115 4006
rect 3122 4004 3230 4020
rect 3237 4004 3243 4006
rect 3251 4004 3266 4020
rect 3332 4014 3351 4017
rect 2973 3992 3071 3994
rect 3098 3992 3266 4004
rect 3281 3994 3297 4008
rect 3332 3995 3354 4014
rect 3364 4008 3380 4009
rect 3363 4006 3380 4008
rect 3364 4001 3380 4006
rect 3354 3994 3360 3995
rect 3363 3994 3392 4001
rect 3281 3993 3392 3994
rect 3281 3992 3398 3993
rect 2957 3984 3008 3992
rect 3055 3984 3089 3992
rect 2957 3972 2982 3984
rect 2989 3972 3008 3984
rect 3062 3982 3089 3984
rect 3098 3982 3319 3992
rect 3354 3989 3360 3992
rect 3062 3978 3319 3982
rect 2957 3964 3008 3972
rect 3055 3964 3319 3978
rect 3363 3984 3398 3992
rect 2909 3916 2928 3950
rect 2973 3956 3002 3964
rect 2973 3950 2990 3956
rect 2973 3948 3007 3950
rect 3055 3948 3071 3964
rect 3072 3954 3280 3964
rect 3281 3954 3297 3964
rect 3345 3960 3360 3975
rect 3363 3972 3364 3984
rect 3371 3972 3398 3984
rect 3363 3964 3398 3972
rect 3363 3963 3392 3964
rect 3083 3950 3297 3954
rect 3098 3948 3297 3950
rect 3332 3950 3345 3960
rect 3363 3950 3380 3963
rect 3332 3948 3380 3950
rect 2974 3944 3007 3948
rect 2970 3942 3007 3944
rect 2970 3941 3037 3942
rect 2970 3936 3001 3941
rect 3007 3936 3037 3941
rect 2970 3932 3037 3936
rect 2943 3929 3037 3932
rect 2943 3922 2992 3929
rect 2943 3916 2973 3922
rect 2992 3917 2997 3922
rect 2909 3900 2989 3916
rect 3001 3908 3037 3929
rect 3098 3924 3287 3948
rect 3332 3947 3379 3948
rect 3345 3942 3379 3947
rect 3113 3921 3287 3924
rect 3106 3918 3287 3921
rect 3315 3941 3379 3942
rect 2909 3898 2928 3900
rect 2943 3898 2977 3900
rect 2909 3882 2989 3898
rect 2909 3876 2928 3882
rect 2625 3850 2728 3860
rect 2579 3848 2728 3850
rect 2749 3848 2784 3860
rect 2418 3846 2580 3848
rect 2430 3826 2449 3846
rect 2464 3844 2494 3846
rect 2313 3818 2354 3826
rect 2436 3822 2449 3826
rect 2501 3830 2580 3846
rect 2612 3846 2784 3848
rect 2612 3830 2691 3846
rect 2698 3844 2728 3846
rect 2276 3808 2305 3818
rect 2319 3808 2348 3818
rect 2363 3808 2393 3822
rect 2436 3808 2479 3822
rect 2501 3818 2691 3830
rect 2756 3826 2762 3846
rect 2486 3808 2516 3818
rect 2517 3808 2675 3818
rect 2679 3808 2709 3818
rect 2713 3808 2743 3822
rect 2771 3808 2784 3846
rect 2856 3860 2885 3876
rect 2899 3860 2928 3876
rect 2943 3866 2973 3882
rect 3001 3860 3007 3908
rect 3010 3902 3029 3908
rect 3044 3902 3074 3910
rect 3010 3894 3074 3902
rect 3010 3878 3090 3894
rect 3106 3887 3168 3918
rect 3184 3887 3246 3918
rect 3315 3916 3364 3941
rect 3379 3916 3409 3932
rect 3278 3902 3308 3910
rect 3315 3908 3425 3916
rect 3278 3894 3323 3902
rect 3010 3876 3029 3878
rect 3044 3876 3090 3878
rect 3010 3860 3090 3876
rect 3117 3874 3152 3887
rect 3193 3884 3230 3887
rect 3193 3882 3235 3884
rect 3122 3871 3152 3874
rect 3131 3867 3138 3871
rect 3138 3866 3139 3867
rect 3097 3860 3107 3866
rect 2856 3852 2891 3860
rect 2856 3826 2857 3852
rect 2864 3826 2891 3852
rect 2799 3808 2829 3822
rect 2856 3818 2891 3826
rect 2893 3852 2934 3860
rect 2893 3826 2908 3852
rect 2915 3826 2934 3852
rect 2998 3848 3029 3860
rect 3044 3848 3147 3860
rect 3159 3850 3185 3876
rect 3200 3871 3230 3882
rect 3262 3878 3324 3894
rect 3262 3876 3308 3878
rect 3262 3860 3324 3876
rect 3336 3860 3342 3908
rect 3345 3900 3425 3908
rect 3345 3898 3364 3900
rect 3379 3898 3413 3900
rect 3345 3882 3425 3898
rect 3345 3860 3364 3882
rect 3379 3866 3409 3882
rect 3437 3876 3443 3950
rect 3446 3876 3465 4020
rect 3480 3876 3486 4020
rect 3495 3950 3508 4020
rect 3560 4016 3582 4020
rect 3553 3994 3582 4008
rect 3635 3994 3651 4008
rect 3689 4004 3695 4006
rect 3702 4004 3810 4020
rect 3817 4004 3823 4006
rect 3831 4004 3846 4020
rect 3912 4014 3931 4017
rect 3553 3992 3651 3994
rect 3678 3992 3846 4004
rect 3861 3994 3877 4008
rect 3912 3995 3934 4014
rect 3944 4008 3960 4009
rect 3943 4006 3960 4008
rect 3944 4001 3960 4006
rect 3934 3994 3940 3995
rect 3943 3994 3972 4001
rect 3861 3993 3972 3994
rect 3861 3992 3978 3993
rect 3537 3984 3588 3992
rect 3635 3984 3669 3992
rect 3537 3972 3562 3984
rect 3569 3972 3588 3984
rect 3642 3982 3669 3984
rect 3678 3982 3899 3992
rect 3934 3989 3940 3992
rect 3642 3978 3899 3982
rect 3537 3964 3588 3972
rect 3635 3964 3899 3978
rect 3943 3984 3978 3992
rect 3489 3916 3508 3950
rect 3553 3956 3582 3964
rect 3553 3950 3570 3956
rect 3553 3948 3587 3950
rect 3635 3948 3651 3964
rect 3652 3954 3860 3964
rect 3861 3954 3877 3964
rect 3925 3960 3940 3975
rect 3943 3972 3944 3984
rect 3951 3972 3978 3984
rect 3943 3964 3978 3972
rect 3943 3963 3972 3964
rect 3663 3950 3877 3954
rect 3678 3948 3877 3950
rect 3912 3950 3925 3960
rect 3943 3950 3960 3963
rect 3912 3948 3960 3950
rect 3554 3944 3587 3948
rect 3550 3942 3587 3944
rect 3550 3941 3617 3942
rect 3550 3936 3581 3941
rect 3587 3936 3617 3941
rect 3550 3932 3617 3936
rect 3523 3929 3617 3932
rect 3523 3922 3572 3929
rect 3523 3916 3553 3922
rect 3572 3917 3577 3922
rect 3489 3900 3569 3916
rect 3581 3908 3617 3929
rect 3678 3924 3867 3948
rect 3912 3947 3959 3948
rect 3925 3942 3959 3947
rect 3693 3921 3867 3924
rect 3686 3918 3867 3921
rect 3895 3941 3959 3942
rect 3489 3898 3508 3900
rect 3523 3898 3557 3900
rect 3489 3882 3569 3898
rect 3489 3876 3508 3882
rect 3205 3850 3308 3860
rect 3159 3848 3308 3850
rect 3329 3848 3364 3860
rect 2998 3846 3160 3848
rect 3010 3826 3029 3846
rect 3044 3844 3074 3846
rect 2893 3818 2934 3826
rect 3016 3822 3029 3826
rect 3081 3830 3160 3846
rect 3192 3846 3364 3848
rect 3192 3830 3271 3846
rect 3278 3844 3308 3846
rect 2856 3808 2885 3818
rect 2899 3808 2928 3818
rect 2943 3808 2973 3822
rect 3016 3808 3059 3822
rect 3081 3818 3271 3830
rect 3336 3826 3342 3846
rect 3066 3808 3096 3818
rect 3097 3808 3255 3818
rect 3259 3808 3289 3818
rect 3293 3808 3323 3822
rect 3351 3808 3364 3846
rect 3436 3860 3465 3876
rect 3479 3860 3508 3876
rect 3523 3866 3553 3882
rect 3581 3860 3587 3908
rect 3590 3902 3609 3908
rect 3624 3902 3654 3910
rect 3590 3894 3654 3902
rect 3590 3878 3670 3894
rect 3686 3887 3748 3918
rect 3764 3887 3826 3918
rect 3895 3916 3944 3941
rect 3959 3916 3989 3932
rect 3858 3902 3888 3910
rect 3895 3908 4005 3916
rect 3858 3894 3903 3902
rect 3590 3876 3609 3878
rect 3624 3876 3670 3878
rect 3590 3860 3670 3876
rect 3697 3874 3732 3887
rect 3773 3884 3810 3887
rect 3773 3882 3815 3884
rect 3702 3871 3732 3874
rect 3711 3867 3718 3871
rect 3718 3866 3719 3867
rect 3677 3860 3687 3866
rect 3436 3852 3471 3860
rect 3436 3826 3437 3852
rect 3444 3826 3471 3852
rect 3379 3808 3409 3822
rect 3436 3818 3471 3826
rect 3473 3852 3514 3860
rect 3473 3826 3488 3852
rect 3495 3826 3514 3852
rect 3578 3848 3609 3860
rect 3624 3848 3727 3860
rect 3739 3850 3765 3876
rect 3780 3871 3810 3882
rect 3842 3878 3904 3894
rect 3842 3876 3888 3878
rect 3842 3860 3904 3876
rect 3916 3860 3922 3908
rect 3925 3900 4005 3908
rect 3925 3898 3944 3900
rect 3959 3898 3993 3900
rect 3925 3882 4005 3898
rect 3925 3860 3944 3882
rect 3959 3866 3989 3882
rect 4017 3876 4023 3950
rect 4026 3876 4045 4020
rect 4060 3876 4066 4020
rect 4075 3950 4088 4020
rect 4140 4016 4162 4020
rect 4133 3994 4162 4008
rect 4215 3994 4231 4008
rect 4269 4004 4275 4006
rect 4282 4004 4390 4020
rect 4397 4004 4403 4006
rect 4411 4004 4426 4020
rect 4492 4014 4511 4017
rect 4133 3992 4231 3994
rect 4258 3992 4426 4004
rect 4441 3994 4457 4008
rect 4492 3995 4514 4014
rect 4524 4008 4540 4009
rect 4523 4006 4540 4008
rect 4524 4001 4540 4006
rect 4514 3994 4520 3995
rect 4523 3994 4552 4001
rect 4441 3993 4552 3994
rect 4441 3992 4558 3993
rect 4117 3984 4168 3992
rect 4215 3984 4249 3992
rect 4117 3972 4142 3984
rect 4149 3972 4168 3984
rect 4222 3982 4249 3984
rect 4258 3982 4479 3992
rect 4514 3989 4520 3992
rect 4222 3978 4479 3982
rect 4117 3964 4168 3972
rect 4215 3964 4479 3978
rect 4523 3984 4558 3992
rect 4069 3916 4088 3950
rect 4133 3956 4162 3964
rect 4133 3950 4150 3956
rect 4133 3948 4167 3950
rect 4215 3948 4231 3964
rect 4232 3954 4440 3964
rect 4441 3954 4457 3964
rect 4505 3960 4520 3975
rect 4523 3972 4524 3984
rect 4531 3972 4558 3984
rect 4523 3964 4558 3972
rect 4523 3963 4552 3964
rect 4243 3950 4457 3954
rect 4258 3948 4457 3950
rect 4492 3950 4505 3960
rect 4523 3950 4540 3963
rect 4492 3948 4540 3950
rect 4134 3944 4167 3948
rect 4130 3942 4167 3944
rect 4130 3941 4197 3942
rect 4130 3936 4161 3941
rect 4167 3936 4197 3941
rect 4130 3932 4197 3936
rect 4103 3929 4197 3932
rect 4103 3922 4152 3929
rect 4103 3916 4133 3922
rect 4152 3917 4157 3922
rect 4069 3900 4149 3916
rect 4161 3908 4197 3929
rect 4258 3924 4447 3948
rect 4492 3947 4539 3948
rect 4505 3942 4539 3947
rect 4273 3921 4447 3924
rect 4266 3918 4447 3921
rect 4475 3941 4539 3942
rect 4069 3898 4088 3900
rect 4103 3898 4137 3900
rect 4069 3882 4149 3898
rect 4069 3876 4088 3882
rect 3785 3850 3888 3860
rect 3739 3848 3888 3850
rect 3909 3848 3944 3860
rect 3578 3846 3740 3848
rect 3590 3826 3609 3846
rect 3624 3844 3654 3846
rect 3473 3818 3514 3826
rect 3596 3822 3609 3826
rect 3661 3830 3740 3846
rect 3772 3846 3944 3848
rect 3772 3830 3851 3846
rect 3858 3844 3888 3846
rect 3436 3808 3465 3818
rect 3479 3808 3508 3818
rect 3523 3808 3553 3822
rect 3596 3808 3639 3822
rect 3661 3818 3851 3830
rect 3916 3826 3922 3846
rect 3646 3808 3676 3818
rect 3677 3808 3835 3818
rect 3839 3808 3869 3818
rect 3873 3808 3903 3822
rect 3931 3808 3944 3846
rect 4016 3860 4045 3876
rect 4059 3860 4088 3876
rect 4103 3866 4133 3882
rect 4161 3860 4167 3908
rect 4170 3902 4189 3908
rect 4204 3902 4234 3910
rect 4170 3894 4234 3902
rect 4170 3878 4250 3894
rect 4266 3887 4328 3918
rect 4344 3887 4406 3918
rect 4475 3916 4524 3941
rect 4539 3916 4569 3932
rect 4438 3902 4468 3910
rect 4475 3908 4585 3916
rect 4438 3894 4483 3902
rect 4170 3876 4189 3878
rect 4204 3876 4250 3878
rect 4170 3860 4250 3876
rect 4277 3874 4312 3887
rect 4353 3884 4390 3887
rect 4353 3882 4395 3884
rect 4282 3871 4312 3874
rect 4291 3867 4298 3871
rect 4298 3866 4299 3867
rect 4257 3860 4267 3866
rect 4016 3852 4051 3860
rect 4016 3826 4017 3852
rect 4024 3826 4051 3852
rect 3959 3808 3989 3822
rect 4016 3818 4051 3826
rect 4053 3852 4094 3860
rect 4053 3826 4068 3852
rect 4075 3826 4094 3852
rect 4158 3848 4189 3860
rect 4204 3848 4307 3860
rect 4319 3850 4345 3876
rect 4360 3871 4390 3882
rect 4422 3878 4484 3894
rect 4422 3876 4468 3878
rect 4422 3860 4484 3876
rect 4496 3860 4502 3908
rect 4505 3900 4585 3908
rect 4505 3898 4524 3900
rect 4539 3898 4573 3900
rect 4505 3882 4585 3898
rect 4505 3860 4524 3882
rect 4539 3866 4569 3882
rect 4597 3876 4603 3950
rect 4606 3876 4625 4020
rect 4640 3876 4646 4020
rect 4655 3950 4668 4020
rect 4720 4016 4742 4020
rect 4713 3994 4742 4008
rect 4795 3994 4811 4008
rect 4849 4004 4855 4006
rect 4862 4004 4970 4020
rect 4977 4004 4983 4006
rect 4991 4004 5006 4020
rect 5072 4014 5091 4017
rect 4713 3992 4811 3994
rect 4838 3992 5006 4004
rect 5021 3994 5037 4008
rect 5072 3995 5094 4014
rect 5104 4008 5120 4009
rect 5103 4006 5120 4008
rect 5104 4001 5120 4006
rect 5094 3994 5100 3995
rect 5103 3994 5132 4001
rect 5021 3993 5132 3994
rect 5021 3992 5138 3993
rect 4697 3984 4748 3992
rect 4795 3984 4829 3992
rect 4697 3972 4722 3984
rect 4729 3972 4748 3984
rect 4802 3982 4829 3984
rect 4838 3982 5059 3992
rect 5094 3989 5100 3992
rect 4802 3978 5059 3982
rect 4697 3964 4748 3972
rect 4795 3964 5059 3978
rect 5103 3984 5138 3992
rect 4649 3916 4668 3950
rect 4713 3956 4742 3964
rect 4713 3950 4730 3956
rect 4713 3948 4747 3950
rect 4795 3948 4811 3964
rect 4812 3954 5020 3964
rect 5021 3954 5037 3964
rect 5085 3960 5100 3975
rect 5103 3972 5104 3984
rect 5111 3972 5138 3984
rect 5103 3964 5138 3972
rect 5103 3963 5132 3964
rect 4823 3950 5037 3954
rect 4838 3948 5037 3950
rect 5072 3950 5085 3960
rect 5103 3950 5120 3963
rect 5072 3948 5120 3950
rect 4714 3944 4747 3948
rect 4710 3942 4747 3944
rect 4710 3941 4777 3942
rect 4710 3936 4741 3941
rect 4747 3936 4777 3941
rect 4710 3932 4777 3936
rect 4683 3929 4777 3932
rect 4683 3922 4732 3929
rect 4683 3916 4713 3922
rect 4732 3917 4737 3922
rect 4649 3900 4729 3916
rect 4741 3908 4777 3929
rect 4838 3924 5027 3948
rect 5072 3947 5119 3948
rect 5085 3942 5119 3947
rect 4853 3921 5027 3924
rect 4846 3918 5027 3921
rect 5055 3941 5119 3942
rect 4649 3898 4668 3900
rect 4683 3898 4717 3900
rect 4649 3882 4729 3898
rect 4649 3876 4668 3882
rect 4365 3850 4468 3860
rect 4319 3848 4468 3850
rect 4489 3848 4524 3860
rect 4158 3846 4320 3848
rect 4170 3826 4189 3846
rect 4204 3844 4234 3846
rect 4053 3818 4094 3826
rect 4176 3822 4189 3826
rect 4241 3830 4320 3846
rect 4352 3846 4524 3848
rect 4352 3830 4431 3846
rect 4438 3844 4468 3846
rect 4016 3808 4045 3818
rect 4059 3808 4088 3818
rect 4103 3808 4133 3822
rect 4176 3808 4219 3822
rect 4241 3818 4431 3830
rect 4496 3826 4502 3846
rect 4226 3808 4256 3818
rect 4257 3808 4415 3818
rect 4419 3808 4449 3818
rect 4453 3808 4483 3822
rect 4511 3808 4524 3846
rect 4596 3860 4625 3876
rect 4639 3860 4668 3876
rect 4683 3866 4713 3882
rect 4741 3860 4747 3908
rect 4750 3902 4769 3908
rect 4784 3902 4814 3910
rect 4750 3894 4814 3902
rect 4750 3878 4830 3894
rect 4846 3887 4908 3918
rect 4924 3887 4986 3918
rect 5055 3916 5104 3941
rect 5119 3916 5149 3932
rect 5018 3902 5048 3910
rect 5055 3908 5165 3916
rect 5018 3894 5063 3902
rect 4750 3876 4769 3878
rect 4784 3876 4830 3878
rect 4750 3860 4830 3876
rect 4857 3874 4892 3887
rect 4933 3884 4970 3887
rect 4933 3882 4975 3884
rect 4862 3871 4892 3874
rect 4871 3867 4878 3871
rect 4878 3866 4879 3867
rect 4837 3860 4847 3866
rect 4596 3852 4631 3860
rect 4596 3826 4597 3852
rect 4604 3826 4631 3852
rect 4539 3808 4569 3822
rect 4596 3818 4631 3826
rect 4633 3852 4674 3860
rect 4633 3826 4648 3852
rect 4655 3826 4674 3852
rect 4738 3848 4769 3860
rect 4784 3848 4887 3860
rect 4899 3850 4925 3876
rect 4940 3871 4970 3882
rect 5002 3878 5064 3894
rect 5002 3876 5048 3878
rect 5002 3860 5064 3876
rect 5076 3860 5082 3908
rect 5085 3900 5165 3908
rect 5085 3898 5104 3900
rect 5119 3898 5153 3900
rect 5085 3882 5165 3898
rect 5085 3860 5104 3882
rect 5119 3866 5149 3882
rect 5177 3876 5183 3950
rect 5186 3876 5205 4020
rect 5220 3876 5226 4020
rect 5235 3950 5248 4020
rect 5300 4016 5322 4020
rect 5293 3994 5322 4008
rect 5375 3994 5391 4008
rect 5429 4004 5435 4006
rect 5442 4004 5550 4020
rect 5557 4004 5563 4006
rect 5571 4004 5586 4020
rect 5652 4014 5671 4017
rect 5293 3992 5391 3994
rect 5418 3992 5586 4004
rect 5601 3994 5617 4008
rect 5652 3995 5674 4014
rect 5684 4008 5700 4009
rect 5683 4006 5700 4008
rect 5684 4001 5700 4006
rect 5674 3994 5680 3995
rect 5683 3994 5712 4001
rect 5601 3993 5712 3994
rect 5601 3992 5718 3993
rect 5277 3984 5328 3992
rect 5375 3984 5409 3992
rect 5277 3972 5302 3984
rect 5309 3972 5328 3984
rect 5382 3982 5409 3984
rect 5418 3982 5639 3992
rect 5674 3989 5680 3992
rect 5382 3978 5639 3982
rect 5277 3964 5328 3972
rect 5375 3964 5639 3978
rect 5683 3984 5718 3992
rect 5229 3916 5248 3950
rect 5293 3956 5322 3964
rect 5293 3950 5310 3956
rect 5293 3948 5327 3950
rect 5375 3948 5391 3964
rect 5392 3954 5600 3964
rect 5601 3954 5617 3964
rect 5665 3960 5680 3975
rect 5683 3972 5684 3984
rect 5691 3972 5718 3984
rect 5683 3964 5718 3972
rect 5683 3963 5712 3964
rect 5403 3950 5617 3954
rect 5418 3948 5617 3950
rect 5652 3950 5665 3960
rect 5683 3950 5700 3963
rect 5652 3948 5700 3950
rect 5294 3944 5327 3948
rect 5290 3942 5327 3944
rect 5290 3941 5357 3942
rect 5290 3936 5321 3941
rect 5327 3936 5357 3941
rect 5290 3932 5357 3936
rect 5263 3929 5357 3932
rect 5263 3922 5312 3929
rect 5263 3916 5293 3922
rect 5312 3917 5317 3922
rect 5229 3900 5309 3916
rect 5321 3908 5357 3929
rect 5418 3924 5607 3948
rect 5652 3947 5699 3948
rect 5665 3942 5699 3947
rect 5433 3921 5607 3924
rect 5426 3918 5607 3921
rect 5635 3941 5699 3942
rect 5229 3898 5248 3900
rect 5263 3898 5297 3900
rect 5229 3882 5309 3898
rect 5229 3876 5248 3882
rect 4945 3850 5048 3860
rect 4899 3848 5048 3850
rect 5069 3848 5104 3860
rect 4738 3846 4900 3848
rect 4750 3826 4769 3846
rect 4784 3844 4814 3846
rect 4633 3818 4674 3826
rect 4756 3822 4769 3826
rect 4821 3830 4900 3846
rect 4932 3846 5104 3848
rect 4932 3830 5011 3846
rect 5018 3844 5048 3846
rect 4596 3808 4625 3818
rect 4639 3808 4668 3818
rect 4683 3808 4713 3822
rect 4756 3808 4799 3822
rect 4821 3818 5011 3830
rect 5076 3826 5082 3846
rect 4806 3808 4836 3818
rect 4837 3808 4995 3818
rect 4999 3808 5029 3818
rect 5033 3808 5063 3822
rect 5091 3808 5104 3846
rect 5176 3860 5205 3876
rect 5219 3860 5248 3876
rect 5263 3866 5293 3882
rect 5321 3860 5327 3908
rect 5330 3902 5349 3908
rect 5364 3902 5394 3910
rect 5330 3894 5394 3902
rect 5330 3878 5410 3894
rect 5426 3887 5488 3918
rect 5504 3887 5566 3918
rect 5635 3916 5684 3941
rect 5699 3916 5729 3932
rect 5598 3902 5628 3910
rect 5635 3908 5745 3916
rect 5598 3894 5643 3902
rect 5330 3876 5349 3878
rect 5364 3876 5410 3878
rect 5330 3860 5410 3876
rect 5437 3874 5472 3887
rect 5513 3884 5550 3887
rect 5513 3882 5555 3884
rect 5442 3871 5472 3874
rect 5451 3867 5458 3871
rect 5458 3866 5459 3867
rect 5417 3860 5427 3866
rect 5176 3852 5211 3860
rect 5176 3826 5177 3852
rect 5184 3826 5211 3852
rect 5119 3808 5149 3822
rect 5176 3818 5211 3826
rect 5213 3852 5254 3860
rect 5213 3826 5228 3852
rect 5235 3826 5254 3852
rect 5318 3848 5349 3860
rect 5364 3848 5467 3860
rect 5479 3850 5505 3876
rect 5520 3871 5550 3882
rect 5582 3878 5644 3894
rect 5582 3876 5628 3878
rect 5582 3860 5644 3876
rect 5656 3860 5662 3908
rect 5665 3900 5745 3908
rect 5665 3898 5684 3900
rect 5699 3898 5733 3900
rect 5665 3882 5745 3898
rect 5665 3860 5684 3882
rect 5699 3866 5729 3882
rect 5757 3876 5763 3950
rect 5766 3876 5785 4020
rect 5800 3876 5806 4020
rect 5815 3950 5828 4020
rect 5880 4016 5902 4020
rect 5873 3994 5902 4008
rect 5955 3994 5971 4008
rect 6009 4004 6015 4006
rect 6022 4004 6130 4020
rect 6137 4004 6143 4006
rect 6151 4004 6166 4020
rect 6232 4014 6251 4017
rect 5873 3992 5971 3994
rect 5998 3992 6166 4004
rect 6181 3994 6197 4008
rect 6232 3995 6254 4014
rect 6264 4008 6280 4009
rect 6263 4006 6280 4008
rect 6264 4001 6280 4006
rect 6254 3994 6260 3995
rect 6263 3994 6292 4001
rect 6181 3993 6292 3994
rect 6181 3992 6298 3993
rect 5857 3984 5908 3992
rect 5955 3984 5989 3992
rect 5857 3972 5882 3984
rect 5889 3972 5908 3984
rect 5962 3982 5989 3984
rect 5998 3982 6219 3992
rect 6254 3989 6260 3992
rect 5962 3978 6219 3982
rect 5857 3964 5908 3972
rect 5955 3964 6219 3978
rect 6263 3984 6298 3992
rect 5809 3916 5828 3950
rect 5873 3956 5902 3964
rect 5873 3950 5890 3956
rect 5873 3948 5907 3950
rect 5955 3948 5971 3964
rect 5972 3954 6180 3964
rect 6181 3954 6197 3964
rect 6245 3960 6260 3975
rect 6263 3972 6264 3984
rect 6271 3972 6298 3984
rect 6263 3964 6298 3972
rect 6263 3963 6292 3964
rect 5983 3950 6197 3954
rect 5998 3948 6197 3950
rect 6232 3950 6245 3960
rect 6263 3950 6280 3963
rect 6232 3948 6280 3950
rect 5874 3944 5907 3948
rect 5870 3942 5907 3944
rect 5870 3941 5937 3942
rect 5870 3936 5901 3941
rect 5907 3936 5937 3941
rect 5870 3932 5937 3936
rect 5843 3929 5937 3932
rect 5843 3922 5892 3929
rect 5843 3916 5873 3922
rect 5892 3917 5897 3922
rect 5809 3900 5889 3916
rect 5901 3908 5937 3929
rect 5998 3924 6187 3948
rect 6232 3947 6279 3948
rect 6245 3942 6279 3947
rect 6013 3921 6187 3924
rect 6006 3918 6187 3921
rect 6215 3941 6279 3942
rect 5809 3898 5828 3900
rect 5843 3898 5877 3900
rect 5809 3882 5889 3898
rect 5809 3876 5828 3882
rect 5525 3850 5628 3860
rect 5479 3848 5628 3850
rect 5649 3848 5684 3860
rect 5318 3846 5480 3848
rect 5330 3826 5349 3846
rect 5364 3844 5394 3846
rect 5213 3818 5254 3826
rect 5336 3822 5349 3826
rect 5401 3830 5480 3846
rect 5512 3846 5684 3848
rect 5512 3830 5591 3846
rect 5598 3844 5628 3846
rect 5176 3808 5205 3818
rect 5219 3808 5248 3818
rect 5263 3808 5293 3822
rect 5336 3808 5379 3822
rect 5401 3818 5591 3830
rect 5656 3826 5662 3846
rect 5386 3808 5416 3818
rect 5417 3808 5575 3818
rect 5579 3808 5609 3818
rect 5613 3808 5643 3822
rect 5671 3808 5684 3846
rect 5756 3860 5785 3876
rect 5799 3860 5828 3876
rect 5843 3866 5873 3882
rect 5901 3860 5907 3908
rect 5910 3902 5929 3908
rect 5944 3902 5974 3910
rect 5910 3894 5974 3902
rect 5910 3878 5990 3894
rect 6006 3887 6068 3918
rect 6084 3887 6146 3918
rect 6215 3916 6264 3941
rect 6279 3916 6309 3932
rect 6178 3902 6208 3910
rect 6215 3908 6325 3916
rect 6178 3894 6223 3902
rect 5910 3876 5929 3878
rect 5944 3876 5990 3878
rect 5910 3860 5990 3876
rect 6017 3874 6052 3887
rect 6093 3884 6130 3887
rect 6093 3882 6135 3884
rect 6022 3871 6052 3874
rect 6031 3867 6038 3871
rect 6038 3866 6039 3867
rect 5997 3860 6007 3866
rect 5756 3852 5791 3860
rect 5756 3826 5757 3852
rect 5764 3826 5791 3852
rect 5699 3808 5729 3822
rect 5756 3818 5791 3826
rect 5793 3852 5834 3860
rect 5793 3826 5808 3852
rect 5815 3826 5834 3852
rect 5898 3848 5929 3860
rect 5944 3848 6047 3860
rect 6059 3850 6085 3876
rect 6100 3871 6130 3882
rect 6162 3878 6224 3894
rect 6162 3876 6208 3878
rect 6162 3860 6224 3876
rect 6236 3860 6242 3908
rect 6245 3900 6325 3908
rect 6245 3898 6264 3900
rect 6279 3898 6313 3900
rect 6245 3882 6325 3898
rect 6245 3860 6264 3882
rect 6279 3866 6309 3882
rect 6337 3876 6343 3950
rect 6346 3876 6365 4020
rect 6380 3876 6386 4020
rect 6395 3950 6408 4020
rect 6460 4016 6482 4020
rect 6453 3994 6482 4008
rect 6535 3994 6551 4008
rect 6589 4004 6595 4006
rect 6602 4004 6710 4020
rect 6717 4004 6723 4006
rect 6731 4004 6746 4020
rect 6812 4014 6831 4017
rect 6453 3992 6551 3994
rect 6578 3992 6746 4004
rect 6761 3994 6777 4008
rect 6812 3995 6834 4014
rect 6844 4008 6860 4009
rect 6843 4006 6860 4008
rect 6844 4001 6860 4006
rect 6834 3994 6840 3995
rect 6843 3994 6872 4001
rect 6761 3993 6872 3994
rect 6761 3992 6878 3993
rect 6437 3984 6488 3992
rect 6535 3984 6569 3992
rect 6437 3972 6462 3984
rect 6469 3972 6488 3984
rect 6542 3982 6569 3984
rect 6578 3982 6799 3992
rect 6834 3989 6840 3992
rect 6542 3978 6799 3982
rect 6437 3964 6488 3972
rect 6535 3964 6799 3978
rect 6843 3984 6878 3992
rect 6389 3916 6408 3950
rect 6453 3956 6482 3964
rect 6453 3950 6470 3956
rect 6453 3948 6487 3950
rect 6535 3948 6551 3964
rect 6552 3954 6760 3964
rect 6761 3954 6777 3964
rect 6825 3960 6840 3975
rect 6843 3972 6844 3984
rect 6851 3972 6878 3984
rect 6843 3964 6878 3972
rect 6843 3963 6872 3964
rect 6563 3950 6777 3954
rect 6578 3948 6777 3950
rect 6812 3950 6825 3960
rect 6843 3950 6860 3963
rect 6812 3948 6860 3950
rect 6454 3944 6487 3948
rect 6450 3942 6487 3944
rect 6450 3941 6517 3942
rect 6450 3936 6481 3941
rect 6487 3936 6517 3941
rect 6450 3932 6517 3936
rect 6423 3929 6517 3932
rect 6423 3922 6472 3929
rect 6423 3916 6453 3922
rect 6472 3917 6477 3922
rect 6389 3900 6469 3916
rect 6481 3908 6517 3929
rect 6578 3924 6767 3948
rect 6812 3947 6859 3948
rect 6825 3942 6859 3947
rect 6593 3921 6767 3924
rect 6586 3918 6767 3921
rect 6795 3941 6859 3942
rect 6389 3898 6408 3900
rect 6423 3898 6457 3900
rect 6389 3882 6469 3898
rect 6389 3876 6408 3882
rect 6105 3850 6208 3860
rect 6059 3848 6208 3850
rect 6229 3848 6264 3860
rect 5898 3846 6060 3848
rect 5910 3826 5929 3846
rect 5944 3844 5974 3846
rect 5793 3818 5834 3826
rect 5916 3822 5929 3826
rect 5981 3830 6060 3846
rect 6092 3846 6264 3848
rect 6092 3830 6171 3846
rect 6178 3844 6208 3846
rect 5756 3808 5785 3818
rect 5799 3808 5828 3818
rect 5843 3808 5873 3822
rect 5916 3808 5959 3822
rect 5981 3818 6171 3830
rect 6236 3826 6242 3846
rect 5966 3808 5996 3818
rect 5997 3808 6155 3818
rect 6159 3808 6189 3818
rect 6193 3808 6223 3822
rect 6251 3808 6264 3846
rect 6336 3860 6365 3876
rect 6379 3860 6408 3876
rect 6423 3866 6453 3882
rect 6481 3860 6487 3908
rect 6490 3902 6509 3908
rect 6524 3902 6554 3910
rect 6490 3894 6554 3902
rect 6490 3878 6570 3894
rect 6586 3887 6648 3918
rect 6664 3887 6726 3918
rect 6795 3916 6844 3941
rect 6859 3916 6889 3932
rect 6758 3902 6788 3910
rect 6795 3908 6905 3916
rect 6758 3894 6803 3902
rect 6490 3876 6509 3878
rect 6524 3876 6570 3878
rect 6490 3860 6570 3876
rect 6597 3874 6632 3887
rect 6673 3884 6710 3887
rect 6673 3882 6715 3884
rect 6602 3871 6632 3874
rect 6611 3867 6618 3871
rect 6618 3866 6619 3867
rect 6577 3860 6587 3866
rect 6336 3852 6371 3860
rect 6336 3826 6337 3852
rect 6344 3826 6371 3852
rect 6279 3808 6309 3822
rect 6336 3818 6371 3826
rect 6373 3852 6414 3860
rect 6373 3826 6388 3852
rect 6395 3826 6414 3852
rect 6478 3848 6509 3860
rect 6524 3848 6627 3860
rect 6639 3850 6665 3876
rect 6680 3871 6710 3882
rect 6742 3878 6804 3894
rect 6742 3876 6788 3878
rect 6742 3860 6804 3876
rect 6816 3860 6822 3908
rect 6825 3900 6905 3908
rect 6825 3898 6844 3900
rect 6859 3898 6893 3900
rect 6825 3882 6905 3898
rect 6825 3860 6844 3882
rect 6859 3866 6889 3882
rect 6917 3876 6923 3950
rect 6926 3876 6945 4020
rect 6960 3876 6966 4020
rect 6975 3950 6988 4020
rect 7040 4016 7062 4020
rect 7033 3994 7062 4008
rect 7115 3994 7131 4008
rect 7169 4004 7175 4006
rect 7182 4004 7290 4020
rect 7297 4004 7303 4006
rect 7311 4004 7326 4020
rect 7392 4014 7411 4017
rect 7033 3992 7131 3994
rect 7158 3992 7326 4004
rect 7341 3994 7357 4008
rect 7392 3995 7414 4014
rect 7424 4008 7440 4009
rect 7423 4006 7440 4008
rect 7424 4001 7440 4006
rect 7414 3994 7420 3995
rect 7423 3994 7452 4001
rect 7341 3993 7452 3994
rect 7341 3992 7458 3993
rect 7017 3984 7068 3992
rect 7115 3984 7149 3992
rect 7017 3972 7042 3984
rect 7049 3972 7068 3984
rect 7122 3982 7149 3984
rect 7158 3982 7379 3992
rect 7414 3989 7420 3992
rect 7122 3978 7379 3982
rect 7017 3964 7068 3972
rect 7115 3964 7379 3978
rect 7423 3984 7458 3992
rect 6969 3916 6988 3950
rect 7033 3956 7062 3964
rect 7033 3950 7050 3956
rect 7033 3948 7067 3950
rect 7115 3948 7131 3964
rect 7132 3954 7340 3964
rect 7341 3954 7357 3964
rect 7405 3960 7420 3975
rect 7423 3972 7424 3984
rect 7431 3972 7458 3984
rect 7423 3964 7458 3972
rect 7423 3963 7452 3964
rect 7143 3950 7357 3954
rect 7158 3948 7357 3950
rect 7392 3950 7405 3960
rect 7423 3950 7440 3963
rect 7392 3948 7440 3950
rect 7034 3944 7067 3948
rect 7030 3942 7067 3944
rect 7030 3941 7097 3942
rect 7030 3936 7061 3941
rect 7067 3936 7097 3941
rect 7030 3932 7097 3936
rect 7003 3929 7097 3932
rect 7003 3922 7052 3929
rect 7003 3916 7033 3922
rect 7052 3917 7057 3922
rect 6969 3900 7049 3916
rect 7061 3908 7097 3929
rect 7158 3924 7347 3948
rect 7392 3947 7439 3948
rect 7405 3942 7439 3947
rect 7173 3921 7347 3924
rect 7166 3918 7347 3921
rect 7375 3941 7439 3942
rect 6969 3898 6988 3900
rect 7003 3898 7037 3900
rect 6969 3882 7049 3898
rect 6969 3876 6988 3882
rect 6685 3850 6788 3860
rect 6639 3848 6788 3850
rect 6809 3848 6844 3860
rect 6478 3846 6640 3848
rect 6490 3826 6509 3846
rect 6524 3844 6554 3846
rect 6373 3818 6414 3826
rect 6496 3822 6509 3826
rect 6561 3830 6640 3846
rect 6672 3846 6844 3848
rect 6672 3830 6751 3846
rect 6758 3844 6788 3846
rect 6336 3808 6365 3818
rect 6379 3808 6408 3818
rect 6423 3808 6453 3822
rect 6496 3808 6539 3822
rect 6561 3818 6751 3830
rect 6816 3826 6822 3846
rect 6546 3808 6576 3818
rect 6577 3808 6735 3818
rect 6739 3808 6769 3818
rect 6773 3808 6803 3822
rect 6831 3808 6844 3846
rect 6916 3860 6945 3876
rect 6959 3860 6988 3876
rect 7003 3866 7033 3882
rect 7061 3860 7067 3908
rect 7070 3902 7089 3908
rect 7104 3902 7134 3910
rect 7070 3894 7134 3902
rect 7070 3878 7150 3894
rect 7166 3887 7228 3918
rect 7244 3887 7306 3918
rect 7375 3916 7424 3941
rect 7439 3916 7469 3932
rect 7338 3902 7368 3910
rect 7375 3908 7485 3916
rect 7338 3894 7383 3902
rect 7070 3876 7089 3878
rect 7104 3876 7150 3878
rect 7070 3860 7150 3876
rect 7177 3874 7212 3887
rect 7253 3884 7290 3887
rect 7253 3882 7295 3884
rect 7182 3871 7212 3874
rect 7191 3867 7198 3871
rect 7198 3866 7199 3867
rect 7157 3860 7167 3866
rect 6916 3852 6951 3860
rect 6916 3826 6917 3852
rect 6924 3826 6951 3852
rect 6859 3808 6889 3822
rect 6916 3818 6951 3826
rect 6953 3852 6994 3860
rect 6953 3826 6968 3852
rect 6975 3826 6994 3852
rect 7058 3848 7089 3860
rect 7104 3848 7207 3860
rect 7219 3850 7245 3876
rect 7260 3871 7290 3882
rect 7322 3878 7384 3894
rect 7322 3876 7368 3878
rect 7322 3860 7384 3876
rect 7396 3860 7402 3908
rect 7405 3900 7485 3908
rect 7405 3898 7424 3900
rect 7439 3898 7473 3900
rect 7405 3882 7485 3898
rect 7405 3860 7424 3882
rect 7439 3866 7469 3882
rect 7497 3876 7503 3950
rect 7506 3876 7525 4020
rect 7540 3876 7546 4020
rect 7555 3950 7568 4020
rect 7620 4016 7642 4020
rect 7613 3994 7642 4008
rect 7695 3994 7711 4008
rect 7749 4004 7755 4006
rect 7762 4004 7870 4020
rect 7877 4004 7883 4006
rect 7891 4004 7906 4020
rect 7972 4014 7991 4017
rect 7613 3992 7711 3994
rect 7738 3992 7906 4004
rect 7921 3994 7937 4008
rect 7972 3995 7994 4014
rect 8004 4008 8020 4009
rect 8003 4006 8020 4008
rect 8004 4001 8020 4006
rect 7994 3994 8000 3995
rect 8003 3994 8032 4001
rect 7921 3993 8032 3994
rect 7921 3992 8038 3993
rect 7597 3984 7648 3992
rect 7695 3984 7729 3992
rect 7597 3972 7622 3984
rect 7629 3972 7648 3984
rect 7702 3982 7729 3984
rect 7738 3982 7959 3992
rect 7994 3989 8000 3992
rect 7702 3978 7959 3982
rect 7597 3964 7648 3972
rect 7695 3964 7959 3978
rect 8003 3984 8038 3992
rect 7549 3916 7568 3950
rect 7613 3956 7642 3964
rect 7613 3950 7630 3956
rect 7613 3948 7647 3950
rect 7695 3948 7711 3964
rect 7712 3954 7920 3964
rect 7921 3954 7937 3964
rect 7985 3960 8000 3975
rect 8003 3972 8004 3984
rect 8011 3972 8038 3984
rect 8003 3964 8038 3972
rect 8003 3963 8032 3964
rect 7723 3950 7937 3954
rect 7738 3948 7937 3950
rect 7972 3950 7985 3960
rect 8003 3950 8020 3963
rect 7972 3948 8020 3950
rect 7614 3944 7647 3948
rect 7610 3942 7647 3944
rect 7610 3941 7677 3942
rect 7610 3936 7641 3941
rect 7647 3936 7677 3941
rect 7610 3932 7677 3936
rect 7583 3929 7677 3932
rect 7583 3922 7632 3929
rect 7583 3916 7613 3922
rect 7632 3917 7637 3922
rect 7549 3900 7629 3916
rect 7641 3908 7677 3929
rect 7738 3924 7927 3948
rect 7972 3947 8019 3948
rect 7985 3942 8019 3947
rect 7753 3921 7927 3924
rect 7746 3918 7927 3921
rect 7955 3941 8019 3942
rect 7549 3898 7568 3900
rect 7583 3898 7617 3900
rect 7549 3882 7629 3898
rect 7549 3876 7568 3882
rect 7265 3850 7368 3860
rect 7219 3848 7368 3850
rect 7389 3848 7424 3860
rect 7058 3846 7220 3848
rect 7070 3826 7089 3846
rect 7104 3844 7134 3846
rect 6953 3818 6994 3826
rect 7076 3822 7089 3826
rect 7141 3830 7220 3846
rect 7252 3846 7424 3848
rect 7252 3830 7331 3846
rect 7338 3844 7368 3846
rect 6916 3808 6945 3818
rect 6959 3808 6988 3818
rect 7003 3808 7033 3822
rect 7076 3808 7119 3822
rect 7141 3818 7331 3830
rect 7396 3826 7402 3846
rect 7126 3808 7156 3818
rect 7157 3808 7315 3818
rect 7319 3808 7349 3818
rect 7353 3808 7383 3822
rect 7411 3808 7424 3846
rect 7496 3860 7525 3876
rect 7539 3860 7568 3876
rect 7583 3866 7613 3882
rect 7641 3860 7647 3908
rect 7650 3902 7669 3908
rect 7684 3902 7714 3910
rect 7650 3894 7714 3902
rect 7650 3878 7730 3894
rect 7746 3887 7808 3918
rect 7824 3887 7886 3918
rect 7955 3916 8004 3941
rect 8019 3916 8049 3932
rect 7918 3902 7948 3910
rect 7955 3908 8065 3916
rect 7918 3894 7963 3902
rect 7650 3876 7669 3878
rect 7684 3876 7730 3878
rect 7650 3860 7730 3876
rect 7757 3874 7792 3887
rect 7833 3884 7870 3887
rect 7833 3882 7875 3884
rect 7762 3871 7792 3874
rect 7771 3867 7778 3871
rect 7778 3866 7779 3867
rect 7737 3860 7747 3866
rect 7496 3852 7531 3860
rect 7496 3826 7497 3852
rect 7504 3826 7531 3852
rect 7439 3808 7469 3822
rect 7496 3818 7531 3826
rect 7533 3852 7574 3860
rect 7533 3826 7548 3852
rect 7555 3826 7574 3852
rect 7638 3848 7669 3860
rect 7684 3848 7787 3860
rect 7799 3850 7825 3876
rect 7840 3871 7870 3882
rect 7902 3878 7964 3894
rect 7902 3876 7948 3878
rect 7902 3860 7964 3876
rect 7976 3860 7982 3908
rect 7985 3900 8065 3908
rect 7985 3898 8004 3900
rect 8019 3898 8053 3900
rect 7985 3882 8065 3898
rect 7985 3860 8004 3882
rect 8019 3866 8049 3882
rect 8077 3876 8083 3950
rect 8086 3876 8105 4020
rect 8120 3876 8126 4020
rect 8135 3950 8148 4020
rect 8200 4016 8222 4020
rect 8193 3994 8222 4008
rect 8275 3994 8291 4008
rect 8329 4004 8335 4006
rect 8342 4004 8450 4020
rect 8457 4004 8463 4006
rect 8471 4004 8486 4020
rect 8552 4014 8571 4017
rect 8193 3992 8291 3994
rect 8318 3992 8486 4004
rect 8501 3994 8517 4008
rect 8552 3995 8574 4014
rect 8584 4008 8600 4009
rect 8583 4006 8600 4008
rect 8584 4001 8600 4006
rect 8574 3994 8580 3995
rect 8583 3994 8612 4001
rect 8501 3993 8612 3994
rect 8501 3992 8618 3993
rect 8177 3984 8228 3992
rect 8275 3984 8309 3992
rect 8177 3972 8202 3984
rect 8209 3972 8228 3984
rect 8282 3982 8309 3984
rect 8318 3982 8539 3992
rect 8574 3989 8580 3992
rect 8282 3978 8539 3982
rect 8177 3964 8228 3972
rect 8275 3964 8539 3978
rect 8583 3984 8618 3992
rect 8129 3916 8148 3950
rect 8193 3956 8222 3964
rect 8193 3950 8210 3956
rect 8193 3948 8227 3950
rect 8275 3948 8291 3964
rect 8292 3954 8500 3964
rect 8501 3954 8517 3964
rect 8565 3960 8580 3975
rect 8583 3972 8584 3984
rect 8591 3972 8618 3984
rect 8583 3964 8618 3972
rect 8583 3963 8612 3964
rect 8303 3950 8517 3954
rect 8318 3948 8517 3950
rect 8552 3950 8565 3960
rect 8583 3950 8600 3963
rect 8552 3948 8600 3950
rect 8194 3944 8227 3948
rect 8190 3942 8227 3944
rect 8190 3941 8257 3942
rect 8190 3936 8221 3941
rect 8227 3936 8257 3941
rect 8190 3932 8257 3936
rect 8163 3929 8257 3932
rect 8163 3922 8212 3929
rect 8163 3916 8193 3922
rect 8212 3917 8217 3922
rect 8129 3900 8209 3916
rect 8221 3908 8257 3929
rect 8318 3924 8507 3948
rect 8552 3947 8599 3948
rect 8565 3942 8599 3947
rect 8333 3921 8507 3924
rect 8326 3918 8507 3921
rect 8535 3941 8599 3942
rect 8129 3898 8148 3900
rect 8163 3898 8197 3900
rect 8129 3882 8209 3898
rect 8129 3876 8148 3882
rect 7845 3850 7948 3860
rect 7799 3848 7948 3850
rect 7969 3848 8004 3860
rect 7638 3846 7800 3848
rect 7650 3826 7669 3846
rect 7684 3844 7714 3846
rect 7533 3818 7574 3826
rect 7656 3822 7669 3826
rect 7721 3830 7800 3846
rect 7832 3846 8004 3848
rect 7832 3830 7911 3846
rect 7918 3844 7948 3846
rect 7496 3808 7525 3818
rect 7539 3808 7568 3818
rect 7583 3808 7613 3822
rect 7656 3808 7699 3822
rect 7721 3818 7911 3830
rect 7976 3826 7982 3846
rect 7706 3808 7736 3818
rect 7737 3808 7895 3818
rect 7899 3808 7929 3818
rect 7933 3808 7963 3822
rect 7991 3808 8004 3846
rect 8076 3860 8105 3876
rect 8119 3860 8148 3876
rect 8163 3866 8193 3882
rect 8221 3860 8227 3908
rect 8230 3902 8249 3908
rect 8264 3902 8294 3910
rect 8230 3894 8294 3902
rect 8230 3878 8310 3894
rect 8326 3887 8388 3918
rect 8404 3887 8466 3918
rect 8535 3916 8584 3941
rect 8599 3916 8629 3932
rect 8498 3902 8528 3910
rect 8535 3908 8645 3916
rect 8498 3894 8543 3902
rect 8230 3876 8249 3878
rect 8264 3876 8310 3878
rect 8230 3860 8310 3876
rect 8337 3874 8372 3887
rect 8413 3884 8450 3887
rect 8413 3882 8455 3884
rect 8342 3871 8372 3874
rect 8351 3867 8358 3871
rect 8358 3866 8359 3867
rect 8317 3860 8327 3866
rect 8076 3852 8111 3860
rect 8076 3826 8077 3852
rect 8084 3826 8111 3852
rect 8019 3808 8049 3822
rect 8076 3818 8111 3826
rect 8113 3852 8154 3860
rect 8113 3826 8128 3852
rect 8135 3826 8154 3852
rect 8218 3848 8249 3860
rect 8264 3848 8367 3860
rect 8379 3850 8405 3876
rect 8420 3871 8450 3882
rect 8482 3878 8544 3894
rect 8482 3876 8528 3878
rect 8482 3860 8544 3876
rect 8556 3860 8562 3908
rect 8565 3900 8645 3908
rect 8565 3898 8584 3900
rect 8599 3898 8633 3900
rect 8565 3882 8645 3898
rect 8565 3860 8584 3882
rect 8599 3866 8629 3882
rect 8657 3876 8663 3950
rect 8666 3876 8685 4020
rect 8700 3876 8706 4020
rect 8715 3950 8728 4020
rect 8780 4016 8802 4020
rect 8773 3994 8802 4008
rect 8855 3994 8871 4008
rect 8909 4004 8915 4006
rect 8922 4004 9030 4020
rect 9037 4004 9043 4006
rect 9051 4004 9066 4020
rect 9132 4014 9151 4017
rect 8773 3992 8871 3994
rect 8898 3992 9066 4004
rect 9081 3994 9097 4008
rect 9132 3995 9154 4014
rect 9164 4008 9180 4009
rect 9163 4006 9180 4008
rect 9164 4001 9180 4006
rect 9154 3994 9160 3995
rect 9163 3994 9192 4001
rect 9081 3993 9192 3994
rect 9081 3992 9198 3993
rect 8757 3984 8808 3992
rect 8855 3984 8889 3992
rect 8757 3972 8782 3984
rect 8789 3972 8808 3984
rect 8862 3982 8889 3984
rect 8898 3982 9119 3992
rect 9154 3989 9160 3992
rect 8862 3978 9119 3982
rect 8757 3964 8808 3972
rect 8855 3964 9119 3978
rect 9163 3984 9198 3992
rect 8709 3916 8728 3950
rect 8773 3956 8802 3964
rect 8773 3950 8790 3956
rect 8773 3948 8807 3950
rect 8855 3948 8871 3964
rect 8872 3954 9080 3964
rect 9081 3954 9097 3964
rect 9145 3960 9160 3975
rect 9163 3972 9164 3984
rect 9171 3972 9198 3984
rect 9163 3964 9198 3972
rect 9163 3963 9192 3964
rect 8883 3950 9097 3954
rect 8898 3948 9097 3950
rect 9132 3950 9145 3960
rect 9163 3950 9180 3963
rect 9132 3948 9180 3950
rect 8774 3944 8807 3948
rect 8770 3942 8807 3944
rect 8770 3941 8837 3942
rect 8770 3936 8801 3941
rect 8807 3936 8837 3941
rect 8770 3932 8837 3936
rect 8743 3929 8837 3932
rect 8743 3922 8792 3929
rect 8743 3916 8773 3922
rect 8792 3917 8797 3922
rect 8709 3900 8789 3916
rect 8801 3908 8837 3929
rect 8898 3924 9087 3948
rect 9132 3947 9179 3948
rect 9145 3942 9179 3947
rect 8913 3921 9087 3924
rect 8906 3918 9087 3921
rect 9115 3941 9179 3942
rect 8709 3898 8728 3900
rect 8743 3898 8777 3900
rect 8709 3882 8789 3898
rect 8709 3876 8728 3882
rect 8425 3850 8528 3860
rect 8379 3848 8528 3850
rect 8549 3848 8584 3860
rect 8218 3846 8380 3848
rect 8230 3826 8249 3846
rect 8264 3844 8294 3846
rect 8113 3818 8154 3826
rect 8236 3822 8249 3826
rect 8301 3830 8380 3846
rect 8412 3846 8584 3848
rect 8412 3830 8491 3846
rect 8498 3844 8528 3846
rect 8076 3808 8105 3818
rect 8119 3808 8148 3818
rect 8163 3808 8193 3822
rect 8236 3808 8279 3822
rect 8301 3818 8491 3830
rect 8556 3826 8562 3846
rect 8286 3808 8316 3818
rect 8317 3808 8475 3818
rect 8479 3808 8509 3818
rect 8513 3808 8543 3822
rect 8571 3808 8584 3846
rect 8656 3860 8685 3876
rect 8699 3860 8728 3876
rect 8743 3866 8773 3882
rect 8801 3860 8807 3908
rect 8810 3902 8829 3908
rect 8844 3902 8874 3910
rect 8810 3894 8874 3902
rect 8810 3878 8890 3894
rect 8906 3887 8968 3918
rect 8984 3887 9046 3918
rect 9115 3916 9164 3941
rect 9179 3916 9209 3932
rect 9078 3902 9108 3910
rect 9115 3908 9225 3916
rect 9078 3894 9123 3902
rect 8810 3876 8829 3878
rect 8844 3876 8890 3878
rect 8810 3860 8890 3876
rect 8917 3874 8952 3887
rect 8993 3884 9030 3887
rect 8993 3882 9035 3884
rect 8922 3871 8952 3874
rect 8931 3867 8938 3871
rect 8938 3866 8939 3867
rect 8897 3860 8907 3866
rect 8656 3852 8691 3860
rect 8656 3826 8657 3852
rect 8664 3826 8691 3852
rect 8599 3808 8629 3822
rect 8656 3818 8691 3826
rect 8693 3852 8734 3860
rect 8693 3826 8708 3852
rect 8715 3826 8734 3852
rect 8798 3848 8829 3860
rect 8844 3848 8947 3860
rect 8959 3850 8985 3876
rect 9000 3871 9030 3882
rect 9062 3878 9124 3894
rect 9062 3876 9108 3878
rect 9062 3860 9124 3876
rect 9136 3860 9142 3908
rect 9145 3900 9225 3908
rect 9145 3898 9164 3900
rect 9179 3898 9213 3900
rect 9145 3882 9225 3898
rect 9145 3860 9164 3882
rect 9179 3866 9209 3882
rect 9237 3876 9243 3950
rect 9246 3876 9265 4020
rect 9280 3876 9286 4020
rect 9295 3950 9308 4020
rect 9360 4016 9382 4020
rect 9353 3994 9382 4008
rect 9435 3994 9451 4008
rect 9489 4004 9495 4006
rect 9502 4004 9610 4020
rect 9617 4004 9623 4006
rect 9631 4004 9646 4020
rect 9712 4014 9731 4017
rect 9353 3992 9451 3994
rect 9478 3992 9646 4004
rect 9661 3994 9677 4008
rect 9712 3995 9734 4014
rect 9744 4008 9760 4009
rect 9743 4006 9760 4008
rect 9744 4001 9760 4006
rect 9734 3994 9740 3995
rect 9743 3994 9772 4001
rect 9661 3993 9772 3994
rect 9661 3992 9778 3993
rect 9337 3984 9388 3992
rect 9435 3984 9469 3992
rect 9337 3972 9362 3984
rect 9369 3972 9388 3984
rect 9442 3982 9469 3984
rect 9478 3982 9699 3992
rect 9734 3989 9740 3992
rect 9442 3978 9699 3982
rect 9337 3964 9388 3972
rect 9435 3964 9699 3978
rect 9743 3984 9778 3992
rect 9289 3916 9308 3950
rect 9353 3956 9382 3964
rect 9353 3950 9370 3956
rect 9353 3948 9387 3950
rect 9435 3948 9451 3964
rect 9452 3954 9660 3964
rect 9661 3954 9677 3964
rect 9725 3960 9740 3975
rect 9743 3972 9744 3984
rect 9751 3972 9778 3984
rect 9743 3964 9778 3972
rect 9743 3963 9772 3964
rect 9463 3950 9677 3954
rect 9478 3948 9677 3950
rect 9712 3950 9725 3960
rect 9743 3950 9760 3963
rect 9712 3948 9760 3950
rect 9354 3944 9387 3948
rect 9350 3942 9387 3944
rect 9350 3941 9417 3942
rect 9350 3936 9381 3941
rect 9387 3936 9417 3941
rect 9350 3932 9417 3936
rect 9323 3929 9417 3932
rect 9323 3922 9372 3929
rect 9323 3916 9353 3922
rect 9372 3917 9377 3922
rect 9289 3900 9369 3916
rect 9381 3908 9417 3929
rect 9478 3924 9667 3948
rect 9712 3947 9759 3948
rect 9725 3942 9759 3947
rect 9493 3921 9667 3924
rect 9486 3918 9667 3921
rect 9695 3941 9759 3942
rect 9289 3898 9308 3900
rect 9323 3898 9357 3900
rect 9289 3882 9369 3898
rect 9289 3876 9308 3882
rect 9005 3850 9108 3860
rect 8959 3848 9108 3850
rect 9129 3848 9164 3860
rect 8798 3846 8960 3848
rect 8810 3826 8829 3846
rect 8844 3844 8874 3846
rect 8693 3818 8734 3826
rect 8816 3822 8829 3826
rect 8881 3830 8960 3846
rect 8992 3846 9164 3848
rect 8992 3830 9071 3846
rect 9078 3844 9108 3846
rect 8656 3808 8685 3818
rect 8699 3808 8728 3818
rect 8743 3808 8773 3822
rect 8816 3808 8859 3822
rect 8881 3818 9071 3830
rect 9136 3826 9142 3846
rect 8866 3808 8896 3818
rect 8897 3808 9055 3818
rect 9059 3808 9089 3818
rect 9093 3808 9123 3822
rect 9151 3808 9164 3846
rect 9236 3860 9265 3876
rect 9279 3860 9308 3876
rect 9323 3866 9353 3882
rect 9381 3860 9387 3908
rect 9390 3902 9409 3908
rect 9424 3902 9454 3910
rect 9390 3894 9454 3902
rect 9390 3878 9470 3894
rect 9486 3887 9548 3918
rect 9564 3887 9626 3918
rect 9695 3916 9744 3941
rect 9759 3916 9789 3932
rect 9658 3902 9688 3910
rect 9695 3908 9805 3916
rect 9658 3894 9703 3902
rect 9390 3876 9409 3878
rect 9424 3876 9470 3878
rect 9390 3860 9470 3876
rect 9497 3874 9532 3887
rect 9573 3884 9610 3887
rect 9573 3882 9615 3884
rect 9502 3871 9532 3874
rect 9511 3867 9518 3871
rect 9518 3866 9519 3867
rect 9477 3860 9487 3866
rect 9236 3852 9271 3860
rect 9236 3826 9237 3852
rect 9244 3826 9271 3852
rect 9179 3808 9209 3822
rect 9236 3818 9271 3826
rect 9273 3852 9314 3860
rect 9273 3826 9288 3852
rect 9295 3826 9314 3852
rect 9378 3848 9409 3860
rect 9424 3848 9527 3860
rect 9539 3850 9565 3876
rect 9580 3871 9610 3882
rect 9642 3878 9704 3894
rect 9642 3876 9688 3878
rect 9642 3860 9704 3876
rect 9716 3860 9722 3908
rect 9725 3900 9805 3908
rect 9725 3898 9744 3900
rect 9759 3898 9793 3900
rect 9725 3882 9805 3898
rect 9725 3860 9744 3882
rect 9759 3866 9789 3882
rect 9817 3876 9823 3950
rect 9826 3876 9845 4020
rect 9860 3876 9866 4020
rect 9875 3950 9888 4020
rect 9940 4016 9962 4020
rect 9933 3994 9962 4008
rect 10015 3994 10031 4008
rect 10069 4004 10075 4006
rect 10082 4004 10190 4020
rect 10197 4004 10203 4006
rect 10211 4004 10226 4020
rect 10292 4014 10311 4017
rect 9933 3992 10031 3994
rect 10058 3992 10226 4004
rect 10241 3994 10257 4008
rect 10292 3995 10314 4014
rect 10324 4008 10340 4009
rect 10323 4006 10340 4008
rect 10324 4001 10340 4006
rect 10314 3994 10320 3995
rect 10323 3994 10352 4001
rect 10241 3993 10352 3994
rect 10241 3992 10358 3993
rect 9917 3984 9968 3992
rect 10015 3984 10049 3992
rect 9917 3972 9942 3984
rect 9949 3972 9968 3984
rect 10022 3982 10049 3984
rect 10058 3982 10279 3992
rect 10314 3989 10320 3992
rect 10022 3978 10279 3982
rect 9917 3964 9968 3972
rect 10015 3964 10279 3978
rect 10323 3984 10358 3992
rect 9869 3916 9888 3950
rect 9933 3956 9962 3964
rect 9933 3950 9950 3956
rect 9933 3948 9967 3950
rect 10015 3948 10031 3964
rect 10032 3954 10240 3964
rect 10241 3954 10257 3964
rect 10305 3960 10320 3975
rect 10323 3972 10324 3984
rect 10331 3972 10358 3984
rect 10323 3964 10358 3972
rect 10323 3963 10352 3964
rect 10043 3950 10257 3954
rect 10058 3948 10257 3950
rect 10292 3950 10305 3960
rect 10323 3950 10340 3963
rect 10292 3948 10340 3950
rect 9934 3944 9967 3948
rect 9930 3942 9967 3944
rect 9930 3941 9997 3942
rect 9930 3936 9961 3941
rect 9967 3936 9997 3941
rect 9930 3932 9997 3936
rect 9903 3929 9997 3932
rect 9903 3922 9952 3929
rect 9903 3916 9933 3922
rect 9952 3917 9957 3922
rect 9869 3900 9949 3916
rect 9961 3908 9997 3929
rect 10058 3924 10247 3948
rect 10292 3947 10339 3948
rect 10305 3942 10339 3947
rect 10073 3921 10247 3924
rect 10066 3918 10247 3921
rect 10275 3941 10339 3942
rect 9869 3898 9888 3900
rect 9903 3898 9937 3900
rect 9869 3882 9949 3898
rect 9869 3876 9888 3882
rect 9585 3850 9688 3860
rect 9539 3848 9688 3850
rect 9709 3848 9744 3860
rect 9378 3846 9540 3848
rect 9390 3826 9409 3846
rect 9424 3844 9454 3846
rect 9273 3818 9314 3826
rect 9396 3822 9409 3826
rect 9461 3830 9540 3846
rect 9572 3846 9744 3848
rect 9572 3830 9651 3846
rect 9658 3844 9688 3846
rect 9236 3808 9265 3818
rect 9279 3808 9308 3818
rect 9323 3808 9353 3822
rect 9396 3808 9439 3822
rect 9461 3818 9651 3830
rect 9716 3826 9722 3846
rect 9446 3808 9476 3818
rect 9477 3808 9635 3818
rect 9639 3808 9669 3818
rect 9673 3808 9703 3822
rect 9731 3808 9744 3846
rect 9816 3860 9845 3876
rect 9859 3860 9888 3876
rect 9903 3866 9933 3882
rect 9961 3860 9967 3908
rect 9970 3902 9989 3908
rect 10004 3902 10034 3910
rect 9970 3894 10034 3902
rect 9970 3878 10050 3894
rect 10066 3887 10128 3918
rect 10144 3887 10206 3918
rect 10275 3916 10324 3941
rect 10339 3916 10369 3932
rect 10238 3902 10268 3910
rect 10275 3908 10385 3916
rect 10238 3894 10283 3902
rect 9970 3876 9989 3878
rect 10004 3876 10050 3878
rect 9970 3860 10050 3876
rect 10077 3874 10112 3887
rect 10153 3884 10190 3887
rect 10153 3882 10195 3884
rect 10082 3871 10112 3874
rect 10091 3867 10098 3871
rect 10098 3866 10099 3867
rect 10057 3860 10067 3866
rect 9816 3852 9851 3860
rect 9816 3826 9817 3852
rect 9824 3826 9851 3852
rect 9759 3808 9789 3822
rect 9816 3818 9851 3826
rect 9853 3852 9894 3860
rect 9853 3826 9868 3852
rect 9875 3826 9894 3852
rect 9958 3848 9989 3860
rect 10004 3848 10107 3860
rect 10119 3850 10145 3876
rect 10160 3871 10190 3882
rect 10222 3878 10284 3894
rect 10222 3876 10268 3878
rect 10222 3860 10284 3876
rect 10296 3860 10302 3908
rect 10305 3900 10385 3908
rect 10305 3898 10324 3900
rect 10339 3898 10373 3900
rect 10305 3882 10385 3898
rect 10305 3860 10324 3882
rect 10339 3866 10369 3882
rect 10397 3876 10403 3950
rect 10406 3876 10425 4020
rect 10440 3876 10446 4020
rect 10455 3950 10468 4020
rect 10520 4016 10542 4020
rect 10513 3994 10542 4008
rect 10595 3994 10611 4008
rect 10649 4004 10655 4006
rect 10662 4004 10770 4020
rect 10777 4004 10783 4006
rect 10791 4004 10806 4020
rect 10872 4014 10891 4017
rect 10513 3992 10611 3994
rect 10638 3992 10806 4004
rect 10821 3994 10837 4008
rect 10872 3995 10894 4014
rect 10904 4008 10920 4009
rect 10903 4006 10920 4008
rect 10904 4001 10920 4006
rect 10894 3994 10900 3995
rect 10903 3994 10932 4001
rect 10821 3993 10932 3994
rect 10821 3992 10938 3993
rect 10497 3984 10548 3992
rect 10595 3984 10629 3992
rect 10497 3972 10522 3984
rect 10529 3972 10548 3984
rect 10602 3982 10629 3984
rect 10638 3982 10859 3992
rect 10894 3989 10900 3992
rect 10602 3978 10859 3982
rect 10497 3964 10548 3972
rect 10595 3964 10859 3978
rect 10903 3984 10938 3992
rect 10449 3916 10468 3950
rect 10513 3956 10542 3964
rect 10513 3950 10530 3956
rect 10513 3948 10547 3950
rect 10595 3948 10611 3964
rect 10612 3954 10820 3964
rect 10821 3954 10837 3964
rect 10885 3960 10900 3975
rect 10903 3972 10904 3984
rect 10911 3972 10938 3984
rect 10903 3964 10938 3972
rect 10903 3963 10932 3964
rect 10623 3950 10837 3954
rect 10638 3948 10837 3950
rect 10872 3950 10885 3960
rect 10903 3950 10920 3963
rect 10872 3948 10920 3950
rect 10514 3944 10547 3948
rect 10510 3942 10547 3944
rect 10510 3941 10577 3942
rect 10510 3936 10541 3941
rect 10547 3936 10577 3941
rect 10510 3932 10577 3936
rect 10483 3929 10577 3932
rect 10483 3922 10532 3929
rect 10483 3916 10513 3922
rect 10532 3917 10537 3922
rect 10449 3900 10529 3916
rect 10541 3908 10577 3929
rect 10638 3924 10827 3948
rect 10872 3947 10919 3948
rect 10885 3942 10919 3947
rect 10653 3921 10827 3924
rect 10646 3918 10827 3921
rect 10855 3941 10919 3942
rect 10449 3898 10468 3900
rect 10483 3898 10517 3900
rect 10449 3882 10529 3898
rect 10449 3876 10468 3882
rect 10165 3850 10268 3860
rect 10119 3848 10268 3850
rect 10289 3848 10324 3860
rect 9958 3846 10120 3848
rect 9970 3826 9989 3846
rect 10004 3844 10034 3846
rect 9853 3818 9894 3826
rect 9976 3822 9989 3826
rect 10041 3830 10120 3846
rect 10152 3846 10324 3848
rect 10152 3830 10231 3846
rect 10238 3844 10268 3846
rect 9816 3808 9845 3818
rect 9859 3808 9888 3818
rect 9903 3808 9933 3822
rect 9976 3808 10019 3822
rect 10041 3818 10231 3830
rect 10296 3826 10302 3846
rect 10026 3808 10056 3818
rect 10057 3808 10215 3818
rect 10219 3808 10249 3818
rect 10253 3808 10283 3822
rect 10311 3808 10324 3846
rect 10396 3860 10425 3876
rect 10439 3860 10468 3876
rect 10483 3866 10513 3882
rect 10541 3860 10547 3908
rect 10550 3902 10569 3908
rect 10584 3902 10614 3910
rect 10550 3894 10614 3902
rect 10550 3878 10630 3894
rect 10646 3887 10708 3918
rect 10724 3887 10786 3918
rect 10855 3916 10904 3941
rect 10919 3916 10949 3932
rect 10818 3902 10848 3910
rect 10855 3908 10965 3916
rect 10818 3894 10863 3902
rect 10550 3876 10569 3878
rect 10584 3876 10630 3878
rect 10550 3860 10630 3876
rect 10657 3874 10692 3887
rect 10733 3884 10770 3887
rect 10733 3882 10775 3884
rect 10662 3871 10692 3874
rect 10671 3867 10678 3871
rect 10678 3866 10679 3867
rect 10637 3860 10647 3866
rect 10396 3852 10431 3860
rect 10396 3826 10397 3852
rect 10404 3826 10431 3852
rect 10339 3808 10369 3822
rect 10396 3818 10431 3826
rect 10433 3852 10474 3860
rect 10433 3826 10448 3852
rect 10455 3826 10474 3852
rect 10538 3848 10569 3860
rect 10584 3848 10687 3860
rect 10699 3850 10725 3876
rect 10740 3871 10770 3882
rect 10802 3878 10864 3894
rect 10802 3876 10848 3878
rect 10802 3860 10864 3876
rect 10876 3860 10882 3908
rect 10885 3900 10965 3908
rect 10885 3898 10904 3900
rect 10919 3898 10953 3900
rect 10885 3882 10965 3898
rect 10885 3860 10904 3882
rect 10919 3866 10949 3882
rect 10977 3876 10983 3950
rect 10986 3876 11005 4020
rect 11020 3876 11026 4020
rect 11035 3950 11048 4020
rect 11100 4016 11122 4020
rect 11093 3994 11122 4008
rect 11175 3994 11191 4008
rect 11229 4004 11235 4006
rect 11242 4004 11350 4020
rect 11357 4004 11363 4006
rect 11371 4004 11386 4020
rect 11452 4014 11471 4017
rect 11093 3992 11191 3994
rect 11218 3992 11386 4004
rect 11401 3994 11417 4008
rect 11452 3995 11474 4014
rect 11484 4008 11500 4009
rect 11483 4006 11500 4008
rect 11484 4001 11500 4006
rect 11474 3994 11480 3995
rect 11483 3994 11512 4001
rect 11401 3993 11512 3994
rect 11401 3992 11518 3993
rect 11077 3984 11128 3992
rect 11175 3984 11209 3992
rect 11077 3972 11102 3984
rect 11109 3972 11128 3984
rect 11182 3982 11209 3984
rect 11218 3982 11439 3992
rect 11474 3989 11480 3992
rect 11182 3978 11439 3982
rect 11077 3964 11128 3972
rect 11175 3964 11439 3978
rect 11483 3984 11518 3992
rect 11029 3916 11048 3950
rect 11093 3956 11122 3964
rect 11093 3950 11110 3956
rect 11093 3948 11127 3950
rect 11175 3948 11191 3964
rect 11192 3954 11400 3964
rect 11401 3954 11417 3964
rect 11465 3960 11480 3975
rect 11483 3972 11484 3984
rect 11491 3972 11518 3984
rect 11483 3964 11518 3972
rect 11483 3963 11512 3964
rect 11203 3950 11417 3954
rect 11218 3948 11417 3950
rect 11452 3950 11465 3960
rect 11483 3950 11500 3963
rect 11452 3948 11500 3950
rect 11094 3944 11127 3948
rect 11090 3942 11127 3944
rect 11090 3941 11157 3942
rect 11090 3936 11121 3941
rect 11127 3936 11157 3941
rect 11090 3932 11157 3936
rect 11063 3929 11157 3932
rect 11063 3922 11112 3929
rect 11063 3916 11093 3922
rect 11112 3917 11117 3922
rect 11029 3900 11109 3916
rect 11121 3908 11157 3929
rect 11218 3924 11407 3948
rect 11452 3947 11499 3948
rect 11465 3942 11499 3947
rect 11233 3921 11407 3924
rect 11226 3918 11407 3921
rect 11435 3941 11499 3942
rect 11029 3898 11048 3900
rect 11063 3898 11097 3900
rect 11029 3882 11109 3898
rect 11029 3876 11048 3882
rect 10745 3850 10848 3860
rect 10699 3848 10848 3850
rect 10869 3848 10904 3860
rect 10538 3846 10700 3848
rect 10550 3826 10569 3846
rect 10584 3844 10614 3846
rect 10433 3818 10474 3826
rect 10556 3822 10569 3826
rect 10621 3830 10700 3846
rect 10732 3846 10904 3848
rect 10732 3830 10811 3846
rect 10818 3844 10848 3846
rect 10396 3808 10425 3818
rect 10439 3808 10468 3818
rect 10483 3808 10513 3822
rect 10556 3808 10599 3822
rect 10621 3818 10811 3830
rect 10876 3826 10882 3846
rect 10606 3808 10636 3818
rect 10637 3808 10795 3818
rect 10799 3808 10829 3818
rect 10833 3808 10863 3822
rect 10891 3808 10904 3846
rect 10976 3860 11005 3876
rect 11019 3860 11048 3876
rect 11063 3866 11093 3882
rect 11121 3860 11127 3908
rect 11130 3902 11149 3908
rect 11164 3902 11194 3910
rect 11130 3894 11194 3902
rect 11130 3878 11210 3894
rect 11226 3887 11288 3918
rect 11304 3887 11366 3918
rect 11435 3916 11484 3941
rect 11499 3916 11529 3932
rect 11398 3902 11428 3910
rect 11435 3908 11545 3916
rect 11398 3894 11443 3902
rect 11130 3876 11149 3878
rect 11164 3876 11210 3878
rect 11130 3860 11210 3876
rect 11237 3874 11272 3887
rect 11313 3884 11350 3887
rect 11313 3882 11355 3884
rect 11242 3871 11272 3874
rect 11251 3867 11258 3871
rect 11258 3866 11259 3867
rect 11217 3860 11227 3866
rect 10976 3852 11011 3860
rect 10976 3826 10977 3852
rect 10984 3826 11011 3852
rect 10919 3808 10949 3822
rect 10976 3818 11011 3826
rect 11013 3852 11054 3860
rect 11013 3826 11028 3852
rect 11035 3826 11054 3852
rect 11118 3848 11149 3860
rect 11164 3848 11267 3860
rect 11279 3850 11305 3876
rect 11320 3871 11350 3882
rect 11382 3878 11444 3894
rect 11382 3876 11428 3878
rect 11382 3860 11444 3876
rect 11456 3860 11462 3908
rect 11465 3900 11545 3908
rect 11465 3898 11484 3900
rect 11499 3898 11533 3900
rect 11465 3882 11545 3898
rect 11465 3860 11484 3882
rect 11499 3866 11529 3882
rect 11557 3876 11563 3950
rect 11566 3876 11585 4020
rect 11600 3876 11606 4020
rect 11615 3950 11628 4020
rect 11680 4016 11702 4020
rect 11673 3994 11702 4008
rect 11755 3994 11771 4008
rect 11809 4004 11815 4006
rect 11822 4004 11930 4020
rect 11937 4004 11943 4006
rect 11951 4004 11966 4020
rect 12032 4014 12051 4017
rect 11673 3992 11771 3994
rect 11798 3992 11966 4004
rect 11981 3994 11997 4008
rect 12032 3995 12054 4014
rect 12064 4008 12080 4009
rect 12063 4006 12080 4008
rect 12064 4001 12080 4006
rect 12054 3994 12060 3995
rect 12063 3994 12092 4001
rect 11981 3993 12092 3994
rect 11981 3992 12098 3993
rect 11657 3984 11708 3992
rect 11755 3984 11789 3992
rect 11657 3972 11682 3984
rect 11689 3972 11708 3984
rect 11762 3982 11789 3984
rect 11798 3982 12019 3992
rect 12054 3989 12060 3992
rect 11762 3978 12019 3982
rect 11657 3964 11708 3972
rect 11755 3964 12019 3978
rect 12063 3984 12098 3992
rect 11609 3916 11628 3950
rect 11673 3956 11702 3964
rect 11673 3950 11690 3956
rect 11673 3948 11707 3950
rect 11755 3948 11771 3964
rect 11772 3954 11980 3964
rect 11981 3954 11997 3964
rect 12045 3960 12060 3975
rect 12063 3972 12064 3984
rect 12071 3972 12098 3984
rect 12063 3964 12098 3972
rect 12063 3963 12092 3964
rect 11783 3950 11997 3954
rect 11798 3948 11997 3950
rect 12032 3950 12045 3960
rect 12063 3950 12080 3963
rect 12032 3948 12080 3950
rect 11674 3944 11707 3948
rect 11670 3942 11707 3944
rect 11670 3941 11737 3942
rect 11670 3936 11701 3941
rect 11707 3936 11737 3941
rect 11670 3932 11737 3936
rect 11643 3929 11737 3932
rect 11643 3922 11692 3929
rect 11643 3916 11673 3922
rect 11692 3917 11697 3922
rect 11609 3900 11689 3916
rect 11701 3908 11737 3929
rect 11798 3924 11987 3948
rect 12032 3947 12079 3948
rect 12045 3942 12079 3947
rect 11813 3921 11987 3924
rect 11806 3918 11987 3921
rect 12015 3941 12079 3942
rect 11609 3898 11628 3900
rect 11643 3898 11677 3900
rect 11609 3882 11689 3898
rect 11609 3876 11628 3882
rect 11325 3850 11428 3860
rect 11279 3848 11428 3850
rect 11449 3848 11484 3860
rect 11118 3846 11280 3848
rect 11130 3826 11149 3846
rect 11164 3844 11194 3846
rect 11013 3818 11054 3826
rect 11136 3822 11149 3826
rect 11201 3830 11280 3846
rect 11312 3846 11484 3848
rect 11312 3830 11391 3846
rect 11398 3844 11428 3846
rect 10976 3808 11005 3818
rect 11019 3808 11048 3818
rect 11063 3808 11093 3822
rect 11136 3808 11179 3822
rect 11201 3818 11391 3830
rect 11456 3826 11462 3846
rect 11186 3808 11216 3818
rect 11217 3808 11375 3818
rect 11379 3808 11409 3818
rect 11413 3808 11443 3822
rect 11471 3808 11484 3846
rect 11556 3860 11585 3876
rect 11599 3860 11628 3876
rect 11643 3866 11673 3882
rect 11701 3860 11707 3908
rect 11710 3902 11729 3908
rect 11744 3902 11774 3910
rect 11710 3894 11774 3902
rect 11710 3878 11790 3894
rect 11806 3887 11868 3918
rect 11884 3887 11946 3918
rect 12015 3916 12064 3941
rect 12079 3916 12109 3932
rect 11978 3902 12008 3910
rect 12015 3908 12125 3916
rect 11978 3894 12023 3902
rect 11710 3876 11729 3878
rect 11744 3876 11790 3878
rect 11710 3860 11790 3876
rect 11817 3874 11852 3887
rect 11893 3884 11930 3887
rect 11893 3882 11935 3884
rect 11822 3871 11852 3874
rect 11831 3867 11838 3871
rect 11838 3866 11839 3867
rect 11797 3860 11807 3866
rect 11556 3852 11591 3860
rect 11556 3826 11557 3852
rect 11564 3826 11591 3852
rect 11499 3808 11529 3822
rect 11556 3818 11591 3826
rect 11593 3852 11634 3860
rect 11593 3826 11608 3852
rect 11615 3826 11634 3852
rect 11698 3848 11729 3860
rect 11744 3848 11847 3860
rect 11859 3850 11885 3876
rect 11900 3871 11930 3882
rect 11962 3878 12024 3894
rect 11962 3876 12008 3878
rect 11962 3860 12024 3876
rect 12036 3860 12042 3908
rect 12045 3900 12125 3908
rect 12045 3898 12064 3900
rect 12079 3898 12113 3900
rect 12045 3882 12125 3898
rect 12045 3860 12064 3882
rect 12079 3866 12109 3882
rect 12137 3876 12143 3950
rect 12146 3876 12165 4020
rect 12180 3876 12186 4020
rect 12195 3950 12208 4020
rect 12260 4016 12282 4020
rect 12253 3994 12282 4008
rect 12335 3994 12351 4008
rect 12389 4004 12395 4006
rect 12402 4004 12510 4020
rect 12517 4004 12523 4006
rect 12531 4004 12546 4020
rect 12612 4014 12631 4017
rect 12253 3992 12351 3994
rect 12378 3992 12546 4004
rect 12561 3994 12577 4008
rect 12612 3995 12634 4014
rect 12644 4008 12660 4009
rect 12643 4006 12660 4008
rect 12644 4001 12660 4006
rect 12634 3994 12640 3995
rect 12643 3994 12672 4001
rect 12561 3993 12672 3994
rect 12561 3992 12678 3993
rect 12237 3984 12288 3992
rect 12335 3984 12369 3992
rect 12237 3972 12262 3984
rect 12269 3972 12288 3984
rect 12342 3982 12369 3984
rect 12378 3982 12599 3992
rect 12634 3989 12640 3992
rect 12342 3978 12599 3982
rect 12237 3964 12288 3972
rect 12335 3964 12599 3978
rect 12643 3984 12678 3992
rect 12189 3916 12208 3950
rect 12253 3956 12282 3964
rect 12253 3950 12270 3956
rect 12253 3948 12287 3950
rect 12335 3948 12351 3964
rect 12352 3954 12560 3964
rect 12561 3954 12577 3964
rect 12625 3960 12640 3975
rect 12643 3972 12644 3984
rect 12651 3972 12678 3984
rect 12643 3964 12678 3972
rect 12643 3963 12672 3964
rect 12363 3950 12577 3954
rect 12378 3948 12577 3950
rect 12612 3950 12625 3960
rect 12643 3950 12660 3963
rect 12612 3948 12660 3950
rect 12254 3944 12287 3948
rect 12250 3942 12287 3944
rect 12250 3941 12317 3942
rect 12250 3936 12281 3941
rect 12287 3936 12317 3941
rect 12250 3932 12317 3936
rect 12223 3929 12317 3932
rect 12223 3922 12272 3929
rect 12223 3916 12253 3922
rect 12272 3917 12277 3922
rect 12189 3900 12269 3916
rect 12281 3908 12317 3929
rect 12378 3924 12567 3948
rect 12612 3947 12659 3948
rect 12625 3942 12659 3947
rect 12393 3921 12567 3924
rect 12386 3918 12567 3921
rect 12595 3941 12659 3942
rect 12189 3898 12208 3900
rect 12223 3898 12257 3900
rect 12189 3882 12269 3898
rect 12189 3876 12208 3882
rect 11905 3850 12008 3860
rect 11859 3848 12008 3850
rect 12029 3848 12064 3860
rect 11698 3846 11860 3848
rect 11710 3826 11729 3846
rect 11744 3844 11774 3846
rect 11593 3818 11634 3826
rect 11716 3822 11729 3826
rect 11781 3830 11860 3846
rect 11892 3846 12064 3848
rect 11892 3830 11971 3846
rect 11978 3844 12008 3846
rect 11556 3808 11585 3818
rect 11599 3808 11628 3818
rect 11643 3808 11673 3822
rect 11716 3808 11759 3822
rect 11781 3818 11971 3830
rect 12036 3826 12042 3846
rect 11766 3808 11796 3818
rect 11797 3808 11955 3818
rect 11959 3808 11989 3818
rect 11993 3808 12023 3822
rect 12051 3808 12064 3846
rect 12136 3860 12165 3876
rect 12179 3860 12208 3876
rect 12223 3866 12253 3882
rect 12281 3860 12287 3908
rect 12290 3902 12309 3908
rect 12324 3902 12354 3910
rect 12290 3894 12354 3902
rect 12290 3878 12370 3894
rect 12386 3887 12448 3918
rect 12464 3887 12526 3918
rect 12595 3916 12644 3941
rect 12659 3916 12689 3932
rect 12558 3902 12588 3910
rect 12595 3908 12705 3916
rect 12558 3894 12603 3902
rect 12290 3876 12309 3878
rect 12324 3876 12370 3878
rect 12290 3860 12370 3876
rect 12397 3874 12432 3887
rect 12473 3884 12510 3887
rect 12473 3882 12515 3884
rect 12402 3871 12432 3874
rect 12411 3867 12418 3871
rect 12418 3866 12419 3867
rect 12377 3860 12387 3866
rect 12136 3852 12171 3860
rect 12136 3826 12137 3852
rect 12144 3826 12171 3852
rect 12079 3808 12109 3822
rect 12136 3818 12171 3826
rect 12173 3852 12214 3860
rect 12173 3826 12188 3852
rect 12195 3826 12214 3852
rect 12278 3848 12309 3860
rect 12324 3848 12427 3860
rect 12439 3850 12465 3876
rect 12480 3871 12510 3882
rect 12542 3878 12604 3894
rect 12542 3876 12588 3878
rect 12542 3860 12604 3876
rect 12616 3860 12622 3908
rect 12625 3900 12705 3908
rect 12625 3898 12644 3900
rect 12659 3898 12693 3900
rect 12625 3882 12705 3898
rect 12625 3860 12644 3882
rect 12659 3866 12689 3882
rect 12717 3876 12723 3950
rect 12726 3876 12745 4020
rect 12760 3876 12766 4020
rect 12775 3950 12788 4020
rect 12840 4016 12862 4020
rect 12833 3994 12862 4008
rect 12915 3994 12931 4008
rect 12969 4004 12975 4006
rect 12982 4004 13090 4020
rect 13097 4004 13103 4006
rect 13111 4004 13126 4020
rect 13192 4014 13211 4017
rect 12833 3992 12931 3994
rect 12958 3992 13126 4004
rect 13141 3994 13157 4008
rect 13192 3995 13214 4014
rect 13224 4008 13240 4009
rect 13223 4006 13240 4008
rect 13224 4001 13240 4006
rect 13214 3994 13220 3995
rect 13223 3994 13252 4001
rect 13141 3993 13252 3994
rect 13141 3992 13258 3993
rect 12817 3984 12868 3992
rect 12915 3984 12949 3992
rect 12817 3972 12842 3984
rect 12849 3972 12868 3984
rect 12922 3982 12949 3984
rect 12958 3982 13179 3992
rect 13214 3989 13220 3992
rect 12922 3978 13179 3982
rect 12817 3964 12868 3972
rect 12915 3964 13179 3978
rect 13223 3984 13258 3992
rect 12769 3916 12788 3950
rect 12833 3956 12862 3964
rect 12833 3950 12850 3956
rect 12833 3948 12867 3950
rect 12915 3948 12931 3964
rect 12932 3954 13140 3964
rect 13141 3954 13157 3964
rect 13205 3960 13220 3975
rect 13223 3972 13224 3984
rect 13231 3972 13258 3984
rect 13223 3964 13258 3972
rect 13223 3963 13252 3964
rect 12943 3950 13157 3954
rect 12958 3948 13157 3950
rect 13192 3950 13205 3960
rect 13223 3950 13240 3963
rect 13192 3948 13240 3950
rect 12834 3944 12867 3948
rect 12830 3942 12867 3944
rect 12830 3941 12897 3942
rect 12830 3936 12861 3941
rect 12867 3936 12897 3941
rect 12830 3932 12897 3936
rect 12803 3929 12897 3932
rect 12803 3922 12852 3929
rect 12803 3916 12833 3922
rect 12852 3917 12857 3922
rect 12769 3900 12849 3916
rect 12861 3908 12897 3929
rect 12958 3924 13147 3948
rect 13192 3947 13239 3948
rect 13205 3942 13239 3947
rect 12973 3921 13147 3924
rect 12966 3918 13147 3921
rect 13175 3941 13239 3942
rect 12769 3898 12788 3900
rect 12803 3898 12837 3900
rect 12769 3882 12849 3898
rect 12769 3876 12788 3882
rect 12485 3850 12588 3860
rect 12439 3848 12588 3850
rect 12609 3848 12644 3860
rect 12278 3846 12440 3848
rect 12290 3826 12309 3846
rect 12324 3844 12354 3846
rect 12173 3818 12214 3826
rect 12296 3822 12309 3826
rect 12361 3830 12440 3846
rect 12472 3846 12644 3848
rect 12472 3830 12551 3846
rect 12558 3844 12588 3846
rect 12136 3808 12165 3818
rect 12179 3808 12208 3818
rect 12223 3808 12253 3822
rect 12296 3808 12339 3822
rect 12361 3818 12551 3830
rect 12616 3826 12622 3846
rect 12346 3808 12376 3818
rect 12377 3808 12535 3818
rect 12539 3808 12569 3818
rect 12573 3808 12603 3822
rect 12631 3808 12644 3846
rect 12716 3860 12745 3876
rect 12759 3860 12788 3876
rect 12803 3866 12833 3882
rect 12861 3860 12867 3908
rect 12870 3902 12889 3908
rect 12904 3902 12934 3910
rect 12870 3894 12934 3902
rect 12870 3878 12950 3894
rect 12966 3887 13028 3918
rect 13044 3887 13106 3918
rect 13175 3916 13224 3941
rect 13239 3916 13269 3932
rect 13138 3902 13168 3910
rect 13175 3908 13285 3916
rect 13138 3894 13183 3902
rect 12870 3876 12889 3878
rect 12904 3876 12950 3878
rect 12870 3860 12950 3876
rect 12977 3874 13012 3887
rect 13053 3884 13090 3887
rect 13053 3882 13095 3884
rect 12982 3871 13012 3874
rect 12991 3867 12998 3871
rect 12998 3866 12999 3867
rect 12957 3860 12967 3866
rect 12716 3852 12751 3860
rect 12716 3826 12717 3852
rect 12724 3826 12751 3852
rect 12659 3808 12689 3822
rect 12716 3818 12751 3826
rect 12753 3852 12794 3860
rect 12753 3826 12768 3852
rect 12775 3826 12794 3852
rect 12858 3848 12889 3860
rect 12904 3848 13007 3860
rect 13019 3850 13045 3876
rect 13060 3871 13090 3882
rect 13122 3878 13184 3894
rect 13122 3876 13168 3878
rect 13122 3860 13184 3876
rect 13196 3860 13202 3908
rect 13205 3900 13285 3908
rect 13205 3898 13224 3900
rect 13239 3898 13273 3900
rect 13205 3882 13285 3898
rect 13205 3860 13224 3882
rect 13239 3866 13269 3882
rect 13297 3876 13303 3950
rect 13306 3876 13325 4020
rect 13340 3876 13346 4020
rect 13355 3950 13368 4020
rect 13420 4016 13442 4020
rect 13413 3994 13442 4008
rect 13495 3994 13511 4008
rect 13549 4004 13555 4006
rect 13562 4004 13670 4020
rect 13677 4004 13683 4006
rect 13691 4004 13706 4020
rect 13772 4014 13791 4017
rect 13413 3992 13511 3994
rect 13538 3992 13706 4004
rect 13721 3994 13737 4008
rect 13772 3995 13794 4014
rect 13804 4008 13820 4009
rect 13803 4006 13820 4008
rect 13804 4001 13820 4006
rect 13794 3994 13800 3995
rect 13803 3994 13832 4001
rect 13721 3993 13832 3994
rect 13721 3992 13838 3993
rect 13397 3984 13448 3992
rect 13495 3984 13529 3992
rect 13397 3972 13422 3984
rect 13429 3972 13448 3984
rect 13502 3982 13529 3984
rect 13538 3982 13759 3992
rect 13794 3989 13800 3992
rect 13502 3978 13759 3982
rect 13397 3964 13448 3972
rect 13495 3964 13759 3978
rect 13803 3984 13838 3992
rect 13349 3916 13368 3950
rect 13413 3956 13442 3964
rect 13413 3950 13430 3956
rect 13413 3948 13447 3950
rect 13495 3948 13511 3964
rect 13512 3954 13720 3964
rect 13721 3954 13737 3964
rect 13785 3960 13800 3975
rect 13803 3972 13804 3984
rect 13811 3972 13838 3984
rect 13803 3964 13838 3972
rect 13803 3963 13832 3964
rect 13523 3950 13737 3954
rect 13538 3948 13737 3950
rect 13772 3950 13785 3960
rect 13803 3950 13820 3963
rect 13772 3948 13820 3950
rect 13414 3944 13447 3948
rect 13410 3942 13447 3944
rect 13410 3941 13477 3942
rect 13410 3936 13441 3941
rect 13447 3936 13477 3941
rect 13410 3932 13477 3936
rect 13383 3929 13477 3932
rect 13383 3922 13432 3929
rect 13383 3916 13413 3922
rect 13432 3917 13437 3922
rect 13349 3900 13429 3916
rect 13441 3908 13477 3929
rect 13538 3924 13727 3948
rect 13772 3947 13819 3948
rect 13785 3942 13819 3947
rect 13553 3921 13727 3924
rect 13546 3918 13727 3921
rect 13755 3941 13819 3942
rect 13349 3898 13368 3900
rect 13383 3898 13417 3900
rect 13349 3882 13429 3898
rect 13349 3876 13368 3882
rect 13065 3850 13168 3860
rect 13019 3848 13168 3850
rect 13189 3848 13224 3860
rect 12858 3846 13020 3848
rect 12870 3826 12889 3846
rect 12904 3844 12934 3846
rect 12753 3818 12794 3826
rect 12876 3822 12889 3826
rect 12941 3830 13020 3846
rect 13052 3846 13224 3848
rect 13052 3830 13131 3846
rect 13138 3844 13168 3846
rect 12716 3808 12745 3818
rect 12759 3808 12788 3818
rect 12803 3808 12833 3822
rect 12876 3808 12919 3822
rect 12941 3818 13131 3830
rect 13196 3826 13202 3846
rect 12926 3808 12956 3818
rect 12957 3808 13115 3818
rect 13119 3808 13149 3818
rect 13153 3808 13183 3822
rect 13211 3808 13224 3846
rect 13296 3860 13325 3876
rect 13339 3860 13368 3876
rect 13383 3866 13413 3882
rect 13441 3860 13447 3908
rect 13450 3902 13469 3908
rect 13484 3902 13514 3910
rect 13450 3894 13514 3902
rect 13450 3878 13530 3894
rect 13546 3887 13608 3918
rect 13624 3887 13686 3918
rect 13755 3916 13804 3941
rect 13819 3916 13849 3932
rect 13718 3902 13748 3910
rect 13755 3908 13865 3916
rect 13718 3894 13763 3902
rect 13450 3876 13469 3878
rect 13484 3876 13530 3878
rect 13450 3860 13530 3876
rect 13557 3874 13592 3887
rect 13633 3884 13670 3887
rect 13633 3882 13675 3884
rect 13562 3871 13592 3874
rect 13571 3867 13578 3871
rect 13578 3866 13579 3867
rect 13537 3860 13547 3866
rect 13296 3852 13331 3860
rect 13296 3826 13297 3852
rect 13304 3826 13331 3852
rect 13239 3808 13269 3822
rect 13296 3818 13331 3826
rect 13333 3852 13374 3860
rect 13333 3826 13348 3852
rect 13355 3826 13374 3852
rect 13438 3848 13469 3860
rect 13484 3848 13587 3860
rect 13599 3850 13625 3876
rect 13640 3871 13670 3882
rect 13702 3878 13764 3894
rect 13702 3876 13748 3878
rect 13702 3860 13764 3876
rect 13776 3860 13782 3908
rect 13785 3900 13865 3908
rect 13785 3898 13804 3900
rect 13819 3898 13853 3900
rect 13785 3882 13865 3898
rect 13785 3860 13804 3882
rect 13819 3866 13849 3882
rect 13877 3876 13883 3950
rect 13886 3876 13905 4020
rect 13920 3876 13926 4020
rect 13935 3950 13948 4020
rect 14000 4016 14022 4020
rect 13993 3994 14022 4008
rect 14075 3994 14091 4008
rect 14129 4004 14135 4006
rect 14142 4004 14250 4020
rect 14257 4004 14263 4006
rect 14271 4004 14286 4020
rect 14352 4014 14371 4017
rect 13993 3992 14091 3994
rect 14118 3992 14286 4004
rect 14301 3994 14317 4008
rect 14352 3995 14374 4014
rect 14384 4008 14400 4009
rect 14383 4006 14400 4008
rect 14384 4001 14400 4006
rect 14374 3994 14380 3995
rect 14383 3994 14412 4001
rect 14301 3993 14412 3994
rect 14301 3992 14418 3993
rect 13977 3984 14028 3992
rect 14075 3984 14109 3992
rect 13977 3972 14002 3984
rect 14009 3972 14028 3984
rect 14082 3982 14109 3984
rect 14118 3982 14339 3992
rect 14374 3989 14380 3992
rect 14082 3978 14339 3982
rect 13977 3964 14028 3972
rect 14075 3964 14339 3978
rect 14383 3984 14418 3992
rect 13929 3916 13948 3950
rect 13993 3956 14022 3964
rect 13993 3950 14010 3956
rect 13993 3948 14027 3950
rect 14075 3948 14091 3964
rect 14092 3954 14300 3964
rect 14301 3954 14317 3964
rect 14365 3960 14380 3975
rect 14383 3972 14384 3984
rect 14391 3972 14418 3984
rect 14383 3964 14418 3972
rect 14383 3963 14412 3964
rect 14103 3950 14317 3954
rect 14118 3948 14317 3950
rect 14352 3950 14365 3960
rect 14383 3950 14400 3963
rect 14352 3948 14400 3950
rect 13994 3944 14027 3948
rect 13990 3942 14027 3944
rect 13990 3941 14057 3942
rect 13990 3936 14021 3941
rect 14027 3936 14057 3941
rect 13990 3932 14057 3936
rect 13963 3929 14057 3932
rect 13963 3922 14012 3929
rect 13963 3916 13993 3922
rect 14012 3917 14017 3922
rect 13929 3900 14009 3916
rect 14021 3908 14057 3929
rect 14118 3924 14307 3948
rect 14352 3947 14399 3948
rect 14365 3942 14399 3947
rect 14133 3921 14307 3924
rect 14126 3918 14307 3921
rect 14335 3941 14399 3942
rect 13929 3898 13948 3900
rect 13963 3898 13997 3900
rect 13929 3882 14009 3898
rect 13929 3876 13948 3882
rect 13645 3850 13748 3860
rect 13599 3848 13748 3850
rect 13769 3848 13804 3860
rect 13438 3846 13600 3848
rect 13450 3826 13469 3846
rect 13484 3844 13514 3846
rect 13333 3818 13374 3826
rect 13456 3822 13469 3826
rect 13521 3830 13600 3846
rect 13632 3846 13804 3848
rect 13632 3830 13711 3846
rect 13718 3844 13748 3846
rect 13296 3808 13325 3818
rect 13339 3808 13368 3818
rect 13383 3808 13413 3822
rect 13456 3808 13499 3822
rect 13521 3818 13711 3830
rect 13776 3826 13782 3846
rect 13506 3808 13536 3818
rect 13537 3808 13695 3818
rect 13699 3808 13729 3818
rect 13733 3808 13763 3822
rect 13791 3808 13804 3846
rect 13876 3860 13905 3876
rect 13919 3860 13948 3876
rect 13963 3866 13993 3882
rect 14021 3860 14027 3908
rect 14030 3902 14049 3908
rect 14064 3902 14094 3910
rect 14030 3894 14094 3902
rect 14030 3878 14110 3894
rect 14126 3887 14188 3918
rect 14204 3887 14266 3918
rect 14335 3916 14384 3941
rect 14399 3916 14429 3932
rect 14298 3902 14328 3910
rect 14335 3908 14445 3916
rect 14298 3894 14343 3902
rect 14030 3876 14049 3878
rect 14064 3876 14110 3878
rect 14030 3860 14110 3876
rect 14137 3874 14172 3887
rect 14213 3884 14250 3887
rect 14213 3882 14255 3884
rect 14142 3871 14172 3874
rect 14151 3867 14158 3871
rect 14158 3866 14159 3867
rect 14117 3860 14127 3866
rect 13876 3852 13911 3860
rect 13876 3826 13877 3852
rect 13884 3826 13911 3852
rect 13819 3808 13849 3822
rect 13876 3818 13911 3826
rect 13913 3852 13954 3860
rect 13913 3826 13928 3852
rect 13935 3826 13954 3852
rect 14018 3848 14049 3860
rect 14064 3848 14167 3860
rect 14179 3850 14205 3876
rect 14220 3871 14250 3882
rect 14282 3878 14344 3894
rect 14282 3876 14328 3878
rect 14282 3860 14344 3876
rect 14356 3860 14362 3908
rect 14365 3900 14445 3908
rect 14365 3898 14384 3900
rect 14399 3898 14433 3900
rect 14365 3882 14445 3898
rect 14365 3860 14384 3882
rect 14399 3866 14429 3882
rect 14457 3876 14463 3950
rect 14466 3876 14485 4020
rect 14500 3876 14506 4020
rect 14515 3950 14528 4020
rect 14580 4016 14602 4020
rect 14573 3994 14602 4008
rect 14655 3994 14671 4008
rect 14709 4004 14715 4006
rect 14722 4004 14830 4020
rect 14837 4004 14843 4006
rect 14851 4004 14866 4020
rect 14932 4014 14951 4017
rect 14573 3992 14671 3994
rect 14698 3992 14866 4004
rect 14881 3994 14897 4008
rect 14932 3995 14954 4014
rect 14964 4008 14980 4009
rect 14963 4006 14980 4008
rect 14964 4001 14980 4006
rect 14954 3994 14960 3995
rect 14963 3994 14992 4001
rect 14881 3993 14992 3994
rect 14881 3992 14998 3993
rect 14557 3984 14608 3992
rect 14655 3984 14689 3992
rect 14557 3972 14582 3984
rect 14589 3972 14608 3984
rect 14662 3982 14689 3984
rect 14698 3982 14919 3992
rect 14954 3989 14960 3992
rect 14662 3978 14919 3982
rect 14557 3964 14608 3972
rect 14655 3964 14919 3978
rect 14963 3984 14998 3992
rect 14509 3916 14528 3950
rect 14573 3956 14602 3964
rect 14573 3950 14590 3956
rect 14573 3948 14607 3950
rect 14655 3948 14671 3964
rect 14672 3954 14880 3964
rect 14881 3954 14897 3964
rect 14945 3960 14960 3975
rect 14963 3972 14964 3984
rect 14971 3972 14998 3984
rect 14963 3964 14998 3972
rect 14963 3963 14992 3964
rect 14683 3950 14897 3954
rect 14698 3948 14897 3950
rect 14932 3950 14945 3960
rect 14963 3950 14980 3963
rect 14932 3948 14980 3950
rect 14574 3944 14607 3948
rect 14570 3942 14607 3944
rect 14570 3941 14637 3942
rect 14570 3936 14601 3941
rect 14607 3936 14637 3941
rect 14570 3932 14637 3936
rect 14543 3929 14637 3932
rect 14543 3922 14592 3929
rect 14543 3916 14573 3922
rect 14592 3917 14597 3922
rect 14509 3900 14589 3916
rect 14601 3908 14637 3929
rect 14698 3924 14887 3948
rect 14932 3947 14979 3948
rect 14945 3942 14979 3947
rect 14713 3921 14887 3924
rect 14706 3918 14887 3921
rect 14915 3941 14979 3942
rect 14509 3898 14528 3900
rect 14543 3898 14577 3900
rect 14509 3882 14589 3898
rect 14509 3876 14528 3882
rect 14225 3850 14328 3860
rect 14179 3848 14328 3850
rect 14349 3848 14384 3860
rect 14018 3846 14180 3848
rect 14030 3826 14049 3846
rect 14064 3844 14094 3846
rect 13913 3818 13954 3826
rect 14036 3822 14049 3826
rect 14101 3830 14180 3846
rect 14212 3846 14384 3848
rect 14212 3830 14291 3846
rect 14298 3844 14328 3846
rect 13876 3808 13905 3818
rect 13919 3808 13948 3818
rect 13963 3808 13993 3822
rect 14036 3808 14079 3822
rect 14101 3818 14291 3830
rect 14356 3826 14362 3846
rect 14086 3808 14116 3818
rect 14117 3808 14275 3818
rect 14279 3808 14309 3818
rect 14313 3808 14343 3822
rect 14371 3808 14384 3846
rect 14456 3860 14485 3876
rect 14499 3860 14528 3876
rect 14543 3866 14573 3882
rect 14601 3860 14607 3908
rect 14610 3902 14629 3908
rect 14644 3902 14674 3910
rect 14610 3894 14674 3902
rect 14610 3878 14690 3894
rect 14706 3887 14768 3918
rect 14784 3887 14846 3918
rect 14915 3916 14964 3941
rect 14979 3916 15009 3932
rect 14878 3902 14908 3910
rect 14915 3908 15025 3916
rect 14878 3894 14923 3902
rect 14610 3876 14629 3878
rect 14644 3876 14690 3878
rect 14610 3860 14690 3876
rect 14717 3874 14752 3887
rect 14793 3884 14830 3887
rect 14793 3882 14835 3884
rect 14722 3871 14752 3874
rect 14731 3867 14738 3871
rect 14738 3866 14739 3867
rect 14697 3860 14707 3866
rect 14456 3852 14491 3860
rect 14456 3826 14457 3852
rect 14464 3826 14491 3852
rect 14399 3808 14429 3822
rect 14456 3818 14491 3826
rect 14493 3852 14534 3860
rect 14493 3826 14508 3852
rect 14515 3826 14534 3852
rect 14598 3848 14629 3860
rect 14644 3848 14747 3860
rect 14759 3850 14785 3876
rect 14800 3871 14830 3882
rect 14862 3878 14924 3894
rect 14862 3876 14908 3878
rect 14862 3860 14924 3876
rect 14936 3860 14942 3908
rect 14945 3900 15025 3908
rect 14945 3898 14964 3900
rect 14979 3898 15013 3900
rect 14945 3882 15025 3898
rect 14945 3860 14964 3882
rect 14979 3866 15009 3882
rect 15037 3876 15043 3950
rect 15046 3876 15065 4020
rect 15080 3876 15086 4020
rect 15095 3950 15108 4020
rect 15160 4016 15182 4020
rect 15153 3994 15182 4008
rect 15235 3994 15251 4008
rect 15289 4004 15295 4006
rect 15302 4004 15410 4020
rect 15417 4004 15423 4006
rect 15431 4004 15446 4020
rect 15512 4014 15531 4017
rect 15153 3992 15251 3994
rect 15278 3992 15446 4004
rect 15461 3994 15477 4008
rect 15512 3995 15534 4014
rect 15544 4008 15560 4009
rect 15543 4006 15560 4008
rect 15544 4001 15560 4006
rect 15534 3994 15540 3995
rect 15543 3994 15572 4001
rect 15461 3993 15572 3994
rect 15461 3992 15578 3993
rect 15137 3984 15188 3992
rect 15235 3984 15269 3992
rect 15137 3972 15162 3984
rect 15169 3972 15188 3984
rect 15242 3982 15269 3984
rect 15278 3982 15499 3992
rect 15534 3989 15540 3992
rect 15242 3978 15499 3982
rect 15137 3964 15188 3972
rect 15235 3964 15499 3978
rect 15543 3984 15578 3992
rect 15089 3916 15108 3950
rect 15153 3956 15182 3964
rect 15153 3950 15170 3956
rect 15153 3948 15187 3950
rect 15235 3948 15251 3964
rect 15252 3954 15460 3964
rect 15461 3954 15477 3964
rect 15525 3960 15540 3975
rect 15543 3972 15544 3984
rect 15551 3972 15578 3984
rect 15543 3964 15578 3972
rect 15543 3963 15572 3964
rect 15263 3950 15477 3954
rect 15278 3948 15477 3950
rect 15512 3950 15525 3960
rect 15543 3950 15560 3963
rect 15512 3948 15560 3950
rect 15154 3944 15187 3948
rect 15150 3942 15187 3944
rect 15150 3941 15217 3942
rect 15150 3936 15181 3941
rect 15187 3936 15217 3941
rect 15150 3932 15217 3936
rect 15123 3929 15217 3932
rect 15123 3922 15172 3929
rect 15123 3916 15153 3922
rect 15172 3917 15177 3922
rect 15089 3900 15169 3916
rect 15181 3908 15217 3929
rect 15278 3924 15467 3948
rect 15512 3947 15559 3948
rect 15525 3942 15559 3947
rect 15293 3921 15467 3924
rect 15286 3918 15467 3921
rect 15495 3941 15559 3942
rect 15089 3898 15108 3900
rect 15123 3898 15157 3900
rect 15089 3882 15169 3898
rect 15089 3876 15108 3882
rect 14805 3850 14908 3860
rect 14759 3848 14908 3850
rect 14929 3848 14964 3860
rect 14598 3846 14760 3848
rect 14610 3826 14629 3846
rect 14644 3844 14674 3846
rect 14493 3818 14534 3826
rect 14616 3822 14629 3826
rect 14681 3830 14760 3846
rect 14792 3846 14964 3848
rect 14792 3830 14871 3846
rect 14878 3844 14908 3846
rect 14456 3808 14485 3818
rect 14499 3808 14528 3818
rect 14543 3808 14573 3822
rect 14616 3808 14659 3822
rect 14681 3818 14871 3830
rect 14936 3826 14942 3846
rect 14666 3808 14696 3818
rect 14697 3808 14855 3818
rect 14859 3808 14889 3818
rect 14893 3808 14923 3822
rect 14951 3808 14964 3846
rect 15036 3860 15065 3876
rect 15079 3860 15108 3876
rect 15123 3866 15153 3882
rect 15181 3860 15187 3908
rect 15190 3902 15209 3908
rect 15224 3902 15254 3910
rect 15190 3894 15254 3902
rect 15190 3878 15270 3894
rect 15286 3887 15348 3918
rect 15364 3887 15426 3918
rect 15495 3916 15544 3941
rect 15559 3916 15589 3932
rect 15458 3902 15488 3910
rect 15495 3908 15605 3916
rect 15458 3894 15503 3902
rect 15190 3876 15209 3878
rect 15224 3876 15270 3878
rect 15190 3860 15270 3876
rect 15297 3874 15332 3887
rect 15373 3884 15410 3887
rect 15373 3882 15415 3884
rect 15302 3871 15332 3874
rect 15311 3867 15318 3871
rect 15318 3866 15319 3867
rect 15277 3860 15287 3866
rect 15036 3852 15071 3860
rect 15036 3826 15037 3852
rect 15044 3826 15071 3852
rect 14979 3808 15009 3822
rect 15036 3818 15071 3826
rect 15073 3852 15114 3860
rect 15073 3826 15088 3852
rect 15095 3826 15114 3852
rect 15178 3848 15209 3860
rect 15224 3848 15327 3860
rect 15339 3850 15365 3876
rect 15380 3871 15410 3882
rect 15442 3878 15504 3894
rect 15442 3876 15488 3878
rect 15442 3860 15504 3876
rect 15516 3860 15522 3908
rect 15525 3900 15605 3908
rect 15525 3898 15544 3900
rect 15559 3898 15593 3900
rect 15525 3882 15605 3898
rect 15525 3860 15544 3882
rect 15559 3866 15589 3882
rect 15617 3876 15623 3950
rect 15626 3876 15645 4020
rect 15660 3876 15666 4020
rect 15675 3950 15688 4020
rect 15740 4016 15762 4020
rect 15733 3994 15762 4008
rect 15815 3994 15831 4008
rect 15869 4004 15875 4006
rect 15882 4004 15990 4020
rect 15997 4004 16003 4006
rect 16011 4004 16026 4020
rect 16092 4014 16111 4017
rect 15733 3992 15831 3994
rect 15858 3992 16026 4004
rect 16041 3994 16057 4008
rect 16092 3995 16114 4014
rect 16124 4008 16140 4009
rect 16123 4006 16140 4008
rect 16124 4001 16140 4006
rect 16114 3994 16120 3995
rect 16123 3994 16152 4001
rect 16041 3993 16152 3994
rect 16041 3992 16158 3993
rect 15717 3984 15768 3992
rect 15815 3984 15849 3992
rect 15717 3972 15742 3984
rect 15749 3972 15768 3984
rect 15822 3982 15849 3984
rect 15858 3982 16079 3992
rect 16114 3989 16120 3992
rect 15822 3978 16079 3982
rect 15717 3964 15768 3972
rect 15815 3964 16079 3978
rect 16123 3984 16158 3992
rect 15669 3916 15688 3950
rect 15733 3956 15762 3964
rect 15733 3950 15750 3956
rect 15733 3948 15767 3950
rect 15815 3948 15831 3964
rect 15832 3954 16040 3964
rect 16041 3954 16057 3964
rect 16105 3960 16120 3975
rect 16123 3972 16124 3984
rect 16131 3972 16158 3984
rect 16123 3964 16158 3972
rect 16123 3963 16152 3964
rect 15843 3950 16057 3954
rect 15858 3948 16057 3950
rect 16092 3950 16105 3960
rect 16123 3950 16140 3963
rect 16092 3948 16140 3950
rect 15734 3944 15767 3948
rect 15730 3942 15767 3944
rect 15730 3941 15797 3942
rect 15730 3936 15761 3941
rect 15767 3936 15797 3941
rect 15730 3932 15797 3936
rect 15703 3929 15797 3932
rect 15703 3922 15752 3929
rect 15703 3916 15733 3922
rect 15752 3917 15757 3922
rect 15669 3900 15749 3916
rect 15761 3908 15797 3929
rect 15858 3924 16047 3948
rect 16092 3947 16139 3948
rect 16105 3942 16139 3947
rect 15873 3921 16047 3924
rect 15866 3918 16047 3921
rect 16075 3941 16139 3942
rect 15669 3898 15688 3900
rect 15703 3898 15737 3900
rect 15669 3882 15749 3898
rect 15669 3876 15688 3882
rect 15385 3850 15488 3860
rect 15339 3848 15488 3850
rect 15509 3848 15544 3860
rect 15178 3846 15340 3848
rect 15190 3826 15209 3846
rect 15224 3844 15254 3846
rect 15073 3818 15114 3826
rect 15196 3822 15209 3826
rect 15261 3830 15340 3846
rect 15372 3846 15544 3848
rect 15372 3830 15451 3846
rect 15458 3844 15488 3846
rect 15036 3808 15065 3818
rect 15079 3808 15108 3818
rect 15123 3808 15153 3822
rect 15196 3808 15239 3822
rect 15261 3818 15451 3830
rect 15516 3826 15522 3846
rect 15246 3808 15276 3818
rect 15277 3808 15435 3818
rect 15439 3808 15469 3818
rect 15473 3808 15503 3822
rect 15531 3808 15544 3846
rect 15616 3860 15645 3876
rect 15659 3860 15688 3876
rect 15703 3866 15733 3882
rect 15761 3860 15767 3908
rect 15770 3902 15789 3908
rect 15804 3902 15834 3910
rect 15770 3894 15834 3902
rect 15770 3878 15850 3894
rect 15866 3887 15928 3918
rect 15944 3887 16006 3918
rect 16075 3916 16124 3941
rect 16139 3916 16169 3932
rect 16038 3902 16068 3910
rect 16075 3908 16185 3916
rect 16038 3894 16083 3902
rect 15770 3876 15789 3878
rect 15804 3876 15850 3878
rect 15770 3860 15850 3876
rect 15877 3874 15912 3887
rect 15953 3884 15990 3887
rect 15953 3882 15995 3884
rect 15882 3871 15912 3874
rect 15891 3867 15898 3871
rect 15898 3866 15899 3867
rect 15857 3860 15867 3866
rect 15616 3852 15651 3860
rect 15616 3826 15617 3852
rect 15624 3826 15651 3852
rect 15559 3808 15589 3822
rect 15616 3818 15651 3826
rect 15653 3852 15694 3860
rect 15653 3826 15668 3852
rect 15675 3826 15694 3852
rect 15758 3848 15789 3860
rect 15804 3848 15907 3860
rect 15919 3850 15945 3876
rect 15960 3871 15990 3882
rect 16022 3878 16084 3894
rect 16022 3876 16068 3878
rect 16022 3860 16084 3876
rect 16096 3860 16102 3908
rect 16105 3900 16185 3908
rect 16105 3898 16124 3900
rect 16139 3898 16173 3900
rect 16105 3882 16185 3898
rect 16105 3860 16124 3882
rect 16139 3866 16169 3882
rect 16197 3876 16203 3950
rect 16206 3876 16225 4020
rect 16240 3876 16246 4020
rect 16255 3950 16268 4020
rect 16320 4016 16342 4020
rect 16313 3994 16342 4008
rect 16395 3994 16411 4008
rect 16449 4004 16455 4006
rect 16462 4004 16570 4020
rect 16577 4004 16583 4006
rect 16591 4004 16606 4020
rect 16672 4014 16691 4017
rect 16313 3992 16411 3994
rect 16438 3992 16606 4004
rect 16621 3994 16637 4008
rect 16672 3995 16694 4014
rect 16704 4008 16720 4009
rect 16703 4006 16720 4008
rect 16704 4001 16720 4006
rect 16694 3994 16700 3995
rect 16703 3994 16732 4001
rect 16621 3993 16732 3994
rect 16621 3992 16738 3993
rect 16297 3984 16348 3992
rect 16395 3984 16429 3992
rect 16297 3972 16322 3984
rect 16329 3972 16348 3984
rect 16402 3982 16429 3984
rect 16438 3982 16659 3992
rect 16694 3989 16700 3992
rect 16402 3978 16659 3982
rect 16297 3964 16348 3972
rect 16395 3964 16659 3978
rect 16703 3984 16738 3992
rect 16249 3916 16268 3950
rect 16313 3956 16342 3964
rect 16313 3950 16330 3956
rect 16313 3948 16347 3950
rect 16395 3948 16411 3964
rect 16412 3954 16620 3964
rect 16621 3954 16637 3964
rect 16685 3960 16700 3975
rect 16703 3972 16704 3984
rect 16711 3972 16738 3984
rect 16703 3964 16738 3972
rect 16703 3963 16732 3964
rect 16423 3950 16637 3954
rect 16438 3948 16637 3950
rect 16672 3950 16685 3960
rect 16703 3950 16720 3963
rect 16672 3948 16720 3950
rect 16314 3944 16347 3948
rect 16310 3942 16347 3944
rect 16310 3941 16377 3942
rect 16310 3936 16341 3941
rect 16347 3936 16377 3941
rect 16310 3932 16377 3936
rect 16283 3929 16377 3932
rect 16283 3922 16332 3929
rect 16283 3916 16313 3922
rect 16332 3917 16337 3922
rect 16249 3900 16329 3916
rect 16341 3908 16377 3929
rect 16438 3924 16627 3948
rect 16672 3947 16719 3948
rect 16685 3942 16719 3947
rect 16453 3921 16627 3924
rect 16446 3918 16627 3921
rect 16655 3941 16719 3942
rect 16249 3898 16268 3900
rect 16283 3898 16317 3900
rect 16249 3882 16329 3898
rect 16249 3876 16268 3882
rect 15965 3850 16068 3860
rect 15919 3848 16068 3850
rect 16089 3848 16124 3860
rect 15758 3846 15920 3848
rect 15770 3826 15789 3846
rect 15804 3844 15834 3846
rect 15653 3818 15694 3826
rect 15776 3822 15789 3826
rect 15841 3830 15920 3846
rect 15952 3846 16124 3848
rect 15952 3830 16031 3846
rect 16038 3844 16068 3846
rect 15616 3808 15645 3818
rect 15659 3808 15688 3818
rect 15703 3808 15733 3822
rect 15776 3808 15819 3822
rect 15841 3818 16031 3830
rect 16096 3826 16102 3846
rect 15826 3808 15856 3818
rect 15857 3808 16015 3818
rect 16019 3808 16049 3818
rect 16053 3808 16083 3822
rect 16111 3808 16124 3846
rect 16196 3860 16225 3876
rect 16239 3860 16268 3876
rect 16283 3866 16313 3882
rect 16341 3860 16347 3908
rect 16350 3902 16369 3908
rect 16384 3902 16414 3910
rect 16350 3894 16414 3902
rect 16350 3878 16430 3894
rect 16446 3887 16508 3918
rect 16524 3887 16586 3918
rect 16655 3916 16704 3941
rect 16719 3916 16749 3932
rect 16618 3902 16648 3910
rect 16655 3908 16765 3916
rect 16618 3894 16663 3902
rect 16350 3876 16369 3878
rect 16384 3876 16430 3878
rect 16350 3860 16430 3876
rect 16457 3874 16492 3887
rect 16533 3884 16570 3887
rect 16533 3882 16575 3884
rect 16462 3871 16492 3874
rect 16471 3867 16478 3871
rect 16478 3866 16479 3867
rect 16437 3860 16447 3866
rect 16196 3852 16231 3860
rect 16196 3826 16197 3852
rect 16204 3826 16231 3852
rect 16139 3808 16169 3822
rect 16196 3818 16231 3826
rect 16233 3852 16274 3860
rect 16233 3826 16248 3852
rect 16255 3826 16274 3852
rect 16338 3848 16369 3860
rect 16384 3848 16487 3860
rect 16499 3850 16525 3876
rect 16540 3871 16570 3882
rect 16602 3878 16664 3894
rect 16602 3876 16648 3878
rect 16602 3860 16664 3876
rect 16676 3860 16682 3908
rect 16685 3900 16765 3908
rect 16685 3898 16704 3900
rect 16719 3898 16753 3900
rect 16685 3882 16765 3898
rect 16685 3860 16704 3882
rect 16719 3866 16749 3882
rect 16777 3876 16783 3950
rect 16786 3876 16805 4020
rect 16820 3876 16826 4020
rect 16835 3950 16848 4020
rect 16900 4016 16922 4020
rect 16893 3994 16922 4008
rect 16975 3994 16991 4008
rect 17029 4004 17035 4006
rect 17042 4004 17150 4020
rect 17157 4004 17163 4006
rect 17171 4004 17186 4020
rect 17252 4014 17271 4017
rect 16893 3992 16991 3994
rect 17018 3992 17186 4004
rect 17201 3994 17217 4008
rect 17252 3995 17274 4014
rect 17284 4008 17300 4009
rect 17283 4006 17300 4008
rect 17284 4001 17300 4006
rect 17274 3994 17280 3995
rect 17283 3994 17312 4001
rect 17201 3993 17312 3994
rect 17201 3992 17318 3993
rect 16877 3984 16928 3992
rect 16975 3984 17009 3992
rect 16877 3972 16902 3984
rect 16909 3972 16928 3984
rect 16982 3982 17009 3984
rect 17018 3982 17239 3992
rect 17274 3989 17280 3992
rect 16982 3978 17239 3982
rect 16877 3964 16928 3972
rect 16975 3964 17239 3978
rect 17283 3984 17318 3992
rect 16829 3916 16848 3950
rect 16893 3956 16922 3964
rect 16893 3950 16910 3956
rect 16893 3948 16927 3950
rect 16975 3948 16991 3964
rect 16992 3954 17200 3964
rect 17201 3954 17217 3964
rect 17265 3960 17280 3975
rect 17283 3972 17284 3984
rect 17291 3972 17318 3984
rect 17283 3964 17318 3972
rect 17283 3963 17312 3964
rect 17003 3950 17217 3954
rect 17018 3948 17217 3950
rect 17252 3950 17265 3960
rect 17283 3950 17300 3963
rect 17252 3948 17300 3950
rect 16894 3944 16927 3948
rect 16890 3942 16927 3944
rect 16890 3941 16957 3942
rect 16890 3936 16921 3941
rect 16927 3936 16957 3941
rect 16890 3932 16957 3936
rect 16863 3929 16957 3932
rect 16863 3922 16912 3929
rect 16863 3916 16893 3922
rect 16912 3917 16917 3922
rect 16829 3900 16909 3916
rect 16921 3908 16957 3929
rect 17018 3924 17207 3948
rect 17252 3947 17299 3948
rect 17265 3942 17299 3947
rect 17033 3921 17207 3924
rect 17026 3918 17207 3921
rect 17235 3941 17299 3942
rect 16829 3898 16848 3900
rect 16863 3898 16897 3900
rect 16829 3882 16909 3898
rect 16829 3876 16848 3882
rect 16545 3850 16648 3860
rect 16499 3848 16648 3850
rect 16669 3848 16704 3860
rect 16338 3846 16500 3848
rect 16350 3826 16369 3846
rect 16384 3844 16414 3846
rect 16233 3818 16274 3826
rect 16356 3822 16369 3826
rect 16421 3830 16500 3846
rect 16532 3846 16704 3848
rect 16532 3830 16611 3846
rect 16618 3844 16648 3846
rect 16196 3808 16225 3818
rect 16239 3808 16268 3818
rect 16283 3808 16313 3822
rect 16356 3808 16399 3822
rect 16421 3818 16611 3830
rect 16676 3826 16682 3846
rect 16406 3808 16436 3818
rect 16437 3808 16595 3818
rect 16599 3808 16629 3818
rect 16633 3808 16663 3822
rect 16691 3808 16704 3846
rect 16776 3860 16805 3876
rect 16819 3860 16848 3876
rect 16863 3866 16893 3882
rect 16921 3860 16927 3908
rect 16930 3902 16949 3908
rect 16964 3902 16994 3910
rect 16930 3894 16994 3902
rect 16930 3878 17010 3894
rect 17026 3887 17088 3918
rect 17104 3887 17166 3918
rect 17235 3916 17284 3941
rect 17299 3916 17329 3932
rect 17198 3902 17228 3910
rect 17235 3908 17345 3916
rect 17198 3894 17243 3902
rect 16930 3876 16949 3878
rect 16964 3876 17010 3878
rect 16930 3860 17010 3876
rect 17037 3874 17072 3887
rect 17113 3884 17150 3887
rect 17113 3882 17155 3884
rect 17042 3871 17072 3874
rect 17051 3867 17058 3871
rect 17058 3866 17059 3867
rect 17017 3860 17027 3866
rect 16776 3852 16811 3860
rect 16776 3826 16777 3852
rect 16784 3826 16811 3852
rect 16719 3808 16749 3822
rect 16776 3818 16811 3826
rect 16813 3852 16854 3860
rect 16813 3826 16828 3852
rect 16835 3826 16854 3852
rect 16918 3848 16949 3860
rect 16964 3848 17067 3860
rect 17079 3850 17105 3876
rect 17120 3871 17150 3882
rect 17182 3878 17244 3894
rect 17182 3876 17228 3878
rect 17182 3860 17244 3876
rect 17256 3860 17262 3908
rect 17265 3900 17345 3908
rect 17265 3898 17284 3900
rect 17299 3898 17333 3900
rect 17265 3882 17345 3898
rect 17265 3860 17284 3882
rect 17299 3866 17329 3882
rect 17357 3876 17363 3950
rect 17366 3876 17385 4020
rect 17400 3876 17406 4020
rect 17415 3950 17428 4020
rect 17480 4016 17502 4020
rect 17473 3994 17502 4008
rect 17555 3994 17571 4008
rect 17609 4004 17615 4006
rect 17622 4004 17730 4020
rect 17737 4004 17743 4006
rect 17751 4004 17766 4020
rect 17832 4014 17851 4017
rect 17473 3992 17571 3994
rect 17598 3992 17766 4004
rect 17781 3994 17797 4008
rect 17832 3995 17854 4014
rect 17864 4008 17880 4009
rect 17863 4006 17880 4008
rect 17864 4001 17880 4006
rect 17854 3994 17860 3995
rect 17863 3994 17892 4001
rect 17781 3993 17892 3994
rect 17781 3992 17898 3993
rect 17457 3984 17508 3992
rect 17555 3984 17589 3992
rect 17457 3972 17482 3984
rect 17489 3972 17508 3984
rect 17562 3982 17589 3984
rect 17598 3982 17819 3992
rect 17854 3989 17860 3992
rect 17562 3978 17819 3982
rect 17457 3964 17508 3972
rect 17555 3964 17819 3978
rect 17863 3984 17898 3992
rect 17409 3916 17428 3950
rect 17473 3956 17502 3964
rect 17473 3950 17490 3956
rect 17473 3948 17507 3950
rect 17555 3948 17571 3964
rect 17572 3954 17780 3964
rect 17781 3954 17797 3964
rect 17845 3960 17860 3975
rect 17863 3972 17864 3984
rect 17871 3972 17898 3984
rect 17863 3964 17898 3972
rect 17863 3963 17892 3964
rect 17583 3950 17797 3954
rect 17598 3948 17797 3950
rect 17832 3950 17845 3960
rect 17863 3950 17880 3963
rect 17832 3948 17880 3950
rect 17474 3944 17507 3948
rect 17470 3942 17507 3944
rect 17470 3941 17537 3942
rect 17470 3936 17501 3941
rect 17507 3936 17537 3941
rect 17470 3932 17537 3936
rect 17443 3929 17537 3932
rect 17443 3922 17492 3929
rect 17443 3916 17473 3922
rect 17492 3917 17497 3922
rect 17409 3900 17489 3916
rect 17501 3908 17537 3929
rect 17598 3924 17787 3948
rect 17832 3947 17879 3948
rect 17845 3942 17879 3947
rect 17613 3921 17787 3924
rect 17606 3918 17787 3921
rect 17815 3941 17879 3942
rect 17409 3898 17428 3900
rect 17443 3898 17477 3900
rect 17409 3882 17489 3898
rect 17409 3876 17428 3882
rect 17125 3850 17228 3860
rect 17079 3848 17228 3850
rect 17249 3848 17284 3860
rect 16918 3846 17080 3848
rect 16930 3826 16949 3846
rect 16964 3844 16994 3846
rect 16813 3818 16854 3826
rect 16936 3822 16949 3826
rect 17001 3830 17080 3846
rect 17112 3846 17284 3848
rect 17112 3830 17191 3846
rect 17198 3844 17228 3846
rect 16776 3808 16805 3818
rect 16819 3808 16848 3818
rect 16863 3808 16893 3822
rect 16936 3808 16979 3822
rect 17001 3818 17191 3830
rect 17256 3826 17262 3846
rect 16986 3808 17016 3818
rect 17017 3808 17175 3818
rect 17179 3808 17209 3818
rect 17213 3808 17243 3822
rect 17271 3808 17284 3846
rect 17356 3860 17385 3876
rect 17399 3860 17428 3876
rect 17443 3866 17473 3882
rect 17501 3860 17507 3908
rect 17510 3902 17529 3908
rect 17544 3902 17574 3910
rect 17510 3894 17574 3902
rect 17510 3878 17590 3894
rect 17606 3887 17668 3918
rect 17684 3887 17746 3918
rect 17815 3916 17864 3941
rect 17879 3916 17909 3932
rect 17778 3902 17808 3910
rect 17815 3908 17925 3916
rect 17778 3894 17823 3902
rect 17510 3876 17529 3878
rect 17544 3876 17590 3878
rect 17510 3860 17590 3876
rect 17617 3874 17652 3887
rect 17693 3884 17730 3887
rect 17693 3882 17735 3884
rect 17622 3871 17652 3874
rect 17631 3867 17638 3871
rect 17638 3866 17639 3867
rect 17597 3860 17607 3866
rect 17356 3852 17391 3860
rect 17356 3826 17357 3852
rect 17364 3826 17391 3852
rect 17299 3808 17329 3822
rect 17356 3818 17391 3826
rect 17393 3852 17434 3860
rect 17393 3826 17408 3852
rect 17415 3826 17434 3852
rect 17498 3848 17529 3860
rect 17544 3848 17647 3860
rect 17659 3850 17685 3876
rect 17700 3871 17730 3882
rect 17762 3878 17824 3894
rect 17762 3876 17808 3878
rect 17762 3860 17824 3876
rect 17836 3860 17842 3908
rect 17845 3900 17925 3908
rect 17845 3898 17864 3900
rect 17879 3898 17913 3900
rect 17845 3882 17925 3898
rect 17845 3860 17864 3882
rect 17879 3866 17909 3882
rect 17937 3876 17943 3950
rect 17946 3876 17965 4020
rect 17980 3876 17986 4020
rect 17995 3950 18008 4020
rect 18060 4016 18082 4020
rect 18053 3994 18082 4008
rect 18135 3994 18151 4008
rect 18189 4004 18195 4006
rect 18202 4004 18310 4020
rect 18317 4004 18323 4006
rect 18331 4004 18346 4020
rect 18412 4014 18431 4017
rect 18053 3992 18151 3994
rect 18178 3992 18346 4004
rect 18361 3994 18377 4008
rect 18412 3995 18434 4014
rect 18444 4008 18460 4009
rect 18443 4006 18460 4008
rect 18444 4001 18460 4006
rect 18434 3994 18440 3995
rect 18443 3994 18472 4001
rect 18361 3993 18472 3994
rect 18361 3992 18478 3993
rect 18037 3984 18088 3992
rect 18135 3984 18169 3992
rect 18037 3972 18062 3984
rect 18069 3972 18088 3984
rect 18142 3982 18169 3984
rect 18178 3982 18399 3992
rect 18434 3989 18440 3992
rect 18142 3978 18399 3982
rect 18037 3964 18088 3972
rect 18135 3964 18399 3978
rect 18443 3984 18478 3992
rect 17989 3916 18008 3950
rect 18053 3956 18082 3964
rect 18053 3950 18070 3956
rect 18053 3948 18087 3950
rect 18135 3948 18151 3964
rect 18152 3954 18360 3964
rect 18361 3954 18377 3964
rect 18425 3960 18440 3975
rect 18443 3972 18444 3984
rect 18451 3972 18478 3984
rect 18443 3964 18478 3972
rect 18443 3963 18472 3964
rect 18163 3950 18377 3954
rect 18178 3948 18377 3950
rect 18412 3950 18425 3960
rect 18443 3950 18460 3963
rect 18412 3948 18460 3950
rect 18054 3944 18087 3948
rect 18050 3942 18087 3944
rect 18050 3941 18117 3942
rect 18050 3936 18081 3941
rect 18087 3936 18117 3941
rect 18050 3932 18117 3936
rect 18023 3929 18117 3932
rect 18023 3922 18072 3929
rect 18023 3916 18053 3922
rect 18072 3917 18077 3922
rect 17989 3900 18069 3916
rect 18081 3908 18117 3929
rect 18178 3924 18367 3948
rect 18412 3947 18459 3948
rect 18425 3942 18459 3947
rect 18193 3921 18367 3924
rect 18186 3918 18367 3921
rect 18395 3941 18459 3942
rect 17989 3898 18008 3900
rect 18023 3898 18057 3900
rect 17989 3882 18069 3898
rect 17989 3876 18008 3882
rect 17705 3850 17808 3860
rect 17659 3848 17808 3850
rect 17829 3848 17864 3860
rect 17498 3846 17660 3848
rect 17510 3826 17529 3846
rect 17544 3844 17574 3846
rect 17393 3818 17434 3826
rect 17516 3822 17529 3826
rect 17581 3830 17660 3846
rect 17692 3846 17864 3848
rect 17692 3830 17771 3846
rect 17778 3844 17808 3846
rect 17356 3808 17385 3818
rect 17399 3808 17428 3818
rect 17443 3808 17473 3822
rect 17516 3808 17559 3822
rect 17581 3818 17771 3830
rect 17836 3826 17842 3846
rect 17566 3808 17596 3818
rect 17597 3808 17755 3818
rect 17759 3808 17789 3818
rect 17793 3808 17823 3822
rect 17851 3808 17864 3846
rect 17936 3860 17965 3876
rect 17979 3860 18008 3876
rect 18023 3866 18053 3882
rect 18081 3860 18087 3908
rect 18090 3902 18109 3908
rect 18124 3902 18154 3910
rect 18090 3894 18154 3902
rect 18090 3878 18170 3894
rect 18186 3887 18248 3918
rect 18264 3887 18326 3918
rect 18395 3916 18444 3941
rect 18459 3916 18489 3932
rect 18358 3902 18388 3910
rect 18395 3908 18505 3916
rect 18358 3894 18403 3902
rect 18090 3876 18109 3878
rect 18124 3876 18170 3878
rect 18090 3860 18170 3876
rect 18197 3874 18232 3887
rect 18273 3884 18310 3887
rect 18273 3882 18315 3884
rect 18202 3871 18232 3874
rect 18211 3867 18218 3871
rect 18218 3866 18219 3867
rect 18177 3860 18187 3866
rect 17936 3852 17971 3860
rect 17936 3826 17937 3852
rect 17944 3826 17971 3852
rect 17879 3808 17909 3822
rect 17936 3818 17971 3826
rect 17973 3852 18014 3860
rect 17973 3826 17988 3852
rect 17995 3826 18014 3852
rect 18078 3848 18109 3860
rect 18124 3848 18227 3860
rect 18239 3850 18265 3876
rect 18280 3871 18310 3882
rect 18342 3878 18404 3894
rect 18342 3876 18388 3878
rect 18342 3860 18404 3876
rect 18416 3860 18422 3908
rect 18425 3900 18505 3908
rect 18425 3898 18444 3900
rect 18459 3898 18493 3900
rect 18425 3882 18505 3898
rect 18425 3860 18444 3882
rect 18459 3866 18489 3882
rect 18517 3876 18523 3950
rect 18532 3876 18545 4020
rect 18285 3850 18388 3860
rect 18239 3848 18388 3850
rect 18409 3848 18444 3860
rect 18078 3846 18240 3848
rect 18090 3826 18109 3846
rect 18124 3844 18154 3846
rect 17973 3818 18014 3826
rect 18096 3822 18109 3826
rect 18161 3830 18240 3846
rect 18272 3846 18444 3848
rect 18272 3830 18351 3846
rect 18358 3844 18388 3846
rect 17936 3808 17965 3818
rect 17979 3808 18008 3818
rect 18023 3808 18053 3822
rect 18096 3808 18139 3822
rect 18161 3818 18351 3830
rect 18416 3826 18422 3846
rect 18146 3808 18176 3818
rect 18177 3808 18335 3818
rect 18339 3808 18369 3818
rect 18373 3808 18403 3822
rect 18431 3808 18444 3846
rect 18516 3860 18545 3876
rect 18516 3852 18551 3860
rect 18516 3826 18517 3852
rect 18524 3826 18551 3852
rect 18459 3808 18489 3822
rect 18516 3818 18551 3826
rect 18516 3808 18545 3818
rect -1 3802 18545 3808
rect 0 3794 18545 3802
rect 15 3764 28 3794
rect 43 3780 73 3794
rect 116 3780 159 3794
rect 166 3780 386 3794
rect 393 3780 423 3794
rect 83 3766 98 3778
rect 117 3766 130 3780
rect 198 3776 351 3780
rect 80 3764 102 3766
rect 180 3764 372 3776
rect 451 3764 464 3794
rect 479 3780 509 3794
rect 546 3764 565 3794
rect 580 3764 586 3794
rect 595 3764 608 3794
rect 623 3780 653 3794
rect 696 3780 739 3794
rect 746 3780 966 3794
rect 973 3780 1003 3794
rect 663 3766 678 3778
rect 697 3766 710 3780
rect 778 3776 931 3780
rect 660 3764 682 3766
rect 760 3764 952 3776
rect 1031 3764 1044 3794
rect 1059 3780 1089 3794
rect 1126 3764 1145 3794
rect 1160 3764 1166 3794
rect 1175 3764 1188 3794
rect 1203 3780 1233 3794
rect 1276 3780 1319 3794
rect 1326 3780 1546 3794
rect 1553 3780 1583 3794
rect 1243 3766 1258 3778
rect 1277 3766 1290 3780
rect 1358 3776 1511 3780
rect 1240 3764 1262 3766
rect 1340 3764 1532 3776
rect 1611 3764 1624 3794
rect 1639 3780 1669 3794
rect 1706 3764 1725 3794
rect 1740 3764 1746 3794
rect 1755 3764 1768 3794
rect 1783 3780 1813 3794
rect 1856 3780 1899 3794
rect 1906 3780 2126 3794
rect 2133 3780 2163 3794
rect 1823 3766 1838 3778
rect 1857 3766 1870 3780
rect 1938 3776 2091 3780
rect 1820 3764 1842 3766
rect 1920 3764 2112 3776
rect 2191 3764 2204 3794
rect 2219 3780 2249 3794
rect 2286 3764 2305 3794
rect 2320 3764 2326 3794
rect 2335 3764 2348 3794
rect 2363 3780 2393 3794
rect 2436 3780 2479 3794
rect 2486 3780 2706 3794
rect 2713 3780 2743 3794
rect 2403 3766 2418 3778
rect 2437 3766 2450 3780
rect 2518 3776 2671 3780
rect 2400 3764 2422 3766
rect 2500 3764 2692 3776
rect 2771 3764 2784 3794
rect 2799 3780 2829 3794
rect 2866 3764 2885 3794
rect 2900 3764 2906 3794
rect 2915 3764 2928 3794
rect 2943 3780 2973 3794
rect 3016 3780 3059 3794
rect 3066 3780 3286 3794
rect 3293 3780 3323 3794
rect 2983 3766 2998 3778
rect 3017 3766 3030 3780
rect 3098 3776 3251 3780
rect 2980 3764 3002 3766
rect 3080 3764 3272 3776
rect 3351 3764 3364 3794
rect 3379 3780 3409 3794
rect 3446 3764 3465 3794
rect 3480 3764 3486 3794
rect 3495 3764 3508 3794
rect 3523 3780 3553 3794
rect 3596 3780 3639 3794
rect 3646 3780 3866 3794
rect 3873 3780 3903 3794
rect 3563 3766 3578 3778
rect 3597 3766 3610 3780
rect 3678 3776 3831 3780
rect 3560 3764 3582 3766
rect 3660 3764 3852 3776
rect 3931 3764 3944 3794
rect 3959 3780 3989 3794
rect 4026 3764 4045 3794
rect 4060 3764 4066 3794
rect 4075 3764 4088 3794
rect 4103 3780 4133 3794
rect 4176 3780 4219 3794
rect 4226 3780 4446 3794
rect 4453 3780 4483 3794
rect 4143 3766 4158 3778
rect 4177 3766 4190 3780
rect 4258 3776 4411 3780
rect 4140 3764 4162 3766
rect 4240 3764 4432 3776
rect 4511 3764 4524 3794
rect 4539 3780 4569 3794
rect 4606 3764 4625 3794
rect 4640 3764 4646 3794
rect 4655 3764 4668 3794
rect 4683 3780 4713 3794
rect 4756 3780 4799 3794
rect 4806 3780 5026 3794
rect 5033 3780 5063 3794
rect 4723 3766 4738 3778
rect 4757 3766 4770 3780
rect 4838 3776 4991 3780
rect 4720 3764 4742 3766
rect 4820 3764 5012 3776
rect 5091 3764 5104 3794
rect 5119 3780 5149 3794
rect 5186 3764 5205 3794
rect 5220 3764 5226 3794
rect 5235 3764 5248 3794
rect 5263 3780 5293 3794
rect 5336 3780 5379 3794
rect 5386 3780 5606 3794
rect 5613 3780 5643 3794
rect 5303 3766 5318 3778
rect 5337 3766 5350 3780
rect 5418 3776 5571 3780
rect 5300 3764 5322 3766
rect 5400 3764 5592 3776
rect 5671 3764 5684 3794
rect 5699 3780 5729 3794
rect 5766 3764 5785 3794
rect 5800 3764 5806 3794
rect 5815 3764 5828 3794
rect 5843 3780 5873 3794
rect 5916 3780 5959 3794
rect 5966 3780 6186 3794
rect 6193 3780 6223 3794
rect 5883 3766 5898 3778
rect 5917 3766 5930 3780
rect 5998 3776 6151 3780
rect 5880 3764 5902 3766
rect 5980 3764 6172 3776
rect 6251 3764 6264 3794
rect 6279 3780 6309 3794
rect 6346 3764 6365 3794
rect 6380 3764 6386 3794
rect 6395 3764 6408 3794
rect 6423 3780 6453 3794
rect 6496 3780 6539 3794
rect 6546 3780 6766 3794
rect 6773 3780 6803 3794
rect 6463 3766 6478 3778
rect 6497 3766 6510 3780
rect 6578 3776 6731 3780
rect 6460 3764 6482 3766
rect 6560 3764 6752 3776
rect 6831 3764 6844 3794
rect 6859 3780 6889 3794
rect 6926 3764 6945 3794
rect 6960 3764 6966 3794
rect 6975 3764 6988 3794
rect 7003 3780 7033 3794
rect 7076 3780 7119 3794
rect 7126 3780 7346 3794
rect 7353 3780 7383 3794
rect 7043 3766 7058 3778
rect 7077 3766 7090 3780
rect 7158 3776 7311 3780
rect 7040 3764 7062 3766
rect 7140 3764 7332 3776
rect 7411 3764 7424 3794
rect 7439 3780 7469 3794
rect 7506 3764 7525 3794
rect 7540 3764 7546 3794
rect 7555 3764 7568 3794
rect 7583 3780 7613 3794
rect 7656 3780 7699 3794
rect 7706 3780 7926 3794
rect 7933 3780 7963 3794
rect 7623 3766 7638 3778
rect 7657 3766 7670 3780
rect 7738 3776 7891 3780
rect 7620 3764 7642 3766
rect 7720 3764 7912 3776
rect 7991 3764 8004 3794
rect 8019 3780 8049 3794
rect 8086 3764 8105 3794
rect 8120 3764 8126 3794
rect 8135 3764 8148 3794
rect 8163 3780 8193 3794
rect 8236 3780 8279 3794
rect 8286 3780 8506 3794
rect 8513 3780 8543 3794
rect 8203 3766 8218 3778
rect 8237 3766 8250 3780
rect 8318 3776 8471 3780
rect 8200 3764 8222 3766
rect 8300 3764 8492 3776
rect 8571 3764 8584 3794
rect 8599 3780 8629 3794
rect 8666 3764 8685 3794
rect 8700 3764 8706 3794
rect 8715 3764 8728 3794
rect 8743 3780 8773 3794
rect 8816 3780 8859 3794
rect 8866 3780 9086 3794
rect 9093 3780 9123 3794
rect 8783 3766 8798 3778
rect 8817 3766 8830 3780
rect 8898 3776 9051 3780
rect 8780 3764 8802 3766
rect 8880 3764 9072 3776
rect 9151 3764 9164 3794
rect 9179 3780 9209 3794
rect 9246 3764 9265 3794
rect 9280 3764 9286 3794
rect 9295 3764 9308 3794
rect 9323 3780 9353 3794
rect 9396 3780 9439 3794
rect 9446 3780 9666 3794
rect 9673 3780 9703 3794
rect 9363 3766 9378 3778
rect 9397 3766 9410 3780
rect 9478 3776 9631 3780
rect 9360 3764 9382 3766
rect 9460 3764 9652 3776
rect 9731 3764 9744 3794
rect 9759 3780 9789 3794
rect 9826 3764 9845 3794
rect 9860 3764 9866 3794
rect 9875 3764 9888 3794
rect 9903 3780 9933 3794
rect 9976 3780 10019 3794
rect 10026 3780 10246 3794
rect 10253 3780 10283 3794
rect 9943 3766 9958 3778
rect 9977 3766 9990 3780
rect 10058 3776 10211 3780
rect 9940 3764 9962 3766
rect 10040 3764 10232 3776
rect 10311 3764 10324 3794
rect 10339 3780 10369 3794
rect 10406 3764 10425 3794
rect 10440 3764 10446 3794
rect 10455 3764 10468 3794
rect 10483 3780 10513 3794
rect 10556 3780 10599 3794
rect 10606 3780 10826 3794
rect 10833 3780 10863 3794
rect 10523 3766 10538 3778
rect 10557 3766 10570 3780
rect 10638 3776 10791 3780
rect 10520 3764 10542 3766
rect 10620 3764 10812 3776
rect 10891 3764 10904 3794
rect 10919 3780 10949 3794
rect 10986 3764 11005 3794
rect 11020 3764 11026 3794
rect 11035 3764 11048 3794
rect 11063 3780 11093 3794
rect 11136 3780 11179 3794
rect 11186 3780 11406 3794
rect 11413 3780 11443 3794
rect 11103 3766 11118 3778
rect 11137 3766 11150 3780
rect 11218 3776 11371 3780
rect 11100 3764 11122 3766
rect 11200 3764 11392 3776
rect 11471 3764 11484 3794
rect 11499 3780 11529 3794
rect 11566 3764 11585 3794
rect 11600 3764 11606 3794
rect 11615 3764 11628 3794
rect 11643 3780 11673 3794
rect 11716 3780 11759 3794
rect 11766 3780 11986 3794
rect 11993 3780 12023 3794
rect 11683 3766 11698 3778
rect 11717 3766 11730 3780
rect 11798 3776 11951 3780
rect 11680 3764 11702 3766
rect 11780 3764 11972 3776
rect 12051 3764 12064 3794
rect 12079 3780 12109 3794
rect 12146 3764 12165 3794
rect 12180 3764 12186 3794
rect 12195 3764 12208 3794
rect 12223 3780 12253 3794
rect 12296 3780 12339 3794
rect 12346 3780 12566 3794
rect 12573 3780 12603 3794
rect 12263 3766 12278 3778
rect 12297 3766 12310 3780
rect 12378 3776 12531 3780
rect 12260 3764 12282 3766
rect 12360 3764 12552 3776
rect 12631 3764 12644 3794
rect 12659 3780 12689 3794
rect 12726 3764 12745 3794
rect 12760 3764 12766 3794
rect 12775 3764 12788 3794
rect 12803 3780 12833 3794
rect 12876 3780 12919 3794
rect 12926 3780 13146 3794
rect 13153 3780 13183 3794
rect 12843 3766 12858 3778
rect 12877 3766 12890 3780
rect 12958 3776 13111 3780
rect 12840 3764 12862 3766
rect 12940 3764 13132 3776
rect 13211 3764 13224 3794
rect 13239 3780 13269 3794
rect 13306 3764 13325 3794
rect 13340 3764 13346 3794
rect 13355 3764 13368 3794
rect 13383 3780 13413 3794
rect 13456 3780 13499 3794
rect 13506 3780 13726 3794
rect 13733 3780 13763 3794
rect 13423 3766 13438 3778
rect 13457 3766 13470 3780
rect 13538 3776 13691 3780
rect 13420 3764 13442 3766
rect 13520 3764 13712 3776
rect 13791 3764 13804 3794
rect 13819 3780 13849 3794
rect 13886 3764 13905 3794
rect 13920 3764 13926 3794
rect 13935 3764 13948 3794
rect 13963 3780 13993 3794
rect 14036 3780 14079 3794
rect 14086 3780 14306 3794
rect 14313 3780 14343 3794
rect 14003 3766 14018 3778
rect 14037 3766 14050 3780
rect 14118 3776 14271 3780
rect 14000 3764 14022 3766
rect 14100 3764 14292 3776
rect 14371 3764 14384 3794
rect 14399 3780 14429 3794
rect 14466 3764 14485 3794
rect 14500 3764 14506 3794
rect 14515 3764 14528 3794
rect 14543 3780 14573 3794
rect 14616 3780 14659 3794
rect 14666 3780 14886 3794
rect 14893 3780 14923 3794
rect 14583 3766 14598 3778
rect 14617 3766 14630 3780
rect 14698 3776 14851 3780
rect 14580 3764 14602 3766
rect 14680 3764 14872 3776
rect 14951 3764 14964 3794
rect 14979 3780 15009 3794
rect 15046 3764 15065 3794
rect 15080 3764 15086 3794
rect 15095 3764 15108 3794
rect 15123 3780 15153 3794
rect 15196 3780 15239 3794
rect 15246 3780 15466 3794
rect 15473 3780 15503 3794
rect 15163 3766 15178 3778
rect 15197 3766 15210 3780
rect 15278 3776 15431 3780
rect 15160 3764 15182 3766
rect 15260 3764 15452 3776
rect 15531 3764 15544 3794
rect 15559 3780 15589 3794
rect 15626 3764 15645 3794
rect 15660 3764 15666 3794
rect 15675 3764 15688 3794
rect 15703 3780 15733 3794
rect 15776 3780 15819 3794
rect 15826 3780 16046 3794
rect 16053 3780 16083 3794
rect 15743 3766 15758 3778
rect 15777 3766 15790 3780
rect 15858 3776 16011 3780
rect 15740 3764 15762 3766
rect 15840 3764 16032 3776
rect 16111 3764 16124 3794
rect 16139 3780 16169 3794
rect 16206 3764 16225 3794
rect 16240 3764 16246 3794
rect 16255 3764 16268 3794
rect 16283 3780 16313 3794
rect 16356 3780 16399 3794
rect 16406 3780 16626 3794
rect 16633 3780 16663 3794
rect 16323 3766 16338 3778
rect 16357 3766 16370 3780
rect 16438 3776 16591 3780
rect 16320 3764 16342 3766
rect 16420 3764 16612 3776
rect 16691 3764 16704 3794
rect 16719 3780 16749 3794
rect 16786 3764 16805 3794
rect 16820 3764 16826 3794
rect 16835 3764 16848 3794
rect 16863 3780 16893 3794
rect 16936 3780 16979 3794
rect 16986 3780 17206 3794
rect 17213 3780 17243 3794
rect 16903 3766 16918 3778
rect 16937 3766 16950 3780
rect 17018 3776 17171 3780
rect 16900 3764 16922 3766
rect 17000 3764 17192 3776
rect 17271 3764 17284 3794
rect 17299 3780 17329 3794
rect 17366 3764 17385 3794
rect 17400 3764 17406 3794
rect 17415 3764 17428 3794
rect 17443 3780 17473 3794
rect 17516 3780 17559 3794
rect 17566 3780 17786 3794
rect 17793 3780 17823 3794
rect 17483 3766 17498 3778
rect 17517 3766 17530 3780
rect 17598 3776 17751 3780
rect 17480 3764 17502 3766
rect 17580 3764 17772 3776
rect 17851 3764 17864 3794
rect 17879 3780 17909 3794
rect 17946 3764 17965 3794
rect 17980 3764 17986 3794
rect 17995 3764 18008 3794
rect 18023 3780 18053 3794
rect 18096 3780 18139 3794
rect 18146 3780 18366 3794
rect 18373 3780 18403 3794
rect 18063 3766 18078 3778
rect 18097 3766 18110 3780
rect 18178 3776 18331 3780
rect 18060 3764 18082 3766
rect 18160 3764 18352 3776
rect 18431 3764 18444 3794
rect 18459 3780 18489 3794
rect 18532 3764 18545 3794
rect 0 3750 18545 3764
rect 15 3680 28 3750
rect 80 3746 102 3750
rect 73 3724 102 3738
rect 155 3724 171 3738
rect 209 3734 215 3736
rect 222 3734 330 3750
rect 337 3734 343 3736
rect 351 3734 366 3750
rect 432 3744 451 3747
rect 73 3722 171 3724
rect 198 3722 366 3734
rect 381 3724 397 3738
rect 432 3725 454 3744
rect 464 3738 480 3739
rect 463 3736 480 3738
rect 464 3731 480 3736
rect 454 3724 460 3725
rect 463 3724 492 3731
rect 381 3723 492 3724
rect 381 3722 498 3723
rect 57 3714 108 3722
rect 155 3714 189 3722
rect 57 3702 82 3714
rect 89 3702 108 3714
rect 162 3712 189 3714
rect 198 3712 419 3722
rect 454 3719 460 3722
rect 162 3708 419 3712
rect 57 3694 108 3702
rect 155 3694 419 3708
rect 463 3714 498 3722
rect 9 3646 28 3680
rect 73 3686 102 3694
rect 73 3680 90 3686
rect 73 3678 107 3680
rect 155 3678 171 3694
rect 172 3684 380 3694
rect 381 3684 397 3694
rect 445 3690 460 3705
rect 463 3702 464 3714
rect 471 3702 498 3714
rect 463 3694 498 3702
rect 463 3693 492 3694
rect 183 3680 397 3684
rect 198 3678 397 3680
rect 432 3680 445 3690
rect 463 3680 480 3693
rect 432 3678 480 3680
rect 74 3674 107 3678
rect 70 3672 107 3674
rect 70 3671 137 3672
rect 70 3666 101 3671
rect 107 3666 137 3671
rect 70 3662 137 3666
rect 43 3659 137 3662
rect 43 3652 92 3659
rect 43 3646 73 3652
rect 92 3647 97 3652
rect 9 3630 89 3646
rect 101 3638 137 3659
rect 198 3654 387 3678
rect 432 3677 479 3678
rect 445 3672 479 3677
rect 213 3651 387 3654
rect 206 3648 387 3651
rect 415 3671 479 3672
rect 9 3628 28 3630
rect 43 3628 77 3630
rect 9 3612 89 3628
rect 9 3606 28 3612
rect -1 3590 28 3606
rect 43 3596 73 3612
rect 101 3590 107 3638
rect 110 3632 129 3638
rect 144 3632 174 3640
rect 110 3624 174 3632
rect 110 3608 190 3624
rect 206 3617 268 3648
rect 284 3617 346 3648
rect 415 3646 464 3671
rect 479 3646 509 3662
rect 378 3632 408 3640
rect 415 3638 525 3646
rect 378 3624 423 3632
rect 110 3606 129 3608
rect 144 3606 190 3608
rect 110 3590 190 3606
rect 217 3604 252 3617
rect 293 3614 330 3617
rect 293 3612 335 3614
rect 222 3601 252 3604
rect 231 3597 238 3601
rect 238 3596 239 3597
rect 197 3590 207 3596
rect -7 3582 34 3590
rect -7 3556 8 3582
rect 15 3556 34 3582
rect 98 3578 129 3590
rect 144 3578 247 3590
rect 259 3580 285 3606
rect 300 3601 330 3612
rect 362 3608 424 3624
rect 362 3606 408 3608
rect 362 3590 424 3606
rect 436 3590 442 3638
rect 445 3630 525 3638
rect 445 3628 464 3630
rect 479 3628 513 3630
rect 445 3612 525 3628
rect 445 3590 464 3612
rect 479 3596 509 3612
rect 537 3606 543 3680
rect 546 3606 565 3750
rect 580 3606 586 3750
rect 595 3680 608 3750
rect 660 3746 682 3750
rect 653 3724 682 3738
rect 735 3724 751 3738
rect 789 3734 795 3736
rect 802 3734 910 3750
rect 917 3734 923 3736
rect 931 3734 946 3750
rect 1012 3744 1031 3747
rect 653 3722 751 3724
rect 778 3722 946 3734
rect 961 3724 977 3738
rect 1012 3725 1034 3744
rect 1044 3738 1060 3739
rect 1043 3736 1060 3738
rect 1044 3731 1060 3736
rect 1034 3724 1040 3725
rect 1043 3724 1072 3731
rect 961 3723 1072 3724
rect 961 3722 1078 3723
rect 637 3714 688 3722
rect 735 3714 769 3722
rect 637 3702 662 3714
rect 669 3702 688 3714
rect 742 3712 769 3714
rect 778 3712 999 3722
rect 1034 3719 1040 3722
rect 742 3708 999 3712
rect 637 3694 688 3702
rect 735 3694 999 3708
rect 1043 3714 1078 3722
rect 589 3646 608 3680
rect 653 3686 682 3694
rect 653 3680 670 3686
rect 653 3678 687 3680
rect 735 3678 751 3694
rect 752 3684 960 3694
rect 961 3684 977 3694
rect 1025 3690 1040 3705
rect 1043 3702 1044 3714
rect 1051 3702 1078 3714
rect 1043 3694 1078 3702
rect 1043 3693 1072 3694
rect 763 3680 977 3684
rect 778 3678 977 3680
rect 1012 3680 1025 3690
rect 1043 3680 1060 3693
rect 1012 3678 1060 3680
rect 654 3674 687 3678
rect 650 3672 687 3674
rect 650 3671 717 3672
rect 650 3666 681 3671
rect 687 3666 717 3671
rect 650 3662 717 3666
rect 623 3659 717 3662
rect 623 3652 672 3659
rect 623 3646 653 3652
rect 672 3647 677 3652
rect 589 3630 669 3646
rect 681 3638 717 3659
rect 778 3654 967 3678
rect 1012 3677 1059 3678
rect 1025 3672 1059 3677
rect 793 3651 967 3654
rect 786 3648 967 3651
rect 995 3671 1059 3672
rect 589 3628 608 3630
rect 623 3628 657 3630
rect 589 3612 669 3628
rect 589 3606 608 3612
rect 305 3580 408 3590
rect 259 3578 408 3580
rect 429 3578 464 3590
rect 98 3576 260 3578
rect 110 3556 129 3576
rect 144 3574 174 3576
rect -7 3548 34 3556
rect 116 3552 129 3556
rect 181 3560 260 3576
rect 292 3576 464 3578
rect 292 3560 371 3576
rect 378 3574 408 3576
rect -1 3538 28 3548
rect 43 3538 73 3552
rect 116 3538 159 3552
rect 181 3548 371 3560
rect 436 3556 442 3576
rect 166 3538 196 3548
rect 197 3538 355 3548
rect 359 3538 389 3548
rect 393 3538 423 3552
rect 451 3538 464 3576
rect 536 3590 565 3606
rect 579 3590 608 3606
rect 623 3596 653 3612
rect 681 3590 687 3638
rect 690 3632 709 3638
rect 724 3632 754 3640
rect 690 3624 754 3632
rect 690 3608 770 3624
rect 786 3617 848 3648
rect 864 3617 926 3648
rect 995 3646 1044 3671
rect 1059 3646 1089 3662
rect 958 3632 988 3640
rect 995 3638 1105 3646
rect 958 3624 1003 3632
rect 690 3606 709 3608
rect 724 3606 770 3608
rect 690 3590 770 3606
rect 797 3604 832 3617
rect 873 3614 910 3617
rect 873 3612 915 3614
rect 802 3601 832 3604
rect 811 3597 818 3601
rect 818 3596 819 3597
rect 777 3590 787 3596
rect 536 3582 571 3590
rect 536 3556 537 3582
rect 544 3556 571 3582
rect 479 3538 509 3552
rect 536 3548 571 3556
rect 573 3582 614 3590
rect 573 3556 588 3582
rect 595 3556 614 3582
rect 678 3578 709 3590
rect 724 3578 827 3590
rect 839 3580 865 3606
rect 880 3601 910 3612
rect 942 3608 1004 3624
rect 942 3606 988 3608
rect 942 3590 1004 3606
rect 1016 3590 1022 3638
rect 1025 3630 1105 3638
rect 1025 3628 1044 3630
rect 1059 3628 1093 3630
rect 1025 3612 1105 3628
rect 1025 3590 1044 3612
rect 1059 3596 1089 3612
rect 1117 3606 1123 3680
rect 1126 3606 1145 3750
rect 1160 3606 1166 3750
rect 1175 3680 1188 3750
rect 1240 3746 1262 3750
rect 1233 3724 1262 3738
rect 1315 3724 1331 3738
rect 1369 3734 1375 3736
rect 1382 3734 1490 3750
rect 1497 3734 1503 3736
rect 1511 3734 1526 3750
rect 1592 3744 1611 3747
rect 1233 3722 1331 3724
rect 1358 3722 1526 3734
rect 1541 3724 1557 3738
rect 1592 3725 1614 3744
rect 1624 3738 1640 3739
rect 1623 3736 1640 3738
rect 1624 3731 1640 3736
rect 1614 3724 1620 3725
rect 1623 3724 1652 3731
rect 1541 3723 1652 3724
rect 1541 3722 1658 3723
rect 1217 3714 1268 3722
rect 1315 3714 1349 3722
rect 1217 3702 1242 3714
rect 1249 3702 1268 3714
rect 1322 3712 1349 3714
rect 1358 3712 1579 3722
rect 1614 3719 1620 3722
rect 1322 3708 1579 3712
rect 1217 3694 1268 3702
rect 1315 3694 1579 3708
rect 1623 3714 1658 3722
rect 1169 3646 1188 3680
rect 1233 3686 1262 3694
rect 1233 3680 1250 3686
rect 1233 3678 1267 3680
rect 1315 3678 1331 3694
rect 1332 3684 1540 3694
rect 1541 3684 1557 3694
rect 1605 3690 1620 3705
rect 1623 3702 1624 3714
rect 1631 3702 1658 3714
rect 1623 3694 1658 3702
rect 1623 3693 1652 3694
rect 1343 3680 1557 3684
rect 1358 3678 1557 3680
rect 1592 3680 1605 3690
rect 1623 3680 1640 3693
rect 1592 3678 1640 3680
rect 1234 3674 1267 3678
rect 1230 3672 1267 3674
rect 1230 3671 1297 3672
rect 1230 3666 1261 3671
rect 1267 3666 1297 3671
rect 1230 3662 1297 3666
rect 1203 3659 1297 3662
rect 1203 3652 1252 3659
rect 1203 3646 1233 3652
rect 1252 3647 1257 3652
rect 1169 3630 1249 3646
rect 1261 3638 1297 3659
rect 1358 3654 1547 3678
rect 1592 3677 1639 3678
rect 1605 3672 1639 3677
rect 1373 3651 1547 3654
rect 1366 3648 1547 3651
rect 1575 3671 1639 3672
rect 1169 3628 1188 3630
rect 1203 3628 1237 3630
rect 1169 3612 1249 3628
rect 1169 3606 1188 3612
rect 885 3580 988 3590
rect 839 3578 988 3580
rect 1009 3578 1044 3590
rect 678 3576 840 3578
rect 690 3556 709 3576
rect 724 3574 754 3576
rect 573 3548 614 3556
rect 696 3552 709 3556
rect 761 3560 840 3576
rect 872 3576 1044 3578
rect 872 3560 951 3576
rect 958 3574 988 3576
rect 536 3538 565 3548
rect 579 3538 608 3548
rect 623 3538 653 3552
rect 696 3538 739 3552
rect 761 3548 951 3560
rect 1016 3556 1022 3576
rect 746 3538 776 3548
rect 777 3538 935 3548
rect 939 3538 969 3548
rect 973 3538 1003 3552
rect 1031 3538 1044 3576
rect 1116 3590 1145 3606
rect 1159 3590 1188 3606
rect 1203 3596 1233 3612
rect 1261 3590 1267 3638
rect 1270 3632 1289 3638
rect 1304 3632 1334 3640
rect 1270 3624 1334 3632
rect 1270 3608 1350 3624
rect 1366 3617 1428 3648
rect 1444 3617 1506 3648
rect 1575 3646 1624 3671
rect 1639 3646 1669 3662
rect 1538 3632 1568 3640
rect 1575 3638 1685 3646
rect 1538 3624 1583 3632
rect 1270 3606 1289 3608
rect 1304 3606 1350 3608
rect 1270 3590 1350 3606
rect 1377 3604 1412 3617
rect 1453 3614 1490 3617
rect 1453 3612 1495 3614
rect 1382 3601 1412 3604
rect 1391 3597 1398 3601
rect 1398 3596 1399 3597
rect 1357 3590 1367 3596
rect 1116 3582 1151 3590
rect 1116 3556 1117 3582
rect 1124 3556 1151 3582
rect 1059 3538 1089 3552
rect 1116 3548 1151 3556
rect 1153 3582 1194 3590
rect 1153 3556 1168 3582
rect 1175 3556 1194 3582
rect 1258 3578 1289 3590
rect 1304 3578 1407 3590
rect 1419 3580 1445 3606
rect 1460 3601 1490 3612
rect 1522 3608 1584 3624
rect 1522 3606 1568 3608
rect 1522 3590 1584 3606
rect 1596 3590 1602 3638
rect 1605 3630 1685 3638
rect 1605 3628 1624 3630
rect 1639 3628 1673 3630
rect 1605 3612 1685 3628
rect 1605 3590 1624 3612
rect 1639 3596 1669 3612
rect 1697 3606 1703 3680
rect 1706 3606 1725 3750
rect 1740 3606 1746 3750
rect 1755 3680 1768 3750
rect 1820 3746 1842 3750
rect 1813 3724 1842 3738
rect 1895 3724 1911 3738
rect 1949 3734 1955 3736
rect 1962 3734 2070 3750
rect 2077 3734 2083 3736
rect 2091 3734 2106 3750
rect 2172 3744 2191 3747
rect 1813 3722 1911 3724
rect 1938 3722 2106 3734
rect 2121 3724 2137 3738
rect 2172 3725 2194 3744
rect 2204 3738 2220 3739
rect 2203 3736 2220 3738
rect 2204 3731 2220 3736
rect 2194 3724 2200 3725
rect 2203 3724 2232 3731
rect 2121 3723 2232 3724
rect 2121 3722 2238 3723
rect 1797 3714 1848 3722
rect 1895 3714 1929 3722
rect 1797 3702 1822 3714
rect 1829 3702 1848 3714
rect 1902 3712 1929 3714
rect 1938 3712 2159 3722
rect 2194 3719 2200 3722
rect 1902 3708 2159 3712
rect 1797 3694 1848 3702
rect 1895 3694 2159 3708
rect 2203 3714 2238 3722
rect 1749 3646 1768 3680
rect 1813 3686 1842 3694
rect 1813 3680 1830 3686
rect 1813 3678 1847 3680
rect 1895 3678 1911 3694
rect 1912 3684 2120 3694
rect 2121 3684 2137 3694
rect 2185 3690 2200 3705
rect 2203 3702 2204 3714
rect 2211 3702 2238 3714
rect 2203 3694 2238 3702
rect 2203 3693 2232 3694
rect 1923 3680 2137 3684
rect 1938 3678 2137 3680
rect 2172 3680 2185 3690
rect 2203 3680 2220 3693
rect 2172 3678 2220 3680
rect 1814 3674 1847 3678
rect 1810 3672 1847 3674
rect 1810 3671 1877 3672
rect 1810 3666 1841 3671
rect 1847 3666 1877 3671
rect 1810 3662 1877 3666
rect 1783 3659 1877 3662
rect 1783 3652 1832 3659
rect 1783 3646 1813 3652
rect 1832 3647 1837 3652
rect 1749 3630 1829 3646
rect 1841 3638 1877 3659
rect 1938 3654 2127 3678
rect 2172 3677 2219 3678
rect 2185 3672 2219 3677
rect 1953 3651 2127 3654
rect 1946 3648 2127 3651
rect 2155 3671 2219 3672
rect 1749 3628 1768 3630
rect 1783 3628 1817 3630
rect 1749 3612 1829 3628
rect 1749 3606 1768 3612
rect 1465 3580 1568 3590
rect 1419 3578 1568 3580
rect 1589 3578 1624 3590
rect 1258 3576 1420 3578
rect 1270 3556 1289 3576
rect 1304 3574 1334 3576
rect 1153 3548 1194 3556
rect 1276 3552 1289 3556
rect 1341 3560 1420 3576
rect 1452 3576 1624 3578
rect 1452 3560 1531 3576
rect 1538 3574 1568 3576
rect 1116 3538 1145 3548
rect 1159 3538 1188 3548
rect 1203 3538 1233 3552
rect 1276 3538 1319 3552
rect 1341 3548 1531 3560
rect 1596 3556 1602 3576
rect 1326 3538 1356 3548
rect 1357 3538 1515 3548
rect 1519 3538 1549 3548
rect 1553 3538 1583 3552
rect 1611 3538 1624 3576
rect 1696 3590 1725 3606
rect 1739 3590 1768 3606
rect 1783 3596 1813 3612
rect 1841 3590 1847 3638
rect 1850 3632 1869 3638
rect 1884 3632 1914 3640
rect 1850 3624 1914 3632
rect 1850 3608 1930 3624
rect 1946 3617 2008 3648
rect 2024 3617 2086 3648
rect 2155 3646 2204 3671
rect 2219 3646 2249 3662
rect 2118 3632 2148 3640
rect 2155 3638 2265 3646
rect 2118 3624 2163 3632
rect 1850 3606 1869 3608
rect 1884 3606 1930 3608
rect 1850 3590 1930 3606
rect 1957 3604 1992 3617
rect 2033 3614 2070 3617
rect 2033 3612 2075 3614
rect 1962 3601 1992 3604
rect 1971 3597 1978 3601
rect 1978 3596 1979 3597
rect 1937 3590 1947 3596
rect 1696 3582 1731 3590
rect 1696 3556 1697 3582
rect 1704 3556 1731 3582
rect 1639 3538 1669 3552
rect 1696 3548 1731 3556
rect 1733 3582 1774 3590
rect 1733 3556 1748 3582
rect 1755 3556 1774 3582
rect 1838 3578 1869 3590
rect 1884 3578 1987 3590
rect 1999 3580 2025 3606
rect 2040 3601 2070 3612
rect 2102 3608 2164 3624
rect 2102 3606 2148 3608
rect 2102 3590 2164 3606
rect 2176 3590 2182 3638
rect 2185 3630 2265 3638
rect 2185 3628 2204 3630
rect 2219 3628 2253 3630
rect 2185 3612 2265 3628
rect 2185 3590 2204 3612
rect 2219 3596 2249 3612
rect 2277 3606 2283 3680
rect 2286 3606 2305 3750
rect 2320 3606 2326 3750
rect 2335 3680 2348 3750
rect 2400 3746 2422 3750
rect 2393 3724 2422 3738
rect 2475 3724 2491 3738
rect 2529 3734 2535 3736
rect 2542 3734 2650 3750
rect 2657 3734 2663 3736
rect 2671 3734 2686 3750
rect 2752 3744 2771 3747
rect 2393 3722 2491 3724
rect 2518 3722 2686 3734
rect 2701 3724 2717 3738
rect 2752 3725 2774 3744
rect 2784 3738 2800 3739
rect 2783 3736 2800 3738
rect 2784 3731 2800 3736
rect 2774 3724 2780 3725
rect 2783 3724 2812 3731
rect 2701 3723 2812 3724
rect 2701 3722 2818 3723
rect 2377 3714 2428 3722
rect 2475 3714 2509 3722
rect 2377 3702 2402 3714
rect 2409 3702 2428 3714
rect 2482 3712 2509 3714
rect 2518 3712 2739 3722
rect 2774 3719 2780 3722
rect 2482 3708 2739 3712
rect 2377 3694 2428 3702
rect 2475 3694 2739 3708
rect 2783 3714 2818 3722
rect 2329 3646 2348 3680
rect 2393 3686 2422 3694
rect 2393 3680 2410 3686
rect 2393 3678 2427 3680
rect 2475 3678 2491 3694
rect 2492 3684 2700 3694
rect 2701 3684 2717 3694
rect 2765 3690 2780 3705
rect 2783 3702 2784 3714
rect 2791 3702 2818 3714
rect 2783 3694 2818 3702
rect 2783 3693 2812 3694
rect 2503 3680 2717 3684
rect 2518 3678 2717 3680
rect 2752 3680 2765 3690
rect 2783 3680 2800 3693
rect 2752 3678 2800 3680
rect 2394 3674 2427 3678
rect 2390 3672 2427 3674
rect 2390 3671 2457 3672
rect 2390 3666 2421 3671
rect 2427 3666 2457 3671
rect 2390 3662 2457 3666
rect 2363 3659 2457 3662
rect 2363 3652 2412 3659
rect 2363 3646 2393 3652
rect 2412 3647 2417 3652
rect 2329 3630 2409 3646
rect 2421 3638 2457 3659
rect 2518 3654 2707 3678
rect 2752 3677 2799 3678
rect 2765 3672 2799 3677
rect 2533 3651 2707 3654
rect 2526 3648 2707 3651
rect 2735 3671 2799 3672
rect 2329 3628 2348 3630
rect 2363 3628 2397 3630
rect 2329 3612 2409 3628
rect 2329 3606 2348 3612
rect 2045 3580 2148 3590
rect 1999 3578 2148 3580
rect 2169 3578 2204 3590
rect 1838 3576 2000 3578
rect 1850 3556 1869 3576
rect 1884 3574 1914 3576
rect 1733 3548 1774 3556
rect 1856 3552 1869 3556
rect 1921 3560 2000 3576
rect 2032 3576 2204 3578
rect 2032 3560 2111 3576
rect 2118 3574 2148 3576
rect 1696 3538 1725 3548
rect 1739 3538 1768 3548
rect 1783 3538 1813 3552
rect 1856 3538 1899 3552
rect 1921 3548 2111 3560
rect 2176 3556 2182 3576
rect 1906 3538 1936 3548
rect 1937 3538 2095 3548
rect 2099 3538 2129 3548
rect 2133 3538 2163 3552
rect 2191 3538 2204 3576
rect 2276 3590 2305 3606
rect 2319 3590 2348 3606
rect 2363 3596 2393 3612
rect 2421 3590 2427 3638
rect 2430 3632 2449 3638
rect 2464 3632 2494 3640
rect 2430 3624 2494 3632
rect 2430 3608 2510 3624
rect 2526 3617 2588 3648
rect 2604 3617 2666 3648
rect 2735 3646 2784 3671
rect 2799 3646 2829 3662
rect 2698 3632 2728 3640
rect 2735 3638 2845 3646
rect 2698 3624 2743 3632
rect 2430 3606 2449 3608
rect 2464 3606 2510 3608
rect 2430 3590 2510 3606
rect 2537 3604 2572 3617
rect 2613 3614 2650 3617
rect 2613 3612 2655 3614
rect 2542 3601 2572 3604
rect 2551 3597 2558 3601
rect 2558 3596 2559 3597
rect 2517 3590 2527 3596
rect 2276 3582 2311 3590
rect 2276 3556 2277 3582
rect 2284 3556 2311 3582
rect 2219 3538 2249 3552
rect 2276 3548 2311 3556
rect 2313 3582 2354 3590
rect 2313 3556 2328 3582
rect 2335 3556 2354 3582
rect 2418 3578 2449 3590
rect 2464 3578 2567 3590
rect 2579 3580 2605 3606
rect 2620 3601 2650 3612
rect 2682 3608 2744 3624
rect 2682 3606 2728 3608
rect 2682 3590 2744 3606
rect 2756 3590 2762 3638
rect 2765 3630 2845 3638
rect 2765 3628 2784 3630
rect 2799 3628 2833 3630
rect 2765 3612 2845 3628
rect 2765 3590 2784 3612
rect 2799 3596 2829 3612
rect 2857 3606 2863 3680
rect 2866 3606 2885 3750
rect 2900 3606 2906 3750
rect 2915 3680 2928 3750
rect 2980 3746 3002 3750
rect 2973 3724 3002 3738
rect 3055 3724 3071 3738
rect 3109 3734 3115 3736
rect 3122 3734 3230 3750
rect 3237 3734 3243 3736
rect 3251 3734 3266 3750
rect 3332 3744 3351 3747
rect 2973 3722 3071 3724
rect 3098 3722 3266 3734
rect 3281 3724 3297 3738
rect 3332 3725 3354 3744
rect 3364 3738 3380 3739
rect 3363 3736 3380 3738
rect 3364 3731 3380 3736
rect 3354 3724 3360 3725
rect 3363 3724 3392 3731
rect 3281 3723 3392 3724
rect 3281 3722 3398 3723
rect 2957 3714 3008 3722
rect 3055 3714 3089 3722
rect 2957 3702 2982 3714
rect 2989 3702 3008 3714
rect 3062 3712 3089 3714
rect 3098 3712 3319 3722
rect 3354 3719 3360 3722
rect 3062 3708 3319 3712
rect 2957 3694 3008 3702
rect 3055 3694 3319 3708
rect 3363 3714 3398 3722
rect 2909 3646 2928 3680
rect 2973 3686 3002 3694
rect 2973 3680 2990 3686
rect 2973 3678 3007 3680
rect 3055 3678 3071 3694
rect 3072 3684 3280 3694
rect 3281 3684 3297 3694
rect 3345 3690 3360 3705
rect 3363 3702 3364 3714
rect 3371 3702 3398 3714
rect 3363 3694 3398 3702
rect 3363 3693 3392 3694
rect 3083 3680 3297 3684
rect 3098 3678 3297 3680
rect 3332 3680 3345 3690
rect 3363 3680 3380 3693
rect 3332 3678 3380 3680
rect 2974 3674 3007 3678
rect 2970 3672 3007 3674
rect 2970 3671 3037 3672
rect 2970 3666 3001 3671
rect 3007 3666 3037 3671
rect 2970 3662 3037 3666
rect 2943 3659 3037 3662
rect 2943 3652 2992 3659
rect 2943 3646 2973 3652
rect 2992 3647 2997 3652
rect 2909 3630 2989 3646
rect 3001 3638 3037 3659
rect 3098 3654 3287 3678
rect 3332 3677 3379 3678
rect 3345 3672 3379 3677
rect 3113 3651 3287 3654
rect 3106 3648 3287 3651
rect 3315 3671 3379 3672
rect 2909 3628 2928 3630
rect 2943 3628 2977 3630
rect 2909 3612 2989 3628
rect 2909 3606 2928 3612
rect 2625 3580 2728 3590
rect 2579 3578 2728 3580
rect 2749 3578 2784 3590
rect 2418 3576 2580 3578
rect 2430 3556 2449 3576
rect 2464 3574 2494 3576
rect 2313 3548 2354 3556
rect 2436 3552 2449 3556
rect 2501 3560 2580 3576
rect 2612 3576 2784 3578
rect 2612 3560 2691 3576
rect 2698 3574 2728 3576
rect 2276 3538 2305 3548
rect 2319 3538 2348 3548
rect 2363 3538 2393 3552
rect 2436 3538 2479 3552
rect 2501 3548 2691 3560
rect 2756 3556 2762 3576
rect 2486 3538 2516 3548
rect 2517 3538 2675 3548
rect 2679 3538 2709 3548
rect 2713 3538 2743 3552
rect 2771 3538 2784 3576
rect 2856 3590 2885 3606
rect 2899 3590 2928 3606
rect 2943 3596 2973 3612
rect 3001 3590 3007 3638
rect 3010 3632 3029 3638
rect 3044 3632 3074 3640
rect 3010 3624 3074 3632
rect 3010 3608 3090 3624
rect 3106 3617 3168 3648
rect 3184 3617 3246 3648
rect 3315 3646 3364 3671
rect 3379 3646 3409 3662
rect 3278 3632 3308 3640
rect 3315 3638 3425 3646
rect 3278 3624 3323 3632
rect 3010 3606 3029 3608
rect 3044 3606 3090 3608
rect 3010 3590 3090 3606
rect 3117 3604 3152 3617
rect 3193 3614 3230 3617
rect 3193 3612 3235 3614
rect 3122 3601 3152 3604
rect 3131 3597 3138 3601
rect 3138 3596 3139 3597
rect 3097 3590 3107 3596
rect 2856 3582 2891 3590
rect 2856 3556 2857 3582
rect 2864 3556 2891 3582
rect 2799 3538 2829 3552
rect 2856 3548 2891 3556
rect 2893 3582 2934 3590
rect 2893 3556 2908 3582
rect 2915 3556 2934 3582
rect 2998 3578 3029 3590
rect 3044 3578 3147 3590
rect 3159 3580 3185 3606
rect 3200 3601 3230 3612
rect 3262 3608 3324 3624
rect 3262 3606 3308 3608
rect 3262 3590 3324 3606
rect 3336 3590 3342 3638
rect 3345 3630 3425 3638
rect 3345 3628 3364 3630
rect 3379 3628 3413 3630
rect 3345 3612 3425 3628
rect 3345 3590 3364 3612
rect 3379 3596 3409 3612
rect 3437 3606 3443 3680
rect 3446 3606 3465 3750
rect 3480 3606 3486 3750
rect 3495 3680 3508 3750
rect 3560 3746 3582 3750
rect 3553 3724 3582 3738
rect 3635 3724 3651 3738
rect 3689 3734 3695 3736
rect 3702 3734 3810 3750
rect 3817 3734 3823 3736
rect 3831 3734 3846 3750
rect 3912 3744 3931 3747
rect 3553 3722 3651 3724
rect 3678 3722 3846 3734
rect 3861 3724 3877 3738
rect 3912 3725 3934 3744
rect 3944 3738 3960 3739
rect 3943 3736 3960 3738
rect 3944 3731 3960 3736
rect 3934 3724 3940 3725
rect 3943 3724 3972 3731
rect 3861 3723 3972 3724
rect 3861 3722 3978 3723
rect 3537 3714 3588 3722
rect 3635 3714 3669 3722
rect 3537 3702 3562 3714
rect 3569 3702 3588 3714
rect 3642 3712 3669 3714
rect 3678 3712 3899 3722
rect 3934 3719 3940 3722
rect 3642 3708 3899 3712
rect 3537 3694 3588 3702
rect 3635 3694 3899 3708
rect 3943 3714 3978 3722
rect 3489 3646 3508 3680
rect 3553 3686 3582 3694
rect 3553 3680 3570 3686
rect 3553 3678 3587 3680
rect 3635 3678 3651 3694
rect 3652 3684 3860 3694
rect 3861 3684 3877 3694
rect 3925 3690 3940 3705
rect 3943 3702 3944 3714
rect 3951 3702 3978 3714
rect 3943 3694 3978 3702
rect 3943 3693 3972 3694
rect 3663 3680 3877 3684
rect 3678 3678 3877 3680
rect 3912 3680 3925 3690
rect 3943 3680 3960 3693
rect 3912 3678 3960 3680
rect 3554 3674 3587 3678
rect 3550 3672 3587 3674
rect 3550 3671 3617 3672
rect 3550 3666 3581 3671
rect 3587 3666 3617 3671
rect 3550 3662 3617 3666
rect 3523 3659 3617 3662
rect 3523 3652 3572 3659
rect 3523 3646 3553 3652
rect 3572 3647 3577 3652
rect 3489 3630 3569 3646
rect 3581 3638 3617 3659
rect 3678 3654 3867 3678
rect 3912 3677 3959 3678
rect 3925 3672 3959 3677
rect 3693 3651 3867 3654
rect 3686 3648 3867 3651
rect 3895 3671 3959 3672
rect 3489 3628 3508 3630
rect 3523 3628 3557 3630
rect 3489 3612 3569 3628
rect 3489 3606 3508 3612
rect 3205 3580 3308 3590
rect 3159 3578 3308 3580
rect 3329 3578 3364 3590
rect 2998 3576 3160 3578
rect 3010 3556 3029 3576
rect 3044 3574 3074 3576
rect 2893 3548 2934 3556
rect 3016 3552 3029 3556
rect 3081 3560 3160 3576
rect 3192 3576 3364 3578
rect 3192 3560 3271 3576
rect 3278 3574 3308 3576
rect 2856 3538 2885 3548
rect 2899 3538 2928 3548
rect 2943 3538 2973 3552
rect 3016 3538 3059 3552
rect 3081 3548 3271 3560
rect 3336 3556 3342 3576
rect 3066 3538 3096 3548
rect 3097 3538 3255 3548
rect 3259 3538 3289 3548
rect 3293 3538 3323 3552
rect 3351 3538 3364 3576
rect 3436 3590 3465 3606
rect 3479 3590 3508 3606
rect 3523 3596 3553 3612
rect 3581 3590 3587 3638
rect 3590 3632 3609 3638
rect 3624 3632 3654 3640
rect 3590 3624 3654 3632
rect 3590 3608 3670 3624
rect 3686 3617 3748 3648
rect 3764 3617 3826 3648
rect 3895 3646 3944 3671
rect 3959 3646 3989 3662
rect 3858 3632 3888 3640
rect 3895 3638 4005 3646
rect 3858 3624 3903 3632
rect 3590 3606 3609 3608
rect 3624 3606 3670 3608
rect 3590 3590 3670 3606
rect 3697 3604 3732 3617
rect 3773 3614 3810 3617
rect 3773 3612 3815 3614
rect 3702 3601 3732 3604
rect 3711 3597 3718 3601
rect 3718 3596 3719 3597
rect 3677 3590 3687 3596
rect 3436 3582 3471 3590
rect 3436 3556 3437 3582
rect 3444 3556 3471 3582
rect 3379 3538 3409 3552
rect 3436 3548 3471 3556
rect 3473 3582 3514 3590
rect 3473 3556 3488 3582
rect 3495 3556 3514 3582
rect 3578 3578 3609 3590
rect 3624 3578 3727 3590
rect 3739 3580 3765 3606
rect 3780 3601 3810 3612
rect 3842 3608 3904 3624
rect 3842 3606 3888 3608
rect 3842 3590 3904 3606
rect 3916 3590 3922 3638
rect 3925 3630 4005 3638
rect 3925 3628 3944 3630
rect 3959 3628 3993 3630
rect 3925 3612 4005 3628
rect 3925 3590 3944 3612
rect 3959 3596 3989 3612
rect 4017 3606 4023 3680
rect 4026 3606 4045 3750
rect 4060 3606 4066 3750
rect 4075 3680 4088 3750
rect 4140 3746 4162 3750
rect 4133 3724 4162 3738
rect 4215 3724 4231 3738
rect 4269 3734 4275 3736
rect 4282 3734 4390 3750
rect 4397 3734 4403 3736
rect 4411 3734 4426 3750
rect 4492 3744 4511 3747
rect 4133 3722 4231 3724
rect 4258 3722 4426 3734
rect 4441 3724 4457 3738
rect 4492 3725 4514 3744
rect 4524 3738 4540 3739
rect 4523 3736 4540 3738
rect 4524 3731 4540 3736
rect 4514 3724 4520 3725
rect 4523 3724 4552 3731
rect 4441 3723 4552 3724
rect 4441 3722 4558 3723
rect 4117 3714 4168 3722
rect 4215 3714 4249 3722
rect 4117 3702 4142 3714
rect 4149 3702 4168 3714
rect 4222 3712 4249 3714
rect 4258 3712 4479 3722
rect 4514 3719 4520 3722
rect 4222 3708 4479 3712
rect 4117 3694 4168 3702
rect 4215 3694 4479 3708
rect 4523 3714 4558 3722
rect 4069 3646 4088 3680
rect 4133 3686 4162 3694
rect 4133 3680 4150 3686
rect 4133 3678 4167 3680
rect 4215 3678 4231 3694
rect 4232 3684 4440 3694
rect 4441 3684 4457 3694
rect 4505 3690 4520 3705
rect 4523 3702 4524 3714
rect 4531 3702 4558 3714
rect 4523 3694 4558 3702
rect 4523 3693 4552 3694
rect 4243 3680 4457 3684
rect 4258 3678 4457 3680
rect 4492 3680 4505 3690
rect 4523 3680 4540 3693
rect 4492 3678 4540 3680
rect 4134 3674 4167 3678
rect 4130 3672 4167 3674
rect 4130 3671 4197 3672
rect 4130 3666 4161 3671
rect 4167 3666 4197 3671
rect 4130 3662 4197 3666
rect 4103 3659 4197 3662
rect 4103 3652 4152 3659
rect 4103 3646 4133 3652
rect 4152 3647 4157 3652
rect 4069 3630 4149 3646
rect 4161 3638 4197 3659
rect 4258 3654 4447 3678
rect 4492 3677 4539 3678
rect 4505 3672 4539 3677
rect 4273 3651 4447 3654
rect 4266 3648 4447 3651
rect 4475 3671 4539 3672
rect 4069 3628 4088 3630
rect 4103 3628 4137 3630
rect 4069 3612 4149 3628
rect 4069 3606 4088 3612
rect 3785 3580 3888 3590
rect 3739 3578 3888 3580
rect 3909 3578 3944 3590
rect 3578 3576 3740 3578
rect 3590 3556 3609 3576
rect 3624 3574 3654 3576
rect 3473 3548 3514 3556
rect 3596 3552 3609 3556
rect 3661 3560 3740 3576
rect 3772 3576 3944 3578
rect 3772 3560 3851 3576
rect 3858 3574 3888 3576
rect 3436 3538 3465 3548
rect 3479 3538 3508 3548
rect 3523 3538 3553 3552
rect 3596 3538 3639 3552
rect 3661 3548 3851 3560
rect 3916 3556 3922 3576
rect 3646 3538 3676 3548
rect 3677 3538 3835 3548
rect 3839 3538 3869 3548
rect 3873 3538 3903 3552
rect 3931 3538 3944 3576
rect 4016 3590 4045 3606
rect 4059 3590 4088 3606
rect 4103 3596 4133 3612
rect 4161 3590 4167 3638
rect 4170 3632 4189 3638
rect 4204 3632 4234 3640
rect 4170 3624 4234 3632
rect 4170 3608 4250 3624
rect 4266 3617 4328 3648
rect 4344 3617 4406 3648
rect 4475 3646 4524 3671
rect 4539 3646 4569 3662
rect 4438 3632 4468 3640
rect 4475 3638 4585 3646
rect 4438 3624 4483 3632
rect 4170 3606 4189 3608
rect 4204 3606 4250 3608
rect 4170 3590 4250 3606
rect 4277 3604 4312 3617
rect 4353 3614 4390 3617
rect 4353 3612 4395 3614
rect 4282 3601 4312 3604
rect 4291 3597 4298 3601
rect 4298 3596 4299 3597
rect 4257 3590 4267 3596
rect 4016 3582 4051 3590
rect 4016 3556 4017 3582
rect 4024 3556 4051 3582
rect 3959 3538 3989 3552
rect 4016 3548 4051 3556
rect 4053 3582 4094 3590
rect 4053 3556 4068 3582
rect 4075 3556 4094 3582
rect 4158 3578 4189 3590
rect 4204 3578 4307 3590
rect 4319 3580 4345 3606
rect 4360 3601 4390 3612
rect 4422 3608 4484 3624
rect 4422 3606 4468 3608
rect 4422 3590 4484 3606
rect 4496 3590 4502 3638
rect 4505 3630 4585 3638
rect 4505 3628 4524 3630
rect 4539 3628 4573 3630
rect 4505 3612 4585 3628
rect 4505 3590 4524 3612
rect 4539 3596 4569 3612
rect 4597 3606 4603 3680
rect 4606 3606 4625 3750
rect 4640 3606 4646 3750
rect 4655 3680 4668 3750
rect 4720 3746 4742 3750
rect 4713 3724 4742 3738
rect 4795 3724 4811 3738
rect 4849 3734 4855 3736
rect 4862 3734 4970 3750
rect 4977 3734 4983 3736
rect 4991 3734 5006 3750
rect 5072 3744 5091 3747
rect 4713 3722 4811 3724
rect 4838 3722 5006 3734
rect 5021 3724 5037 3738
rect 5072 3725 5094 3744
rect 5104 3738 5120 3739
rect 5103 3736 5120 3738
rect 5104 3731 5120 3736
rect 5094 3724 5100 3725
rect 5103 3724 5132 3731
rect 5021 3723 5132 3724
rect 5021 3722 5138 3723
rect 4697 3714 4748 3722
rect 4795 3714 4829 3722
rect 4697 3702 4722 3714
rect 4729 3702 4748 3714
rect 4802 3712 4829 3714
rect 4838 3712 5059 3722
rect 5094 3719 5100 3722
rect 4802 3708 5059 3712
rect 4697 3694 4748 3702
rect 4795 3694 5059 3708
rect 5103 3714 5138 3722
rect 4649 3646 4668 3680
rect 4713 3686 4742 3694
rect 4713 3680 4730 3686
rect 4713 3678 4747 3680
rect 4795 3678 4811 3694
rect 4812 3684 5020 3694
rect 5021 3684 5037 3694
rect 5085 3690 5100 3705
rect 5103 3702 5104 3714
rect 5111 3702 5138 3714
rect 5103 3694 5138 3702
rect 5103 3693 5132 3694
rect 4823 3680 5037 3684
rect 4838 3678 5037 3680
rect 5072 3680 5085 3690
rect 5103 3680 5120 3693
rect 5072 3678 5120 3680
rect 4714 3674 4747 3678
rect 4710 3672 4747 3674
rect 4710 3671 4777 3672
rect 4710 3666 4741 3671
rect 4747 3666 4777 3671
rect 4710 3662 4777 3666
rect 4683 3659 4777 3662
rect 4683 3652 4732 3659
rect 4683 3646 4713 3652
rect 4732 3647 4737 3652
rect 4649 3630 4729 3646
rect 4741 3638 4777 3659
rect 4838 3654 5027 3678
rect 5072 3677 5119 3678
rect 5085 3672 5119 3677
rect 4853 3651 5027 3654
rect 4846 3648 5027 3651
rect 5055 3671 5119 3672
rect 4649 3628 4668 3630
rect 4683 3628 4717 3630
rect 4649 3612 4729 3628
rect 4649 3606 4668 3612
rect 4365 3580 4468 3590
rect 4319 3578 4468 3580
rect 4489 3578 4524 3590
rect 4158 3576 4320 3578
rect 4170 3556 4189 3576
rect 4204 3574 4234 3576
rect 4053 3548 4094 3556
rect 4176 3552 4189 3556
rect 4241 3560 4320 3576
rect 4352 3576 4524 3578
rect 4352 3560 4431 3576
rect 4438 3574 4468 3576
rect 4016 3538 4045 3548
rect 4059 3538 4088 3548
rect 4103 3538 4133 3552
rect 4176 3538 4219 3552
rect 4241 3548 4431 3560
rect 4496 3556 4502 3576
rect 4226 3538 4256 3548
rect 4257 3538 4415 3548
rect 4419 3538 4449 3548
rect 4453 3538 4483 3552
rect 4511 3538 4524 3576
rect 4596 3590 4625 3606
rect 4639 3590 4668 3606
rect 4683 3596 4713 3612
rect 4741 3590 4747 3638
rect 4750 3632 4769 3638
rect 4784 3632 4814 3640
rect 4750 3624 4814 3632
rect 4750 3608 4830 3624
rect 4846 3617 4908 3648
rect 4924 3617 4986 3648
rect 5055 3646 5104 3671
rect 5119 3646 5149 3662
rect 5018 3632 5048 3640
rect 5055 3638 5165 3646
rect 5018 3624 5063 3632
rect 4750 3606 4769 3608
rect 4784 3606 4830 3608
rect 4750 3590 4830 3606
rect 4857 3604 4892 3617
rect 4933 3614 4970 3617
rect 4933 3612 4975 3614
rect 4862 3601 4892 3604
rect 4871 3597 4878 3601
rect 4878 3596 4879 3597
rect 4837 3590 4847 3596
rect 4596 3582 4631 3590
rect 4596 3556 4597 3582
rect 4604 3556 4631 3582
rect 4539 3538 4569 3552
rect 4596 3548 4631 3556
rect 4633 3582 4674 3590
rect 4633 3556 4648 3582
rect 4655 3556 4674 3582
rect 4738 3578 4769 3590
rect 4784 3578 4887 3590
rect 4899 3580 4925 3606
rect 4940 3601 4970 3612
rect 5002 3608 5064 3624
rect 5002 3606 5048 3608
rect 5002 3590 5064 3606
rect 5076 3590 5082 3638
rect 5085 3630 5165 3638
rect 5085 3628 5104 3630
rect 5119 3628 5153 3630
rect 5085 3612 5165 3628
rect 5085 3590 5104 3612
rect 5119 3596 5149 3612
rect 5177 3606 5183 3680
rect 5186 3606 5205 3750
rect 5220 3606 5226 3750
rect 5235 3680 5248 3750
rect 5300 3746 5322 3750
rect 5293 3724 5322 3738
rect 5375 3724 5391 3738
rect 5429 3734 5435 3736
rect 5442 3734 5550 3750
rect 5557 3734 5563 3736
rect 5571 3734 5586 3750
rect 5652 3744 5671 3747
rect 5293 3722 5391 3724
rect 5418 3722 5586 3734
rect 5601 3724 5617 3738
rect 5652 3725 5674 3744
rect 5684 3738 5700 3739
rect 5683 3736 5700 3738
rect 5684 3731 5700 3736
rect 5674 3724 5680 3725
rect 5683 3724 5712 3731
rect 5601 3723 5712 3724
rect 5601 3722 5718 3723
rect 5277 3714 5328 3722
rect 5375 3714 5409 3722
rect 5277 3702 5302 3714
rect 5309 3702 5328 3714
rect 5382 3712 5409 3714
rect 5418 3712 5639 3722
rect 5674 3719 5680 3722
rect 5382 3708 5639 3712
rect 5277 3694 5328 3702
rect 5375 3694 5639 3708
rect 5683 3714 5718 3722
rect 5229 3646 5248 3680
rect 5293 3686 5322 3694
rect 5293 3680 5310 3686
rect 5293 3678 5327 3680
rect 5375 3678 5391 3694
rect 5392 3684 5600 3694
rect 5601 3684 5617 3694
rect 5665 3690 5680 3705
rect 5683 3702 5684 3714
rect 5691 3702 5718 3714
rect 5683 3694 5718 3702
rect 5683 3693 5712 3694
rect 5403 3680 5617 3684
rect 5418 3678 5617 3680
rect 5652 3680 5665 3690
rect 5683 3680 5700 3693
rect 5652 3678 5700 3680
rect 5294 3674 5327 3678
rect 5290 3672 5327 3674
rect 5290 3671 5357 3672
rect 5290 3666 5321 3671
rect 5327 3666 5357 3671
rect 5290 3662 5357 3666
rect 5263 3659 5357 3662
rect 5263 3652 5312 3659
rect 5263 3646 5293 3652
rect 5312 3647 5317 3652
rect 5229 3630 5309 3646
rect 5321 3638 5357 3659
rect 5418 3654 5607 3678
rect 5652 3677 5699 3678
rect 5665 3672 5699 3677
rect 5433 3651 5607 3654
rect 5426 3648 5607 3651
rect 5635 3671 5699 3672
rect 5229 3628 5248 3630
rect 5263 3628 5297 3630
rect 5229 3612 5309 3628
rect 5229 3606 5248 3612
rect 4945 3580 5048 3590
rect 4899 3578 5048 3580
rect 5069 3578 5104 3590
rect 4738 3576 4900 3578
rect 4750 3556 4769 3576
rect 4784 3574 4814 3576
rect 4633 3548 4674 3556
rect 4756 3552 4769 3556
rect 4821 3560 4900 3576
rect 4932 3576 5104 3578
rect 4932 3560 5011 3576
rect 5018 3574 5048 3576
rect 4596 3538 4625 3548
rect 4639 3538 4668 3548
rect 4683 3538 4713 3552
rect 4756 3538 4799 3552
rect 4821 3548 5011 3560
rect 5076 3556 5082 3576
rect 4806 3538 4836 3548
rect 4837 3538 4995 3548
rect 4999 3538 5029 3548
rect 5033 3538 5063 3552
rect 5091 3538 5104 3576
rect 5176 3590 5205 3606
rect 5219 3590 5248 3606
rect 5263 3596 5293 3612
rect 5321 3590 5327 3638
rect 5330 3632 5349 3638
rect 5364 3632 5394 3640
rect 5330 3624 5394 3632
rect 5330 3608 5410 3624
rect 5426 3617 5488 3648
rect 5504 3617 5566 3648
rect 5635 3646 5684 3671
rect 5699 3646 5729 3662
rect 5598 3632 5628 3640
rect 5635 3638 5745 3646
rect 5598 3624 5643 3632
rect 5330 3606 5349 3608
rect 5364 3606 5410 3608
rect 5330 3590 5410 3606
rect 5437 3604 5472 3617
rect 5513 3614 5550 3617
rect 5513 3612 5555 3614
rect 5442 3601 5472 3604
rect 5451 3597 5458 3601
rect 5458 3596 5459 3597
rect 5417 3590 5427 3596
rect 5176 3582 5211 3590
rect 5176 3556 5177 3582
rect 5184 3556 5211 3582
rect 5119 3538 5149 3552
rect 5176 3548 5211 3556
rect 5213 3582 5254 3590
rect 5213 3556 5228 3582
rect 5235 3556 5254 3582
rect 5318 3578 5349 3590
rect 5364 3578 5467 3590
rect 5479 3580 5505 3606
rect 5520 3601 5550 3612
rect 5582 3608 5644 3624
rect 5582 3606 5628 3608
rect 5582 3590 5644 3606
rect 5656 3590 5662 3638
rect 5665 3630 5745 3638
rect 5665 3628 5684 3630
rect 5699 3628 5733 3630
rect 5665 3612 5745 3628
rect 5665 3590 5684 3612
rect 5699 3596 5729 3612
rect 5757 3606 5763 3680
rect 5766 3606 5785 3750
rect 5800 3606 5806 3750
rect 5815 3680 5828 3750
rect 5880 3746 5902 3750
rect 5873 3724 5902 3738
rect 5955 3724 5971 3738
rect 6009 3734 6015 3736
rect 6022 3734 6130 3750
rect 6137 3734 6143 3736
rect 6151 3734 6166 3750
rect 6232 3744 6251 3747
rect 5873 3722 5971 3724
rect 5998 3722 6166 3734
rect 6181 3724 6197 3738
rect 6232 3725 6254 3744
rect 6264 3738 6280 3739
rect 6263 3736 6280 3738
rect 6264 3731 6280 3736
rect 6254 3724 6260 3725
rect 6263 3724 6292 3731
rect 6181 3723 6292 3724
rect 6181 3722 6298 3723
rect 5857 3714 5908 3722
rect 5955 3714 5989 3722
rect 5857 3702 5882 3714
rect 5889 3702 5908 3714
rect 5962 3712 5989 3714
rect 5998 3712 6219 3722
rect 6254 3719 6260 3722
rect 5962 3708 6219 3712
rect 5857 3694 5908 3702
rect 5955 3694 6219 3708
rect 6263 3714 6298 3722
rect 5809 3646 5828 3680
rect 5873 3686 5902 3694
rect 5873 3680 5890 3686
rect 5873 3678 5907 3680
rect 5955 3678 5971 3694
rect 5972 3684 6180 3694
rect 6181 3684 6197 3694
rect 6245 3690 6260 3705
rect 6263 3702 6264 3714
rect 6271 3702 6298 3714
rect 6263 3694 6298 3702
rect 6263 3693 6292 3694
rect 5983 3680 6197 3684
rect 5998 3678 6197 3680
rect 6232 3680 6245 3690
rect 6263 3680 6280 3693
rect 6232 3678 6280 3680
rect 5874 3674 5907 3678
rect 5870 3672 5907 3674
rect 5870 3671 5937 3672
rect 5870 3666 5901 3671
rect 5907 3666 5937 3671
rect 5870 3662 5937 3666
rect 5843 3659 5937 3662
rect 5843 3652 5892 3659
rect 5843 3646 5873 3652
rect 5892 3647 5897 3652
rect 5809 3630 5889 3646
rect 5901 3638 5937 3659
rect 5998 3654 6187 3678
rect 6232 3677 6279 3678
rect 6245 3672 6279 3677
rect 6013 3651 6187 3654
rect 6006 3648 6187 3651
rect 6215 3671 6279 3672
rect 5809 3628 5828 3630
rect 5843 3628 5877 3630
rect 5809 3612 5889 3628
rect 5809 3606 5828 3612
rect 5525 3580 5628 3590
rect 5479 3578 5628 3580
rect 5649 3578 5684 3590
rect 5318 3576 5480 3578
rect 5330 3556 5349 3576
rect 5364 3574 5394 3576
rect 5213 3548 5254 3556
rect 5336 3552 5349 3556
rect 5401 3560 5480 3576
rect 5512 3576 5684 3578
rect 5512 3560 5591 3576
rect 5598 3574 5628 3576
rect 5176 3538 5205 3548
rect 5219 3538 5248 3548
rect 5263 3538 5293 3552
rect 5336 3538 5379 3552
rect 5401 3548 5591 3560
rect 5656 3556 5662 3576
rect 5386 3538 5416 3548
rect 5417 3538 5575 3548
rect 5579 3538 5609 3548
rect 5613 3538 5643 3552
rect 5671 3538 5684 3576
rect 5756 3590 5785 3606
rect 5799 3590 5828 3606
rect 5843 3596 5873 3612
rect 5901 3590 5907 3638
rect 5910 3632 5929 3638
rect 5944 3632 5974 3640
rect 5910 3624 5974 3632
rect 5910 3608 5990 3624
rect 6006 3617 6068 3648
rect 6084 3617 6146 3648
rect 6215 3646 6264 3671
rect 6279 3646 6309 3662
rect 6178 3632 6208 3640
rect 6215 3638 6325 3646
rect 6178 3624 6223 3632
rect 5910 3606 5929 3608
rect 5944 3606 5990 3608
rect 5910 3590 5990 3606
rect 6017 3604 6052 3617
rect 6093 3614 6130 3617
rect 6093 3612 6135 3614
rect 6022 3601 6052 3604
rect 6031 3597 6038 3601
rect 6038 3596 6039 3597
rect 5997 3590 6007 3596
rect 5756 3582 5791 3590
rect 5756 3556 5757 3582
rect 5764 3556 5791 3582
rect 5699 3538 5729 3552
rect 5756 3548 5791 3556
rect 5793 3582 5834 3590
rect 5793 3556 5808 3582
rect 5815 3556 5834 3582
rect 5898 3578 5929 3590
rect 5944 3578 6047 3590
rect 6059 3580 6085 3606
rect 6100 3601 6130 3612
rect 6162 3608 6224 3624
rect 6162 3606 6208 3608
rect 6162 3590 6224 3606
rect 6236 3590 6242 3638
rect 6245 3630 6325 3638
rect 6245 3628 6264 3630
rect 6279 3628 6313 3630
rect 6245 3612 6325 3628
rect 6245 3590 6264 3612
rect 6279 3596 6309 3612
rect 6337 3606 6343 3680
rect 6346 3606 6365 3750
rect 6380 3606 6386 3750
rect 6395 3680 6408 3750
rect 6460 3746 6482 3750
rect 6453 3724 6482 3738
rect 6535 3724 6551 3738
rect 6589 3734 6595 3736
rect 6602 3734 6710 3750
rect 6717 3734 6723 3736
rect 6731 3734 6746 3750
rect 6812 3744 6831 3747
rect 6453 3722 6551 3724
rect 6578 3722 6746 3734
rect 6761 3724 6777 3738
rect 6812 3725 6834 3744
rect 6844 3738 6860 3739
rect 6843 3736 6860 3738
rect 6844 3731 6860 3736
rect 6834 3724 6840 3725
rect 6843 3724 6872 3731
rect 6761 3723 6872 3724
rect 6761 3722 6878 3723
rect 6437 3714 6488 3722
rect 6535 3714 6569 3722
rect 6437 3702 6462 3714
rect 6469 3702 6488 3714
rect 6542 3712 6569 3714
rect 6578 3712 6799 3722
rect 6834 3719 6840 3722
rect 6542 3708 6799 3712
rect 6437 3694 6488 3702
rect 6535 3694 6799 3708
rect 6843 3714 6878 3722
rect 6389 3646 6408 3680
rect 6453 3686 6482 3694
rect 6453 3680 6470 3686
rect 6453 3678 6487 3680
rect 6535 3678 6551 3694
rect 6552 3684 6760 3694
rect 6761 3684 6777 3694
rect 6825 3690 6840 3705
rect 6843 3702 6844 3714
rect 6851 3702 6878 3714
rect 6843 3694 6878 3702
rect 6843 3693 6872 3694
rect 6563 3680 6777 3684
rect 6578 3678 6777 3680
rect 6812 3680 6825 3690
rect 6843 3680 6860 3693
rect 6812 3678 6860 3680
rect 6454 3674 6487 3678
rect 6450 3672 6487 3674
rect 6450 3671 6517 3672
rect 6450 3666 6481 3671
rect 6487 3666 6517 3671
rect 6450 3662 6517 3666
rect 6423 3659 6517 3662
rect 6423 3652 6472 3659
rect 6423 3646 6453 3652
rect 6472 3647 6477 3652
rect 6389 3630 6469 3646
rect 6481 3638 6517 3659
rect 6578 3654 6767 3678
rect 6812 3677 6859 3678
rect 6825 3672 6859 3677
rect 6593 3651 6767 3654
rect 6586 3648 6767 3651
rect 6795 3671 6859 3672
rect 6389 3628 6408 3630
rect 6423 3628 6457 3630
rect 6389 3612 6469 3628
rect 6389 3606 6408 3612
rect 6105 3580 6208 3590
rect 6059 3578 6208 3580
rect 6229 3578 6264 3590
rect 5898 3576 6060 3578
rect 5910 3556 5929 3576
rect 5944 3574 5974 3576
rect 5793 3548 5834 3556
rect 5916 3552 5929 3556
rect 5981 3560 6060 3576
rect 6092 3576 6264 3578
rect 6092 3560 6171 3576
rect 6178 3574 6208 3576
rect 5756 3538 5785 3548
rect 5799 3538 5828 3548
rect 5843 3538 5873 3552
rect 5916 3538 5959 3552
rect 5981 3548 6171 3560
rect 6236 3556 6242 3576
rect 5966 3538 5996 3548
rect 5997 3538 6155 3548
rect 6159 3538 6189 3548
rect 6193 3538 6223 3552
rect 6251 3538 6264 3576
rect 6336 3590 6365 3606
rect 6379 3590 6408 3606
rect 6423 3596 6453 3612
rect 6481 3590 6487 3638
rect 6490 3632 6509 3638
rect 6524 3632 6554 3640
rect 6490 3624 6554 3632
rect 6490 3608 6570 3624
rect 6586 3617 6648 3648
rect 6664 3617 6726 3648
rect 6795 3646 6844 3671
rect 6859 3646 6889 3662
rect 6758 3632 6788 3640
rect 6795 3638 6905 3646
rect 6758 3624 6803 3632
rect 6490 3606 6509 3608
rect 6524 3606 6570 3608
rect 6490 3590 6570 3606
rect 6597 3604 6632 3617
rect 6673 3614 6710 3617
rect 6673 3612 6715 3614
rect 6602 3601 6632 3604
rect 6611 3597 6618 3601
rect 6618 3596 6619 3597
rect 6577 3590 6587 3596
rect 6336 3582 6371 3590
rect 6336 3556 6337 3582
rect 6344 3556 6371 3582
rect 6279 3538 6309 3552
rect 6336 3548 6371 3556
rect 6373 3582 6414 3590
rect 6373 3556 6388 3582
rect 6395 3556 6414 3582
rect 6478 3578 6509 3590
rect 6524 3578 6627 3590
rect 6639 3580 6665 3606
rect 6680 3601 6710 3612
rect 6742 3608 6804 3624
rect 6742 3606 6788 3608
rect 6742 3590 6804 3606
rect 6816 3590 6822 3638
rect 6825 3630 6905 3638
rect 6825 3628 6844 3630
rect 6859 3628 6893 3630
rect 6825 3612 6905 3628
rect 6825 3590 6844 3612
rect 6859 3596 6889 3612
rect 6917 3606 6923 3680
rect 6926 3606 6945 3750
rect 6960 3606 6966 3750
rect 6975 3680 6988 3750
rect 7040 3746 7062 3750
rect 7033 3724 7062 3738
rect 7115 3724 7131 3738
rect 7169 3734 7175 3736
rect 7182 3734 7290 3750
rect 7297 3734 7303 3736
rect 7311 3734 7326 3750
rect 7392 3744 7411 3747
rect 7033 3722 7131 3724
rect 7158 3722 7326 3734
rect 7341 3724 7357 3738
rect 7392 3725 7414 3744
rect 7424 3738 7440 3739
rect 7423 3736 7440 3738
rect 7424 3731 7440 3736
rect 7414 3724 7420 3725
rect 7423 3724 7452 3731
rect 7341 3723 7452 3724
rect 7341 3722 7458 3723
rect 7017 3714 7068 3722
rect 7115 3714 7149 3722
rect 7017 3702 7042 3714
rect 7049 3702 7068 3714
rect 7122 3712 7149 3714
rect 7158 3712 7379 3722
rect 7414 3719 7420 3722
rect 7122 3708 7379 3712
rect 7017 3694 7068 3702
rect 7115 3694 7379 3708
rect 7423 3714 7458 3722
rect 6969 3646 6988 3680
rect 7033 3686 7062 3694
rect 7033 3680 7050 3686
rect 7033 3678 7067 3680
rect 7115 3678 7131 3694
rect 7132 3684 7340 3694
rect 7341 3684 7357 3694
rect 7405 3690 7420 3705
rect 7423 3702 7424 3714
rect 7431 3702 7458 3714
rect 7423 3694 7458 3702
rect 7423 3693 7452 3694
rect 7143 3680 7357 3684
rect 7158 3678 7357 3680
rect 7392 3680 7405 3690
rect 7423 3680 7440 3693
rect 7392 3678 7440 3680
rect 7034 3674 7067 3678
rect 7030 3672 7067 3674
rect 7030 3671 7097 3672
rect 7030 3666 7061 3671
rect 7067 3666 7097 3671
rect 7030 3662 7097 3666
rect 7003 3659 7097 3662
rect 7003 3652 7052 3659
rect 7003 3646 7033 3652
rect 7052 3647 7057 3652
rect 6969 3630 7049 3646
rect 7061 3638 7097 3659
rect 7158 3654 7347 3678
rect 7392 3677 7439 3678
rect 7405 3672 7439 3677
rect 7173 3651 7347 3654
rect 7166 3648 7347 3651
rect 7375 3671 7439 3672
rect 6969 3628 6988 3630
rect 7003 3628 7037 3630
rect 6969 3612 7049 3628
rect 6969 3606 6988 3612
rect 6685 3580 6788 3590
rect 6639 3578 6788 3580
rect 6809 3578 6844 3590
rect 6478 3576 6640 3578
rect 6490 3556 6509 3576
rect 6524 3574 6554 3576
rect 6373 3548 6414 3556
rect 6496 3552 6509 3556
rect 6561 3560 6640 3576
rect 6672 3576 6844 3578
rect 6672 3560 6751 3576
rect 6758 3574 6788 3576
rect 6336 3538 6365 3548
rect 6379 3538 6408 3548
rect 6423 3538 6453 3552
rect 6496 3538 6539 3552
rect 6561 3548 6751 3560
rect 6816 3556 6822 3576
rect 6546 3538 6576 3548
rect 6577 3538 6735 3548
rect 6739 3538 6769 3548
rect 6773 3538 6803 3552
rect 6831 3538 6844 3576
rect 6916 3590 6945 3606
rect 6959 3590 6988 3606
rect 7003 3596 7033 3612
rect 7061 3590 7067 3638
rect 7070 3632 7089 3638
rect 7104 3632 7134 3640
rect 7070 3624 7134 3632
rect 7070 3608 7150 3624
rect 7166 3617 7228 3648
rect 7244 3617 7306 3648
rect 7375 3646 7424 3671
rect 7439 3646 7469 3662
rect 7338 3632 7368 3640
rect 7375 3638 7485 3646
rect 7338 3624 7383 3632
rect 7070 3606 7089 3608
rect 7104 3606 7150 3608
rect 7070 3590 7150 3606
rect 7177 3604 7212 3617
rect 7253 3614 7290 3617
rect 7253 3612 7295 3614
rect 7182 3601 7212 3604
rect 7191 3597 7198 3601
rect 7198 3596 7199 3597
rect 7157 3590 7167 3596
rect 6916 3582 6951 3590
rect 6916 3556 6917 3582
rect 6924 3556 6951 3582
rect 6859 3538 6889 3552
rect 6916 3548 6951 3556
rect 6953 3582 6994 3590
rect 6953 3556 6968 3582
rect 6975 3556 6994 3582
rect 7058 3578 7089 3590
rect 7104 3578 7207 3590
rect 7219 3580 7245 3606
rect 7260 3601 7290 3612
rect 7322 3608 7384 3624
rect 7322 3606 7368 3608
rect 7322 3590 7384 3606
rect 7396 3590 7402 3638
rect 7405 3630 7485 3638
rect 7405 3628 7424 3630
rect 7439 3628 7473 3630
rect 7405 3612 7485 3628
rect 7405 3590 7424 3612
rect 7439 3596 7469 3612
rect 7497 3606 7503 3680
rect 7506 3606 7525 3750
rect 7540 3606 7546 3750
rect 7555 3680 7568 3750
rect 7620 3746 7642 3750
rect 7613 3724 7642 3738
rect 7695 3724 7711 3738
rect 7749 3734 7755 3736
rect 7762 3734 7870 3750
rect 7877 3734 7883 3736
rect 7891 3734 7906 3750
rect 7972 3744 7991 3747
rect 7613 3722 7711 3724
rect 7738 3722 7906 3734
rect 7921 3724 7937 3738
rect 7972 3725 7994 3744
rect 8004 3738 8020 3739
rect 8003 3736 8020 3738
rect 8004 3731 8020 3736
rect 7994 3724 8000 3725
rect 8003 3724 8032 3731
rect 7921 3723 8032 3724
rect 7921 3722 8038 3723
rect 7597 3714 7648 3722
rect 7695 3714 7729 3722
rect 7597 3702 7622 3714
rect 7629 3702 7648 3714
rect 7702 3712 7729 3714
rect 7738 3712 7959 3722
rect 7994 3719 8000 3722
rect 7702 3708 7959 3712
rect 7597 3694 7648 3702
rect 7695 3694 7959 3708
rect 8003 3714 8038 3722
rect 7549 3646 7568 3680
rect 7613 3686 7642 3694
rect 7613 3680 7630 3686
rect 7613 3678 7647 3680
rect 7695 3678 7711 3694
rect 7712 3684 7920 3694
rect 7921 3684 7937 3694
rect 7985 3690 8000 3705
rect 8003 3702 8004 3714
rect 8011 3702 8038 3714
rect 8003 3694 8038 3702
rect 8003 3693 8032 3694
rect 7723 3680 7937 3684
rect 7738 3678 7937 3680
rect 7972 3680 7985 3690
rect 8003 3680 8020 3693
rect 7972 3678 8020 3680
rect 7614 3674 7647 3678
rect 7610 3672 7647 3674
rect 7610 3671 7677 3672
rect 7610 3666 7641 3671
rect 7647 3666 7677 3671
rect 7610 3662 7677 3666
rect 7583 3659 7677 3662
rect 7583 3652 7632 3659
rect 7583 3646 7613 3652
rect 7632 3647 7637 3652
rect 7549 3630 7629 3646
rect 7641 3638 7677 3659
rect 7738 3654 7927 3678
rect 7972 3677 8019 3678
rect 7985 3672 8019 3677
rect 7753 3651 7927 3654
rect 7746 3648 7927 3651
rect 7955 3671 8019 3672
rect 7549 3628 7568 3630
rect 7583 3628 7617 3630
rect 7549 3612 7629 3628
rect 7549 3606 7568 3612
rect 7265 3580 7368 3590
rect 7219 3578 7368 3580
rect 7389 3578 7424 3590
rect 7058 3576 7220 3578
rect 7070 3556 7089 3576
rect 7104 3574 7134 3576
rect 6953 3548 6994 3556
rect 7076 3552 7089 3556
rect 7141 3560 7220 3576
rect 7252 3576 7424 3578
rect 7252 3560 7331 3576
rect 7338 3574 7368 3576
rect 6916 3538 6945 3548
rect 6959 3538 6988 3548
rect 7003 3538 7033 3552
rect 7076 3538 7119 3552
rect 7141 3548 7331 3560
rect 7396 3556 7402 3576
rect 7126 3538 7156 3548
rect 7157 3538 7315 3548
rect 7319 3538 7349 3548
rect 7353 3538 7383 3552
rect 7411 3538 7424 3576
rect 7496 3590 7525 3606
rect 7539 3590 7568 3606
rect 7583 3596 7613 3612
rect 7641 3590 7647 3638
rect 7650 3632 7669 3638
rect 7684 3632 7714 3640
rect 7650 3624 7714 3632
rect 7650 3608 7730 3624
rect 7746 3617 7808 3648
rect 7824 3617 7886 3648
rect 7955 3646 8004 3671
rect 8019 3646 8049 3662
rect 7918 3632 7948 3640
rect 7955 3638 8065 3646
rect 7918 3624 7963 3632
rect 7650 3606 7669 3608
rect 7684 3606 7730 3608
rect 7650 3590 7730 3606
rect 7757 3604 7792 3617
rect 7833 3614 7870 3617
rect 7833 3612 7875 3614
rect 7762 3601 7792 3604
rect 7771 3597 7778 3601
rect 7778 3596 7779 3597
rect 7737 3590 7747 3596
rect 7496 3582 7531 3590
rect 7496 3556 7497 3582
rect 7504 3556 7531 3582
rect 7439 3538 7469 3552
rect 7496 3548 7531 3556
rect 7533 3582 7574 3590
rect 7533 3556 7548 3582
rect 7555 3556 7574 3582
rect 7638 3578 7669 3590
rect 7684 3578 7787 3590
rect 7799 3580 7825 3606
rect 7840 3601 7870 3612
rect 7902 3608 7964 3624
rect 7902 3606 7948 3608
rect 7902 3590 7964 3606
rect 7976 3590 7982 3638
rect 7985 3630 8065 3638
rect 7985 3628 8004 3630
rect 8019 3628 8053 3630
rect 7985 3612 8065 3628
rect 7985 3590 8004 3612
rect 8019 3596 8049 3612
rect 8077 3606 8083 3680
rect 8086 3606 8105 3750
rect 8120 3606 8126 3750
rect 8135 3680 8148 3750
rect 8200 3746 8222 3750
rect 8193 3724 8222 3738
rect 8275 3724 8291 3738
rect 8329 3734 8335 3736
rect 8342 3734 8450 3750
rect 8457 3734 8463 3736
rect 8471 3734 8486 3750
rect 8552 3744 8571 3747
rect 8193 3722 8291 3724
rect 8318 3722 8486 3734
rect 8501 3724 8517 3738
rect 8552 3725 8574 3744
rect 8584 3738 8600 3739
rect 8583 3736 8600 3738
rect 8584 3731 8600 3736
rect 8574 3724 8580 3725
rect 8583 3724 8612 3731
rect 8501 3723 8612 3724
rect 8501 3722 8618 3723
rect 8177 3714 8228 3722
rect 8275 3714 8309 3722
rect 8177 3702 8202 3714
rect 8209 3702 8228 3714
rect 8282 3712 8309 3714
rect 8318 3712 8539 3722
rect 8574 3719 8580 3722
rect 8282 3708 8539 3712
rect 8177 3694 8228 3702
rect 8275 3694 8539 3708
rect 8583 3714 8618 3722
rect 8129 3646 8148 3680
rect 8193 3686 8222 3694
rect 8193 3680 8210 3686
rect 8193 3678 8227 3680
rect 8275 3678 8291 3694
rect 8292 3684 8500 3694
rect 8501 3684 8517 3694
rect 8565 3690 8580 3705
rect 8583 3702 8584 3714
rect 8591 3702 8618 3714
rect 8583 3694 8618 3702
rect 8583 3693 8612 3694
rect 8303 3680 8517 3684
rect 8318 3678 8517 3680
rect 8552 3680 8565 3690
rect 8583 3680 8600 3693
rect 8552 3678 8600 3680
rect 8194 3674 8227 3678
rect 8190 3672 8227 3674
rect 8190 3671 8257 3672
rect 8190 3666 8221 3671
rect 8227 3666 8257 3671
rect 8190 3662 8257 3666
rect 8163 3659 8257 3662
rect 8163 3652 8212 3659
rect 8163 3646 8193 3652
rect 8212 3647 8217 3652
rect 8129 3630 8209 3646
rect 8221 3638 8257 3659
rect 8318 3654 8507 3678
rect 8552 3677 8599 3678
rect 8565 3672 8599 3677
rect 8333 3651 8507 3654
rect 8326 3648 8507 3651
rect 8535 3671 8599 3672
rect 8129 3628 8148 3630
rect 8163 3628 8197 3630
rect 8129 3612 8209 3628
rect 8129 3606 8148 3612
rect 7845 3580 7948 3590
rect 7799 3578 7948 3580
rect 7969 3578 8004 3590
rect 7638 3576 7800 3578
rect 7650 3556 7669 3576
rect 7684 3574 7714 3576
rect 7533 3548 7574 3556
rect 7656 3552 7669 3556
rect 7721 3560 7800 3576
rect 7832 3576 8004 3578
rect 7832 3560 7911 3576
rect 7918 3574 7948 3576
rect 7496 3538 7525 3548
rect 7539 3538 7568 3548
rect 7583 3538 7613 3552
rect 7656 3538 7699 3552
rect 7721 3548 7911 3560
rect 7976 3556 7982 3576
rect 7706 3538 7736 3548
rect 7737 3538 7895 3548
rect 7899 3538 7929 3548
rect 7933 3538 7963 3552
rect 7991 3538 8004 3576
rect 8076 3590 8105 3606
rect 8119 3590 8148 3606
rect 8163 3596 8193 3612
rect 8221 3590 8227 3638
rect 8230 3632 8249 3638
rect 8264 3632 8294 3640
rect 8230 3624 8294 3632
rect 8230 3608 8310 3624
rect 8326 3617 8388 3648
rect 8404 3617 8466 3648
rect 8535 3646 8584 3671
rect 8599 3646 8629 3662
rect 8498 3632 8528 3640
rect 8535 3638 8645 3646
rect 8498 3624 8543 3632
rect 8230 3606 8249 3608
rect 8264 3606 8310 3608
rect 8230 3590 8310 3606
rect 8337 3604 8372 3617
rect 8413 3614 8450 3617
rect 8413 3612 8455 3614
rect 8342 3601 8372 3604
rect 8351 3597 8358 3601
rect 8358 3596 8359 3597
rect 8317 3590 8327 3596
rect 8076 3582 8111 3590
rect 8076 3556 8077 3582
rect 8084 3556 8111 3582
rect 8019 3538 8049 3552
rect 8076 3548 8111 3556
rect 8113 3582 8154 3590
rect 8113 3556 8128 3582
rect 8135 3556 8154 3582
rect 8218 3578 8249 3590
rect 8264 3578 8367 3590
rect 8379 3580 8405 3606
rect 8420 3601 8450 3612
rect 8482 3608 8544 3624
rect 8482 3606 8528 3608
rect 8482 3590 8544 3606
rect 8556 3590 8562 3638
rect 8565 3630 8645 3638
rect 8565 3628 8584 3630
rect 8599 3628 8633 3630
rect 8565 3612 8645 3628
rect 8565 3590 8584 3612
rect 8599 3596 8629 3612
rect 8657 3606 8663 3680
rect 8666 3606 8685 3750
rect 8700 3606 8706 3750
rect 8715 3680 8728 3750
rect 8780 3746 8802 3750
rect 8773 3724 8802 3738
rect 8855 3724 8871 3738
rect 8909 3734 8915 3736
rect 8922 3734 9030 3750
rect 9037 3734 9043 3736
rect 9051 3734 9066 3750
rect 9132 3744 9151 3747
rect 8773 3722 8871 3724
rect 8898 3722 9066 3734
rect 9081 3724 9097 3738
rect 9132 3725 9154 3744
rect 9164 3738 9180 3739
rect 9163 3736 9180 3738
rect 9164 3731 9180 3736
rect 9154 3724 9160 3725
rect 9163 3724 9192 3731
rect 9081 3723 9192 3724
rect 9081 3722 9198 3723
rect 8757 3714 8808 3722
rect 8855 3714 8889 3722
rect 8757 3702 8782 3714
rect 8789 3702 8808 3714
rect 8862 3712 8889 3714
rect 8898 3712 9119 3722
rect 9154 3719 9160 3722
rect 8862 3708 9119 3712
rect 8757 3694 8808 3702
rect 8855 3694 9119 3708
rect 9163 3714 9198 3722
rect 8709 3646 8728 3680
rect 8773 3686 8802 3694
rect 8773 3680 8790 3686
rect 8773 3678 8807 3680
rect 8855 3678 8871 3694
rect 8872 3684 9080 3694
rect 9081 3684 9097 3694
rect 9145 3690 9160 3705
rect 9163 3702 9164 3714
rect 9171 3702 9198 3714
rect 9163 3694 9198 3702
rect 9163 3693 9192 3694
rect 8883 3680 9097 3684
rect 8898 3678 9097 3680
rect 9132 3680 9145 3690
rect 9163 3680 9180 3693
rect 9132 3678 9180 3680
rect 8774 3674 8807 3678
rect 8770 3672 8807 3674
rect 8770 3671 8837 3672
rect 8770 3666 8801 3671
rect 8807 3666 8837 3671
rect 8770 3662 8837 3666
rect 8743 3659 8837 3662
rect 8743 3652 8792 3659
rect 8743 3646 8773 3652
rect 8792 3647 8797 3652
rect 8709 3630 8789 3646
rect 8801 3638 8837 3659
rect 8898 3654 9087 3678
rect 9132 3677 9179 3678
rect 9145 3672 9179 3677
rect 8913 3651 9087 3654
rect 8906 3648 9087 3651
rect 9115 3671 9179 3672
rect 8709 3628 8728 3630
rect 8743 3628 8777 3630
rect 8709 3612 8789 3628
rect 8709 3606 8728 3612
rect 8425 3580 8528 3590
rect 8379 3578 8528 3580
rect 8549 3578 8584 3590
rect 8218 3576 8380 3578
rect 8230 3556 8249 3576
rect 8264 3574 8294 3576
rect 8113 3548 8154 3556
rect 8236 3552 8249 3556
rect 8301 3560 8380 3576
rect 8412 3576 8584 3578
rect 8412 3560 8491 3576
rect 8498 3574 8528 3576
rect 8076 3538 8105 3548
rect 8119 3538 8148 3548
rect 8163 3538 8193 3552
rect 8236 3538 8279 3552
rect 8301 3548 8491 3560
rect 8556 3556 8562 3576
rect 8286 3538 8316 3548
rect 8317 3538 8475 3548
rect 8479 3538 8509 3548
rect 8513 3538 8543 3552
rect 8571 3538 8584 3576
rect 8656 3590 8685 3606
rect 8699 3590 8728 3606
rect 8743 3596 8773 3612
rect 8801 3590 8807 3638
rect 8810 3632 8829 3638
rect 8844 3632 8874 3640
rect 8810 3624 8874 3632
rect 8810 3608 8890 3624
rect 8906 3617 8968 3648
rect 8984 3617 9046 3648
rect 9115 3646 9164 3671
rect 9179 3646 9209 3662
rect 9078 3632 9108 3640
rect 9115 3638 9225 3646
rect 9078 3624 9123 3632
rect 8810 3606 8829 3608
rect 8844 3606 8890 3608
rect 8810 3590 8890 3606
rect 8917 3604 8952 3617
rect 8993 3614 9030 3617
rect 8993 3612 9035 3614
rect 8922 3601 8952 3604
rect 8931 3597 8938 3601
rect 8938 3596 8939 3597
rect 8897 3590 8907 3596
rect 8656 3582 8691 3590
rect 8656 3556 8657 3582
rect 8664 3556 8691 3582
rect 8599 3538 8629 3552
rect 8656 3548 8691 3556
rect 8693 3582 8734 3590
rect 8693 3556 8708 3582
rect 8715 3556 8734 3582
rect 8798 3578 8829 3590
rect 8844 3578 8947 3590
rect 8959 3580 8985 3606
rect 9000 3601 9030 3612
rect 9062 3608 9124 3624
rect 9062 3606 9108 3608
rect 9062 3590 9124 3606
rect 9136 3590 9142 3638
rect 9145 3630 9225 3638
rect 9145 3628 9164 3630
rect 9179 3628 9213 3630
rect 9145 3612 9225 3628
rect 9145 3590 9164 3612
rect 9179 3596 9209 3612
rect 9237 3606 9243 3680
rect 9246 3606 9265 3750
rect 9280 3606 9286 3750
rect 9295 3680 9308 3750
rect 9360 3746 9382 3750
rect 9353 3724 9382 3738
rect 9435 3724 9451 3738
rect 9489 3734 9495 3736
rect 9502 3734 9610 3750
rect 9617 3734 9623 3736
rect 9631 3734 9646 3750
rect 9712 3744 9731 3747
rect 9353 3722 9451 3724
rect 9478 3722 9646 3734
rect 9661 3724 9677 3738
rect 9712 3725 9734 3744
rect 9744 3738 9760 3739
rect 9743 3736 9760 3738
rect 9744 3731 9760 3736
rect 9734 3724 9740 3725
rect 9743 3724 9772 3731
rect 9661 3723 9772 3724
rect 9661 3722 9778 3723
rect 9337 3714 9388 3722
rect 9435 3714 9469 3722
rect 9337 3702 9362 3714
rect 9369 3702 9388 3714
rect 9442 3712 9469 3714
rect 9478 3712 9699 3722
rect 9734 3719 9740 3722
rect 9442 3708 9699 3712
rect 9337 3694 9388 3702
rect 9435 3694 9699 3708
rect 9743 3714 9778 3722
rect 9289 3646 9308 3680
rect 9353 3686 9382 3694
rect 9353 3680 9370 3686
rect 9353 3678 9387 3680
rect 9435 3678 9451 3694
rect 9452 3684 9660 3694
rect 9661 3684 9677 3694
rect 9725 3690 9740 3705
rect 9743 3702 9744 3714
rect 9751 3702 9778 3714
rect 9743 3694 9778 3702
rect 9743 3693 9772 3694
rect 9463 3680 9677 3684
rect 9478 3678 9677 3680
rect 9712 3680 9725 3690
rect 9743 3680 9760 3693
rect 9712 3678 9760 3680
rect 9354 3674 9387 3678
rect 9350 3672 9387 3674
rect 9350 3671 9417 3672
rect 9350 3666 9381 3671
rect 9387 3666 9417 3671
rect 9350 3662 9417 3666
rect 9323 3659 9417 3662
rect 9323 3652 9372 3659
rect 9323 3646 9353 3652
rect 9372 3647 9377 3652
rect 9289 3630 9369 3646
rect 9381 3638 9417 3659
rect 9478 3654 9667 3678
rect 9712 3677 9759 3678
rect 9725 3672 9759 3677
rect 9493 3651 9667 3654
rect 9486 3648 9667 3651
rect 9695 3671 9759 3672
rect 9289 3628 9308 3630
rect 9323 3628 9357 3630
rect 9289 3612 9369 3628
rect 9289 3606 9308 3612
rect 9005 3580 9108 3590
rect 8959 3578 9108 3580
rect 9129 3578 9164 3590
rect 8798 3576 8960 3578
rect 8810 3556 8829 3576
rect 8844 3574 8874 3576
rect 8693 3548 8734 3556
rect 8816 3552 8829 3556
rect 8881 3560 8960 3576
rect 8992 3576 9164 3578
rect 8992 3560 9071 3576
rect 9078 3574 9108 3576
rect 8656 3538 8685 3548
rect 8699 3538 8728 3548
rect 8743 3538 8773 3552
rect 8816 3538 8859 3552
rect 8881 3548 9071 3560
rect 9136 3556 9142 3576
rect 8866 3538 8896 3548
rect 8897 3538 9055 3548
rect 9059 3538 9089 3548
rect 9093 3538 9123 3552
rect 9151 3538 9164 3576
rect 9236 3590 9265 3606
rect 9279 3590 9308 3606
rect 9323 3596 9353 3612
rect 9381 3590 9387 3638
rect 9390 3632 9409 3638
rect 9424 3632 9454 3640
rect 9390 3624 9454 3632
rect 9390 3608 9470 3624
rect 9486 3617 9548 3648
rect 9564 3617 9626 3648
rect 9695 3646 9744 3671
rect 9759 3646 9789 3662
rect 9658 3632 9688 3640
rect 9695 3638 9805 3646
rect 9658 3624 9703 3632
rect 9390 3606 9409 3608
rect 9424 3606 9470 3608
rect 9390 3590 9470 3606
rect 9497 3604 9532 3617
rect 9573 3614 9610 3617
rect 9573 3612 9615 3614
rect 9502 3601 9532 3604
rect 9511 3597 9518 3601
rect 9518 3596 9519 3597
rect 9477 3590 9487 3596
rect 9236 3582 9271 3590
rect 9236 3556 9237 3582
rect 9244 3556 9271 3582
rect 9179 3538 9209 3552
rect 9236 3548 9271 3556
rect 9273 3582 9314 3590
rect 9273 3556 9288 3582
rect 9295 3556 9314 3582
rect 9378 3578 9409 3590
rect 9424 3578 9527 3590
rect 9539 3580 9565 3606
rect 9580 3601 9610 3612
rect 9642 3608 9704 3624
rect 9642 3606 9688 3608
rect 9642 3590 9704 3606
rect 9716 3590 9722 3638
rect 9725 3630 9805 3638
rect 9725 3628 9744 3630
rect 9759 3628 9793 3630
rect 9725 3612 9805 3628
rect 9725 3590 9744 3612
rect 9759 3596 9789 3612
rect 9817 3606 9823 3680
rect 9826 3606 9845 3750
rect 9860 3606 9866 3750
rect 9875 3680 9888 3750
rect 9940 3746 9962 3750
rect 9933 3724 9962 3738
rect 10015 3724 10031 3738
rect 10069 3734 10075 3736
rect 10082 3734 10190 3750
rect 10197 3734 10203 3736
rect 10211 3734 10226 3750
rect 10292 3744 10311 3747
rect 9933 3722 10031 3724
rect 10058 3722 10226 3734
rect 10241 3724 10257 3738
rect 10292 3725 10314 3744
rect 10324 3738 10340 3739
rect 10323 3736 10340 3738
rect 10324 3731 10340 3736
rect 10314 3724 10320 3725
rect 10323 3724 10352 3731
rect 10241 3723 10352 3724
rect 10241 3722 10358 3723
rect 9917 3714 9968 3722
rect 10015 3714 10049 3722
rect 9917 3702 9942 3714
rect 9949 3702 9968 3714
rect 10022 3712 10049 3714
rect 10058 3712 10279 3722
rect 10314 3719 10320 3722
rect 10022 3708 10279 3712
rect 9917 3694 9968 3702
rect 10015 3694 10279 3708
rect 10323 3714 10358 3722
rect 9869 3646 9888 3680
rect 9933 3686 9962 3694
rect 9933 3680 9950 3686
rect 9933 3678 9967 3680
rect 10015 3678 10031 3694
rect 10032 3684 10240 3694
rect 10241 3684 10257 3694
rect 10305 3690 10320 3705
rect 10323 3702 10324 3714
rect 10331 3702 10358 3714
rect 10323 3694 10358 3702
rect 10323 3693 10352 3694
rect 10043 3680 10257 3684
rect 10058 3678 10257 3680
rect 10292 3680 10305 3690
rect 10323 3680 10340 3693
rect 10292 3678 10340 3680
rect 9934 3674 9967 3678
rect 9930 3672 9967 3674
rect 9930 3671 9997 3672
rect 9930 3666 9961 3671
rect 9967 3666 9997 3671
rect 9930 3662 9997 3666
rect 9903 3659 9997 3662
rect 9903 3652 9952 3659
rect 9903 3646 9933 3652
rect 9952 3647 9957 3652
rect 9869 3630 9949 3646
rect 9961 3638 9997 3659
rect 10058 3654 10247 3678
rect 10292 3677 10339 3678
rect 10305 3672 10339 3677
rect 10073 3651 10247 3654
rect 10066 3648 10247 3651
rect 10275 3671 10339 3672
rect 9869 3628 9888 3630
rect 9903 3628 9937 3630
rect 9869 3612 9949 3628
rect 9869 3606 9888 3612
rect 9585 3580 9688 3590
rect 9539 3578 9688 3580
rect 9709 3578 9744 3590
rect 9378 3576 9540 3578
rect 9390 3556 9409 3576
rect 9424 3574 9454 3576
rect 9273 3548 9314 3556
rect 9396 3552 9409 3556
rect 9461 3560 9540 3576
rect 9572 3576 9744 3578
rect 9572 3560 9651 3576
rect 9658 3574 9688 3576
rect 9236 3538 9265 3548
rect 9279 3538 9308 3548
rect 9323 3538 9353 3552
rect 9396 3538 9439 3552
rect 9461 3548 9651 3560
rect 9716 3556 9722 3576
rect 9446 3538 9476 3548
rect 9477 3538 9635 3548
rect 9639 3538 9669 3548
rect 9673 3538 9703 3552
rect 9731 3538 9744 3576
rect 9816 3590 9845 3606
rect 9859 3590 9888 3606
rect 9903 3596 9933 3612
rect 9961 3590 9967 3638
rect 9970 3632 9989 3638
rect 10004 3632 10034 3640
rect 9970 3624 10034 3632
rect 9970 3608 10050 3624
rect 10066 3617 10128 3648
rect 10144 3617 10206 3648
rect 10275 3646 10324 3671
rect 10339 3646 10369 3662
rect 10238 3632 10268 3640
rect 10275 3638 10385 3646
rect 10238 3624 10283 3632
rect 9970 3606 9989 3608
rect 10004 3606 10050 3608
rect 9970 3590 10050 3606
rect 10077 3604 10112 3617
rect 10153 3614 10190 3617
rect 10153 3612 10195 3614
rect 10082 3601 10112 3604
rect 10091 3597 10098 3601
rect 10098 3596 10099 3597
rect 10057 3590 10067 3596
rect 9816 3582 9851 3590
rect 9816 3556 9817 3582
rect 9824 3556 9851 3582
rect 9759 3538 9789 3552
rect 9816 3548 9851 3556
rect 9853 3582 9894 3590
rect 9853 3556 9868 3582
rect 9875 3556 9894 3582
rect 9958 3578 9989 3590
rect 10004 3578 10107 3590
rect 10119 3580 10145 3606
rect 10160 3601 10190 3612
rect 10222 3608 10284 3624
rect 10222 3606 10268 3608
rect 10222 3590 10284 3606
rect 10296 3590 10302 3638
rect 10305 3630 10385 3638
rect 10305 3628 10324 3630
rect 10339 3628 10373 3630
rect 10305 3612 10385 3628
rect 10305 3590 10324 3612
rect 10339 3596 10369 3612
rect 10397 3606 10403 3680
rect 10406 3606 10425 3750
rect 10440 3606 10446 3750
rect 10455 3680 10468 3750
rect 10520 3746 10542 3750
rect 10513 3724 10542 3738
rect 10595 3724 10611 3738
rect 10649 3734 10655 3736
rect 10662 3734 10770 3750
rect 10777 3734 10783 3736
rect 10791 3734 10806 3750
rect 10872 3744 10891 3747
rect 10513 3722 10611 3724
rect 10638 3722 10806 3734
rect 10821 3724 10837 3738
rect 10872 3725 10894 3744
rect 10904 3738 10920 3739
rect 10903 3736 10920 3738
rect 10904 3731 10920 3736
rect 10894 3724 10900 3725
rect 10903 3724 10932 3731
rect 10821 3723 10932 3724
rect 10821 3722 10938 3723
rect 10497 3714 10548 3722
rect 10595 3714 10629 3722
rect 10497 3702 10522 3714
rect 10529 3702 10548 3714
rect 10602 3712 10629 3714
rect 10638 3712 10859 3722
rect 10894 3719 10900 3722
rect 10602 3708 10859 3712
rect 10497 3694 10548 3702
rect 10595 3694 10859 3708
rect 10903 3714 10938 3722
rect 10449 3646 10468 3680
rect 10513 3686 10542 3694
rect 10513 3680 10530 3686
rect 10513 3678 10547 3680
rect 10595 3678 10611 3694
rect 10612 3684 10820 3694
rect 10821 3684 10837 3694
rect 10885 3690 10900 3705
rect 10903 3702 10904 3714
rect 10911 3702 10938 3714
rect 10903 3694 10938 3702
rect 10903 3693 10932 3694
rect 10623 3680 10837 3684
rect 10638 3678 10837 3680
rect 10872 3680 10885 3690
rect 10903 3680 10920 3693
rect 10872 3678 10920 3680
rect 10514 3674 10547 3678
rect 10510 3672 10547 3674
rect 10510 3671 10577 3672
rect 10510 3666 10541 3671
rect 10547 3666 10577 3671
rect 10510 3662 10577 3666
rect 10483 3659 10577 3662
rect 10483 3652 10532 3659
rect 10483 3646 10513 3652
rect 10532 3647 10537 3652
rect 10449 3630 10529 3646
rect 10541 3638 10577 3659
rect 10638 3654 10827 3678
rect 10872 3677 10919 3678
rect 10885 3672 10919 3677
rect 10653 3651 10827 3654
rect 10646 3648 10827 3651
rect 10855 3671 10919 3672
rect 10449 3628 10468 3630
rect 10483 3628 10517 3630
rect 10449 3612 10529 3628
rect 10449 3606 10468 3612
rect 10165 3580 10268 3590
rect 10119 3578 10268 3580
rect 10289 3578 10324 3590
rect 9958 3576 10120 3578
rect 9970 3556 9989 3576
rect 10004 3574 10034 3576
rect 9853 3548 9894 3556
rect 9976 3552 9989 3556
rect 10041 3560 10120 3576
rect 10152 3576 10324 3578
rect 10152 3560 10231 3576
rect 10238 3574 10268 3576
rect 9816 3538 9845 3548
rect 9859 3538 9888 3548
rect 9903 3538 9933 3552
rect 9976 3538 10019 3552
rect 10041 3548 10231 3560
rect 10296 3556 10302 3576
rect 10026 3538 10056 3548
rect 10057 3538 10215 3548
rect 10219 3538 10249 3548
rect 10253 3538 10283 3552
rect 10311 3538 10324 3576
rect 10396 3590 10425 3606
rect 10439 3590 10468 3606
rect 10483 3596 10513 3612
rect 10541 3590 10547 3638
rect 10550 3632 10569 3638
rect 10584 3632 10614 3640
rect 10550 3624 10614 3632
rect 10550 3608 10630 3624
rect 10646 3617 10708 3648
rect 10724 3617 10786 3648
rect 10855 3646 10904 3671
rect 10919 3646 10949 3662
rect 10818 3632 10848 3640
rect 10855 3638 10965 3646
rect 10818 3624 10863 3632
rect 10550 3606 10569 3608
rect 10584 3606 10630 3608
rect 10550 3590 10630 3606
rect 10657 3604 10692 3617
rect 10733 3614 10770 3617
rect 10733 3612 10775 3614
rect 10662 3601 10692 3604
rect 10671 3597 10678 3601
rect 10678 3596 10679 3597
rect 10637 3590 10647 3596
rect 10396 3582 10431 3590
rect 10396 3556 10397 3582
rect 10404 3556 10431 3582
rect 10339 3538 10369 3552
rect 10396 3548 10431 3556
rect 10433 3582 10474 3590
rect 10433 3556 10448 3582
rect 10455 3556 10474 3582
rect 10538 3578 10569 3590
rect 10584 3578 10687 3590
rect 10699 3580 10725 3606
rect 10740 3601 10770 3612
rect 10802 3608 10864 3624
rect 10802 3606 10848 3608
rect 10802 3590 10864 3606
rect 10876 3590 10882 3638
rect 10885 3630 10965 3638
rect 10885 3628 10904 3630
rect 10919 3628 10953 3630
rect 10885 3612 10965 3628
rect 10885 3590 10904 3612
rect 10919 3596 10949 3612
rect 10977 3606 10983 3680
rect 10986 3606 11005 3750
rect 11020 3606 11026 3750
rect 11035 3680 11048 3750
rect 11100 3746 11122 3750
rect 11093 3724 11122 3738
rect 11175 3724 11191 3738
rect 11229 3734 11235 3736
rect 11242 3734 11350 3750
rect 11357 3734 11363 3736
rect 11371 3734 11386 3750
rect 11452 3744 11471 3747
rect 11093 3722 11191 3724
rect 11218 3722 11386 3734
rect 11401 3724 11417 3738
rect 11452 3725 11474 3744
rect 11484 3738 11500 3739
rect 11483 3736 11500 3738
rect 11484 3731 11500 3736
rect 11474 3724 11480 3725
rect 11483 3724 11512 3731
rect 11401 3723 11512 3724
rect 11401 3722 11518 3723
rect 11077 3714 11128 3722
rect 11175 3714 11209 3722
rect 11077 3702 11102 3714
rect 11109 3702 11128 3714
rect 11182 3712 11209 3714
rect 11218 3712 11439 3722
rect 11474 3719 11480 3722
rect 11182 3708 11439 3712
rect 11077 3694 11128 3702
rect 11175 3694 11439 3708
rect 11483 3714 11518 3722
rect 11029 3646 11048 3680
rect 11093 3686 11122 3694
rect 11093 3680 11110 3686
rect 11093 3678 11127 3680
rect 11175 3678 11191 3694
rect 11192 3684 11400 3694
rect 11401 3684 11417 3694
rect 11465 3690 11480 3705
rect 11483 3702 11484 3714
rect 11491 3702 11518 3714
rect 11483 3694 11518 3702
rect 11483 3693 11512 3694
rect 11203 3680 11417 3684
rect 11218 3678 11417 3680
rect 11452 3680 11465 3690
rect 11483 3680 11500 3693
rect 11452 3678 11500 3680
rect 11094 3674 11127 3678
rect 11090 3672 11127 3674
rect 11090 3671 11157 3672
rect 11090 3666 11121 3671
rect 11127 3666 11157 3671
rect 11090 3662 11157 3666
rect 11063 3659 11157 3662
rect 11063 3652 11112 3659
rect 11063 3646 11093 3652
rect 11112 3647 11117 3652
rect 11029 3630 11109 3646
rect 11121 3638 11157 3659
rect 11218 3654 11407 3678
rect 11452 3677 11499 3678
rect 11465 3672 11499 3677
rect 11233 3651 11407 3654
rect 11226 3648 11407 3651
rect 11435 3671 11499 3672
rect 11029 3628 11048 3630
rect 11063 3628 11097 3630
rect 11029 3612 11109 3628
rect 11029 3606 11048 3612
rect 10745 3580 10848 3590
rect 10699 3578 10848 3580
rect 10869 3578 10904 3590
rect 10538 3576 10700 3578
rect 10550 3556 10569 3576
rect 10584 3574 10614 3576
rect 10433 3548 10474 3556
rect 10556 3552 10569 3556
rect 10621 3560 10700 3576
rect 10732 3576 10904 3578
rect 10732 3560 10811 3576
rect 10818 3574 10848 3576
rect 10396 3538 10425 3548
rect 10439 3538 10468 3548
rect 10483 3538 10513 3552
rect 10556 3538 10599 3552
rect 10621 3548 10811 3560
rect 10876 3556 10882 3576
rect 10606 3538 10636 3548
rect 10637 3538 10795 3548
rect 10799 3538 10829 3548
rect 10833 3538 10863 3552
rect 10891 3538 10904 3576
rect 10976 3590 11005 3606
rect 11019 3590 11048 3606
rect 11063 3596 11093 3612
rect 11121 3590 11127 3638
rect 11130 3632 11149 3638
rect 11164 3632 11194 3640
rect 11130 3624 11194 3632
rect 11130 3608 11210 3624
rect 11226 3617 11288 3648
rect 11304 3617 11366 3648
rect 11435 3646 11484 3671
rect 11499 3646 11529 3662
rect 11398 3632 11428 3640
rect 11435 3638 11545 3646
rect 11398 3624 11443 3632
rect 11130 3606 11149 3608
rect 11164 3606 11210 3608
rect 11130 3590 11210 3606
rect 11237 3604 11272 3617
rect 11313 3614 11350 3617
rect 11313 3612 11355 3614
rect 11242 3601 11272 3604
rect 11251 3597 11258 3601
rect 11258 3596 11259 3597
rect 11217 3590 11227 3596
rect 10976 3582 11011 3590
rect 10976 3556 10977 3582
rect 10984 3556 11011 3582
rect 10919 3538 10949 3552
rect 10976 3548 11011 3556
rect 11013 3582 11054 3590
rect 11013 3556 11028 3582
rect 11035 3556 11054 3582
rect 11118 3578 11149 3590
rect 11164 3578 11267 3590
rect 11279 3580 11305 3606
rect 11320 3601 11350 3612
rect 11382 3608 11444 3624
rect 11382 3606 11428 3608
rect 11382 3590 11444 3606
rect 11456 3590 11462 3638
rect 11465 3630 11545 3638
rect 11465 3628 11484 3630
rect 11499 3628 11533 3630
rect 11465 3612 11545 3628
rect 11465 3590 11484 3612
rect 11499 3596 11529 3612
rect 11557 3606 11563 3680
rect 11566 3606 11585 3750
rect 11600 3606 11606 3750
rect 11615 3680 11628 3750
rect 11680 3746 11702 3750
rect 11673 3724 11702 3738
rect 11755 3724 11771 3738
rect 11809 3734 11815 3736
rect 11822 3734 11930 3750
rect 11937 3734 11943 3736
rect 11951 3734 11966 3750
rect 12032 3744 12051 3747
rect 11673 3722 11771 3724
rect 11798 3722 11966 3734
rect 11981 3724 11997 3738
rect 12032 3725 12054 3744
rect 12064 3738 12080 3739
rect 12063 3736 12080 3738
rect 12064 3731 12080 3736
rect 12054 3724 12060 3725
rect 12063 3724 12092 3731
rect 11981 3723 12092 3724
rect 11981 3722 12098 3723
rect 11657 3714 11708 3722
rect 11755 3714 11789 3722
rect 11657 3702 11682 3714
rect 11689 3702 11708 3714
rect 11762 3712 11789 3714
rect 11798 3712 12019 3722
rect 12054 3719 12060 3722
rect 11762 3708 12019 3712
rect 11657 3694 11708 3702
rect 11755 3694 12019 3708
rect 12063 3714 12098 3722
rect 11609 3646 11628 3680
rect 11673 3686 11702 3694
rect 11673 3680 11690 3686
rect 11673 3678 11707 3680
rect 11755 3678 11771 3694
rect 11772 3684 11980 3694
rect 11981 3684 11997 3694
rect 12045 3690 12060 3705
rect 12063 3702 12064 3714
rect 12071 3702 12098 3714
rect 12063 3694 12098 3702
rect 12063 3693 12092 3694
rect 11783 3680 11997 3684
rect 11798 3678 11997 3680
rect 12032 3680 12045 3690
rect 12063 3680 12080 3693
rect 12032 3678 12080 3680
rect 11674 3674 11707 3678
rect 11670 3672 11707 3674
rect 11670 3671 11737 3672
rect 11670 3666 11701 3671
rect 11707 3666 11737 3671
rect 11670 3662 11737 3666
rect 11643 3659 11737 3662
rect 11643 3652 11692 3659
rect 11643 3646 11673 3652
rect 11692 3647 11697 3652
rect 11609 3630 11689 3646
rect 11701 3638 11737 3659
rect 11798 3654 11987 3678
rect 12032 3677 12079 3678
rect 12045 3672 12079 3677
rect 11813 3651 11987 3654
rect 11806 3648 11987 3651
rect 12015 3671 12079 3672
rect 11609 3628 11628 3630
rect 11643 3628 11677 3630
rect 11609 3612 11689 3628
rect 11609 3606 11628 3612
rect 11325 3580 11428 3590
rect 11279 3578 11428 3580
rect 11449 3578 11484 3590
rect 11118 3576 11280 3578
rect 11130 3556 11149 3576
rect 11164 3574 11194 3576
rect 11013 3548 11054 3556
rect 11136 3552 11149 3556
rect 11201 3560 11280 3576
rect 11312 3576 11484 3578
rect 11312 3560 11391 3576
rect 11398 3574 11428 3576
rect 10976 3538 11005 3548
rect 11019 3538 11048 3548
rect 11063 3538 11093 3552
rect 11136 3538 11179 3552
rect 11201 3548 11391 3560
rect 11456 3556 11462 3576
rect 11186 3538 11216 3548
rect 11217 3538 11375 3548
rect 11379 3538 11409 3548
rect 11413 3538 11443 3552
rect 11471 3538 11484 3576
rect 11556 3590 11585 3606
rect 11599 3590 11628 3606
rect 11643 3596 11673 3612
rect 11701 3590 11707 3638
rect 11710 3632 11729 3638
rect 11744 3632 11774 3640
rect 11710 3624 11774 3632
rect 11710 3608 11790 3624
rect 11806 3617 11868 3648
rect 11884 3617 11946 3648
rect 12015 3646 12064 3671
rect 12079 3646 12109 3662
rect 11978 3632 12008 3640
rect 12015 3638 12125 3646
rect 11978 3624 12023 3632
rect 11710 3606 11729 3608
rect 11744 3606 11790 3608
rect 11710 3590 11790 3606
rect 11817 3604 11852 3617
rect 11893 3614 11930 3617
rect 11893 3612 11935 3614
rect 11822 3601 11852 3604
rect 11831 3597 11838 3601
rect 11838 3596 11839 3597
rect 11797 3590 11807 3596
rect 11556 3582 11591 3590
rect 11556 3556 11557 3582
rect 11564 3556 11591 3582
rect 11499 3538 11529 3552
rect 11556 3548 11591 3556
rect 11593 3582 11634 3590
rect 11593 3556 11608 3582
rect 11615 3556 11634 3582
rect 11698 3578 11729 3590
rect 11744 3578 11847 3590
rect 11859 3580 11885 3606
rect 11900 3601 11930 3612
rect 11962 3608 12024 3624
rect 11962 3606 12008 3608
rect 11962 3590 12024 3606
rect 12036 3590 12042 3638
rect 12045 3630 12125 3638
rect 12045 3628 12064 3630
rect 12079 3628 12113 3630
rect 12045 3612 12125 3628
rect 12045 3590 12064 3612
rect 12079 3596 12109 3612
rect 12137 3606 12143 3680
rect 12146 3606 12165 3750
rect 12180 3606 12186 3750
rect 12195 3680 12208 3750
rect 12260 3746 12282 3750
rect 12253 3724 12282 3738
rect 12335 3724 12351 3738
rect 12389 3734 12395 3736
rect 12402 3734 12510 3750
rect 12517 3734 12523 3736
rect 12531 3734 12546 3750
rect 12612 3744 12631 3747
rect 12253 3722 12351 3724
rect 12378 3722 12546 3734
rect 12561 3724 12577 3738
rect 12612 3725 12634 3744
rect 12644 3738 12660 3739
rect 12643 3736 12660 3738
rect 12644 3731 12660 3736
rect 12634 3724 12640 3725
rect 12643 3724 12672 3731
rect 12561 3723 12672 3724
rect 12561 3722 12678 3723
rect 12237 3714 12288 3722
rect 12335 3714 12369 3722
rect 12237 3702 12262 3714
rect 12269 3702 12288 3714
rect 12342 3712 12369 3714
rect 12378 3712 12599 3722
rect 12634 3719 12640 3722
rect 12342 3708 12599 3712
rect 12237 3694 12288 3702
rect 12335 3694 12599 3708
rect 12643 3714 12678 3722
rect 12189 3646 12208 3680
rect 12253 3686 12282 3694
rect 12253 3680 12270 3686
rect 12253 3678 12287 3680
rect 12335 3678 12351 3694
rect 12352 3684 12560 3694
rect 12561 3684 12577 3694
rect 12625 3690 12640 3705
rect 12643 3702 12644 3714
rect 12651 3702 12678 3714
rect 12643 3694 12678 3702
rect 12643 3693 12672 3694
rect 12363 3680 12577 3684
rect 12378 3678 12577 3680
rect 12612 3680 12625 3690
rect 12643 3680 12660 3693
rect 12612 3678 12660 3680
rect 12254 3674 12287 3678
rect 12250 3672 12287 3674
rect 12250 3671 12317 3672
rect 12250 3666 12281 3671
rect 12287 3666 12317 3671
rect 12250 3662 12317 3666
rect 12223 3659 12317 3662
rect 12223 3652 12272 3659
rect 12223 3646 12253 3652
rect 12272 3647 12277 3652
rect 12189 3630 12269 3646
rect 12281 3638 12317 3659
rect 12378 3654 12567 3678
rect 12612 3677 12659 3678
rect 12625 3672 12659 3677
rect 12393 3651 12567 3654
rect 12386 3648 12567 3651
rect 12595 3671 12659 3672
rect 12189 3628 12208 3630
rect 12223 3628 12257 3630
rect 12189 3612 12269 3628
rect 12189 3606 12208 3612
rect 11905 3580 12008 3590
rect 11859 3578 12008 3580
rect 12029 3578 12064 3590
rect 11698 3576 11860 3578
rect 11710 3556 11729 3576
rect 11744 3574 11774 3576
rect 11593 3548 11634 3556
rect 11716 3552 11729 3556
rect 11781 3560 11860 3576
rect 11892 3576 12064 3578
rect 11892 3560 11971 3576
rect 11978 3574 12008 3576
rect 11556 3538 11585 3548
rect 11599 3538 11628 3548
rect 11643 3538 11673 3552
rect 11716 3538 11759 3552
rect 11781 3548 11971 3560
rect 12036 3556 12042 3576
rect 11766 3538 11796 3548
rect 11797 3538 11955 3548
rect 11959 3538 11989 3548
rect 11993 3538 12023 3552
rect 12051 3538 12064 3576
rect 12136 3590 12165 3606
rect 12179 3590 12208 3606
rect 12223 3596 12253 3612
rect 12281 3590 12287 3638
rect 12290 3632 12309 3638
rect 12324 3632 12354 3640
rect 12290 3624 12354 3632
rect 12290 3608 12370 3624
rect 12386 3617 12448 3648
rect 12464 3617 12526 3648
rect 12595 3646 12644 3671
rect 12659 3646 12689 3662
rect 12558 3632 12588 3640
rect 12595 3638 12705 3646
rect 12558 3624 12603 3632
rect 12290 3606 12309 3608
rect 12324 3606 12370 3608
rect 12290 3590 12370 3606
rect 12397 3604 12432 3617
rect 12473 3614 12510 3617
rect 12473 3612 12515 3614
rect 12402 3601 12432 3604
rect 12411 3597 12418 3601
rect 12418 3596 12419 3597
rect 12377 3590 12387 3596
rect 12136 3582 12171 3590
rect 12136 3556 12137 3582
rect 12144 3556 12171 3582
rect 12079 3538 12109 3552
rect 12136 3548 12171 3556
rect 12173 3582 12214 3590
rect 12173 3556 12188 3582
rect 12195 3556 12214 3582
rect 12278 3578 12309 3590
rect 12324 3578 12427 3590
rect 12439 3580 12465 3606
rect 12480 3601 12510 3612
rect 12542 3608 12604 3624
rect 12542 3606 12588 3608
rect 12542 3590 12604 3606
rect 12616 3590 12622 3638
rect 12625 3630 12705 3638
rect 12625 3628 12644 3630
rect 12659 3628 12693 3630
rect 12625 3612 12705 3628
rect 12625 3590 12644 3612
rect 12659 3596 12689 3612
rect 12717 3606 12723 3680
rect 12726 3606 12745 3750
rect 12760 3606 12766 3750
rect 12775 3680 12788 3750
rect 12840 3746 12862 3750
rect 12833 3724 12862 3738
rect 12915 3724 12931 3738
rect 12969 3734 12975 3736
rect 12982 3734 13090 3750
rect 13097 3734 13103 3736
rect 13111 3734 13126 3750
rect 13192 3744 13211 3747
rect 12833 3722 12931 3724
rect 12958 3722 13126 3734
rect 13141 3724 13157 3738
rect 13192 3725 13214 3744
rect 13224 3738 13240 3739
rect 13223 3736 13240 3738
rect 13224 3731 13240 3736
rect 13214 3724 13220 3725
rect 13223 3724 13252 3731
rect 13141 3723 13252 3724
rect 13141 3722 13258 3723
rect 12817 3714 12868 3722
rect 12915 3714 12949 3722
rect 12817 3702 12842 3714
rect 12849 3702 12868 3714
rect 12922 3712 12949 3714
rect 12958 3712 13179 3722
rect 13214 3719 13220 3722
rect 12922 3708 13179 3712
rect 12817 3694 12868 3702
rect 12915 3694 13179 3708
rect 13223 3714 13258 3722
rect 12769 3646 12788 3680
rect 12833 3686 12862 3694
rect 12833 3680 12850 3686
rect 12833 3678 12867 3680
rect 12915 3678 12931 3694
rect 12932 3684 13140 3694
rect 13141 3684 13157 3694
rect 13205 3690 13220 3705
rect 13223 3702 13224 3714
rect 13231 3702 13258 3714
rect 13223 3694 13258 3702
rect 13223 3693 13252 3694
rect 12943 3680 13157 3684
rect 12958 3678 13157 3680
rect 13192 3680 13205 3690
rect 13223 3680 13240 3693
rect 13192 3678 13240 3680
rect 12834 3674 12867 3678
rect 12830 3672 12867 3674
rect 12830 3671 12897 3672
rect 12830 3666 12861 3671
rect 12867 3666 12897 3671
rect 12830 3662 12897 3666
rect 12803 3659 12897 3662
rect 12803 3652 12852 3659
rect 12803 3646 12833 3652
rect 12852 3647 12857 3652
rect 12769 3630 12849 3646
rect 12861 3638 12897 3659
rect 12958 3654 13147 3678
rect 13192 3677 13239 3678
rect 13205 3672 13239 3677
rect 12973 3651 13147 3654
rect 12966 3648 13147 3651
rect 13175 3671 13239 3672
rect 12769 3628 12788 3630
rect 12803 3628 12837 3630
rect 12769 3612 12849 3628
rect 12769 3606 12788 3612
rect 12485 3580 12588 3590
rect 12439 3578 12588 3580
rect 12609 3578 12644 3590
rect 12278 3576 12440 3578
rect 12290 3556 12309 3576
rect 12324 3574 12354 3576
rect 12173 3548 12214 3556
rect 12296 3552 12309 3556
rect 12361 3560 12440 3576
rect 12472 3576 12644 3578
rect 12472 3560 12551 3576
rect 12558 3574 12588 3576
rect 12136 3538 12165 3548
rect 12179 3538 12208 3548
rect 12223 3538 12253 3552
rect 12296 3538 12339 3552
rect 12361 3548 12551 3560
rect 12616 3556 12622 3576
rect 12346 3538 12376 3548
rect 12377 3538 12535 3548
rect 12539 3538 12569 3548
rect 12573 3538 12603 3552
rect 12631 3538 12644 3576
rect 12716 3590 12745 3606
rect 12759 3590 12788 3606
rect 12803 3596 12833 3612
rect 12861 3590 12867 3638
rect 12870 3632 12889 3638
rect 12904 3632 12934 3640
rect 12870 3624 12934 3632
rect 12870 3608 12950 3624
rect 12966 3617 13028 3648
rect 13044 3617 13106 3648
rect 13175 3646 13224 3671
rect 13239 3646 13269 3662
rect 13138 3632 13168 3640
rect 13175 3638 13285 3646
rect 13138 3624 13183 3632
rect 12870 3606 12889 3608
rect 12904 3606 12950 3608
rect 12870 3590 12950 3606
rect 12977 3604 13012 3617
rect 13053 3614 13090 3617
rect 13053 3612 13095 3614
rect 12982 3601 13012 3604
rect 12991 3597 12998 3601
rect 12998 3596 12999 3597
rect 12957 3590 12967 3596
rect 12716 3582 12751 3590
rect 12716 3556 12717 3582
rect 12724 3556 12751 3582
rect 12659 3538 12689 3552
rect 12716 3548 12751 3556
rect 12753 3582 12794 3590
rect 12753 3556 12768 3582
rect 12775 3556 12794 3582
rect 12858 3578 12889 3590
rect 12904 3578 13007 3590
rect 13019 3580 13045 3606
rect 13060 3601 13090 3612
rect 13122 3608 13184 3624
rect 13122 3606 13168 3608
rect 13122 3590 13184 3606
rect 13196 3590 13202 3638
rect 13205 3630 13285 3638
rect 13205 3628 13224 3630
rect 13239 3628 13273 3630
rect 13205 3612 13285 3628
rect 13205 3590 13224 3612
rect 13239 3596 13269 3612
rect 13297 3606 13303 3680
rect 13306 3606 13325 3750
rect 13340 3606 13346 3750
rect 13355 3680 13368 3750
rect 13420 3746 13442 3750
rect 13413 3724 13442 3738
rect 13495 3724 13511 3738
rect 13549 3734 13555 3736
rect 13562 3734 13670 3750
rect 13677 3734 13683 3736
rect 13691 3734 13706 3750
rect 13772 3744 13791 3747
rect 13413 3722 13511 3724
rect 13538 3722 13706 3734
rect 13721 3724 13737 3738
rect 13772 3725 13794 3744
rect 13804 3738 13820 3739
rect 13803 3736 13820 3738
rect 13804 3731 13820 3736
rect 13794 3724 13800 3725
rect 13803 3724 13832 3731
rect 13721 3723 13832 3724
rect 13721 3722 13838 3723
rect 13397 3714 13448 3722
rect 13495 3714 13529 3722
rect 13397 3702 13422 3714
rect 13429 3702 13448 3714
rect 13502 3712 13529 3714
rect 13538 3712 13759 3722
rect 13794 3719 13800 3722
rect 13502 3708 13759 3712
rect 13397 3694 13448 3702
rect 13495 3694 13759 3708
rect 13803 3714 13838 3722
rect 13349 3646 13368 3680
rect 13413 3686 13442 3694
rect 13413 3680 13430 3686
rect 13413 3678 13447 3680
rect 13495 3678 13511 3694
rect 13512 3684 13720 3694
rect 13721 3684 13737 3694
rect 13785 3690 13800 3705
rect 13803 3702 13804 3714
rect 13811 3702 13838 3714
rect 13803 3694 13838 3702
rect 13803 3693 13832 3694
rect 13523 3680 13737 3684
rect 13538 3678 13737 3680
rect 13772 3680 13785 3690
rect 13803 3680 13820 3693
rect 13772 3678 13820 3680
rect 13414 3674 13447 3678
rect 13410 3672 13447 3674
rect 13410 3671 13477 3672
rect 13410 3666 13441 3671
rect 13447 3666 13477 3671
rect 13410 3662 13477 3666
rect 13383 3659 13477 3662
rect 13383 3652 13432 3659
rect 13383 3646 13413 3652
rect 13432 3647 13437 3652
rect 13349 3630 13429 3646
rect 13441 3638 13477 3659
rect 13538 3654 13727 3678
rect 13772 3677 13819 3678
rect 13785 3672 13819 3677
rect 13553 3651 13727 3654
rect 13546 3648 13727 3651
rect 13755 3671 13819 3672
rect 13349 3628 13368 3630
rect 13383 3628 13417 3630
rect 13349 3612 13429 3628
rect 13349 3606 13368 3612
rect 13065 3580 13168 3590
rect 13019 3578 13168 3580
rect 13189 3578 13224 3590
rect 12858 3576 13020 3578
rect 12870 3556 12889 3576
rect 12904 3574 12934 3576
rect 12753 3548 12794 3556
rect 12876 3552 12889 3556
rect 12941 3560 13020 3576
rect 13052 3576 13224 3578
rect 13052 3560 13131 3576
rect 13138 3574 13168 3576
rect 12716 3538 12745 3548
rect 12759 3538 12788 3548
rect 12803 3538 12833 3552
rect 12876 3538 12919 3552
rect 12941 3548 13131 3560
rect 13196 3556 13202 3576
rect 12926 3538 12956 3548
rect 12957 3538 13115 3548
rect 13119 3538 13149 3548
rect 13153 3538 13183 3552
rect 13211 3538 13224 3576
rect 13296 3590 13325 3606
rect 13339 3590 13368 3606
rect 13383 3596 13413 3612
rect 13441 3590 13447 3638
rect 13450 3632 13469 3638
rect 13484 3632 13514 3640
rect 13450 3624 13514 3632
rect 13450 3608 13530 3624
rect 13546 3617 13608 3648
rect 13624 3617 13686 3648
rect 13755 3646 13804 3671
rect 13819 3646 13849 3662
rect 13718 3632 13748 3640
rect 13755 3638 13865 3646
rect 13718 3624 13763 3632
rect 13450 3606 13469 3608
rect 13484 3606 13530 3608
rect 13450 3590 13530 3606
rect 13557 3604 13592 3617
rect 13633 3614 13670 3617
rect 13633 3612 13675 3614
rect 13562 3601 13592 3604
rect 13571 3597 13578 3601
rect 13578 3596 13579 3597
rect 13537 3590 13547 3596
rect 13296 3582 13331 3590
rect 13296 3556 13297 3582
rect 13304 3556 13331 3582
rect 13239 3538 13269 3552
rect 13296 3548 13331 3556
rect 13333 3582 13374 3590
rect 13333 3556 13348 3582
rect 13355 3556 13374 3582
rect 13438 3578 13469 3590
rect 13484 3578 13587 3590
rect 13599 3580 13625 3606
rect 13640 3601 13670 3612
rect 13702 3608 13764 3624
rect 13702 3606 13748 3608
rect 13702 3590 13764 3606
rect 13776 3590 13782 3638
rect 13785 3630 13865 3638
rect 13785 3628 13804 3630
rect 13819 3628 13853 3630
rect 13785 3612 13865 3628
rect 13785 3590 13804 3612
rect 13819 3596 13849 3612
rect 13877 3606 13883 3680
rect 13886 3606 13905 3750
rect 13920 3606 13926 3750
rect 13935 3680 13948 3750
rect 14000 3746 14022 3750
rect 13993 3724 14022 3738
rect 14075 3724 14091 3738
rect 14129 3734 14135 3736
rect 14142 3734 14250 3750
rect 14257 3734 14263 3736
rect 14271 3734 14286 3750
rect 14352 3744 14371 3747
rect 13993 3722 14091 3724
rect 14118 3722 14286 3734
rect 14301 3724 14317 3738
rect 14352 3725 14374 3744
rect 14384 3738 14400 3739
rect 14383 3736 14400 3738
rect 14384 3731 14400 3736
rect 14374 3724 14380 3725
rect 14383 3724 14412 3731
rect 14301 3723 14412 3724
rect 14301 3722 14418 3723
rect 13977 3714 14028 3722
rect 14075 3714 14109 3722
rect 13977 3702 14002 3714
rect 14009 3702 14028 3714
rect 14082 3712 14109 3714
rect 14118 3712 14339 3722
rect 14374 3719 14380 3722
rect 14082 3708 14339 3712
rect 13977 3694 14028 3702
rect 14075 3694 14339 3708
rect 14383 3714 14418 3722
rect 13929 3646 13948 3680
rect 13993 3686 14022 3694
rect 13993 3680 14010 3686
rect 13993 3678 14027 3680
rect 14075 3678 14091 3694
rect 14092 3684 14300 3694
rect 14301 3684 14317 3694
rect 14365 3690 14380 3705
rect 14383 3702 14384 3714
rect 14391 3702 14418 3714
rect 14383 3694 14418 3702
rect 14383 3693 14412 3694
rect 14103 3680 14317 3684
rect 14118 3678 14317 3680
rect 14352 3680 14365 3690
rect 14383 3680 14400 3693
rect 14352 3678 14400 3680
rect 13994 3674 14027 3678
rect 13990 3672 14027 3674
rect 13990 3671 14057 3672
rect 13990 3666 14021 3671
rect 14027 3666 14057 3671
rect 13990 3662 14057 3666
rect 13963 3659 14057 3662
rect 13963 3652 14012 3659
rect 13963 3646 13993 3652
rect 14012 3647 14017 3652
rect 13929 3630 14009 3646
rect 14021 3638 14057 3659
rect 14118 3654 14307 3678
rect 14352 3677 14399 3678
rect 14365 3672 14399 3677
rect 14133 3651 14307 3654
rect 14126 3648 14307 3651
rect 14335 3671 14399 3672
rect 13929 3628 13948 3630
rect 13963 3628 13997 3630
rect 13929 3612 14009 3628
rect 13929 3606 13948 3612
rect 13645 3580 13748 3590
rect 13599 3578 13748 3580
rect 13769 3578 13804 3590
rect 13438 3576 13600 3578
rect 13450 3556 13469 3576
rect 13484 3574 13514 3576
rect 13333 3548 13374 3556
rect 13456 3552 13469 3556
rect 13521 3560 13600 3576
rect 13632 3576 13804 3578
rect 13632 3560 13711 3576
rect 13718 3574 13748 3576
rect 13296 3538 13325 3548
rect 13339 3538 13368 3548
rect 13383 3538 13413 3552
rect 13456 3538 13499 3552
rect 13521 3548 13711 3560
rect 13776 3556 13782 3576
rect 13506 3538 13536 3548
rect 13537 3538 13695 3548
rect 13699 3538 13729 3548
rect 13733 3538 13763 3552
rect 13791 3538 13804 3576
rect 13876 3590 13905 3606
rect 13919 3590 13948 3606
rect 13963 3596 13993 3612
rect 14021 3590 14027 3638
rect 14030 3632 14049 3638
rect 14064 3632 14094 3640
rect 14030 3624 14094 3632
rect 14030 3608 14110 3624
rect 14126 3617 14188 3648
rect 14204 3617 14266 3648
rect 14335 3646 14384 3671
rect 14399 3646 14429 3662
rect 14298 3632 14328 3640
rect 14335 3638 14445 3646
rect 14298 3624 14343 3632
rect 14030 3606 14049 3608
rect 14064 3606 14110 3608
rect 14030 3590 14110 3606
rect 14137 3604 14172 3617
rect 14213 3614 14250 3617
rect 14213 3612 14255 3614
rect 14142 3601 14172 3604
rect 14151 3597 14158 3601
rect 14158 3596 14159 3597
rect 14117 3590 14127 3596
rect 13876 3582 13911 3590
rect 13876 3556 13877 3582
rect 13884 3556 13911 3582
rect 13819 3538 13849 3552
rect 13876 3548 13911 3556
rect 13913 3582 13954 3590
rect 13913 3556 13928 3582
rect 13935 3556 13954 3582
rect 14018 3578 14049 3590
rect 14064 3578 14167 3590
rect 14179 3580 14205 3606
rect 14220 3601 14250 3612
rect 14282 3608 14344 3624
rect 14282 3606 14328 3608
rect 14282 3590 14344 3606
rect 14356 3590 14362 3638
rect 14365 3630 14445 3638
rect 14365 3628 14384 3630
rect 14399 3628 14433 3630
rect 14365 3612 14445 3628
rect 14365 3590 14384 3612
rect 14399 3596 14429 3612
rect 14457 3606 14463 3680
rect 14466 3606 14485 3750
rect 14500 3606 14506 3750
rect 14515 3680 14528 3750
rect 14580 3746 14602 3750
rect 14573 3724 14602 3738
rect 14655 3724 14671 3738
rect 14709 3734 14715 3736
rect 14722 3734 14830 3750
rect 14837 3734 14843 3736
rect 14851 3734 14866 3750
rect 14932 3744 14951 3747
rect 14573 3722 14671 3724
rect 14698 3722 14866 3734
rect 14881 3724 14897 3738
rect 14932 3725 14954 3744
rect 14964 3738 14980 3739
rect 14963 3736 14980 3738
rect 14964 3731 14980 3736
rect 14954 3724 14960 3725
rect 14963 3724 14992 3731
rect 14881 3723 14992 3724
rect 14881 3722 14998 3723
rect 14557 3714 14608 3722
rect 14655 3714 14689 3722
rect 14557 3702 14582 3714
rect 14589 3702 14608 3714
rect 14662 3712 14689 3714
rect 14698 3712 14919 3722
rect 14954 3719 14960 3722
rect 14662 3708 14919 3712
rect 14557 3694 14608 3702
rect 14655 3694 14919 3708
rect 14963 3714 14998 3722
rect 14509 3646 14528 3680
rect 14573 3686 14602 3694
rect 14573 3680 14590 3686
rect 14573 3678 14607 3680
rect 14655 3678 14671 3694
rect 14672 3684 14880 3694
rect 14881 3684 14897 3694
rect 14945 3690 14960 3705
rect 14963 3702 14964 3714
rect 14971 3702 14998 3714
rect 14963 3694 14998 3702
rect 14963 3693 14992 3694
rect 14683 3680 14897 3684
rect 14698 3678 14897 3680
rect 14932 3680 14945 3690
rect 14963 3680 14980 3693
rect 14932 3678 14980 3680
rect 14574 3674 14607 3678
rect 14570 3672 14607 3674
rect 14570 3671 14637 3672
rect 14570 3666 14601 3671
rect 14607 3666 14637 3671
rect 14570 3662 14637 3666
rect 14543 3659 14637 3662
rect 14543 3652 14592 3659
rect 14543 3646 14573 3652
rect 14592 3647 14597 3652
rect 14509 3630 14589 3646
rect 14601 3638 14637 3659
rect 14698 3654 14887 3678
rect 14932 3677 14979 3678
rect 14945 3672 14979 3677
rect 14713 3651 14887 3654
rect 14706 3648 14887 3651
rect 14915 3671 14979 3672
rect 14509 3628 14528 3630
rect 14543 3628 14577 3630
rect 14509 3612 14589 3628
rect 14509 3606 14528 3612
rect 14225 3580 14328 3590
rect 14179 3578 14328 3580
rect 14349 3578 14384 3590
rect 14018 3576 14180 3578
rect 14030 3556 14049 3576
rect 14064 3574 14094 3576
rect 13913 3548 13954 3556
rect 14036 3552 14049 3556
rect 14101 3560 14180 3576
rect 14212 3576 14384 3578
rect 14212 3560 14291 3576
rect 14298 3574 14328 3576
rect 13876 3538 13905 3548
rect 13919 3538 13948 3548
rect 13963 3538 13993 3552
rect 14036 3538 14079 3552
rect 14101 3548 14291 3560
rect 14356 3556 14362 3576
rect 14086 3538 14116 3548
rect 14117 3538 14275 3548
rect 14279 3538 14309 3548
rect 14313 3538 14343 3552
rect 14371 3538 14384 3576
rect 14456 3590 14485 3606
rect 14499 3590 14528 3606
rect 14543 3596 14573 3612
rect 14601 3590 14607 3638
rect 14610 3632 14629 3638
rect 14644 3632 14674 3640
rect 14610 3624 14674 3632
rect 14610 3608 14690 3624
rect 14706 3617 14768 3648
rect 14784 3617 14846 3648
rect 14915 3646 14964 3671
rect 14979 3646 15009 3662
rect 14878 3632 14908 3640
rect 14915 3638 15025 3646
rect 14878 3624 14923 3632
rect 14610 3606 14629 3608
rect 14644 3606 14690 3608
rect 14610 3590 14690 3606
rect 14717 3604 14752 3617
rect 14793 3614 14830 3617
rect 14793 3612 14835 3614
rect 14722 3601 14752 3604
rect 14731 3597 14738 3601
rect 14738 3596 14739 3597
rect 14697 3590 14707 3596
rect 14456 3582 14491 3590
rect 14456 3556 14457 3582
rect 14464 3556 14491 3582
rect 14399 3538 14429 3552
rect 14456 3548 14491 3556
rect 14493 3582 14534 3590
rect 14493 3556 14508 3582
rect 14515 3556 14534 3582
rect 14598 3578 14629 3590
rect 14644 3578 14747 3590
rect 14759 3580 14785 3606
rect 14800 3601 14830 3612
rect 14862 3608 14924 3624
rect 14862 3606 14908 3608
rect 14862 3590 14924 3606
rect 14936 3590 14942 3638
rect 14945 3630 15025 3638
rect 14945 3628 14964 3630
rect 14979 3628 15013 3630
rect 14945 3612 15025 3628
rect 14945 3590 14964 3612
rect 14979 3596 15009 3612
rect 15037 3606 15043 3680
rect 15046 3606 15065 3750
rect 15080 3606 15086 3750
rect 15095 3680 15108 3750
rect 15160 3746 15182 3750
rect 15153 3724 15182 3738
rect 15235 3724 15251 3738
rect 15289 3734 15295 3736
rect 15302 3734 15410 3750
rect 15417 3734 15423 3736
rect 15431 3734 15446 3750
rect 15512 3744 15531 3747
rect 15153 3722 15251 3724
rect 15278 3722 15446 3734
rect 15461 3724 15477 3738
rect 15512 3725 15534 3744
rect 15544 3738 15560 3739
rect 15543 3736 15560 3738
rect 15544 3731 15560 3736
rect 15534 3724 15540 3725
rect 15543 3724 15572 3731
rect 15461 3723 15572 3724
rect 15461 3722 15578 3723
rect 15137 3714 15188 3722
rect 15235 3714 15269 3722
rect 15137 3702 15162 3714
rect 15169 3702 15188 3714
rect 15242 3712 15269 3714
rect 15278 3712 15499 3722
rect 15534 3719 15540 3722
rect 15242 3708 15499 3712
rect 15137 3694 15188 3702
rect 15235 3694 15499 3708
rect 15543 3714 15578 3722
rect 15089 3646 15108 3680
rect 15153 3686 15182 3694
rect 15153 3680 15170 3686
rect 15153 3678 15187 3680
rect 15235 3678 15251 3694
rect 15252 3684 15460 3694
rect 15461 3684 15477 3694
rect 15525 3690 15540 3705
rect 15543 3702 15544 3714
rect 15551 3702 15578 3714
rect 15543 3694 15578 3702
rect 15543 3693 15572 3694
rect 15263 3680 15477 3684
rect 15278 3678 15477 3680
rect 15512 3680 15525 3690
rect 15543 3680 15560 3693
rect 15512 3678 15560 3680
rect 15154 3674 15187 3678
rect 15150 3672 15187 3674
rect 15150 3671 15217 3672
rect 15150 3666 15181 3671
rect 15187 3666 15217 3671
rect 15150 3662 15217 3666
rect 15123 3659 15217 3662
rect 15123 3652 15172 3659
rect 15123 3646 15153 3652
rect 15172 3647 15177 3652
rect 15089 3630 15169 3646
rect 15181 3638 15217 3659
rect 15278 3654 15467 3678
rect 15512 3677 15559 3678
rect 15525 3672 15559 3677
rect 15293 3651 15467 3654
rect 15286 3648 15467 3651
rect 15495 3671 15559 3672
rect 15089 3628 15108 3630
rect 15123 3628 15157 3630
rect 15089 3612 15169 3628
rect 15089 3606 15108 3612
rect 14805 3580 14908 3590
rect 14759 3578 14908 3580
rect 14929 3578 14964 3590
rect 14598 3576 14760 3578
rect 14610 3556 14629 3576
rect 14644 3574 14674 3576
rect 14493 3548 14534 3556
rect 14616 3552 14629 3556
rect 14681 3560 14760 3576
rect 14792 3576 14964 3578
rect 14792 3560 14871 3576
rect 14878 3574 14908 3576
rect 14456 3538 14485 3548
rect 14499 3538 14528 3548
rect 14543 3538 14573 3552
rect 14616 3538 14659 3552
rect 14681 3548 14871 3560
rect 14936 3556 14942 3576
rect 14666 3538 14696 3548
rect 14697 3538 14855 3548
rect 14859 3538 14889 3548
rect 14893 3538 14923 3552
rect 14951 3538 14964 3576
rect 15036 3590 15065 3606
rect 15079 3590 15108 3606
rect 15123 3596 15153 3612
rect 15181 3590 15187 3638
rect 15190 3632 15209 3638
rect 15224 3632 15254 3640
rect 15190 3624 15254 3632
rect 15190 3608 15270 3624
rect 15286 3617 15348 3648
rect 15364 3617 15426 3648
rect 15495 3646 15544 3671
rect 15559 3646 15589 3662
rect 15458 3632 15488 3640
rect 15495 3638 15605 3646
rect 15458 3624 15503 3632
rect 15190 3606 15209 3608
rect 15224 3606 15270 3608
rect 15190 3590 15270 3606
rect 15297 3604 15332 3617
rect 15373 3614 15410 3617
rect 15373 3612 15415 3614
rect 15302 3601 15332 3604
rect 15311 3597 15318 3601
rect 15318 3596 15319 3597
rect 15277 3590 15287 3596
rect 15036 3582 15071 3590
rect 15036 3556 15037 3582
rect 15044 3556 15071 3582
rect 14979 3538 15009 3552
rect 15036 3548 15071 3556
rect 15073 3582 15114 3590
rect 15073 3556 15088 3582
rect 15095 3556 15114 3582
rect 15178 3578 15209 3590
rect 15224 3578 15327 3590
rect 15339 3580 15365 3606
rect 15380 3601 15410 3612
rect 15442 3608 15504 3624
rect 15442 3606 15488 3608
rect 15442 3590 15504 3606
rect 15516 3590 15522 3638
rect 15525 3630 15605 3638
rect 15525 3628 15544 3630
rect 15559 3628 15593 3630
rect 15525 3612 15605 3628
rect 15525 3590 15544 3612
rect 15559 3596 15589 3612
rect 15617 3606 15623 3680
rect 15626 3606 15645 3750
rect 15660 3606 15666 3750
rect 15675 3680 15688 3750
rect 15740 3746 15762 3750
rect 15733 3724 15762 3738
rect 15815 3724 15831 3738
rect 15869 3734 15875 3736
rect 15882 3734 15990 3750
rect 15997 3734 16003 3736
rect 16011 3734 16026 3750
rect 16092 3744 16111 3747
rect 15733 3722 15831 3724
rect 15858 3722 16026 3734
rect 16041 3724 16057 3738
rect 16092 3725 16114 3744
rect 16124 3738 16140 3739
rect 16123 3736 16140 3738
rect 16124 3731 16140 3736
rect 16114 3724 16120 3725
rect 16123 3724 16152 3731
rect 16041 3723 16152 3724
rect 16041 3722 16158 3723
rect 15717 3714 15768 3722
rect 15815 3714 15849 3722
rect 15717 3702 15742 3714
rect 15749 3702 15768 3714
rect 15822 3712 15849 3714
rect 15858 3712 16079 3722
rect 16114 3719 16120 3722
rect 15822 3708 16079 3712
rect 15717 3694 15768 3702
rect 15815 3694 16079 3708
rect 16123 3714 16158 3722
rect 15669 3646 15688 3680
rect 15733 3686 15762 3694
rect 15733 3680 15750 3686
rect 15733 3678 15767 3680
rect 15815 3678 15831 3694
rect 15832 3684 16040 3694
rect 16041 3684 16057 3694
rect 16105 3690 16120 3705
rect 16123 3702 16124 3714
rect 16131 3702 16158 3714
rect 16123 3694 16158 3702
rect 16123 3693 16152 3694
rect 15843 3680 16057 3684
rect 15858 3678 16057 3680
rect 16092 3680 16105 3690
rect 16123 3680 16140 3693
rect 16092 3678 16140 3680
rect 15734 3674 15767 3678
rect 15730 3672 15767 3674
rect 15730 3671 15797 3672
rect 15730 3666 15761 3671
rect 15767 3666 15797 3671
rect 15730 3662 15797 3666
rect 15703 3659 15797 3662
rect 15703 3652 15752 3659
rect 15703 3646 15733 3652
rect 15752 3647 15757 3652
rect 15669 3630 15749 3646
rect 15761 3638 15797 3659
rect 15858 3654 16047 3678
rect 16092 3677 16139 3678
rect 16105 3672 16139 3677
rect 15873 3651 16047 3654
rect 15866 3648 16047 3651
rect 16075 3671 16139 3672
rect 15669 3628 15688 3630
rect 15703 3628 15737 3630
rect 15669 3612 15749 3628
rect 15669 3606 15688 3612
rect 15385 3580 15488 3590
rect 15339 3578 15488 3580
rect 15509 3578 15544 3590
rect 15178 3576 15340 3578
rect 15190 3556 15209 3576
rect 15224 3574 15254 3576
rect 15073 3548 15114 3556
rect 15196 3552 15209 3556
rect 15261 3560 15340 3576
rect 15372 3576 15544 3578
rect 15372 3560 15451 3576
rect 15458 3574 15488 3576
rect 15036 3538 15065 3548
rect 15079 3538 15108 3548
rect 15123 3538 15153 3552
rect 15196 3538 15239 3552
rect 15261 3548 15451 3560
rect 15516 3556 15522 3576
rect 15246 3538 15276 3548
rect 15277 3538 15435 3548
rect 15439 3538 15469 3548
rect 15473 3538 15503 3552
rect 15531 3538 15544 3576
rect 15616 3590 15645 3606
rect 15659 3590 15688 3606
rect 15703 3596 15733 3612
rect 15761 3590 15767 3638
rect 15770 3632 15789 3638
rect 15804 3632 15834 3640
rect 15770 3624 15834 3632
rect 15770 3608 15850 3624
rect 15866 3617 15928 3648
rect 15944 3617 16006 3648
rect 16075 3646 16124 3671
rect 16139 3646 16169 3662
rect 16038 3632 16068 3640
rect 16075 3638 16185 3646
rect 16038 3624 16083 3632
rect 15770 3606 15789 3608
rect 15804 3606 15850 3608
rect 15770 3590 15850 3606
rect 15877 3604 15912 3617
rect 15953 3614 15990 3617
rect 15953 3612 15995 3614
rect 15882 3601 15912 3604
rect 15891 3597 15898 3601
rect 15898 3596 15899 3597
rect 15857 3590 15867 3596
rect 15616 3582 15651 3590
rect 15616 3556 15617 3582
rect 15624 3556 15651 3582
rect 15559 3538 15589 3552
rect 15616 3548 15651 3556
rect 15653 3582 15694 3590
rect 15653 3556 15668 3582
rect 15675 3556 15694 3582
rect 15758 3578 15789 3590
rect 15804 3578 15907 3590
rect 15919 3580 15945 3606
rect 15960 3601 15990 3612
rect 16022 3608 16084 3624
rect 16022 3606 16068 3608
rect 16022 3590 16084 3606
rect 16096 3590 16102 3638
rect 16105 3630 16185 3638
rect 16105 3628 16124 3630
rect 16139 3628 16173 3630
rect 16105 3612 16185 3628
rect 16105 3590 16124 3612
rect 16139 3596 16169 3612
rect 16197 3606 16203 3680
rect 16206 3606 16225 3750
rect 16240 3606 16246 3750
rect 16255 3680 16268 3750
rect 16320 3746 16342 3750
rect 16313 3724 16342 3738
rect 16395 3724 16411 3738
rect 16449 3734 16455 3736
rect 16462 3734 16570 3750
rect 16577 3734 16583 3736
rect 16591 3734 16606 3750
rect 16672 3744 16691 3747
rect 16313 3722 16411 3724
rect 16438 3722 16606 3734
rect 16621 3724 16637 3738
rect 16672 3725 16694 3744
rect 16704 3738 16720 3739
rect 16703 3736 16720 3738
rect 16704 3731 16720 3736
rect 16694 3724 16700 3725
rect 16703 3724 16732 3731
rect 16621 3723 16732 3724
rect 16621 3722 16738 3723
rect 16297 3714 16348 3722
rect 16395 3714 16429 3722
rect 16297 3702 16322 3714
rect 16329 3702 16348 3714
rect 16402 3712 16429 3714
rect 16438 3712 16659 3722
rect 16694 3719 16700 3722
rect 16402 3708 16659 3712
rect 16297 3694 16348 3702
rect 16395 3694 16659 3708
rect 16703 3714 16738 3722
rect 16249 3646 16268 3680
rect 16313 3686 16342 3694
rect 16313 3680 16330 3686
rect 16313 3678 16347 3680
rect 16395 3678 16411 3694
rect 16412 3684 16620 3694
rect 16621 3684 16637 3694
rect 16685 3690 16700 3705
rect 16703 3702 16704 3714
rect 16711 3702 16738 3714
rect 16703 3694 16738 3702
rect 16703 3693 16732 3694
rect 16423 3680 16637 3684
rect 16438 3678 16637 3680
rect 16672 3680 16685 3690
rect 16703 3680 16720 3693
rect 16672 3678 16720 3680
rect 16314 3674 16347 3678
rect 16310 3672 16347 3674
rect 16310 3671 16377 3672
rect 16310 3666 16341 3671
rect 16347 3666 16377 3671
rect 16310 3662 16377 3666
rect 16283 3659 16377 3662
rect 16283 3652 16332 3659
rect 16283 3646 16313 3652
rect 16332 3647 16337 3652
rect 16249 3630 16329 3646
rect 16341 3638 16377 3659
rect 16438 3654 16627 3678
rect 16672 3677 16719 3678
rect 16685 3672 16719 3677
rect 16453 3651 16627 3654
rect 16446 3648 16627 3651
rect 16655 3671 16719 3672
rect 16249 3628 16268 3630
rect 16283 3628 16317 3630
rect 16249 3612 16329 3628
rect 16249 3606 16268 3612
rect 15965 3580 16068 3590
rect 15919 3578 16068 3580
rect 16089 3578 16124 3590
rect 15758 3576 15920 3578
rect 15770 3556 15789 3576
rect 15804 3574 15834 3576
rect 15653 3548 15694 3556
rect 15776 3552 15789 3556
rect 15841 3560 15920 3576
rect 15952 3576 16124 3578
rect 15952 3560 16031 3576
rect 16038 3574 16068 3576
rect 15616 3538 15645 3548
rect 15659 3538 15688 3548
rect 15703 3538 15733 3552
rect 15776 3538 15819 3552
rect 15841 3548 16031 3560
rect 16096 3556 16102 3576
rect 15826 3538 15856 3548
rect 15857 3538 16015 3548
rect 16019 3538 16049 3548
rect 16053 3538 16083 3552
rect 16111 3538 16124 3576
rect 16196 3590 16225 3606
rect 16239 3590 16268 3606
rect 16283 3596 16313 3612
rect 16341 3590 16347 3638
rect 16350 3632 16369 3638
rect 16384 3632 16414 3640
rect 16350 3624 16414 3632
rect 16350 3608 16430 3624
rect 16446 3617 16508 3648
rect 16524 3617 16586 3648
rect 16655 3646 16704 3671
rect 16719 3646 16749 3662
rect 16618 3632 16648 3640
rect 16655 3638 16765 3646
rect 16618 3624 16663 3632
rect 16350 3606 16369 3608
rect 16384 3606 16430 3608
rect 16350 3590 16430 3606
rect 16457 3604 16492 3617
rect 16533 3614 16570 3617
rect 16533 3612 16575 3614
rect 16462 3601 16492 3604
rect 16471 3597 16478 3601
rect 16478 3596 16479 3597
rect 16437 3590 16447 3596
rect 16196 3582 16231 3590
rect 16196 3556 16197 3582
rect 16204 3556 16231 3582
rect 16139 3538 16169 3552
rect 16196 3548 16231 3556
rect 16233 3582 16274 3590
rect 16233 3556 16248 3582
rect 16255 3556 16274 3582
rect 16338 3578 16369 3590
rect 16384 3578 16487 3590
rect 16499 3580 16525 3606
rect 16540 3601 16570 3612
rect 16602 3608 16664 3624
rect 16602 3606 16648 3608
rect 16602 3590 16664 3606
rect 16676 3590 16682 3638
rect 16685 3630 16765 3638
rect 16685 3628 16704 3630
rect 16719 3628 16753 3630
rect 16685 3612 16765 3628
rect 16685 3590 16704 3612
rect 16719 3596 16749 3612
rect 16777 3606 16783 3680
rect 16786 3606 16805 3750
rect 16820 3606 16826 3750
rect 16835 3680 16848 3750
rect 16900 3746 16922 3750
rect 16893 3724 16922 3738
rect 16975 3724 16991 3738
rect 17029 3734 17035 3736
rect 17042 3734 17150 3750
rect 17157 3734 17163 3736
rect 17171 3734 17186 3750
rect 17252 3744 17271 3747
rect 16893 3722 16991 3724
rect 17018 3722 17186 3734
rect 17201 3724 17217 3738
rect 17252 3725 17274 3744
rect 17284 3738 17300 3739
rect 17283 3736 17300 3738
rect 17284 3731 17300 3736
rect 17274 3724 17280 3725
rect 17283 3724 17312 3731
rect 17201 3723 17312 3724
rect 17201 3722 17318 3723
rect 16877 3714 16928 3722
rect 16975 3714 17009 3722
rect 16877 3702 16902 3714
rect 16909 3702 16928 3714
rect 16982 3712 17009 3714
rect 17018 3712 17239 3722
rect 17274 3719 17280 3722
rect 16982 3708 17239 3712
rect 16877 3694 16928 3702
rect 16975 3694 17239 3708
rect 17283 3714 17318 3722
rect 16829 3646 16848 3680
rect 16893 3686 16922 3694
rect 16893 3680 16910 3686
rect 16893 3678 16927 3680
rect 16975 3678 16991 3694
rect 16992 3684 17200 3694
rect 17201 3684 17217 3694
rect 17265 3690 17280 3705
rect 17283 3702 17284 3714
rect 17291 3702 17318 3714
rect 17283 3694 17318 3702
rect 17283 3693 17312 3694
rect 17003 3680 17217 3684
rect 17018 3678 17217 3680
rect 17252 3680 17265 3690
rect 17283 3680 17300 3693
rect 17252 3678 17300 3680
rect 16894 3674 16927 3678
rect 16890 3672 16927 3674
rect 16890 3671 16957 3672
rect 16890 3666 16921 3671
rect 16927 3666 16957 3671
rect 16890 3662 16957 3666
rect 16863 3659 16957 3662
rect 16863 3652 16912 3659
rect 16863 3646 16893 3652
rect 16912 3647 16917 3652
rect 16829 3630 16909 3646
rect 16921 3638 16957 3659
rect 17018 3654 17207 3678
rect 17252 3677 17299 3678
rect 17265 3672 17299 3677
rect 17033 3651 17207 3654
rect 17026 3648 17207 3651
rect 17235 3671 17299 3672
rect 16829 3628 16848 3630
rect 16863 3628 16897 3630
rect 16829 3612 16909 3628
rect 16829 3606 16848 3612
rect 16545 3580 16648 3590
rect 16499 3578 16648 3580
rect 16669 3578 16704 3590
rect 16338 3576 16500 3578
rect 16350 3556 16369 3576
rect 16384 3574 16414 3576
rect 16233 3548 16274 3556
rect 16356 3552 16369 3556
rect 16421 3560 16500 3576
rect 16532 3576 16704 3578
rect 16532 3560 16611 3576
rect 16618 3574 16648 3576
rect 16196 3538 16225 3548
rect 16239 3538 16268 3548
rect 16283 3538 16313 3552
rect 16356 3538 16399 3552
rect 16421 3548 16611 3560
rect 16676 3556 16682 3576
rect 16406 3538 16436 3548
rect 16437 3538 16595 3548
rect 16599 3538 16629 3548
rect 16633 3538 16663 3552
rect 16691 3538 16704 3576
rect 16776 3590 16805 3606
rect 16819 3590 16848 3606
rect 16863 3596 16893 3612
rect 16921 3590 16927 3638
rect 16930 3632 16949 3638
rect 16964 3632 16994 3640
rect 16930 3624 16994 3632
rect 16930 3608 17010 3624
rect 17026 3617 17088 3648
rect 17104 3617 17166 3648
rect 17235 3646 17284 3671
rect 17299 3646 17329 3662
rect 17198 3632 17228 3640
rect 17235 3638 17345 3646
rect 17198 3624 17243 3632
rect 16930 3606 16949 3608
rect 16964 3606 17010 3608
rect 16930 3590 17010 3606
rect 17037 3604 17072 3617
rect 17113 3614 17150 3617
rect 17113 3612 17155 3614
rect 17042 3601 17072 3604
rect 17051 3597 17058 3601
rect 17058 3596 17059 3597
rect 17017 3590 17027 3596
rect 16776 3582 16811 3590
rect 16776 3556 16777 3582
rect 16784 3556 16811 3582
rect 16719 3538 16749 3552
rect 16776 3548 16811 3556
rect 16813 3582 16854 3590
rect 16813 3556 16828 3582
rect 16835 3556 16854 3582
rect 16918 3578 16949 3590
rect 16964 3578 17067 3590
rect 17079 3580 17105 3606
rect 17120 3601 17150 3612
rect 17182 3608 17244 3624
rect 17182 3606 17228 3608
rect 17182 3590 17244 3606
rect 17256 3590 17262 3638
rect 17265 3630 17345 3638
rect 17265 3628 17284 3630
rect 17299 3628 17333 3630
rect 17265 3612 17345 3628
rect 17265 3590 17284 3612
rect 17299 3596 17329 3612
rect 17357 3606 17363 3680
rect 17366 3606 17385 3750
rect 17400 3606 17406 3750
rect 17415 3680 17428 3750
rect 17480 3746 17502 3750
rect 17473 3724 17502 3738
rect 17555 3724 17571 3738
rect 17609 3734 17615 3736
rect 17622 3734 17730 3750
rect 17737 3734 17743 3736
rect 17751 3734 17766 3750
rect 17832 3744 17851 3747
rect 17473 3722 17571 3724
rect 17598 3722 17766 3734
rect 17781 3724 17797 3738
rect 17832 3725 17854 3744
rect 17864 3738 17880 3739
rect 17863 3736 17880 3738
rect 17864 3731 17880 3736
rect 17854 3724 17860 3725
rect 17863 3724 17892 3731
rect 17781 3723 17892 3724
rect 17781 3722 17898 3723
rect 17457 3714 17508 3722
rect 17555 3714 17589 3722
rect 17457 3702 17482 3714
rect 17489 3702 17508 3714
rect 17562 3712 17589 3714
rect 17598 3712 17819 3722
rect 17854 3719 17860 3722
rect 17562 3708 17819 3712
rect 17457 3694 17508 3702
rect 17555 3694 17819 3708
rect 17863 3714 17898 3722
rect 17409 3646 17428 3680
rect 17473 3686 17502 3694
rect 17473 3680 17490 3686
rect 17473 3678 17507 3680
rect 17555 3678 17571 3694
rect 17572 3684 17780 3694
rect 17781 3684 17797 3694
rect 17845 3690 17860 3705
rect 17863 3702 17864 3714
rect 17871 3702 17898 3714
rect 17863 3694 17898 3702
rect 17863 3693 17892 3694
rect 17583 3680 17797 3684
rect 17598 3678 17797 3680
rect 17832 3680 17845 3690
rect 17863 3680 17880 3693
rect 17832 3678 17880 3680
rect 17474 3674 17507 3678
rect 17470 3672 17507 3674
rect 17470 3671 17537 3672
rect 17470 3666 17501 3671
rect 17507 3666 17537 3671
rect 17470 3662 17537 3666
rect 17443 3659 17537 3662
rect 17443 3652 17492 3659
rect 17443 3646 17473 3652
rect 17492 3647 17497 3652
rect 17409 3630 17489 3646
rect 17501 3638 17537 3659
rect 17598 3654 17787 3678
rect 17832 3677 17879 3678
rect 17845 3672 17879 3677
rect 17613 3651 17787 3654
rect 17606 3648 17787 3651
rect 17815 3671 17879 3672
rect 17409 3628 17428 3630
rect 17443 3628 17477 3630
rect 17409 3612 17489 3628
rect 17409 3606 17428 3612
rect 17125 3580 17228 3590
rect 17079 3578 17228 3580
rect 17249 3578 17284 3590
rect 16918 3576 17080 3578
rect 16930 3556 16949 3576
rect 16964 3574 16994 3576
rect 16813 3548 16854 3556
rect 16936 3552 16949 3556
rect 17001 3560 17080 3576
rect 17112 3576 17284 3578
rect 17112 3560 17191 3576
rect 17198 3574 17228 3576
rect 16776 3538 16805 3548
rect 16819 3538 16848 3548
rect 16863 3538 16893 3552
rect 16936 3538 16979 3552
rect 17001 3548 17191 3560
rect 17256 3556 17262 3576
rect 16986 3538 17016 3548
rect 17017 3538 17175 3548
rect 17179 3538 17209 3548
rect 17213 3538 17243 3552
rect 17271 3538 17284 3576
rect 17356 3590 17385 3606
rect 17399 3590 17428 3606
rect 17443 3596 17473 3612
rect 17501 3590 17507 3638
rect 17510 3632 17529 3638
rect 17544 3632 17574 3640
rect 17510 3624 17574 3632
rect 17510 3608 17590 3624
rect 17606 3617 17668 3648
rect 17684 3617 17746 3648
rect 17815 3646 17864 3671
rect 17879 3646 17909 3662
rect 17778 3632 17808 3640
rect 17815 3638 17925 3646
rect 17778 3624 17823 3632
rect 17510 3606 17529 3608
rect 17544 3606 17590 3608
rect 17510 3590 17590 3606
rect 17617 3604 17652 3617
rect 17693 3614 17730 3617
rect 17693 3612 17735 3614
rect 17622 3601 17652 3604
rect 17631 3597 17638 3601
rect 17638 3596 17639 3597
rect 17597 3590 17607 3596
rect 17356 3582 17391 3590
rect 17356 3556 17357 3582
rect 17364 3556 17391 3582
rect 17299 3538 17329 3552
rect 17356 3548 17391 3556
rect 17393 3582 17434 3590
rect 17393 3556 17408 3582
rect 17415 3556 17434 3582
rect 17498 3578 17529 3590
rect 17544 3578 17647 3590
rect 17659 3580 17685 3606
rect 17700 3601 17730 3612
rect 17762 3608 17824 3624
rect 17762 3606 17808 3608
rect 17762 3590 17824 3606
rect 17836 3590 17842 3638
rect 17845 3630 17925 3638
rect 17845 3628 17864 3630
rect 17879 3628 17913 3630
rect 17845 3612 17925 3628
rect 17845 3590 17864 3612
rect 17879 3596 17909 3612
rect 17937 3606 17943 3680
rect 17946 3606 17965 3750
rect 17980 3606 17986 3750
rect 17995 3680 18008 3750
rect 18060 3746 18082 3750
rect 18053 3724 18082 3738
rect 18135 3724 18151 3738
rect 18189 3734 18195 3736
rect 18202 3734 18310 3750
rect 18317 3734 18323 3736
rect 18331 3734 18346 3750
rect 18412 3744 18431 3747
rect 18053 3722 18151 3724
rect 18178 3722 18346 3734
rect 18361 3724 18377 3738
rect 18412 3725 18434 3744
rect 18444 3738 18460 3739
rect 18443 3736 18460 3738
rect 18444 3731 18460 3736
rect 18434 3724 18440 3725
rect 18443 3724 18472 3731
rect 18361 3723 18472 3724
rect 18361 3722 18478 3723
rect 18037 3714 18088 3722
rect 18135 3714 18169 3722
rect 18037 3702 18062 3714
rect 18069 3702 18088 3714
rect 18142 3712 18169 3714
rect 18178 3712 18399 3722
rect 18434 3719 18440 3722
rect 18142 3708 18399 3712
rect 18037 3694 18088 3702
rect 18135 3694 18399 3708
rect 18443 3714 18478 3722
rect 17989 3646 18008 3680
rect 18053 3686 18082 3694
rect 18053 3680 18070 3686
rect 18053 3678 18087 3680
rect 18135 3678 18151 3694
rect 18152 3684 18360 3694
rect 18361 3684 18377 3694
rect 18425 3690 18440 3705
rect 18443 3702 18444 3714
rect 18451 3702 18478 3714
rect 18443 3694 18478 3702
rect 18443 3693 18472 3694
rect 18163 3680 18377 3684
rect 18178 3678 18377 3680
rect 18412 3680 18425 3690
rect 18443 3680 18460 3693
rect 18412 3678 18460 3680
rect 18054 3674 18087 3678
rect 18050 3672 18087 3674
rect 18050 3671 18117 3672
rect 18050 3666 18081 3671
rect 18087 3666 18117 3671
rect 18050 3662 18117 3666
rect 18023 3659 18117 3662
rect 18023 3652 18072 3659
rect 18023 3646 18053 3652
rect 18072 3647 18077 3652
rect 17989 3630 18069 3646
rect 18081 3638 18117 3659
rect 18178 3654 18367 3678
rect 18412 3677 18459 3678
rect 18425 3672 18459 3677
rect 18193 3651 18367 3654
rect 18186 3648 18367 3651
rect 18395 3671 18459 3672
rect 17989 3628 18008 3630
rect 18023 3628 18057 3630
rect 17989 3612 18069 3628
rect 17989 3606 18008 3612
rect 17705 3580 17808 3590
rect 17659 3578 17808 3580
rect 17829 3578 17864 3590
rect 17498 3576 17660 3578
rect 17510 3556 17529 3576
rect 17544 3574 17574 3576
rect 17393 3548 17434 3556
rect 17516 3552 17529 3556
rect 17581 3560 17660 3576
rect 17692 3576 17864 3578
rect 17692 3560 17771 3576
rect 17778 3574 17808 3576
rect 17356 3538 17385 3548
rect 17399 3538 17428 3548
rect 17443 3538 17473 3552
rect 17516 3538 17559 3552
rect 17581 3548 17771 3560
rect 17836 3556 17842 3576
rect 17566 3538 17596 3548
rect 17597 3538 17755 3548
rect 17759 3538 17789 3548
rect 17793 3538 17823 3552
rect 17851 3538 17864 3576
rect 17936 3590 17965 3606
rect 17979 3590 18008 3606
rect 18023 3596 18053 3612
rect 18081 3590 18087 3638
rect 18090 3632 18109 3638
rect 18124 3632 18154 3640
rect 18090 3624 18154 3632
rect 18090 3608 18170 3624
rect 18186 3617 18248 3648
rect 18264 3617 18326 3648
rect 18395 3646 18444 3671
rect 18459 3646 18489 3662
rect 18358 3632 18388 3640
rect 18395 3638 18505 3646
rect 18358 3624 18403 3632
rect 18090 3606 18109 3608
rect 18124 3606 18170 3608
rect 18090 3590 18170 3606
rect 18197 3604 18232 3617
rect 18273 3614 18310 3617
rect 18273 3612 18315 3614
rect 18202 3601 18232 3604
rect 18211 3597 18218 3601
rect 18218 3596 18219 3597
rect 18177 3590 18187 3596
rect 17936 3582 17971 3590
rect 17936 3556 17937 3582
rect 17944 3556 17971 3582
rect 17879 3538 17909 3552
rect 17936 3548 17971 3556
rect 17973 3582 18014 3590
rect 17973 3556 17988 3582
rect 17995 3556 18014 3582
rect 18078 3578 18109 3590
rect 18124 3578 18227 3590
rect 18239 3580 18265 3606
rect 18280 3601 18310 3612
rect 18342 3608 18404 3624
rect 18342 3606 18388 3608
rect 18342 3590 18404 3606
rect 18416 3590 18422 3638
rect 18425 3630 18505 3638
rect 18425 3628 18444 3630
rect 18459 3628 18493 3630
rect 18425 3612 18505 3628
rect 18425 3590 18444 3612
rect 18459 3596 18489 3612
rect 18517 3606 18523 3680
rect 18532 3606 18545 3750
rect 18285 3580 18388 3590
rect 18239 3578 18388 3580
rect 18409 3578 18444 3590
rect 18078 3576 18240 3578
rect 18090 3556 18109 3576
rect 18124 3574 18154 3576
rect 17973 3548 18014 3556
rect 18096 3552 18109 3556
rect 18161 3560 18240 3576
rect 18272 3576 18444 3578
rect 18272 3560 18351 3576
rect 18358 3574 18388 3576
rect 17936 3538 17965 3548
rect 17979 3538 18008 3548
rect 18023 3538 18053 3552
rect 18096 3538 18139 3552
rect 18161 3548 18351 3560
rect 18416 3556 18422 3576
rect 18146 3538 18176 3548
rect 18177 3538 18335 3548
rect 18339 3538 18369 3548
rect 18373 3538 18403 3552
rect 18431 3538 18444 3576
rect 18516 3590 18545 3606
rect 18516 3582 18551 3590
rect 18516 3556 18517 3582
rect 18524 3556 18551 3582
rect 18459 3538 18489 3552
rect 18516 3548 18551 3556
rect 18516 3538 18545 3548
rect -1 3532 18545 3538
rect 0 3524 18545 3532
rect 15 3494 28 3524
rect 43 3510 73 3524
rect 116 3510 159 3524
rect 166 3510 386 3524
rect 393 3510 423 3524
rect 83 3496 98 3508
rect 117 3496 130 3510
rect 198 3506 351 3510
rect 80 3494 102 3496
rect 180 3494 372 3506
rect 451 3494 464 3524
rect 479 3510 509 3524
rect 546 3494 565 3524
rect 580 3494 586 3524
rect 595 3494 608 3524
rect 623 3510 653 3524
rect 696 3510 739 3524
rect 746 3510 966 3524
rect 973 3510 1003 3524
rect 663 3496 678 3508
rect 697 3496 710 3510
rect 778 3506 931 3510
rect 660 3494 682 3496
rect 760 3494 952 3506
rect 1031 3494 1044 3524
rect 1059 3510 1089 3524
rect 1126 3494 1145 3524
rect 1160 3494 1166 3524
rect 1175 3494 1188 3524
rect 1203 3510 1233 3524
rect 1276 3510 1319 3524
rect 1326 3510 1546 3524
rect 1553 3510 1583 3524
rect 1243 3496 1258 3508
rect 1277 3496 1290 3510
rect 1358 3506 1511 3510
rect 1240 3494 1262 3496
rect 1340 3494 1532 3506
rect 1611 3494 1624 3524
rect 1639 3510 1669 3524
rect 1706 3494 1725 3524
rect 1740 3494 1746 3524
rect 1755 3494 1768 3524
rect 1783 3510 1813 3524
rect 1856 3510 1899 3524
rect 1906 3510 2126 3524
rect 2133 3510 2163 3524
rect 1823 3496 1838 3508
rect 1857 3496 1870 3510
rect 1938 3506 2091 3510
rect 1820 3494 1842 3496
rect 1920 3494 2112 3506
rect 2191 3494 2204 3524
rect 2219 3510 2249 3524
rect 2286 3494 2305 3524
rect 2320 3494 2326 3524
rect 2335 3494 2348 3524
rect 2363 3510 2393 3524
rect 2436 3510 2479 3524
rect 2486 3510 2706 3524
rect 2713 3510 2743 3524
rect 2403 3496 2418 3508
rect 2437 3496 2450 3510
rect 2518 3506 2671 3510
rect 2400 3494 2422 3496
rect 2500 3494 2692 3506
rect 2771 3494 2784 3524
rect 2799 3510 2829 3524
rect 2866 3494 2885 3524
rect 2900 3494 2906 3524
rect 2915 3494 2928 3524
rect 2943 3510 2973 3524
rect 3016 3510 3059 3524
rect 3066 3510 3286 3524
rect 3293 3510 3323 3524
rect 2983 3496 2998 3508
rect 3017 3496 3030 3510
rect 3098 3506 3251 3510
rect 2980 3494 3002 3496
rect 3080 3494 3272 3506
rect 3351 3494 3364 3524
rect 3379 3510 3409 3524
rect 3446 3494 3465 3524
rect 3480 3494 3486 3524
rect 3495 3494 3508 3524
rect 3523 3510 3553 3524
rect 3596 3510 3639 3524
rect 3646 3510 3866 3524
rect 3873 3510 3903 3524
rect 3563 3496 3578 3508
rect 3597 3496 3610 3510
rect 3678 3506 3831 3510
rect 3560 3494 3582 3496
rect 3660 3494 3852 3506
rect 3931 3494 3944 3524
rect 3959 3510 3989 3524
rect 4026 3494 4045 3524
rect 4060 3494 4066 3524
rect 4075 3494 4088 3524
rect 4103 3510 4133 3524
rect 4176 3510 4219 3524
rect 4226 3510 4446 3524
rect 4453 3510 4483 3524
rect 4143 3496 4158 3508
rect 4177 3496 4190 3510
rect 4258 3506 4411 3510
rect 4140 3494 4162 3496
rect 4240 3494 4432 3506
rect 4511 3494 4524 3524
rect 4539 3510 4569 3524
rect 4606 3494 4625 3524
rect 4640 3494 4646 3524
rect 4655 3494 4668 3524
rect 4683 3510 4713 3524
rect 4756 3510 4799 3524
rect 4806 3510 5026 3524
rect 5033 3510 5063 3524
rect 4723 3496 4738 3508
rect 4757 3496 4770 3510
rect 4838 3506 4991 3510
rect 4720 3494 4742 3496
rect 4820 3494 5012 3506
rect 5091 3494 5104 3524
rect 5119 3510 5149 3524
rect 5186 3494 5205 3524
rect 5220 3494 5226 3524
rect 5235 3494 5248 3524
rect 5263 3510 5293 3524
rect 5336 3510 5379 3524
rect 5386 3510 5606 3524
rect 5613 3510 5643 3524
rect 5303 3496 5318 3508
rect 5337 3496 5350 3510
rect 5418 3506 5571 3510
rect 5300 3494 5322 3496
rect 5400 3494 5592 3506
rect 5671 3494 5684 3524
rect 5699 3510 5729 3524
rect 5766 3494 5785 3524
rect 5800 3494 5806 3524
rect 5815 3494 5828 3524
rect 5843 3510 5873 3524
rect 5916 3510 5959 3524
rect 5966 3510 6186 3524
rect 6193 3510 6223 3524
rect 5883 3496 5898 3508
rect 5917 3496 5930 3510
rect 5998 3506 6151 3510
rect 5880 3494 5902 3496
rect 5980 3494 6172 3506
rect 6251 3494 6264 3524
rect 6279 3510 6309 3524
rect 6346 3494 6365 3524
rect 6380 3494 6386 3524
rect 6395 3494 6408 3524
rect 6423 3510 6453 3524
rect 6496 3510 6539 3524
rect 6546 3510 6766 3524
rect 6773 3510 6803 3524
rect 6463 3496 6478 3508
rect 6497 3496 6510 3510
rect 6578 3506 6731 3510
rect 6460 3494 6482 3496
rect 6560 3494 6752 3506
rect 6831 3494 6844 3524
rect 6859 3510 6889 3524
rect 6926 3494 6945 3524
rect 6960 3494 6966 3524
rect 6975 3494 6988 3524
rect 7003 3510 7033 3524
rect 7076 3510 7119 3524
rect 7126 3510 7346 3524
rect 7353 3510 7383 3524
rect 7043 3496 7058 3508
rect 7077 3496 7090 3510
rect 7158 3506 7311 3510
rect 7040 3494 7062 3496
rect 7140 3494 7332 3506
rect 7411 3494 7424 3524
rect 7439 3510 7469 3524
rect 7506 3494 7525 3524
rect 7540 3494 7546 3524
rect 7555 3494 7568 3524
rect 7583 3510 7613 3524
rect 7656 3510 7699 3524
rect 7706 3510 7926 3524
rect 7933 3510 7963 3524
rect 7623 3496 7638 3508
rect 7657 3496 7670 3510
rect 7738 3506 7891 3510
rect 7620 3494 7642 3496
rect 7720 3494 7912 3506
rect 7991 3494 8004 3524
rect 8019 3510 8049 3524
rect 8086 3494 8105 3524
rect 8120 3494 8126 3524
rect 8135 3494 8148 3524
rect 8163 3510 8193 3524
rect 8236 3510 8279 3524
rect 8286 3510 8506 3524
rect 8513 3510 8543 3524
rect 8203 3496 8218 3508
rect 8237 3496 8250 3510
rect 8318 3506 8471 3510
rect 8200 3494 8222 3496
rect 8300 3494 8492 3506
rect 8571 3494 8584 3524
rect 8599 3510 8629 3524
rect 8666 3494 8685 3524
rect 8700 3494 8706 3524
rect 8715 3494 8728 3524
rect 8743 3510 8773 3524
rect 8816 3510 8859 3524
rect 8866 3510 9086 3524
rect 9093 3510 9123 3524
rect 8783 3496 8798 3508
rect 8817 3496 8830 3510
rect 8898 3506 9051 3510
rect 8780 3494 8802 3496
rect 8880 3494 9072 3506
rect 9151 3494 9164 3524
rect 9179 3510 9209 3524
rect 9246 3494 9265 3524
rect 9280 3494 9286 3524
rect 9295 3494 9308 3524
rect 9323 3510 9353 3524
rect 9396 3510 9439 3524
rect 9446 3510 9666 3524
rect 9673 3510 9703 3524
rect 9363 3496 9378 3508
rect 9397 3496 9410 3510
rect 9478 3506 9631 3510
rect 9360 3494 9382 3496
rect 9460 3494 9652 3506
rect 9731 3494 9744 3524
rect 9759 3510 9789 3524
rect 9826 3494 9845 3524
rect 9860 3494 9866 3524
rect 9875 3494 9888 3524
rect 9903 3510 9933 3524
rect 9976 3510 10019 3524
rect 10026 3510 10246 3524
rect 10253 3510 10283 3524
rect 9943 3496 9958 3508
rect 9977 3496 9990 3510
rect 10058 3506 10211 3510
rect 9940 3494 9962 3496
rect 10040 3494 10232 3506
rect 10311 3494 10324 3524
rect 10339 3510 10369 3524
rect 10406 3494 10425 3524
rect 10440 3494 10446 3524
rect 10455 3494 10468 3524
rect 10483 3510 10513 3524
rect 10556 3510 10599 3524
rect 10606 3510 10826 3524
rect 10833 3510 10863 3524
rect 10523 3496 10538 3508
rect 10557 3496 10570 3510
rect 10638 3506 10791 3510
rect 10520 3494 10542 3496
rect 10620 3494 10812 3506
rect 10891 3494 10904 3524
rect 10919 3510 10949 3524
rect 10986 3494 11005 3524
rect 11020 3494 11026 3524
rect 11035 3494 11048 3524
rect 11063 3510 11093 3524
rect 11136 3510 11179 3524
rect 11186 3510 11406 3524
rect 11413 3510 11443 3524
rect 11103 3496 11118 3508
rect 11137 3496 11150 3510
rect 11218 3506 11371 3510
rect 11100 3494 11122 3496
rect 11200 3494 11392 3506
rect 11471 3494 11484 3524
rect 11499 3510 11529 3524
rect 11566 3494 11585 3524
rect 11600 3494 11606 3524
rect 11615 3494 11628 3524
rect 11643 3510 11673 3524
rect 11716 3510 11759 3524
rect 11766 3510 11986 3524
rect 11993 3510 12023 3524
rect 11683 3496 11698 3508
rect 11717 3496 11730 3510
rect 11798 3506 11951 3510
rect 11680 3494 11702 3496
rect 11780 3494 11972 3506
rect 12051 3494 12064 3524
rect 12079 3510 12109 3524
rect 12146 3494 12165 3524
rect 12180 3494 12186 3524
rect 12195 3494 12208 3524
rect 12223 3510 12253 3524
rect 12296 3510 12339 3524
rect 12346 3510 12566 3524
rect 12573 3510 12603 3524
rect 12263 3496 12278 3508
rect 12297 3496 12310 3510
rect 12378 3506 12531 3510
rect 12260 3494 12282 3496
rect 12360 3494 12552 3506
rect 12631 3494 12644 3524
rect 12659 3510 12689 3524
rect 12726 3494 12745 3524
rect 12760 3494 12766 3524
rect 12775 3494 12788 3524
rect 12803 3510 12833 3524
rect 12876 3510 12919 3524
rect 12926 3510 13146 3524
rect 13153 3510 13183 3524
rect 12843 3496 12858 3508
rect 12877 3496 12890 3510
rect 12958 3506 13111 3510
rect 12840 3494 12862 3496
rect 12940 3494 13132 3506
rect 13211 3494 13224 3524
rect 13239 3510 13269 3524
rect 13306 3494 13325 3524
rect 13340 3494 13346 3524
rect 13355 3494 13368 3524
rect 13383 3510 13413 3524
rect 13456 3510 13499 3524
rect 13506 3510 13726 3524
rect 13733 3510 13763 3524
rect 13423 3496 13438 3508
rect 13457 3496 13470 3510
rect 13538 3506 13691 3510
rect 13420 3494 13442 3496
rect 13520 3494 13712 3506
rect 13791 3494 13804 3524
rect 13819 3510 13849 3524
rect 13886 3494 13905 3524
rect 13920 3494 13926 3524
rect 13935 3494 13948 3524
rect 13963 3510 13993 3524
rect 14036 3510 14079 3524
rect 14086 3510 14306 3524
rect 14313 3510 14343 3524
rect 14003 3496 14018 3508
rect 14037 3496 14050 3510
rect 14118 3506 14271 3510
rect 14000 3494 14022 3496
rect 14100 3494 14292 3506
rect 14371 3494 14384 3524
rect 14399 3510 14429 3524
rect 14466 3494 14485 3524
rect 14500 3494 14506 3524
rect 14515 3494 14528 3524
rect 14543 3510 14573 3524
rect 14616 3510 14659 3524
rect 14666 3510 14886 3524
rect 14893 3510 14923 3524
rect 14583 3496 14598 3508
rect 14617 3496 14630 3510
rect 14698 3506 14851 3510
rect 14580 3494 14602 3496
rect 14680 3494 14872 3506
rect 14951 3494 14964 3524
rect 14979 3510 15009 3524
rect 15046 3494 15065 3524
rect 15080 3494 15086 3524
rect 15095 3494 15108 3524
rect 15123 3510 15153 3524
rect 15196 3510 15239 3524
rect 15246 3510 15466 3524
rect 15473 3510 15503 3524
rect 15163 3496 15178 3508
rect 15197 3496 15210 3510
rect 15278 3506 15431 3510
rect 15160 3494 15182 3496
rect 15260 3494 15452 3506
rect 15531 3494 15544 3524
rect 15559 3510 15589 3524
rect 15626 3494 15645 3524
rect 15660 3494 15666 3524
rect 15675 3494 15688 3524
rect 15703 3510 15733 3524
rect 15776 3510 15819 3524
rect 15826 3510 16046 3524
rect 16053 3510 16083 3524
rect 15743 3496 15758 3508
rect 15777 3496 15790 3510
rect 15858 3506 16011 3510
rect 15740 3494 15762 3496
rect 15840 3494 16032 3506
rect 16111 3494 16124 3524
rect 16139 3510 16169 3524
rect 16206 3494 16225 3524
rect 16240 3494 16246 3524
rect 16255 3494 16268 3524
rect 16283 3510 16313 3524
rect 16356 3510 16399 3524
rect 16406 3510 16626 3524
rect 16633 3510 16663 3524
rect 16323 3496 16338 3508
rect 16357 3496 16370 3510
rect 16438 3506 16591 3510
rect 16320 3494 16342 3496
rect 16420 3494 16612 3506
rect 16691 3494 16704 3524
rect 16719 3510 16749 3524
rect 16786 3494 16805 3524
rect 16820 3494 16826 3524
rect 16835 3494 16848 3524
rect 16863 3510 16893 3524
rect 16936 3510 16979 3524
rect 16986 3510 17206 3524
rect 17213 3510 17243 3524
rect 16903 3496 16918 3508
rect 16937 3496 16950 3510
rect 17018 3506 17171 3510
rect 16900 3494 16922 3496
rect 17000 3494 17192 3506
rect 17271 3494 17284 3524
rect 17299 3510 17329 3524
rect 17366 3494 17385 3524
rect 17400 3494 17406 3524
rect 17415 3494 17428 3524
rect 17443 3510 17473 3524
rect 17516 3510 17559 3524
rect 17566 3510 17786 3524
rect 17793 3510 17823 3524
rect 17483 3496 17498 3508
rect 17517 3496 17530 3510
rect 17598 3506 17751 3510
rect 17480 3494 17502 3496
rect 17580 3494 17772 3506
rect 17851 3494 17864 3524
rect 17879 3510 17909 3524
rect 17946 3494 17965 3524
rect 17980 3494 17986 3524
rect 17995 3494 18008 3524
rect 18023 3510 18053 3524
rect 18096 3510 18139 3524
rect 18146 3510 18366 3524
rect 18373 3510 18403 3524
rect 18063 3496 18078 3508
rect 18097 3496 18110 3510
rect 18178 3506 18331 3510
rect 18060 3494 18082 3496
rect 18160 3494 18352 3506
rect 18431 3494 18444 3524
rect 18459 3510 18489 3524
rect 18532 3494 18545 3524
rect 0 3480 18545 3494
rect 15 3410 28 3480
rect 80 3476 102 3480
rect 73 3454 102 3468
rect 155 3454 171 3468
rect 209 3464 215 3466
rect 222 3464 330 3480
rect 337 3464 343 3466
rect 351 3464 366 3480
rect 432 3474 451 3477
rect 73 3452 171 3454
rect 198 3452 366 3464
rect 381 3454 397 3468
rect 432 3455 454 3474
rect 464 3468 480 3469
rect 463 3466 480 3468
rect 464 3461 480 3466
rect 454 3454 460 3455
rect 463 3454 492 3461
rect 381 3453 492 3454
rect 381 3452 498 3453
rect 57 3444 108 3452
rect 155 3444 189 3452
rect 57 3432 82 3444
rect 89 3432 108 3444
rect 162 3442 189 3444
rect 198 3442 419 3452
rect 454 3449 460 3452
rect 162 3438 419 3442
rect 57 3424 108 3432
rect 155 3424 419 3438
rect 463 3444 498 3452
rect 9 3376 28 3410
rect 73 3416 102 3424
rect 73 3410 90 3416
rect 73 3408 107 3410
rect 155 3408 171 3424
rect 172 3414 380 3424
rect 381 3414 397 3424
rect 445 3420 460 3435
rect 463 3432 464 3444
rect 471 3432 498 3444
rect 463 3424 498 3432
rect 463 3423 492 3424
rect 183 3410 397 3414
rect 198 3408 397 3410
rect 432 3410 445 3420
rect 463 3410 480 3423
rect 432 3408 480 3410
rect 74 3404 107 3408
rect 70 3402 107 3404
rect 70 3401 137 3402
rect 70 3396 101 3401
rect 107 3396 137 3401
rect 70 3392 137 3396
rect 43 3389 137 3392
rect 43 3382 92 3389
rect 43 3376 73 3382
rect 92 3377 97 3382
rect 9 3360 89 3376
rect 101 3368 137 3389
rect 198 3384 387 3408
rect 432 3407 479 3408
rect 445 3402 479 3407
rect 213 3381 387 3384
rect 206 3378 387 3381
rect 415 3401 479 3402
rect 9 3358 28 3360
rect 43 3358 77 3360
rect 9 3342 89 3358
rect 9 3336 28 3342
rect -1 3320 28 3336
rect 43 3326 73 3342
rect 101 3320 107 3368
rect 110 3362 129 3368
rect 144 3362 174 3370
rect 110 3354 174 3362
rect 110 3338 190 3354
rect 206 3347 268 3378
rect 284 3347 346 3378
rect 415 3376 464 3401
rect 479 3376 509 3392
rect 378 3362 408 3370
rect 415 3368 525 3376
rect 378 3354 423 3362
rect 110 3336 129 3338
rect 144 3336 190 3338
rect 110 3320 190 3336
rect 217 3334 252 3347
rect 293 3344 330 3347
rect 293 3342 335 3344
rect 222 3331 252 3334
rect 231 3327 238 3331
rect 238 3326 239 3327
rect 197 3320 207 3326
rect -7 3312 34 3320
rect -7 3286 8 3312
rect 15 3286 34 3312
rect 98 3308 129 3320
rect 144 3308 247 3320
rect 259 3310 285 3336
rect 300 3331 330 3342
rect 362 3338 424 3354
rect 362 3336 408 3338
rect 362 3320 424 3336
rect 436 3320 442 3368
rect 445 3360 525 3368
rect 445 3358 464 3360
rect 479 3358 513 3360
rect 445 3342 525 3358
rect 445 3320 464 3342
rect 479 3326 509 3342
rect 537 3336 543 3410
rect 546 3336 565 3480
rect 580 3336 586 3480
rect 595 3410 608 3480
rect 660 3476 682 3480
rect 653 3454 682 3468
rect 735 3454 751 3468
rect 789 3464 795 3466
rect 802 3464 910 3480
rect 917 3464 923 3466
rect 931 3464 946 3480
rect 1012 3474 1031 3477
rect 653 3452 751 3454
rect 778 3452 946 3464
rect 961 3454 977 3468
rect 1012 3455 1034 3474
rect 1044 3468 1060 3469
rect 1043 3466 1060 3468
rect 1044 3461 1060 3466
rect 1034 3454 1040 3455
rect 1043 3454 1072 3461
rect 961 3453 1072 3454
rect 961 3452 1078 3453
rect 637 3444 688 3452
rect 735 3444 769 3452
rect 637 3432 662 3444
rect 669 3432 688 3444
rect 742 3442 769 3444
rect 778 3442 999 3452
rect 1034 3449 1040 3452
rect 742 3438 999 3442
rect 637 3424 688 3432
rect 735 3424 999 3438
rect 1043 3444 1078 3452
rect 589 3376 608 3410
rect 653 3416 682 3424
rect 653 3410 670 3416
rect 653 3408 687 3410
rect 735 3408 751 3424
rect 752 3414 960 3424
rect 961 3414 977 3424
rect 1025 3420 1040 3435
rect 1043 3432 1044 3444
rect 1051 3432 1078 3444
rect 1043 3424 1078 3432
rect 1043 3423 1072 3424
rect 763 3410 977 3414
rect 778 3408 977 3410
rect 1012 3410 1025 3420
rect 1043 3410 1060 3423
rect 1012 3408 1060 3410
rect 654 3404 687 3408
rect 650 3402 687 3404
rect 650 3401 717 3402
rect 650 3396 681 3401
rect 687 3396 717 3401
rect 650 3392 717 3396
rect 623 3389 717 3392
rect 623 3382 672 3389
rect 623 3376 653 3382
rect 672 3377 677 3382
rect 589 3360 669 3376
rect 681 3368 717 3389
rect 778 3384 967 3408
rect 1012 3407 1059 3408
rect 1025 3402 1059 3407
rect 793 3381 967 3384
rect 786 3378 967 3381
rect 995 3401 1059 3402
rect 589 3358 608 3360
rect 623 3358 657 3360
rect 589 3342 669 3358
rect 589 3336 608 3342
rect 305 3310 408 3320
rect 259 3308 408 3310
rect 429 3308 464 3320
rect 98 3306 260 3308
rect 110 3286 129 3306
rect 144 3304 174 3306
rect -7 3278 34 3286
rect 116 3282 129 3286
rect 181 3290 260 3306
rect 292 3306 464 3308
rect 292 3290 371 3306
rect 378 3304 408 3306
rect -1 3268 28 3278
rect 43 3268 73 3282
rect 116 3268 159 3282
rect 181 3278 371 3290
rect 436 3286 442 3306
rect 166 3268 196 3278
rect 197 3268 355 3278
rect 359 3268 389 3278
rect 393 3268 423 3282
rect 451 3268 464 3306
rect 536 3320 565 3336
rect 579 3320 608 3336
rect 623 3326 653 3342
rect 681 3320 687 3368
rect 690 3362 709 3368
rect 724 3362 754 3370
rect 690 3354 754 3362
rect 690 3338 770 3354
rect 786 3347 848 3378
rect 864 3347 926 3378
rect 995 3376 1044 3401
rect 1059 3376 1089 3392
rect 958 3362 988 3370
rect 995 3368 1105 3376
rect 958 3354 1003 3362
rect 690 3336 709 3338
rect 724 3336 770 3338
rect 690 3320 770 3336
rect 797 3334 832 3347
rect 873 3344 910 3347
rect 873 3342 915 3344
rect 802 3331 832 3334
rect 811 3327 818 3331
rect 818 3326 819 3327
rect 777 3320 787 3326
rect 536 3312 571 3320
rect 536 3286 537 3312
rect 544 3286 571 3312
rect 479 3268 509 3282
rect 536 3278 571 3286
rect 573 3312 614 3320
rect 573 3286 588 3312
rect 595 3286 614 3312
rect 678 3308 709 3320
rect 724 3308 827 3320
rect 839 3310 865 3336
rect 880 3331 910 3342
rect 942 3338 1004 3354
rect 942 3336 988 3338
rect 942 3320 1004 3336
rect 1016 3320 1022 3368
rect 1025 3360 1105 3368
rect 1025 3358 1044 3360
rect 1059 3358 1093 3360
rect 1025 3342 1105 3358
rect 1025 3320 1044 3342
rect 1059 3326 1089 3342
rect 1117 3336 1123 3410
rect 1126 3336 1145 3480
rect 1160 3336 1166 3480
rect 1175 3410 1188 3480
rect 1240 3476 1262 3480
rect 1233 3454 1262 3468
rect 1315 3454 1331 3468
rect 1369 3464 1375 3466
rect 1382 3464 1490 3480
rect 1497 3464 1503 3466
rect 1511 3464 1526 3480
rect 1592 3474 1611 3477
rect 1233 3452 1331 3454
rect 1358 3452 1526 3464
rect 1541 3454 1557 3468
rect 1592 3455 1614 3474
rect 1624 3468 1640 3469
rect 1623 3466 1640 3468
rect 1624 3461 1640 3466
rect 1614 3454 1620 3455
rect 1623 3454 1652 3461
rect 1541 3453 1652 3454
rect 1541 3452 1658 3453
rect 1217 3444 1268 3452
rect 1315 3444 1349 3452
rect 1217 3432 1242 3444
rect 1249 3432 1268 3444
rect 1322 3442 1349 3444
rect 1358 3442 1579 3452
rect 1614 3449 1620 3452
rect 1322 3438 1579 3442
rect 1217 3424 1268 3432
rect 1315 3424 1579 3438
rect 1623 3444 1658 3452
rect 1169 3376 1188 3410
rect 1233 3416 1262 3424
rect 1233 3410 1250 3416
rect 1233 3408 1267 3410
rect 1315 3408 1331 3424
rect 1332 3414 1540 3424
rect 1541 3414 1557 3424
rect 1605 3420 1620 3435
rect 1623 3432 1624 3444
rect 1631 3432 1658 3444
rect 1623 3424 1658 3432
rect 1623 3423 1652 3424
rect 1343 3410 1557 3414
rect 1358 3408 1557 3410
rect 1592 3410 1605 3420
rect 1623 3410 1640 3423
rect 1592 3408 1640 3410
rect 1234 3404 1267 3408
rect 1230 3402 1267 3404
rect 1230 3401 1297 3402
rect 1230 3396 1261 3401
rect 1267 3396 1297 3401
rect 1230 3392 1297 3396
rect 1203 3389 1297 3392
rect 1203 3382 1252 3389
rect 1203 3376 1233 3382
rect 1252 3377 1257 3382
rect 1169 3360 1249 3376
rect 1261 3368 1297 3389
rect 1358 3384 1547 3408
rect 1592 3407 1639 3408
rect 1605 3402 1639 3407
rect 1373 3381 1547 3384
rect 1366 3378 1547 3381
rect 1575 3401 1639 3402
rect 1169 3358 1188 3360
rect 1203 3358 1237 3360
rect 1169 3342 1249 3358
rect 1169 3336 1188 3342
rect 885 3310 988 3320
rect 839 3308 988 3310
rect 1009 3308 1044 3320
rect 678 3306 840 3308
rect 690 3286 709 3306
rect 724 3304 754 3306
rect 573 3278 614 3286
rect 696 3282 709 3286
rect 761 3290 840 3306
rect 872 3306 1044 3308
rect 872 3290 951 3306
rect 958 3304 988 3306
rect 536 3268 565 3278
rect 579 3268 608 3278
rect 623 3268 653 3282
rect 696 3268 739 3282
rect 761 3278 951 3290
rect 1016 3286 1022 3306
rect 746 3268 776 3278
rect 777 3268 935 3278
rect 939 3268 969 3278
rect 973 3268 1003 3282
rect 1031 3268 1044 3306
rect 1116 3320 1145 3336
rect 1159 3320 1188 3336
rect 1203 3326 1233 3342
rect 1261 3320 1267 3368
rect 1270 3362 1289 3368
rect 1304 3362 1334 3370
rect 1270 3354 1334 3362
rect 1270 3338 1350 3354
rect 1366 3347 1428 3378
rect 1444 3347 1506 3378
rect 1575 3376 1624 3401
rect 1639 3376 1669 3392
rect 1538 3362 1568 3370
rect 1575 3368 1685 3376
rect 1538 3354 1583 3362
rect 1270 3336 1289 3338
rect 1304 3336 1350 3338
rect 1270 3320 1350 3336
rect 1377 3334 1412 3347
rect 1453 3344 1490 3347
rect 1453 3342 1495 3344
rect 1382 3331 1412 3334
rect 1391 3327 1398 3331
rect 1398 3326 1399 3327
rect 1357 3320 1367 3326
rect 1116 3312 1151 3320
rect 1116 3286 1117 3312
rect 1124 3286 1151 3312
rect 1059 3268 1089 3282
rect 1116 3278 1151 3286
rect 1153 3312 1194 3320
rect 1153 3286 1168 3312
rect 1175 3286 1194 3312
rect 1258 3308 1289 3320
rect 1304 3308 1407 3320
rect 1419 3310 1445 3336
rect 1460 3331 1490 3342
rect 1522 3338 1584 3354
rect 1522 3336 1568 3338
rect 1522 3320 1584 3336
rect 1596 3320 1602 3368
rect 1605 3360 1685 3368
rect 1605 3358 1624 3360
rect 1639 3358 1673 3360
rect 1605 3342 1685 3358
rect 1605 3320 1624 3342
rect 1639 3326 1669 3342
rect 1697 3336 1703 3410
rect 1706 3336 1725 3480
rect 1740 3336 1746 3480
rect 1755 3410 1768 3480
rect 1820 3476 1842 3480
rect 1813 3454 1842 3468
rect 1895 3454 1911 3468
rect 1949 3464 1955 3466
rect 1962 3464 2070 3480
rect 2077 3464 2083 3466
rect 2091 3464 2106 3480
rect 2172 3474 2191 3477
rect 1813 3452 1911 3454
rect 1938 3452 2106 3464
rect 2121 3454 2137 3468
rect 2172 3455 2194 3474
rect 2204 3468 2220 3469
rect 2203 3466 2220 3468
rect 2204 3461 2220 3466
rect 2194 3454 2200 3455
rect 2203 3454 2232 3461
rect 2121 3453 2232 3454
rect 2121 3452 2238 3453
rect 1797 3444 1848 3452
rect 1895 3444 1929 3452
rect 1797 3432 1822 3444
rect 1829 3432 1848 3444
rect 1902 3442 1929 3444
rect 1938 3442 2159 3452
rect 2194 3449 2200 3452
rect 1902 3438 2159 3442
rect 1797 3424 1848 3432
rect 1895 3424 2159 3438
rect 2203 3444 2238 3452
rect 1749 3376 1768 3410
rect 1813 3416 1842 3424
rect 1813 3410 1830 3416
rect 1813 3408 1847 3410
rect 1895 3408 1911 3424
rect 1912 3414 2120 3424
rect 2121 3414 2137 3424
rect 2185 3420 2200 3435
rect 2203 3432 2204 3444
rect 2211 3432 2238 3444
rect 2203 3424 2238 3432
rect 2203 3423 2232 3424
rect 1923 3410 2137 3414
rect 1938 3408 2137 3410
rect 2172 3410 2185 3420
rect 2203 3410 2220 3423
rect 2172 3408 2220 3410
rect 1814 3404 1847 3408
rect 1810 3402 1847 3404
rect 1810 3401 1877 3402
rect 1810 3396 1841 3401
rect 1847 3396 1877 3401
rect 1810 3392 1877 3396
rect 1783 3389 1877 3392
rect 1783 3382 1832 3389
rect 1783 3376 1813 3382
rect 1832 3377 1837 3382
rect 1749 3360 1829 3376
rect 1841 3368 1877 3389
rect 1938 3384 2127 3408
rect 2172 3407 2219 3408
rect 2185 3402 2219 3407
rect 1953 3381 2127 3384
rect 1946 3378 2127 3381
rect 2155 3401 2219 3402
rect 1749 3358 1768 3360
rect 1783 3358 1817 3360
rect 1749 3342 1829 3358
rect 1749 3336 1768 3342
rect 1465 3310 1568 3320
rect 1419 3308 1568 3310
rect 1589 3308 1624 3320
rect 1258 3306 1420 3308
rect 1270 3286 1289 3306
rect 1304 3304 1334 3306
rect 1153 3278 1194 3286
rect 1276 3282 1289 3286
rect 1341 3290 1420 3306
rect 1452 3306 1624 3308
rect 1452 3290 1531 3306
rect 1538 3304 1568 3306
rect 1116 3268 1145 3278
rect 1159 3268 1188 3278
rect 1203 3268 1233 3282
rect 1276 3268 1319 3282
rect 1341 3278 1531 3290
rect 1596 3286 1602 3306
rect 1326 3268 1356 3278
rect 1357 3268 1515 3278
rect 1519 3268 1549 3278
rect 1553 3268 1583 3282
rect 1611 3268 1624 3306
rect 1696 3320 1725 3336
rect 1739 3320 1768 3336
rect 1783 3326 1813 3342
rect 1841 3320 1847 3368
rect 1850 3362 1869 3368
rect 1884 3362 1914 3370
rect 1850 3354 1914 3362
rect 1850 3338 1930 3354
rect 1946 3347 2008 3378
rect 2024 3347 2086 3378
rect 2155 3376 2204 3401
rect 2219 3376 2249 3392
rect 2118 3362 2148 3370
rect 2155 3368 2265 3376
rect 2118 3354 2163 3362
rect 1850 3336 1869 3338
rect 1884 3336 1930 3338
rect 1850 3320 1930 3336
rect 1957 3334 1992 3347
rect 2033 3344 2070 3347
rect 2033 3342 2075 3344
rect 1962 3331 1992 3334
rect 1971 3327 1978 3331
rect 1978 3326 1979 3327
rect 1937 3320 1947 3326
rect 1696 3312 1731 3320
rect 1696 3286 1697 3312
rect 1704 3286 1731 3312
rect 1639 3268 1669 3282
rect 1696 3278 1731 3286
rect 1733 3312 1774 3320
rect 1733 3286 1748 3312
rect 1755 3286 1774 3312
rect 1838 3308 1869 3320
rect 1884 3308 1987 3320
rect 1999 3310 2025 3336
rect 2040 3331 2070 3342
rect 2102 3338 2164 3354
rect 2102 3336 2148 3338
rect 2102 3320 2164 3336
rect 2176 3320 2182 3368
rect 2185 3360 2265 3368
rect 2185 3358 2204 3360
rect 2219 3358 2253 3360
rect 2185 3342 2265 3358
rect 2185 3320 2204 3342
rect 2219 3326 2249 3342
rect 2277 3336 2283 3410
rect 2286 3336 2305 3480
rect 2320 3336 2326 3480
rect 2335 3410 2348 3480
rect 2400 3476 2422 3480
rect 2393 3454 2422 3468
rect 2475 3454 2491 3468
rect 2529 3464 2535 3466
rect 2542 3464 2650 3480
rect 2657 3464 2663 3466
rect 2671 3464 2686 3480
rect 2752 3474 2771 3477
rect 2393 3452 2491 3454
rect 2518 3452 2686 3464
rect 2701 3454 2717 3468
rect 2752 3455 2774 3474
rect 2784 3468 2800 3469
rect 2783 3466 2800 3468
rect 2784 3461 2800 3466
rect 2774 3454 2780 3455
rect 2783 3454 2812 3461
rect 2701 3453 2812 3454
rect 2701 3452 2818 3453
rect 2377 3444 2428 3452
rect 2475 3444 2509 3452
rect 2377 3432 2402 3444
rect 2409 3432 2428 3444
rect 2482 3442 2509 3444
rect 2518 3442 2739 3452
rect 2774 3449 2780 3452
rect 2482 3438 2739 3442
rect 2377 3424 2428 3432
rect 2475 3424 2739 3438
rect 2783 3444 2818 3452
rect 2329 3376 2348 3410
rect 2393 3416 2422 3424
rect 2393 3410 2410 3416
rect 2393 3408 2427 3410
rect 2475 3408 2491 3424
rect 2492 3414 2700 3424
rect 2701 3414 2717 3424
rect 2765 3420 2780 3435
rect 2783 3432 2784 3444
rect 2791 3432 2818 3444
rect 2783 3424 2818 3432
rect 2783 3423 2812 3424
rect 2503 3410 2717 3414
rect 2518 3408 2717 3410
rect 2752 3410 2765 3420
rect 2783 3410 2800 3423
rect 2752 3408 2800 3410
rect 2394 3404 2427 3408
rect 2390 3402 2427 3404
rect 2390 3401 2457 3402
rect 2390 3396 2421 3401
rect 2427 3396 2457 3401
rect 2390 3392 2457 3396
rect 2363 3389 2457 3392
rect 2363 3382 2412 3389
rect 2363 3376 2393 3382
rect 2412 3377 2417 3382
rect 2329 3360 2409 3376
rect 2421 3368 2457 3389
rect 2518 3384 2707 3408
rect 2752 3407 2799 3408
rect 2765 3402 2799 3407
rect 2533 3381 2707 3384
rect 2526 3378 2707 3381
rect 2735 3401 2799 3402
rect 2329 3358 2348 3360
rect 2363 3358 2397 3360
rect 2329 3342 2409 3358
rect 2329 3336 2348 3342
rect 2045 3310 2148 3320
rect 1999 3308 2148 3310
rect 2169 3308 2204 3320
rect 1838 3306 2000 3308
rect 1850 3286 1869 3306
rect 1884 3304 1914 3306
rect 1733 3278 1774 3286
rect 1856 3282 1869 3286
rect 1921 3290 2000 3306
rect 2032 3306 2204 3308
rect 2032 3290 2111 3306
rect 2118 3304 2148 3306
rect 1696 3268 1725 3278
rect 1739 3268 1768 3278
rect 1783 3268 1813 3282
rect 1856 3268 1899 3282
rect 1921 3278 2111 3290
rect 2176 3286 2182 3306
rect 1906 3268 1936 3278
rect 1937 3268 2095 3278
rect 2099 3268 2129 3278
rect 2133 3268 2163 3282
rect 2191 3268 2204 3306
rect 2276 3320 2305 3336
rect 2319 3320 2348 3336
rect 2363 3326 2393 3342
rect 2421 3320 2427 3368
rect 2430 3362 2449 3368
rect 2464 3362 2494 3370
rect 2430 3354 2494 3362
rect 2430 3338 2510 3354
rect 2526 3347 2588 3378
rect 2604 3347 2666 3378
rect 2735 3376 2784 3401
rect 2799 3376 2829 3392
rect 2698 3362 2728 3370
rect 2735 3368 2845 3376
rect 2698 3354 2743 3362
rect 2430 3336 2449 3338
rect 2464 3336 2510 3338
rect 2430 3320 2510 3336
rect 2537 3334 2572 3347
rect 2613 3344 2650 3347
rect 2613 3342 2655 3344
rect 2542 3331 2572 3334
rect 2551 3327 2558 3331
rect 2558 3326 2559 3327
rect 2517 3320 2527 3326
rect 2276 3312 2311 3320
rect 2276 3286 2277 3312
rect 2284 3286 2311 3312
rect 2219 3268 2249 3282
rect 2276 3278 2311 3286
rect 2313 3312 2354 3320
rect 2313 3286 2328 3312
rect 2335 3286 2354 3312
rect 2418 3308 2449 3320
rect 2464 3308 2567 3320
rect 2579 3310 2605 3336
rect 2620 3331 2650 3342
rect 2682 3338 2744 3354
rect 2682 3336 2728 3338
rect 2682 3320 2744 3336
rect 2756 3320 2762 3368
rect 2765 3360 2845 3368
rect 2765 3358 2784 3360
rect 2799 3358 2833 3360
rect 2765 3342 2845 3358
rect 2765 3320 2784 3342
rect 2799 3326 2829 3342
rect 2857 3336 2863 3410
rect 2866 3336 2885 3480
rect 2900 3336 2906 3480
rect 2915 3410 2928 3480
rect 2980 3476 3002 3480
rect 2973 3454 3002 3468
rect 3055 3454 3071 3468
rect 3109 3464 3115 3466
rect 3122 3464 3230 3480
rect 3237 3464 3243 3466
rect 3251 3464 3266 3480
rect 3332 3474 3351 3477
rect 2973 3452 3071 3454
rect 3098 3452 3266 3464
rect 3281 3454 3297 3468
rect 3332 3455 3354 3474
rect 3364 3468 3380 3469
rect 3363 3466 3380 3468
rect 3364 3461 3380 3466
rect 3354 3454 3360 3455
rect 3363 3454 3392 3461
rect 3281 3453 3392 3454
rect 3281 3452 3398 3453
rect 2957 3444 3008 3452
rect 3055 3444 3089 3452
rect 2957 3432 2982 3444
rect 2989 3432 3008 3444
rect 3062 3442 3089 3444
rect 3098 3442 3319 3452
rect 3354 3449 3360 3452
rect 3062 3438 3319 3442
rect 2957 3424 3008 3432
rect 3055 3424 3319 3438
rect 3363 3444 3398 3452
rect 2909 3376 2928 3410
rect 2973 3416 3002 3424
rect 2973 3410 2990 3416
rect 2973 3408 3007 3410
rect 3055 3408 3071 3424
rect 3072 3414 3280 3424
rect 3281 3414 3297 3424
rect 3345 3420 3360 3435
rect 3363 3432 3364 3444
rect 3371 3432 3398 3444
rect 3363 3424 3398 3432
rect 3363 3423 3392 3424
rect 3083 3410 3297 3414
rect 3098 3408 3297 3410
rect 3332 3410 3345 3420
rect 3363 3410 3380 3423
rect 3332 3408 3380 3410
rect 2974 3404 3007 3408
rect 2970 3402 3007 3404
rect 2970 3401 3037 3402
rect 2970 3396 3001 3401
rect 3007 3396 3037 3401
rect 2970 3392 3037 3396
rect 2943 3389 3037 3392
rect 2943 3382 2992 3389
rect 2943 3376 2973 3382
rect 2992 3377 2997 3382
rect 2909 3360 2989 3376
rect 3001 3368 3037 3389
rect 3098 3384 3287 3408
rect 3332 3407 3379 3408
rect 3345 3402 3379 3407
rect 3113 3381 3287 3384
rect 3106 3378 3287 3381
rect 3315 3401 3379 3402
rect 2909 3358 2928 3360
rect 2943 3358 2977 3360
rect 2909 3342 2989 3358
rect 2909 3336 2928 3342
rect 2625 3310 2728 3320
rect 2579 3308 2728 3310
rect 2749 3308 2784 3320
rect 2418 3306 2580 3308
rect 2430 3286 2449 3306
rect 2464 3304 2494 3306
rect 2313 3278 2354 3286
rect 2436 3282 2449 3286
rect 2501 3290 2580 3306
rect 2612 3306 2784 3308
rect 2612 3290 2691 3306
rect 2698 3304 2728 3306
rect 2276 3268 2305 3278
rect 2319 3268 2348 3278
rect 2363 3268 2393 3282
rect 2436 3268 2479 3282
rect 2501 3278 2691 3290
rect 2756 3286 2762 3306
rect 2486 3268 2516 3278
rect 2517 3268 2675 3278
rect 2679 3268 2709 3278
rect 2713 3268 2743 3282
rect 2771 3268 2784 3306
rect 2856 3320 2885 3336
rect 2899 3320 2928 3336
rect 2943 3326 2973 3342
rect 3001 3320 3007 3368
rect 3010 3362 3029 3368
rect 3044 3362 3074 3370
rect 3010 3354 3074 3362
rect 3010 3338 3090 3354
rect 3106 3347 3168 3378
rect 3184 3347 3246 3378
rect 3315 3376 3364 3401
rect 3379 3376 3409 3392
rect 3278 3362 3308 3370
rect 3315 3368 3425 3376
rect 3278 3354 3323 3362
rect 3010 3336 3029 3338
rect 3044 3336 3090 3338
rect 3010 3320 3090 3336
rect 3117 3334 3152 3347
rect 3193 3344 3230 3347
rect 3193 3342 3235 3344
rect 3122 3331 3152 3334
rect 3131 3327 3138 3331
rect 3138 3326 3139 3327
rect 3097 3320 3107 3326
rect 2856 3312 2891 3320
rect 2856 3286 2857 3312
rect 2864 3286 2891 3312
rect 2799 3268 2829 3282
rect 2856 3278 2891 3286
rect 2893 3312 2934 3320
rect 2893 3286 2908 3312
rect 2915 3286 2934 3312
rect 2998 3308 3029 3320
rect 3044 3308 3147 3320
rect 3159 3310 3185 3336
rect 3200 3331 3230 3342
rect 3262 3338 3324 3354
rect 3262 3336 3308 3338
rect 3262 3320 3324 3336
rect 3336 3320 3342 3368
rect 3345 3360 3425 3368
rect 3345 3358 3364 3360
rect 3379 3358 3413 3360
rect 3345 3342 3425 3358
rect 3345 3320 3364 3342
rect 3379 3326 3409 3342
rect 3437 3336 3443 3410
rect 3446 3336 3465 3480
rect 3480 3336 3486 3480
rect 3495 3410 3508 3480
rect 3560 3476 3582 3480
rect 3553 3454 3582 3468
rect 3635 3454 3651 3468
rect 3689 3464 3695 3466
rect 3702 3464 3810 3480
rect 3817 3464 3823 3466
rect 3831 3464 3846 3480
rect 3912 3474 3931 3477
rect 3553 3452 3651 3454
rect 3678 3452 3846 3464
rect 3861 3454 3877 3468
rect 3912 3455 3934 3474
rect 3944 3468 3960 3469
rect 3943 3466 3960 3468
rect 3944 3461 3960 3466
rect 3934 3454 3940 3455
rect 3943 3454 3972 3461
rect 3861 3453 3972 3454
rect 3861 3452 3978 3453
rect 3537 3444 3588 3452
rect 3635 3444 3669 3452
rect 3537 3432 3562 3444
rect 3569 3432 3588 3444
rect 3642 3442 3669 3444
rect 3678 3442 3899 3452
rect 3934 3449 3940 3452
rect 3642 3438 3899 3442
rect 3537 3424 3588 3432
rect 3635 3424 3899 3438
rect 3943 3444 3978 3452
rect 3489 3376 3508 3410
rect 3553 3416 3582 3424
rect 3553 3410 3570 3416
rect 3553 3408 3587 3410
rect 3635 3408 3651 3424
rect 3652 3414 3860 3424
rect 3861 3414 3877 3424
rect 3925 3420 3940 3435
rect 3943 3432 3944 3444
rect 3951 3432 3978 3444
rect 3943 3424 3978 3432
rect 3943 3423 3972 3424
rect 3663 3410 3877 3414
rect 3678 3408 3877 3410
rect 3912 3410 3925 3420
rect 3943 3410 3960 3423
rect 3912 3408 3960 3410
rect 3554 3404 3587 3408
rect 3550 3402 3587 3404
rect 3550 3401 3617 3402
rect 3550 3396 3581 3401
rect 3587 3396 3617 3401
rect 3550 3392 3617 3396
rect 3523 3389 3617 3392
rect 3523 3382 3572 3389
rect 3523 3376 3553 3382
rect 3572 3377 3577 3382
rect 3489 3360 3569 3376
rect 3581 3368 3617 3389
rect 3678 3384 3867 3408
rect 3912 3407 3959 3408
rect 3925 3402 3959 3407
rect 3693 3381 3867 3384
rect 3686 3378 3867 3381
rect 3895 3401 3959 3402
rect 3489 3358 3508 3360
rect 3523 3358 3557 3360
rect 3489 3342 3569 3358
rect 3489 3336 3508 3342
rect 3205 3310 3308 3320
rect 3159 3308 3308 3310
rect 3329 3308 3364 3320
rect 2998 3306 3160 3308
rect 3010 3286 3029 3306
rect 3044 3304 3074 3306
rect 2893 3278 2934 3286
rect 3016 3282 3029 3286
rect 3081 3290 3160 3306
rect 3192 3306 3364 3308
rect 3192 3290 3271 3306
rect 3278 3304 3308 3306
rect 2856 3268 2885 3278
rect 2899 3268 2928 3278
rect 2943 3268 2973 3282
rect 3016 3268 3059 3282
rect 3081 3278 3271 3290
rect 3336 3286 3342 3306
rect 3066 3268 3096 3278
rect 3097 3268 3255 3278
rect 3259 3268 3289 3278
rect 3293 3268 3323 3282
rect 3351 3268 3364 3306
rect 3436 3320 3465 3336
rect 3479 3320 3508 3336
rect 3523 3326 3553 3342
rect 3581 3320 3587 3368
rect 3590 3362 3609 3368
rect 3624 3362 3654 3370
rect 3590 3354 3654 3362
rect 3590 3338 3670 3354
rect 3686 3347 3748 3378
rect 3764 3347 3826 3378
rect 3895 3376 3944 3401
rect 3959 3376 3989 3392
rect 3858 3362 3888 3370
rect 3895 3368 4005 3376
rect 3858 3354 3903 3362
rect 3590 3336 3609 3338
rect 3624 3336 3670 3338
rect 3590 3320 3670 3336
rect 3697 3334 3732 3347
rect 3773 3344 3810 3347
rect 3773 3342 3815 3344
rect 3702 3331 3732 3334
rect 3711 3327 3718 3331
rect 3718 3326 3719 3327
rect 3677 3320 3687 3326
rect 3436 3312 3471 3320
rect 3436 3286 3437 3312
rect 3444 3286 3471 3312
rect 3379 3268 3409 3282
rect 3436 3278 3471 3286
rect 3473 3312 3514 3320
rect 3473 3286 3488 3312
rect 3495 3286 3514 3312
rect 3578 3308 3609 3320
rect 3624 3308 3727 3320
rect 3739 3310 3765 3336
rect 3780 3331 3810 3342
rect 3842 3338 3904 3354
rect 3842 3336 3888 3338
rect 3842 3320 3904 3336
rect 3916 3320 3922 3368
rect 3925 3360 4005 3368
rect 3925 3358 3944 3360
rect 3959 3358 3993 3360
rect 3925 3342 4005 3358
rect 3925 3320 3944 3342
rect 3959 3326 3989 3342
rect 4017 3336 4023 3410
rect 4026 3336 4045 3480
rect 4060 3336 4066 3480
rect 4075 3410 4088 3480
rect 4140 3476 4162 3480
rect 4133 3454 4162 3468
rect 4215 3454 4231 3468
rect 4269 3464 4275 3466
rect 4282 3464 4390 3480
rect 4397 3464 4403 3466
rect 4411 3464 4426 3480
rect 4492 3474 4511 3477
rect 4133 3452 4231 3454
rect 4258 3452 4426 3464
rect 4441 3454 4457 3468
rect 4492 3455 4514 3474
rect 4524 3468 4540 3469
rect 4523 3466 4540 3468
rect 4524 3461 4540 3466
rect 4514 3454 4520 3455
rect 4523 3454 4552 3461
rect 4441 3453 4552 3454
rect 4441 3452 4558 3453
rect 4117 3444 4168 3452
rect 4215 3444 4249 3452
rect 4117 3432 4142 3444
rect 4149 3432 4168 3444
rect 4222 3442 4249 3444
rect 4258 3442 4479 3452
rect 4514 3449 4520 3452
rect 4222 3438 4479 3442
rect 4117 3424 4168 3432
rect 4215 3424 4479 3438
rect 4523 3444 4558 3452
rect 4069 3376 4088 3410
rect 4133 3416 4162 3424
rect 4133 3410 4150 3416
rect 4133 3408 4167 3410
rect 4215 3408 4231 3424
rect 4232 3414 4440 3424
rect 4441 3414 4457 3424
rect 4505 3420 4520 3435
rect 4523 3432 4524 3444
rect 4531 3432 4558 3444
rect 4523 3424 4558 3432
rect 4523 3423 4552 3424
rect 4243 3410 4457 3414
rect 4258 3408 4457 3410
rect 4492 3410 4505 3420
rect 4523 3410 4540 3423
rect 4492 3408 4540 3410
rect 4134 3404 4167 3408
rect 4130 3402 4167 3404
rect 4130 3401 4197 3402
rect 4130 3396 4161 3401
rect 4167 3396 4197 3401
rect 4130 3392 4197 3396
rect 4103 3389 4197 3392
rect 4103 3382 4152 3389
rect 4103 3376 4133 3382
rect 4152 3377 4157 3382
rect 4069 3360 4149 3376
rect 4161 3368 4197 3389
rect 4258 3384 4447 3408
rect 4492 3407 4539 3408
rect 4505 3402 4539 3407
rect 4273 3381 4447 3384
rect 4266 3378 4447 3381
rect 4475 3401 4539 3402
rect 4069 3358 4088 3360
rect 4103 3358 4137 3360
rect 4069 3342 4149 3358
rect 4069 3336 4088 3342
rect 3785 3310 3888 3320
rect 3739 3308 3888 3310
rect 3909 3308 3944 3320
rect 3578 3306 3740 3308
rect 3590 3286 3609 3306
rect 3624 3304 3654 3306
rect 3473 3278 3514 3286
rect 3596 3282 3609 3286
rect 3661 3290 3740 3306
rect 3772 3306 3944 3308
rect 3772 3290 3851 3306
rect 3858 3304 3888 3306
rect 3436 3268 3465 3278
rect 3479 3268 3508 3278
rect 3523 3268 3553 3282
rect 3596 3268 3639 3282
rect 3661 3278 3851 3290
rect 3916 3286 3922 3306
rect 3646 3268 3676 3278
rect 3677 3268 3835 3278
rect 3839 3268 3869 3278
rect 3873 3268 3903 3282
rect 3931 3268 3944 3306
rect 4016 3320 4045 3336
rect 4059 3320 4088 3336
rect 4103 3326 4133 3342
rect 4161 3320 4167 3368
rect 4170 3362 4189 3368
rect 4204 3362 4234 3370
rect 4170 3354 4234 3362
rect 4170 3338 4250 3354
rect 4266 3347 4328 3378
rect 4344 3347 4406 3378
rect 4475 3376 4524 3401
rect 4539 3376 4569 3392
rect 4438 3362 4468 3370
rect 4475 3368 4585 3376
rect 4438 3354 4483 3362
rect 4170 3336 4189 3338
rect 4204 3336 4250 3338
rect 4170 3320 4250 3336
rect 4277 3334 4312 3347
rect 4353 3344 4390 3347
rect 4353 3342 4395 3344
rect 4282 3331 4312 3334
rect 4291 3327 4298 3331
rect 4298 3326 4299 3327
rect 4257 3320 4267 3326
rect 4016 3312 4051 3320
rect 4016 3286 4017 3312
rect 4024 3286 4051 3312
rect 3959 3268 3989 3282
rect 4016 3278 4051 3286
rect 4053 3312 4094 3320
rect 4053 3286 4068 3312
rect 4075 3286 4094 3312
rect 4158 3308 4189 3320
rect 4204 3308 4307 3320
rect 4319 3310 4345 3336
rect 4360 3331 4390 3342
rect 4422 3338 4484 3354
rect 4422 3336 4468 3338
rect 4422 3320 4484 3336
rect 4496 3320 4502 3368
rect 4505 3360 4585 3368
rect 4505 3358 4524 3360
rect 4539 3358 4573 3360
rect 4505 3342 4585 3358
rect 4505 3320 4524 3342
rect 4539 3326 4569 3342
rect 4597 3336 4603 3410
rect 4606 3336 4625 3480
rect 4640 3336 4646 3480
rect 4655 3410 4668 3480
rect 4720 3476 4742 3480
rect 4713 3454 4742 3468
rect 4795 3454 4811 3468
rect 4849 3464 4855 3466
rect 4862 3464 4970 3480
rect 4977 3464 4983 3466
rect 4991 3464 5006 3480
rect 5072 3474 5091 3477
rect 4713 3452 4811 3454
rect 4838 3452 5006 3464
rect 5021 3454 5037 3468
rect 5072 3455 5094 3474
rect 5104 3468 5120 3469
rect 5103 3466 5120 3468
rect 5104 3461 5120 3466
rect 5094 3454 5100 3455
rect 5103 3454 5132 3461
rect 5021 3453 5132 3454
rect 5021 3452 5138 3453
rect 4697 3444 4748 3452
rect 4795 3444 4829 3452
rect 4697 3432 4722 3444
rect 4729 3432 4748 3444
rect 4802 3442 4829 3444
rect 4838 3442 5059 3452
rect 5094 3449 5100 3452
rect 4802 3438 5059 3442
rect 4697 3424 4748 3432
rect 4795 3424 5059 3438
rect 5103 3444 5138 3452
rect 4649 3376 4668 3410
rect 4713 3416 4742 3424
rect 4713 3410 4730 3416
rect 4713 3408 4747 3410
rect 4795 3408 4811 3424
rect 4812 3414 5020 3424
rect 5021 3414 5037 3424
rect 5085 3420 5100 3435
rect 5103 3432 5104 3444
rect 5111 3432 5138 3444
rect 5103 3424 5138 3432
rect 5103 3423 5132 3424
rect 4823 3410 5037 3414
rect 4838 3408 5037 3410
rect 5072 3410 5085 3420
rect 5103 3410 5120 3423
rect 5072 3408 5120 3410
rect 4714 3404 4747 3408
rect 4710 3402 4747 3404
rect 4710 3401 4777 3402
rect 4710 3396 4741 3401
rect 4747 3396 4777 3401
rect 4710 3392 4777 3396
rect 4683 3389 4777 3392
rect 4683 3382 4732 3389
rect 4683 3376 4713 3382
rect 4732 3377 4737 3382
rect 4649 3360 4729 3376
rect 4741 3368 4777 3389
rect 4838 3384 5027 3408
rect 5072 3407 5119 3408
rect 5085 3402 5119 3407
rect 4853 3381 5027 3384
rect 4846 3378 5027 3381
rect 5055 3401 5119 3402
rect 4649 3358 4668 3360
rect 4683 3358 4717 3360
rect 4649 3342 4729 3358
rect 4649 3336 4668 3342
rect 4365 3310 4468 3320
rect 4319 3308 4468 3310
rect 4489 3308 4524 3320
rect 4158 3306 4320 3308
rect 4170 3286 4189 3306
rect 4204 3304 4234 3306
rect 4053 3278 4094 3286
rect 4176 3282 4189 3286
rect 4241 3290 4320 3306
rect 4352 3306 4524 3308
rect 4352 3290 4431 3306
rect 4438 3304 4468 3306
rect 4016 3268 4045 3278
rect 4059 3268 4088 3278
rect 4103 3268 4133 3282
rect 4176 3268 4219 3282
rect 4241 3278 4431 3290
rect 4496 3286 4502 3306
rect 4226 3268 4256 3278
rect 4257 3268 4415 3278
rect 4419 3268 4449 3278
rect 4453 3268 4483 3282
rect 4511 3268 4524 3306
rect 4596 3320 4625 3336
rect 4639 3320 4668 3336
rect 4683 3326 4713 3342
rect 4741 3320 4747 3368
rect 4750 3362 4769 3368
rect 4784 3362 4814 3370
rect 4750 3354 4814 3362
rect 4750 3338 4830 3354
rect 4846 3347 4908 3378
rect 4924 3347 4986 3378
rect 5055 3376 5104 3401
rect 5119 3376 5149 3392
rect 5018 3362 5048 3370
rect 5055 3368 5165 3376
rect 5018 3354 5063 3362
rect 4750 3336 4769 3338
rect 4784 3336 4830 3338
rect 4750 3320 4830 3336
rect 4857 3334 4892 3347
rect 4933 3344 4970 3347
rect 4933 3342 4975 3344
rect 4862 3331 4892 3334
rect 4871 3327 4878 3331
rect 4878 3326 4879 3327
rect 4837 3320 4847 3326
rect 4596 3312 4631 3320
rect 4596 3286 4597 3312
rect 4604 3286 4631 3312
rect 4539 3268 4569 3282
rect 4596 3278 4631 3286
rect 4633 3312 4674 3320
rect 4633 3286 4648 3312
rect 4655 3286 4674 3312
rect 4738 3308 4769 3320
rect 4784 3308 4887 3320
rect 4899 3310 4925 3336
rect 4940 3331 4970 3342
rect 5002 3338 5064 3354
rect 5002 3336 5048 3338
rect 5002 3320 5064 3336
rect 5076 3320 5082 3368
rect 5085 3360 5165 3368
rect 5085 3358 5104 3360
rect 5119 3358 5153 3360
rect 5085 3342 5165 3358
rect 5085 3320 5104 3342
rect 5119 3326 5149 3342
rect 5177 3336 5183 3410
rect 5186 3336 5205 3480
rect 5220 3336 5226 3480
rect 5235 3410 5248 3480
rect 5300 3476 5322 3480
rect 5293 3454 5322 3468
rect 5375 3454 5391 3468
rect 5429 3464 5435 3466
rect 5442 3464 5550 3480
rect 5557 3464 5563 3466
rect 5571 3464 5586 3480
rect 5652 3474 5671 3477
rect 5293 3452 5391 3454
rect 5418 3452 5586 3464
rect 5601 3454 5617 3468
rect 5652 3455 5674 3474
rect 5684 3468 5700 3469
rect 5683 3466 5700 3468
rect 5684 3461 5700 3466
rect 5674 3454 5680 3455
rect 5683 3454 5712 3461
rect 5601 3453 5712 3454
rect 5601 3452 5718 3453
rect 5277 3444 5328 3452
rect 5375 3444 5409 3452
rect 5277 3432 5302 3444
rect 5309 3432 5328 3444
rect 5382 3442 5409 3444
rect 5418 3442 5639 3452
rect 5674 3449 5680 3452
rect 5382 3438 5639 3442
rect 5277 3424 5328 3432
rect 5375 3424 5639 3438
rect 5683 3444 5718 3452
rect 5229 3376 5248 3410
rect 5293 3416 5322 3424
rect 5293 3410 5310 3416
rect 5293 3408 5327 3410
rect 5375 3408 5391 3424
rect 5392 3414 5600 3424
rect 5601 3414 5617 3424
rect 5665 3420 5680 3435
rect 5683 3432 5684 3444
rect 5691 3432 5718 3444
rect 5683 3424 5718 3432
rect 5683 3423 5712 3424
rect 5403 3410 5617 3414
rect 5418 3408 5617 3410
rect 5652 3410 5665 3420
rect 5683 3410 5700 3423
rect 5652 3408 5700 3410
rect 5294 3404 5327 3408
rect 5290 3402 5327 3404
rect 5290 3401 5357 3402
rect 5290 3396 5321 3401
rect 5327 3396 5357 3401
rect 5290 3392 5357 3396
rect 5263 3389 5357 3392
rect 5263 3382 5312 3389
rect 5263 3376 5293 3382
rect 5312 3377 5317 3382
rect 5229 3360 5309 3376
rect 5321 3368 5357 3389
rect 5418 3384 5607 3408
rect 5652 3407 5699 3408
rect 5665 3402 5699 3407
rect 5433 3381 5607 3384
rect 5426 3378 5607 3381
rect 5635 3401 5699 3402
rect 5229 3358 5248 3360
rect 5263 3358 5297 3360
rect 5229 3342 5309 3358
rect 5229 3336 5248 3342
rect 4945 3310 5048 3320
rect 4899 3308 5048 3310
rect 5069 3308 5104 3320
rect 4738 3306 4900 3308
rect 4750 3286 4769 3306
rect 4784 3304 4814 3306
rect 4633 3278 4674 3286
rect 4756 3282 4769 3286
rect 4821 3290 4900 3306
rect 4932 3306 5104 3308
rect 4932 3290 5011 3306
rect 5018 3304 5048 3306
rect 4596 3268 4625 3278
rect 4639 3268 4668 3278
rect 4683 3268 4713 3282
rect 4756 3268 4799 3282
rect 4821 3278 5011 3290
rect 5076 3286 5082 3306
rect 4806 3268 4836 3278
rect 4837 3268 4995 3278
rect 4999 3268 5029 3278
rect 5033 3268 5063 3282
rect 5091 3268 5104 3306
rect 5176 3320 5205 3336
rect 5219 3320 5248 3336
rect 5263 3326 5293 3342
rect 5321 3320 5327 3368
rect 5330 3362 5349 3368
rect 5364 3362 5394 3370
rect 5330 3354 5394 3362
rect 5330 3338 5410 3354
rect 5426 3347 5488 3378
rect 5504 3347 5566 3378
rect 5635 3376 5684 3401
rect 5699 3376 5729 3392
rect 5598 3362 5628 3370
rect 5635 3368 5745 3376
rect 5598 3354 5643 3362
rect 5330 3336 5349 3338
rect 5364 3336 5410 3338
rect 5330 3320 5410 3336
rect 5437 3334 5472 3347
rect 5513 3344 5550 3347
rect 5513 3342 5555 3344
rect 5442 3331 5472 3334
rect 5451 3327 5458 3331
rect 5458 3326 5459 3327
rect 5417 3320 5427 3326
rect 5176 3312 5211 3320
rect 5176 3286 5177 3312
rect 5184 3286 5211 3312
rect 5119 3268 5149 3282
rect 5176 3278 5211 3286
rect 5213 3312 5254 3320
rect 5213 3286 5228 3312
rect 5235 3286 5254 3312
rect 5318 3308 5349 3320
rect 5364 3308 5467 3320
rect 5479 3310 5505 3336
rect 5520 3331 5550 3342
rect 5582 3338 5644 3354
rect 5582 3336 5628 3338
rect 5582 3320 5644 3336
rect 5656 3320 5662 3368
rect 5665 3360 5745 3368
rect 5665 3358 5684 3360
rect 5699 3358 5733 3360
rect 5665 3342 5745 3358
rect 5665 3320 5684 3342
rect 5699 3326 5729 3342
rect 5757 3336 5763 3410
rect 5766 3336 5785 3480
rect 5800 3336 5806 3480
rect 5815 3410 5828 3480
rect 5880 3476 5902 3480
rect 5873 3454 5902 3468
rect 5955 3454 5971 3468
rect 6009 3464 6015 3466
rect 6022 3464 6130 3480
rect 6137 3464 6143 3466
rect 6151 3464 6166 3480
rect 6232 3474 6251 3477
rect 5873 3452 5971 3454
rect 5998 3452 6166 3464
rect 6181 3454 6197 3468
rect 6232 3455 6254 3474
rect 6264 3468 6280 3469
rect 6263 3466 6280 3468
rect 6264 3461 6280 3466
rect 6254 3454 6260 3455
rect 6263 3454 6292 3461
rect 6181 3453 6292 3454
rect 6181 3452 6298 3453
rect 5857 3444 5908 3452
rect 5955 3444 5989 3452
rect 5857 3432 5882 3444
rect 5889 3432 5908 3444
rect 5962 3442 5989 3444
rect 5998 3442 6219 3452
rect 6254 3449 6260 3452
rect 5962 3438 6219 3442
rect 5857 3424 5908 3432
rect 5955 3424 6219 3438
rect 6263 3444 6298 3452
rect 5809 3376 5828 3410
rect 5873 3416 5902 3424
rect 5873 3410 5890 3416
rect 5873 3408 5907 3410
rect 5955 3408 5971 3424
rect 5972 3414 6180 3424
rect 6181 3414 6197 3424
rect 6245 3420 6260 3435
rect 6263 3432 6264 3444
rect 6271 3432 6298 3444
rect 6263 3424 6298 3432
rect 6263 3423 6292 3424
rect 5983 3410 6197 3414
rect 5998 3408 6197 3410
rect 6232 3410 6245 3420
rect 6263 3410 6280 3423
rect 6232 3408 6280 3410
rect 5874 3404 5907 3408
rect 5870 3402 5907 3404
rect 5870 3401 5937 3402
rect 5870 3396 5901 3401
rect 5907 3396 5937 3401
rect 5870 3392 5937 3396
rect 5843 3389 5937 3392
rect 5843 3382 5892 3389
rect 5843 3376 5873 3382
rect 5892 3377 5897 3382
rect 5809 3360 5889 3376
rect 5901 3368 5937 3389
rect 5998 3384 6187 3408
rect 6232 3407 6279 3408
rect 6245 3402 6279 3407
rect 6013 3381 6187 3384
rect 6006 3378 6187 3381
rect 6215 3401 6279 3402
rect 5809 3358 5828 3360
rect 5843 3358 5877 3360
rect 5809 3342 5889 3358
rect 5809 3336 5828 3342
rect 5525 3310 5628 3320
rect 5479 3308 5628 3310
rect 5649 3308 5684 3320
rect 5318 3306 5480 3308
rect 5330 3286 5349 3306
rect 5364 3304 5394 3306
rect 5213 3278 5254 3286
rect 5336 3282 5349 3286
rect 5401 3290 5480 3306
rect 5512 3306 5684 3308
rect 5512 3290 5591 3306
rect 5598 3304 5628 3306
rect 5176 3268 5205 3278
rect 5219 3268 5248 3278
rect 5263 3268 5293 3282
rect 5336 3268 5379 3282
rect 5401 3278 5591 3290
rect 5656 3286 5662 3306
rect 5386 3268 5416 3278
rect 5417 3268 5575 3278
rect 5579 3268 5609 3278
rect 5613 3268 5643 3282
rect 5671 3268 5684 3306
rect 5756 3320 5785 3336
rect 5799 3320 5828 3336
rect 5843 3326 5873 3342
rect 5901 3320 5907 3368
rect 5910 3362 5929 3368
rect 5944 3362 5974 3370
rect 5910 3354 5974 3362
rect 5910 3338 5990 3354
rect 6006 3347 6068 3378
rect 6084 3347 6146 3378
rect 6215 3376 6264 3401
rect 6279 3376 6309 3392
rect 6178 3362 6208 3370
rect 6215 3368 6325 3376
rect 6178 3354 6223 3362
rect 5910 3336 5929 3338
rect 5944 3336 5990 3338
rect 5910 3320 5990 3336
rect 6017 3334 6052 3347
rect 6093 3344 6130 3347
rect 6093 3342 6135 3344
rect 6022 3331 6052 3334
rect 6031 3327 6038 3331
rect 6038 3326 6039 3327
rect 5997 3320 6007 3326
rect 5756 3312 5791 3320
rect 5756 3286 5757 3312
rect 5764 3286 5791 3312
rect 5699 3268 5729 3282
rect 5756 3278 5791 3286
rect 5793 3312 5834 3320
rect 5793 3286 5808 3312
rect 5815 3286 5834 3312
rect 5898 3308 5929 3320
rect 5944 3308 6047 3320
rect 6059 3310 6085 3336
rect 6100 3331 6130 3342
rect 6162 3338 6224 3354
rect 6162 3336 6208 3338
rect 6162 3320 6224 3336
rect 6236 3320 6242 3368
rect 6245 3360 6325 3368
rect 6245 3358 6264 3360
rect 6279 3358 6313 3360
rect 6245 3342 6325 3358
rect 6245 3320 6264 3342
rect 6279 3326 6309 3342
rect 6337 3336 6343 3410
rect 6346 3336 6365 3480
rect 6380 3336 6386 3480
rect 6395 3410 6408 3480
rect 6460 3476 6482 3480
rect 6453 3454 6482 3468
rect 6535 3454 6551 3468
rect 6589 3464 6595 3466
rect 6602 3464 6710 3480
rect 6717 3464 6723 3466
rect 6731 3464 6746 3480
rect 6812 3474 6831 3477
rect 6453 3452 6551 3454
rect 6578 3452 6746 3464
rect 6761 3454 6777 3468
rect 6812 3455 6834 3474
rect 6844 3468 6860 3469
rect 6843 3466 6860 3468
rect 6844 3461 6860 3466
rect 6834 3454 6840 3455
rect 6843 3454 6872 3461
rect 6761 3453 6872 3454
rect 6761 3452 6878 3453
rect 6437 3444 6488 3452
rect 6535 3444 6569 3452
rect 6437 3432 6462 3444
rect 6469 3432 6488 3444
rect 6542 3442 6569 3444
rect 6578 3442 6799 3452
rect 6834 3449 6840 3452
rect 6542 3438 6799 3442
rect 6437 3424 6488 3432
rect 6535 3424 6799 3438
rect 6843 3444 6878 3452
rect 6389 3376 6408 3410
rect 6453 3416 6482 3424
rect 6453 3410 6470 3416
rect 6453 3408 6487 3410
rect 6535 3408 6551 3424
rect 6552 3414 6760 3424
rect 6761 3414 6777 3424
rect 6825 3420 6840 3435
rect 6843 3432 6844 3444
rect 6851 3432 6878 3444
rect 6843 3424 6878 3432
rect 6843 3423 6872 3424
rect 6563 3410 6777 3414
rect 6578 3408 6777 3410
rect 6812 3410 6825 3420
rect 6843 3410 6860 3423
rect 6812 3408 6860 3410
rect 6454 3404 6487 3408
rect 6450 3402 6487 3404
rect 6450 3401 6517 3402
rect 6450 3396 6481 3401
rect 6487 3396 6517 3401
rect 6450 3392 6517 3396
rect 6423 3389 6517 3392
rect 6423 3382 6472 3389
rect 6423 3376 6453 3382
rect 6472 3377 6477 3382
rect 6389 3360 6469 3376
rect 6481 3368 6517 3389
rect 6578 3384 6767 3408
rect 6812 3407 6859 3408
rect 6825 3402 6859 3407
rect 6593 3381 6767 3384
rect 6586 3378 6767 3381
rect 6795 3401 6859 3402
rect 6389 3358 6408 3360
rect 6423 3358 6457 3360
rect 6389 3342 6469 3358
rect 6389 3336 6408 3342
rect 6105 3310 6208 3320
rect 6059 3308 6208 3310
rect 6229 3308 6264 3320
rect 5898 3306 6060 3308
rect 5910 3286 5929 3306
rect 5944 3304 5974 3306
rect 5793 3278 5834 3286
rect 5916 3282 5929 3286
rect 5981 3290 6060 3306
rect 6092 3306 6264 3308
rect 6092 3290 6171 3306
rect 6178 3304 6208 3306
rect 5756 3268 5785 3278
rect 5799 3268 5828 3278
rect 5843 3268 5873 3282
rect 5916 3268 5959 3282
rect 5981 3278 6171 3290
rect 6236 3286 6242 3306
rect 5966 3268 5996 3278
rect 5997 3268 6155 3278
rect 6159 3268 6189 3278
rect 6193 3268 6223 3282
rect 6251 3268 6264 3306
rect 6336 3320 6365 3336
rect 6379 3320 6408 3336
rect 6423 3326 6453 3342
rect 6481 3320 6487 3368
rect 6490 3362 6509 3368
rect 6524 3362 6554 3370
rect 6490 3354 6554 3362
rect 6490 3338 6570 3354
rect 6586 3347 6648 3378
rect 6664 3347 6726 3378
rect 6795 3376 6844 3401
rect 6859 3376 6889 3392
rect 6758 3362 6788 3370
rect 6795 3368 6905 3376
rect 6758 3354 6803 3362
rect 6490 3336 6509 3338
rect 6524 3336 6570 3338
rect 6490 3320 6570 3336
rect 6597 3334 6632 3347
rect 6673 3344 6710 3347
rect 6673 3342 6715 3344
rect 6602 3331 6632 3334
rect 6611 3327 6618 3331
rect 6618 3326 6619 3327
rect 6577 3320 6587 3326
rect 6336 3312 6371 3320
rect 6336 3286 6337 3312
rect 6344 3286 6371 3312
rect 6279 3268 6309 3282
rect 6336 3278 6371 3286
rect 6373 3312 6414 3320
rect 6373 3286 6388 3312
rect 6395 3286 6414 3312
rect 6478 3308 6509 3320
rect 6524 3308 6627 3320
rect 6639 3310 6665 3336
rect 6680 3331 6710 3342
rect 6742 3338 6804 3354
rect 6742 3336 6788 3338
rect 6742 3320 6804 3336
rect 6816 3320 6822 3368
rect 6825 3360 6905 3368
rect 6825 3358 6844 3360
rect 6859 3358 6893 3360
rect 6825 3342 6905 3358
rect 6825 3320 6844 3342
rect 6859 3326 6889 3342
rect 6917 3336 6923 3410
rect 6926 3336 6945 3480
rect 6960 3336 6966 3480
rect 6975 3410 6988 3480
rect 7040 3476 7062 3480
rect 7033 3454 7062 3468
rect 7115 3454 7131 3468
rect 7169 3464 7175 3466
rect 7182 3464 7290 3480
rect 7297 3464 7303 3466
rect 7311 3464 7326 3480
rect 7392 3474 7411 3477
rect 7033 3452 7131 3454
rect 7158 3452 7326 3464
rect 7341 3454 7357 3468
rect 7392 3455 7414 3474
rect 7424 3468 7440 3469
rect 7423 3466 7440 3468
rect 7424 3461 7440 3466
rect 7414 3454 7420 3455
rect 7423 3454 7452 3461
rect 7341 3453 7452 3454
rect 7341 3452 7458 3453
rect 7017 3444 7068 3452
rect 7115 3444 7149 3452
rect 7017 3432 7042 3444
rect 7049 3432 7068 3444
rect 7122 3442 7149 3444
rect 7158 3442 7379 3452
rect 7414 3449 7420 3452
rect 7122 3438 7379 3442
rect 7017 3424 7068 3432
rect 7115 3424 7379 3438
rect 7423 3444 7458 3452
rect 6969 3376 6988 3410
rect 7033 3416 7062 3424
rect 7033 3410 7050 3416
rect 7033 3408 7067 3410
rect 7115 3408 7131 3424
rect 7132 3414 7340 3424
rect 7341 3414 7357 3424
rect 7405 3420 7420 3435
rect 7423 3432 7424 3444
rect 7431 3432 7458 3444
rect 7423 3424 7458 3432
rect 7423 3423 7452 3424
rect 7143 3410 7357 3414
rect 7158 3408 7357 3410
rect 7392 3410 7405 3420
rect 7423 3410 7440 3423
rect 7392 3408 7440 3410
rect 7034 3404 7067 3408
rect 7030 3402 7067 3404
rect 7030 3401 7097 3402
rect 7030 3396 7061 3401
rect 7067 3396 7097 3401
rect 7030 3392 7097 3396
rect 7003 3389 7097 3392
rect 7003 3382 7052 3389
rect 7003 3376 7033 3382
rect 7052 3377 7057 3382
rect 6969 3360 7049 3376
rect 7061 3368 7097 3389
rect 7158 3384 7347 3408
rect 7392 3407 7439 3408
rect 7405 3402 7439 3407
rect 7173 3381 7347 3384
rect 7166 3378 7347 3381
rect 7375 3401 7439 3402
rect 6969 3358 6988 3360
rect 7003 3358 7037 3360
rect 6969 3342 7049 3358
rect 6969 3336 6988 3342
rect 6685 3310 6788 3320
rect 6639 3308 6788 3310
rect 6809 3308 6844 3320
rect 6478 3306 6640 3308
rect 6490 3286 6509 3306
rect 6524 3304 6554 3306
rect 6373 3278 6414 3286
rect 6496 3282 6509 3286
rect 6561 3290 6640 3306
rect 6672 3306 6844 3308
rect 6672 3290 6751 3306
rect 6758 3304 6788 3306
rect 6336 3268 6365 3278
rect 6379 3268 6408 3278
rect 6423 3268 6453 3282
rect 6496 3268 6539 3282
rect 6561 3278 6751 3290
rect 6816 3286 6822 3306
rect 6546 3268 6576 3278
rect 6577 3268 6735 3278
rect 6739 3268 6769 3278
rect 6773 3268 6803 3282
rect 6831 3268 6844 3306
rect 6916 3320 6945 3336
rect 6959 3320 6988 3336
rect 7003 3326 7033 3342
rect 7061 3320 7067 3368
rect 7070 3362 7089 3368
rect 7104 3362 7134 3370
rect 7070 3354 7134 3362
rect 7070 3338 7150 3354
rect 7166 3347 7228 3378
rect 7244 3347 7306 3378
rect 7375 3376 7424 3401
rect 7439 3376 7469 3392
rect 7338 3362 7368 3370
rect 7375 3368 7485 3376
rect 7338 3354 7383 3362
rect 7070 3336 7089 3338
rect 7104 3336 7150 3338
rect 7070 3320 7150 3336
rect 7177 3334 7212 3347
rect 7253 3344 7290 3347
rect 7253 3342 7295 3344
rect 7182 3331 7212 3334
rect 7191 3327 7198 3331
rect 7198 3326 7199 3327
rect 7157 3320 7167 3326
rect 6916 3312 6951 3320
rect 6916 3286 6917 3312
rect 6924 3286 6951 3312
rect 6859 3268 6889 3282
rect 6916 3278 6951 3286
rect 6953 3312 6994 3320
rect 6953 3286 6968 3312
rect 6975 3286 6994 3312
rect 7058 3308 7089 3320
rect 7104 3308 7207 3320
rect 7219 3310 7245 3336
rect 7260 3331 7290 3342
rect 7322 3338 7384 3354
rect 7322 3336 7368 3338
rect 7322 3320 7384 3336
rect 7396 3320 7402 3368
rect 7405 3360 7485 3368
rect 7405 3358 7424 3360
rect 7439 3358 7473 3360
rect 7405 3342 7485 3358
rect 7405 3320 7424 3342
rect 7439 3326 7469 3342
rect 7497 3336 7503 3410
rect 7506 3336 7525 3480
rect 7540 3336 7546 3480
rect 7555 3410 7568 3480
rect 7620 3476 7642 3480
rect 7613 3454 7642 3468
rect 7695 3454 7711 3468
rect 7749 3464 7755 3466
rect 7762 3464 7870 3480
rect 7877 3464 7883 3466
rect 7891 3464 7906 3480
rect 7972 3474 7991 3477
rect 7613 3452 7711 3454
rect 7738 3452 7906 3464
rect 7921 3454 7937 3468
rect 7972 3455 7994 3474
rect 8004 3468 8020 3469
rect 8003 3466 8020 3468
rect 8004 3461 8020 3466
rect 7994 3454 8000 3455
rect 8003 3454 8032 3461
rect 7921 3453 8032 3454
rect 7921 3452 8038 3453
rect 7597 3444 7648 3452
rect 7695 3444 7729 3452
rect 7597 3432 7622 3444
rect 7629 3432 7648 3444
rect 7702 3442 7729 3444
rect 7738 3442 7959 3452
rect 7994 3449 8000 3452
rect 7702 3438 7959 3442
rect 7597 3424 7648 3432
rect 7695 3424 7959 3438
rect 8003 3444 8038 3452
rect 7549 3376 7568 3410
rect 7613 3416 7642 3424
rect 7613 3410 7630 3416
rect 7613 3408 7647 3410
rect 7695 3408 7711 3424
rect 7712 3414 7920 3424
rect 7921 3414 7937 3424
rect 7985 3420 8000 3435
rect 8003 3432 8004 3444
rect 8011 3432 8038 3444
rect 8003 3424 8038 3432
rect 8003 3423 8032 3424
rect 7723 3410 7937 3414
rect 7738 3408 7937 3410
rect 7972 3410 7985 3420
rect 8003 3410 8020 3423
rect 7972 3408 8020 3410
rect 7614 3404 7647 3408
rect 7610 3402 7647 3404
rect 7610 3401 7677 3402
rect 7610 3396 7641 3401
rect 7647 3396 7677 3401
rect 7610 3392 7677 3396
rect 7583 3389 7677 3392
rect 7583 3382 7632 3389
rect 7583 3376 7613 3382
rect 7632 3377 7637 3382
rect 7549 3360 7629 3376
rect 7641 3368 7677 3389
rect 7738 3384 7927 3408
rect 7972 3407 8019 3408
rect 7985 3402 8019 3407
rect 7753 3381 7927 3384
rect 7746 3378 7927 3381
rect 7955 3401 8019 3402
rect 7549 3358 7568 3360
rect 7583 3358 7617 3360
rect 7549 3342 7629 3358
rect 7549 3336 7568 3342
rect 7265 3310 7368 3320
rect 7219 3308 7368 3310
rect 7389 3308 7424 3320
rect 7058 3306 7220 3308
rect 7070 3286 7089 3306
rect 7104 3304 7134 3306
rect 6953 3278 6994 3286
rect 7076 3282 7089 3286
rect 7141 3290 7220 3306
rect 7252 3306 7424 3308
rect 7252 3290 7331 3306
rect 7338 3304 7368 3306
rect 6916 3268 6945 3278
rect 6959 3268 6988 3278
rect 7003 3268 7033 3282
rect 7076 3268 7119 3282
rect 7141 3278 7331 3290
rect 7396 3286 7402 3306
rect 7126 3268 7156 3278
rect 7157 3268 7315 3278
rect 7319 3268 7349 3278
rect 7353 3268 7383 3282
rect 7411 3268 7424 3306
rect 7496 3320 7525 3336
rect 7539 3320 7568 3336
rect 7583 3326 7613 3342
rect 7641 3320 7647 3368
rect 7650 3362 7669 3368
rect 7684 3362 7714 3370
rect 7650 3354 7714 3362
rect 7650 3338 7730 3354
rect 7746 3347 7808 3378
rect 7824 3347 7886 3378
rect 7955 3376 8004 3401
rect 8019 3376 8049 3392
rect 7918 3362 7948 3370
rect 7955 3368 8065 3376
rect 7918 3354 7963 3362
rect 7650 3336 7669 3338
rect 7684 3336 7730 3338
rect 7650 3320 7730 3336
rect 7757 3334 7792 3347
rect 7833 3344 7870 3347
rect 7833 3342 7875 3344
rect 7762 3331 7792 3334
rect 7771 3327 7778 3331
rect 7778 3326 7779 3327
rect 7737 3320 7747 3326
rect 7496 3312 7531 3320
rect 7496 3286 7497 3312
rect 7504 3286 7531 3312
rect 7439 3268 7469 3282
rect 7496 3278 7531 3286
rect 7533 3312 7574 3320
rect 7533 3286 7548 3312
rect 7555 3286 7574 3312
rect 7638 3308 7669 3320
rect 7684 3308 7787 3320
rect 7799 3310 7825 3336
rect 7840 3331 7870 3342
rect 7902 3338 7964 3354
rect 7902 3336 7948 3338
rect 7902 3320 7964 3336
rect 7976 3320 7982 3368
rect 7985 3360 8065 3368
rect 7985 3358 8004 3360
rect 8019 3358 8053 3360
rect 7985 3342 8065 3358
rect 7985 3320 8004 3342
rect 8019 3326 8049 3342
rect 8077 3336 8083 3410
rect 8086 3336 8105 3480
rect 8120 3336 8126 3480
rect 8135 3410 8148 3480
rect 8200 3476 8222 3480
rect 8193 3454 8222 3468
rect 8275 3454 8291 3468
rect 8329 3464 8335 3466
rect 8342 3464 8450 3480
rect 8457 3464 8463 3466
rect 8471 3464 8486 3480
rect 8552 3474 8571 3477
rect 8193 3452 8291 3454
rect 8318 3452 8486 3464
rect 8501 3454 8517 3468
rect 8552 3455 8574 3474
rect 8584 3468 8600 3469
rect 8583 3466 8600 3468
rect 8584 3461 8600 3466
rect 8574 3454 8580 3455
rect 8583 3454 8612 3461
rect 8501 3453 8612 3454
rect 8501 3452 8618 3453
rect 8177 3444 8228 3452
rect 8275 3444 8309 3452
rect 8177 3432 8202 3444
rect 8209 3432 8228 3444
rect 8282 3442 8309 3444
rect 8318 3442 8539 3452
rect 8574 3449 8580 3452
rect 8282 3438 8539 3442
rect 8177 3424 8228 3432
rect 8275 3424 8539 3438
rect 8583 3444 8618 3452
rect 8129 3376 8148 3410
rect 8193 3416 8222 3424
rect 8193 3410 8210 3416
rect 8193 3408 8227 3410
rect 8275 3408 8291 3424
rect 8292 3414 8500 3424
rect 8501 3414 8517 3424
rect 8565 3420 8580 3435
rect 8583 3432 8584 3444
rect 8591 3432 8618 3444
rect 8583 3424 8618 3432
rect 8583 3423 8612 3424
rect 8303 3410 8517 3414
rect 8318 3408 8517 3410
rect 8552 3410 8565 3420
rect 8583 3410 8600 3423
rect 8552 3408 8600 3410
rect 8194 3404 8227 3408
rect 8190 3402 8227 3404
rect 8190 3401 8257 3402
rect 8190 3396 8221 3401
rect 8227 3396 8257 3401
rect 8190 3392 8257 3396
rect 8163 3389 8257 3392
rect 8163 3382 8212 3389
rect 8163 3376 8193 3382
rect 8212 3377 8217 3382
rect 8129 3360 8209 3376
rect 8221 3368 8257 3389
rect 8318 3384 8507 3408
rect 8552 3407 8599 3408
rect 8565 3402 8599 3407
rect 8333 3381 8507 3384
rect 8326 3378 8507 3381
rect 8535 3401 8599 3402
rect 8129 3358 8148 3360
rect 8163 3358 8197 3360
rect 8129 3342 8209 3358
rect 8129 3336 8148 3342
rect 7845 3310 7948 3320
rect 7799 3308 7948 3310
rect 7969 3308 8004 3320
rect 7638 3306 7800 3308
rect 7650 3286 7669 3306
rect 7684 3304 7714 3306
rect 7533 3278 7574 3286
rect 7656 3282 7669 3286
rect 7721 3290 7800 3306
rect 7832 3306 8004 3308
rect 7832 3290 7911 3306
rect 7918 3304 7948 3306
rect 7496 3268 7525 3278
rect 7539 3268 7568 3278
rect 7583 3268 7613 3282
rect 7656 3268 7699 3282
rect 7721 3278 7911 3290
rect 7976 3286 7982 3306
rect 7706 3268 7736 3278
rect 7737 3268 7895 3278
rect 7899 3268 7929 3278
rect 7933 3268 7963 3282
rect 7991 3268 8004 3306
rect 8076 3320 8105 3336
rect 8119 3320 8148 3336
rect 8163 3326 8193 3342
rect 8221 3320 8227 3368
rect 8230 3362 8249 3368
rect 8264 3362 8294 3370
rect 8230 3354 8294 3362
rect 8230 3338 8310 3354
rect 8326 3347 8388 3378
rect 8404 3347 8466 3378
rect 8535 3376 8584 3401
rect 8599 3376 8629 3392
rect 8498 3362 8528 3370
rect 8535 3368 8645 3376
rect 8498 3354 8543 3362
rect 8230 3336 8249 3338
rect 8264 3336 8310 3338
rect 8230 3320 8310 3336
rect 8337 3334 8372 3347
rect 8413 3344 8450 3347
rect 8413 3342 8455 3344
rect 8342 3331 8372 3334
rect 8351 3327 8358 3331
rect 8358 3326 8359 3327
rect 8317 3320 8327 3326
rect 8076 3312 8111 3320
rect 8076 3286 8077 3312
rect 8084 3286 8111 3312
rect 8019 3268 8049 3282
rect 8076 3278 8111 3286
rect 8113 3312 8154 3320
rect 8113 3286 8128 3312
rect 8135 3286 8154 3312
rect 8218 3308 8249 3320
rect 8264 3308 8367 3320
rect 8379 3310 8405 3336
rect 8420 3331 8450 3342
rect 8482 3338 8544 3354
rect 8482 3336 8528 3338
rect 8482 3320 8544 3336
rect 8556 3320 8562 3368
rect 8565 3360 8645 3368
rect 8565 3358 8584 3360
rect 8599 3358 8633 3360
rect 8565 3342 8645 3358
rect 8565 3320 8584 3342
rect 8599 3326 8629 3342
rect 8657 3336 8663 3410
rect 8666 3336 8685 3480
rect 8700 3336 8706 3480
rect 8715 3410 8728 3480
rect 8780 3476 8802 3480
rect 8773 3454 8802 3468
rect 8855 3454 8871 3468
rect 8909 3464 8915 3466
rect 8922 3464 9030 3480
rect 9037 3464 9043 3466
rect 9051 3464 9066 3480
rect 9132 3474 9151 3477
rect 8773 3452 8871 3454
rect 8898 3452 9066 3464
rect 9081 3454 9097 3468
rect 9132 3455 9154 3474
rect 9164 3468 9180 3469
rect 9163 3466 9180 3468
rect 9164 3461 9180 3466
rect 9154 3454 9160 3455
rect 9163 3454 9192 3461
rect 9081 3453 9192 3454
rect 9081 3452 9198 3453
rect 8757 3444 8808 3452
rect 8855 3444 8889 3452
rect 8757 3432 8782 3444
rect 8789 3432 8808 3444
rect 8862 3442 8889 3444
rect 8898 3442 9119 3452
rect 9154 3449 9160 3452
rect 8862 3438 9119 3442
rect 8757 3424 8808 3432
rect 8855 3424 9119 3438
rect 9163 3444 9198 3452
rect 8709 3376 8728 3410
rect 8773 3416 8802 3424
rect 8773 3410 8790 3416
rect 8773 3408 8807 3410
rect 8855 3408 8871 3424
rect 8872 3414 9080 3424
rect 9081 3414 9097 3424
rect 9145 3420 9160 3435
rect 9163 3432 9164 3444
rect 9171 3432 9198 3444
rect 9163 3424 9198 3432
rect 9163 3423 9192 3424
rect 8883 3410 9097 3414
rect 8898 3408 9097 3410
rect 9132 3410 9145 3420
rect 9163 3410 9180 3423
rect 9132 3408 9180 3410
rect 8774 3404 8807 3408
rect 8770 3402 8807 3404
rect 8770 3401 8837 3402
rect 8770 3396 8801 3401
rect 8807 3396 8837 3401
rect 8770 3392 8837 3396
rect 8743 3389 8837 3392
rect 8743 3382 8792 3389
rect 8743 3376 8773 3382
rect 8792 3377 8797 3382
rect 8709 3360 8789 3376
rect 8801 3368 8837 3389
rect 8898 3384 9087 3408
rect 9132 3407 9179 3408
rect 9145 3402 9179 3407
rect 8913 3381 9087 3384
rect 8906 3378 9087 3381
rect 9115 3401 9179 3402
rect 8709 3358 8728 3360
rect 8743 3358 8777 3360
rect 8709 3342 8789 3358
rect 8709 3336 8728 3342
rect 8425 3310 8528 3320
rect 8379 3308 8528 3310
rect 8549 3308 8584 3320
rect 8218 3306 8380 3308
rect 8230 3286 8249 3306
rect 8264 3304 8294 3306
rect 8113 3278 8154 3286
rect 8236 3282 8249 3286
rect 8301 3290 8380 3306
rect 8412 3306 8584 3308
rect 8412 3290 8491 3306
rect 8498 3304 8528 3306
rect 8076 3268 8105 3278
rect 8119 3268 8148 3278
rect 8163 3268 8193 3282
rect 8236 3268 8279 3282
rect 8301 3278 8491 3290
rect 8556 3286 8562 3306
rect 8286 3268 8316 3278
rect 8317 3268 8475 3278
rect 8479 3268 8509 3278
rect 8513 3268 8543 3282
rect 8571 3268 8584 3306
rect 8656 3320 8685 3336
rect 8699 3320 8728 3336
rect 8743 3326 8773 3342
rect 8801 3320 8807 3368
rect 8810 3362 8829 3368
rect 8844 3362 8874 3370
rect 8810 3354 8874 3362
rect 8810 3338 8890 3354
rect 8906 3347 8968 3378
rect 8984 3347 9046 3378
rect 9115 3376 9164 3401
rect 9179 3376 9209 3392
rect 9078 3362 9108 3370
rect 9115 3368 9225 3376
rect 9078 3354 9123 3362
rect 8810 3336 8829 3338
rect 8844 3336 8890 3338
rect 8810 3320 8890 3336
rect 8917 3334 8952 3347
rect 8993 3344 9030 3347
rect 8993 3342 9035 3344
rect 8922 3331 8952 3334
rect 8931 3327 8938 3331
rect 8938 3326 8939 3327
rect 8897 3320 8907 3326
rect 8656 3312 8691 3320
rect 8656 3286 8657 3312
rect 8664 3286 8691 3312
rect 8599 3268 8629 3282
rect 8656 3278 8691 3286
rect 8693 3312 8734 3320
rect 8693 3286 8708 3312
rect 8715 3286 8734 3312
rect 8798 3308 8829 3320
rect 8844 3308 8947 3320
rect 8959 3310 8985 3336
rect 9000 3331 9030 3342
rect 9062 3338 9124 3354
rect 9062 3336 9108 3338
rect 9062 3320 9124 3336
rect 9136 3320 9142 3368
rect 9145 3360 9225 3368
rect 9145 3358 9164 3360
rect 9179 3358 9213 3360
rect 9145 3342 9225 3358
rect 9145 3320 9164 3342
rect 9179 3326 9209 3342
rect 9237 3336 9243 3410
rect 9246 3336 9265 3480
rect 9280 3336 9286 3480
rect 9295 3410 9308 3480
rect 9360 3476 9382 3480
rect 9353 3454 9382 3468
rect 9435 3454 9451 3468
rect 9489 3464 9495 3466
rect 9502 3464 9610 3480
rect 9617 3464 9623 3466
rect 9631 3464 9646 3480
rect 9712 3474 9731 3477
rect 9353 3452 9451 3454
rect 9478 3452 9646 3464
rect 9661 3454 9677 3468
rect 9712 3455 9734 3474
rect 9744 3468 9760 3469
rect 9743 3466 9760 3468
rect 9744 3461 9760 3466
rect 9734 3454 9740 3455
rect 9743 3454 9772 3461
rect 9661 3453 9772 3454
rect 9661 3452 9778 3453
rect 9337 3444 9388 3452
rect 9435 3444 9469 3452
rect 9337 3432 9362 3444
rect 9369 3432 9388 3444
rect 9442 3442 9469 3444
rect 9478 3442 9699 3452
rect 9734 3449 9740 3452
rect 9442 3438 9699 3442
rect 9337 3424 9388 3432
rect 9435 3424 9699 3438
rect 9743 3444 9778 3452
rect 9289 3376 9308 3410
rect 9353 3416 9382 3424
rect 9353 3410 9370 3416
rect 9353 3408 9387 3410
rect 9435 3408 9451 3424
rect 9452 3414 9660 3424
rect 9661 3414 9677 3424
rect 9725 3420 9740 3435
rect 9743 3432 9744 3444
rect 9751 3432 9778 3444
rect 9743 3424 9778 3432
rect 9743 3423 9772 3424
rect 9463 3410 9677 3414
rect 9478 3408 9677 3410
rect 9712 3410 9725 3420
rect 9743 3410 9760 3423
rect 9712 3408 9760 3410
rect 9354 3404 9387 3408
rect 9350 3402 9387 3404
rect 9350 3401 9417 3402
rect 9350 3396 9381 3401
rect 9387 3396 9417 3401
rect 9350 3392 9417 3396
rect 9323 3389 9417 3392
rect 9323 3382 9372 3389
rect 9323 3376 9353 3382
rect 9372 3377 9377 3382
rect 9289 3360 9369 3376
rect 9381 3368 9417 3389
rect 9478 3384 9667 3408
rect 9712 3407 9759 3408
rect 9725 3402 9759 3407
rect 9493 3381 9667 3384
rect 9486 3378 9667 3381
rect 9695 3401 9759 3402
rect 9289 3358 9308 3360
rect 9323 3358 9357 3360
rect 9289 3342 9369 3358
rect 9289 3336 9308 3342
rect 9005 3310 9108 3320
rect 8959 3308 9108 3310
rect 9129 3308 9164 3320
rect 8798 3306 8960 3308
rect 8810 3286 8829 3306
rect 8844 3304 8874 3306
rect 8693 3278 8734 3286
rect 8816 3282 8829 3286
rect 8881 3290 8960 3306
rect 8992 3306 9164 3308
rect 8992 3290 9071 3306
rect 9078 3304 9108 3306
rect 8656 3268 8685 3278
rect 8699 3268 8728 3278
rect 8743 3268 8773 3282
rect 8816 3268 8859 3282
rect 8881 3278 9071 3290
rect 9136 3286 9142 3306
rect 8866 3268 8896 3278
rect 8897 3268 9055 3278
rect 9059 3268 9089 3278
rect 9093 3268 9123 3282
rect 9151 3268 9164 3306
rect 9236 3320 9265 3336
rect 9279 3320 9308 3336
rect 9323 3326 9353 3342
rect 9381 3320 9387 3368
rect 9390 3362 9409 3368
rect 9424 3362 9454 3370
rect 9390 3354 9454 3362
rect 9390 3338 9470 3354
rect 9486 3347 9548 3378
rect 9564 3347 9626 3378
rect 9695 3376 9744 3401
rect 9759 3376 9789 3392
rect 9658 3362 9688 3370
rect 9695 3368 9805 3376
rect 9658 3354 9703 3362
rect 9390 3336 9409 3338
rect 9424 3336 9470 3338
rect 9390 3320 9470 3336
rect 9497 3334 9532 3347
rect 9573 3344 9610 3347
rect 9573 3342 9615 3344
rect 9502 3331 9532 3334
rect 9511 3327 9518 3331
rect 9518 3326 9519 3327
rect 9477 3320 9487 3326
rect 9236 3312 9271 3320
rect 9236 3286 9237 3312
rect 9244 3286 9271 3312
rect 9179 3268 9209 3282
rect 9236 3278 9271 3286
rect 9273 3312 9314 3320
rect 9273 3286 9288 3312
rect 9295 3286 9314 3312
rect 9378 3308 9409 3320
rect 9424 3308 9527 3320
rect 9539 3310 9565 3336
rect 9580 3331 9610 3342
rect 9642 3338 9704 3354
rect 9642 3336 9688 3338
rect 9642 3320 9704 3336
rect 9716 3320 9722 3368
rect 9725 3360 9805 3368
rect 9725 3358 9744 3360
rect 9759 3358 9793 3360
rect 9725 3342 9805 3358
rect 9725 3320 9744 3342
rect 9759 3326 9789 3342
rect 9817 3336 9823 3410
rect 9826 3336 9845 3480
rect 9860 3336 9866 3480
rect 9875 3410 9888 3480
rect 9940 3476 9962 3480
rect 9933 3454 9962 3468
rect 10015 3454 10031 3468
rect 10069 3464 10075 3466
rect 10082 3464 10190 3480
rect 10197 3464 10203 3466
rect 10211 3464 10226 3480
rect 10292 3474 10311 3477
rect 9933 3452 10031 3454
rect 10058 3452 10226 3464
rect 10241 3454 10257 3468
rect 10292 3455 10314 3474
rect 10324 3468 10340 3469
rect 10323 3466 10340 3468
rect 10324 3461 10340 3466
rect 10314 3454 10320 3455
rect 10323 3454 10352 3461
rect 10241 3453 10352 3454
rect 10241 3452 10358 3453
rect 9917 3444 9968 3452
rect 10015 3444 10049 3452
rect 9917 3432 9942 3444
rect 9949 3432 9968 3444
rect 10022 3442 10049 3444
rect 10058 3442 10279 3452
rect 10314 3449 10320 3452
rect 10022 3438 10279 3442
rect 9917 3424 9968 3432
rect 10015 3424 10279 3438
rect 10323 3444 10358 3452
rect 9869 3376 9888 3410
rect 9933 3416 9962 3424
rect 9933 3410 9950 3416
rect 9933 3408 9967 3410
rect 10015 3408 10031 3424
rect 10032 3414 10240 3424
rect 10241 3414 10257 3424
rect 10305 3420 10320 3435
rect 10323 3432 10324 3444
rect 10331 3432 10358 3444
rect 10323 3424 10358 3432
rect 10323 3423 10352 3424
rect 10043 3410 10257 3414
rect 10058 3408 10257 3410
rect 10292 3410 10305 3420
rect 10323 3410 10340 3423
rect 10292 3408 10340 3410
rect 9934 3404 9967 3408
rect 9930 3402 9967 3404
rect 9930 3401 9997 3402
rect 9930 3396 9961 3401
rect 9967 3396 9997 3401
rect 9930 3392 9997 3396
rect 9903 3389 9997 3392
rect 9903 3382 9952 3389
rect 9903 3376 9933 3382
rect 9952 3377 9957 3382
rect 9869 3360 9949 3376
rect 9961 3368 9997 3389
rect 10058 3384 10247 3408
rect 10292 3407 10339 3408
rect 10305 3402 10339 3407
rect 10073 3381 10247 3384
rect 10066 3378 10247 3381
rect 10275 3401 10339 3402
rect 9869 3358 9888 3360
rect 9903 3358 9937 3360
rect 9869 3342 9949 3358
rect 9869 3336 9888 3342
rect 9585 3310 9688 3320
rect 9539 3308 9688 3310
rect 9709 3308 9744 3320
rect 9378 3306 9540 3308
rect 9390 3286 9409 3306
rect 9424 3304 9454 3306
rect 9273 3278 9314 3286
rect 9396 3282 9409 3286
rect 9461 3290 9540 3306
rect 9572 3306 9744 3308
rect 9572 3290 9651 3306
rect 9658 3304 9688 3306
rect 9236 3268 9265 3278
rect 9279 3268 9308 3278
rect 9323 3268 9353 3282
rect 9396 3268 9439 3282
rect 9461 3278 9651 3290
rect 9716 3286 9722 3306
rect 9446 3268 9476 3278
rect 9477 3268 9635 3278
rect 9639 3268 9669 3278
rect 9673 3268 9703 3282
rect 9731 3268 9744 3306
rect 9816 3320 9845 3336
rect 9859 3320 9888 3336
rect 9903 3326 9933 3342
rect 9961 3320 9967 3368
rect 9970 3362 9989 3368
rect 10004 3362 10034 3370
rect 9970 3354 10034 3362
rect 9970 3338 10050 3354
rect 10066 3347 10128 3378
rect 10144 3347 10206 3378
rect 10275 3376 10324 3401
rect 10339 3376 10369 3392
rect 10238 3362 10268 3370
rect 10275 3368 10385 3376
rect 10238 3354 10283 3362
rect 9970 3336 9989 3338
rect 10004 3336 10050 3338
rect 9970 3320 10050 3336
rect 10077 3334 10112 3347
rect 10153 3344 10190 3347
rect 10153 3342 10195 3344
rect 10082 3331 10112 3334
rect 10091 3327 10098 3331
rect 10098 3326 10099 3327
rect 10057 3320 10067 3326
rect 9816 3312 9851 3320
rect 9816 3286 9817 3312
rect 9824 3286 9851 3312
rect 9759 3268 9789 3282
rect 9816 3278 9851 3286
rect 9853 3312 9894 3320
rect 9853 3286 9868 3312
rect 9875 3286 9894 3312
rect 9958 3308 9989 3320
rect 10004 3308 10107 3320
rect 10119 3310 10145 3336
rect 10160 3331 10190 3342
rect 10222 3338 10284 3354
rect 10222 3336 10268 3338
rect 10222 3320 10284 3336
rect 10296 3320 10302 3368
rect 10305 3360 10385 3368
rect 10305 3358 10324 3360
rect 10339 3358 10373 3360
rect 10305 3342 10385 3358
rect 10305 3320 10324 3342
rect 10339 3326 10369 3342
rect 10397 3336 10403 3410
rect 10406 3336 10425 3480
rect 10440 3336 10446 3480
rect 10455 3410 10468 3480
rect 10520 3476 10542 3480
rect 10513 3454 10542 3468
rect 10595 3454 10611 3468
rect 10649 3464 10655 3466
rect 10662 3464 10770 3480
rect 10777 3464 10783 3466
rect 10791 3464 10806 3480
rect 10872 3474 10891 3477
rect 10513 3452 10611 3454
rect 10638 3452 10806 3464
rect 10821 3454 10837 3468
rect 10872 3455 10894 3474
rect 10904 3468 10920 3469
rect 10903 3466 10920 3468
rect 10904 3461 10920 3466
rect 10894 3454 10900 3455
rect 10903 3454 10932 3461
rect 10821 3453 10932 3454
rect 10821 3452 10938 3453
rect 10497 3444 10548 3452
rect 10595 3444 10629 3452
rect 10497 3432 10522 3444
rect 10529 3432 10548 3444
rect 10602 3442 10629 3444
rect 10638 3442 10859 3452
rect 10894 3449 10900 3452
rect 10602 3438 10859 3442
rect 10497 3424 10548 3432
rect 10595 3424 10859 3438
rect 10903 3444 10938 3452
rect 10449 3376 10468 3410
rect 10513 3416 10542 3424
rect 10513 3410 10530 3416
rect 10513 3408 10547 3410
rect 10595 3408 10611 3424
rect 10612 3414 10820 3424
rect 10821 3414 10837 3424
rect 10885 3420 10900 3435
rect 10903 3432 10904 3444
rect 10911 3432 10938 3444
rect 10903 3424 10938 3432
rect 10903 3423 10932 3424
rect 10623 3410 10837 3414
rect 10638 3408 10837 3410
rect 10872 3410 10885 3420
rect 10903 3410 10920 3423
rect 10872 3408 10920 3410
rect 10514 3404 10547 3408
rect 10510 3402 10547 3404
rect 10510 3401 10577 3402
rect 10510 3396 10541 3401
rect 10547 3396 10577 3401
rect 10510 3392 10577 3396
rect 10483 3389 10577 3392
rect 10483 3382 10532 3389
rect 10483 3376 10513 3382
rect 10532 3377 10537 3382
rect 10449 3360 10529 3376
rect 10541 3368 10577 3389
rect 10638 3384 10827 3408
rect 10872 3407 10919 3408
rect 10885 3402 10919 3407
rect 10653 3381 10827 3384
rect 10646 3378 10827 3381
rect 10855 3401 10919 3402
rect 10449 3358 10468 3360
rect 10483 3358 10517 3360
rect 10449 3342 10529 3358
rect 10449 3336 10468 3342
rect 10165 3310 10268 3320
rect 10119 3308 10268 3310
rect 10289 3308 10324 3320
rect 9958 3306 10120 3308
rect 9970 3286 9989 3306
rect 10004 3304 10034 3306
rect 9853 3278 9894 3286
rect 9976 3282 9989 3286
rect 10041 3290 10120 3306
rect 10152 3306 10324 3308
rect 10152 3290 10231 3306
rect 10238 3304 10268 3306
rect 9816 3268 9845 3278
rect 9859 3268 9888 3278
rect 9903 3268 9933 3282
rect 9976 3268 10019 3282
rect 10041 3278 10231 3290
rect 10296 3286 10302 3306
rect 10026 3268 10056 3278
rect 10057 3268 10215 3278
rect 10219 3268 10249 3278
rect 10253 3268 10283 3282
rect 10311 3268 10324 3306
rect 10396 3320 10425 3336
rect 10439 3320 10468 3336
rect 10483 3326 10513 3342
rect 10541 3320 10547 3368
rect 10550 3362 10569 3368
rect 10584 3362 10614 3370
rect 10550 3354 10614 3362
rect 10550 3338 10630 3354
rect 10646 3347 10708 3378
rect 10724 3347 10786 3378
rect 10855 3376 10904 3401
rect 10919 3376 10949 3392
rect 10818 3362 10848 3370
rect 10855 3368 10965 3376
rect 10818 3354 10863 3362
rect 10550 3336 10569 3338
rect 10584 3336 10630 3338
rect 10550 3320 10630 3336
rect 10657 3334 10692 3347
rect 10733 3344 10770 3347
rect 10733 3342 10775 3344
rect 10662 3331 10692 3334
rect 10671 3327 10678 3331
rect 10678 3326 10679 3327
rect 10637 3320 10647 3326
rect 10396 3312 10431 3320
rect 10396 3286 10397 3312
rect 10404 3286 10431 3312
rect 10339 3268 10369 3282
rect 10396 3278 10431 3286
rect 10433 3312 10474 3320
rect 10433 3286 10448 3312
rect 10455 3286 10474 3312
rect 10538 3308 10569 3320
rect 10584 3308 10687 3320
rect 10699 3310 10725 3336
rect 10740 3331 10770 3342
rect 10802 3338 10864 3354
rect 10802 3336 10848 3338
rect 10802 3320 10864 3336
rect 10876 3320 10882 3368
rect 10885 3360 10965 3368
rect 10885 3358 10904 3360
rect 10919 3358 10953 3360
rect 10885 3342 10965 3358
rect 10885 3320 10904 3342
rect 10919 3326 10949 3342
rect 10977 3336 10983 3410
rect 10986 3336 11005 3480
rect 11020 3336 11026 3480
rect 11035 3410 11048 3480
rect 11100 3476 11122 3480
rect 11093 3454 11122 3468
rect 11175 3454 11191 3468
rect 11229 3464 11235 3466
rect 11242 3464 11350 3480
rect 11357 3464 11363 3466
rect 11371 3464 11386 3480
rect 11452 3474 11471 3477
rect 11093 3452 11191 3454
rect 11218 3452 11386 3464
rect 11401 3454 11417 3468
rect 11452 3455 11474 3474
rect 11484 3468 11500 3469
rect 11483 3466 11500 3468
rect 11484 3461 11500 3466
rect 11474 3454 11480 3455
rect 11483 3454 11512 3461
rect 11401 3453 11512 3454
rect 11401 3452 11518 3453
rect 11077 3444 11128 3452
rect 11175 3444 11209 3452
rect 11077 3432 11102 3444
rect 11109 3432 11128 3444
rect 11182 3442 11209 3444
rect 11218 3442 11439 3452
rect 11474 3449 11480 3452
rect 11182 3438 11439 3442
rect 11077 3424 11128 3432
rect 11175 3424 11439 3438
rect 11483 3444 11518 3452
rect 11029 3376 11048 3410
rect 11093 3416 11122 3424
rect 11093 3410 11110 3416
rect 11093 3408 11127 3410
rect 11175 3408 11191 3424
rect 11192 3414 11400 3424
rect 11401 3414 11417 3424
rect 11465 3420 11480 3435
rect 11483 3432 11484 3444
rect 11491 3432 11518 3444
rect 11483 3424 11518 3432
rect 11483 3423 11512 3424
rect 11203 3410 11417 3414
rect 11218 3408 11417 3410
rect 11452 3410 11465 3420
rect 11483 3410 11500 3423
rect 11452 3408 11500 3410
rect 11094 3404 11127 3408
rect 11090 3402 11127 3404
rect 11090 3401 11157 3402
rect 11090 3396 11121 3401
rect 11127 3396 11157 3401
rect 11090 3392 11157 3396
rect 11063 3389 11157 3392
rect 11063 3382 11112 3389
rect 11063 3376 11093 3382
rect 11112 3377 11117 3382
rect 11029 3360 11109 3376
rect 11121 3368 11157 3389
rect 11218 3384 11407 3408
rect 11452 3407 11499 3408
rect 11465 3402 11499 3407
rect 11233 3381 11407 3384
rect 11226 3378 11407 3381
rect 11435 3401 11499 3402
rect 11029 3358 11048 3360
rect 11063 3358 11097 3360
rect 11029 3342 11109 3358
rect 11029 3336 11048 3342
rect 10745 3310 10848 3320
rect 10699 3308 10848 3310
rect 10869 3308 10904 3320
rect 10538 3306 10700 3308
rect 10550 3286 10569 3306
rect 10584 3304 10614 3306
rect 10433 3278 10474 3286
rect 10556 3282 10569 3286
rect 10621 3290 10700 3306
rect 10732 3306 10904 3308
rect 10732 3290 10811 3306
rect 10818 3304 10848 3306
rect 10396 3268 10425 3278
rect 10439 3268 10468 3278
rect 10483 3268 10513 3282
rect 10556 3268 10599 3282
rect 10621 3278 10811 3290
rect 10876 3286 10882 3306
rect 10606 3268 10636 3278
rect 10637 3268 10795 3278
rect 10799 3268 10829 3278
rect 10833 3268 10863 3282
rect 10891 3268 10904 3306
rect 10976 3320 11005 3336
rect 11019 3320 11048 3336
rect 11063 3326 11093 3342
rect 11121 3320 11127 3368
rect 11130 3362 11149 3368
rect 11164 3362 11194 3370
rect 11130 3354 11194 3362
rect 11130 3338 11210 3354
rect 11226 3347 11288 3378
rect 11304 3347 11366 3378
rect 11435 3376 11484 3401
rect 11499 3376 11529 3392
rect 11398 3362 11428 3370
rect 11435 3368 11545 3376
rect 11398 3354 11443 3362
rect 11130 3336 11149 3338
rect 11164 3336 11210 3338
rect 11130 3320 11210 3336
rect 11237 3334 11272 3347
rect 11313 3344 11350 3347
rect 11313 3342 11355 3344
rect 11242 3331 11272 3334
rect 11251 3327 11258 3331
rect 11258 3326 11259 3327
rect 11217 3320 11227 3326
rect 10976 3312 11011 3320
rect 10976 3286 10977 3312
rect 10984 3286 11011 3312
rect 10919 3268 10949 3282
rect 10976 3278 11011 3286
rect 11013 3312 11054 3320
rect 11013 3286 11028 3312
rect 11035 3286 11054 3312
rect 11118 3308 11149 3320
rect 11164 3308 11267 3320
rect 11279 3310 11305 3336
rect 11320 3331 11350 3342
rect 11382 3338 11444 3354
rect 11382 3336 11428 3338
rect 11382 3320 11444 3336
rect 11456 3320 11462 3368
rect 11465 3360 11545 3368
rect 11465 3358 11484 3360
rect 11499 3358 11533 3360
rect 11465 3342 11545 3358
rect 11465 3320 11484 3342
rect 11499 3326 11529 3342
rect 11557 3336 11563 3410
rect 11566 3336 11585 3480
rect 11600 3336 11606 3480
rect 11615 3410 11628 3480
rect 11680 3476 11702 3480
rect 11673 3454 11702 3468
rect 11755 3454 11771 3468
rect 11809 3464 11815 3466
rect 11822 3464 11930 3480
rect 11937 3464 11943 3466
rect 11951 3464 11966 3480
rect 12032 3474 12051 3477
rect 11673 3452 11771 3454
rect 11798 3452 11966 3464
rect 11981 3454 11997 3468
rect 12032 3455 12054 3474
rect 12064 3468 12080 3469
rect 12063 3466 12080 3468
rect 12064 3461 12080 3466
rect 12054 3454 12060 3455
rect 12063 3454 12092 3461
rect 11981 3453 12092 3454
rect 11981 3452 12098 3453
rect 11657 3444 11708 3452
rect 11755 3444 11789 3452
rect 11657 3432 11682 3444
rect 11689 3432 11708 3444
rect 11762 3442 11789 3444
rect 11798 3442 12019 3452
rect 12054 3449 12060 3452
rect 11762 3438 12019 3442
rect 11657 3424 11708 3432
rect 11755 3424 12019 3438
rect 12063 3444 12098 3452
rect 11609 3376 11628 3410
rect 11673 3416 11702 3424
rect 11673 3410 11690 3416
rect 11673 3408 11707 3410
rect 11755 3408 11771 3424
rect 11772 3414 11980 3424
rect 11981 3414 11997 3424
rect 12045 3420 12060 3435
rect 12063 3432 12064 3444
rect 12071 3432 12098 3444
rect 12063 3424 12098 3432
rect 12063 3423 12092 3424
rect 11783 3410 11997 3414
rect 11798 3408 11997 3410
rect 12032 3410 12045 3420
rect 12063 3410 12080 3423
rect 12032 3408 12080 3410
rect 11674 3404 11707 3408
rect 11670 3402 11707 3404
rect 11670 3401 11737 3402
rect 11670 3396 11701 3401
rect 11707 3396 11737 3401
rect 11670 3392 11737 3396
rect 11643 3389 11737 3392
rect 11643 3382 11692 3389
rect 11643 3376 11673 3382
rect 11692 3377 11697 3382
rect 11609 3360 11689 3376
rect 11701 3368 11737 3389
rect 11798 3384 11987 3408
rect 12032 3407 12079 3408
rect 12045 3402 12079 3407
rect 11813 3381 11987 3384
rect 11806 3378 11987 3381
rect 12015 3401 12079 3402
rect 11609 3358 11628 3360
rect 11643 3358 11677 3360
rect 11609 3342 11689 3358
rect 11609 3336 11628 3342
rect 11325 3310 11428 3320
rect 11279 3308 11428 3310
rect 11449 3308 11484 3320
rect 11118 3306 11280 3308
rect 11130 3286 11149 3306
rect 11164 3304 11194 3306
rect 11013 3278 11054 3286
rect 11136 3282 11149 3286
rect 11201 3290 11280 3306
rect 11312 3306 11484 3308
rect 11312 3290 11391 3306
rect 11398 3304 11428 3306
rect 10976 3268 11005 3278
rect 11019 3268 11048 3278
rect 11063 3268 11093 3282
rect 11136 3268 11179 3282
rect 11201 3278 11391 3290
rect 11456 3286 11462 3306
rect 11186 3268 11216 3278
rect 11217 3268 11375 3278
rect 11379 3268 11409 3278
rect 11413 3268 11443 3282
rect 11471 3268 11484 3306
rect 11556 3320 11585 3336
rect 11599 3320 11628 3336
rect 11643 3326 11673 3342
rect 11701 3320 11707 3368
rect 11710 3362 11729 3368
rect 11744 3362 11774 3370
rect 11710 3354 11774 3362
rect 11710 3338 11790 3354
rect 11806 3347 11868 3378
rect 11884 3347 11946 3378
rect 12015 3376 12064 3401
rect 12079 3376 12109 3392
rect 11978 3362 12008 3370
rect 12015 3368 12125 3376
rect 11978 3354 12023 3362
rect 11710 3336 11729 3338
rect 11744 3336 11790 3338
rect 11710 3320 11790 3336
rect 11817 3334 11852 3347
rect 11893 3344 11930 3347
rect 11893 3342 11935 3344
rect 11822 3331 11852 3334
rect 11831 3327 11838 3331
rect 11838 3326 11839 3327
rect 11797 3320 11807 3326
rect 11556 3312 11591 3320
rect 11556 3286 11557 3312
rect 11564 3286 11591 3312
rect 11499 3268 11529 3282
rect 11556 3278 11591 3286
rect 11593 3312 11634 3320
rect 11593 3286 11608 3312
rect 11615 3286 11634 3312
rect 11698 3308 11729 3320
rect 11744 3308 11847 3320
rect 11859 3310 11885 3336
rect 11900 3331 11930 3342
rect 11962 3338 12024 3354
rect 11962 3336 12008 3338
rect 11962 3320 12024 3336
rect 12036 3320 12042 3368
rect 12045 3360 12125 3368
rect 12045 3358 12064 3360
rect 12079 3358 12113 3360
rect 12045 3342 12125 3358
rect 12045 3320 12064 3342
rect 12079 3326 12109 3342
rect 12137 3336 12143 3410
rect 12146 3336 12165 3480
rect 12180 3336 12186 3480
rect 12195 3410 12208 3480
rect 12260 3476 12282 3480
rect 12253 3454 12282 3468
rect 12335 3454 12351 3468
rect 12389 3464 12395 3466
rect 12402 3464 12510 3480
rect 12517 3464 12523 3466
rect 12531 3464 12546 3480
rect 12612 3474 12631 3477
rect 12253 3452 12351 3454
rect 12378 3452 12546 3464
rect 12561 3454 12577 3468
rect 12612 3455 12634 3474
rect 12644 3468 12660 3469
rect 12643 3466 12660 3468
rect 12644 3461 12660 3466
rect 12634 3454 12640 3455
rect 12643 3454 12672 3461
rect 12561 3453 12672 3454
rect 12561 3452 12678 3453
rect 12237 3444 12288 3452
rect 12335 3444 12369 3452
rect 12237 3432 12262 3444
rect 12269 3432 12288 3444
rect 12342 3442 12369 3444
rect 12378 3442 12599 3452
rect 12634 3449 12640 3452
rect 12342 3438 12599 3442
rect 12237 3424 12288 3432
rect 12335 3424 12599 3438
rect 12643 3444 12678 3452
rect 12189 3376 12208 3410
rect 12253 3416 12282 3424
rect 12253 3410 12270 3416
rect 12253 3408 12287 3410
rect 12335 3408 12351 3424
rect 12352 3414 12560 3424
rect 12561 3414 12577 3424
rect 12625 3420 12640 3435
rect 12643 3432 12644 3444
rect 12651 3432 12678 3444
rect 12643 3424 12678 3432
rect 12643 3423 12672 3424
rect 12363 3410 12577 3414
rect 12378 3408 12577 3410
rect 12612 3410 12625 3420
rect 12643 3410 12660 3423
rect 12612 3408 12660 3410
rect 12254 3404 12287 3408
rect 12250 3402 12287 3404
rect 12250 3401 12317 3402
rect 12250 3396 12281 3401
rect 12287 3396 12317 3401
rect 12250 3392 12317 3396
rect 12223 3389 12317 3392
rect 12223 3382 12272 3389
rect 12223 3376 12253 3382
rect 12272 3377 12277 3382
rect 12189 3360 12269 3376
rect 12281 3368 12317 3389
rect 12378 3384 12567 3408
rect 12612 3407 12659 3408
rect 12625 3402 12659 3407
rect 12393 3381 12567 3384
rect 12386 3378 12567 3381
rect 12595 3401 12659 3402
rect 12189 3358 12208 3360
rect 12223 3358 12257 3360
rect 12189 3342 12269 3358
rect 12189 3336 12208 3342
rect 11905 3310 12008 3320
rect 11859 3308 12008 3310
rect 12029 3308 12064 3320
rect 11698 3306 11860 3308
rect 11710 3286 11729 3306
rect 11744 3304 11774 3306
rect 11593 3278 11634 3286
rect 11716 3282 11729 3286
rect 11781 3290 11860 3306
rect 11892 3306 12064 3308
rect 11892 3290 11971 3306
rect 11978 3304 12008 3306
rect 11556 3268 11585 3278
rect 11599 3268 11628 3278
rect 11643 3268 11673 3282
rect 11716 3268 11759 3282
rect 11781 3278 11971 3290
rect 12036 3286 12042 3306
rect 11766 3268 11796 3278
rect 11797 3268 11955 3278
rect 11959 3268 11989 3278
rect 11993 3268 12023 3282
rect 12051 3268 12064 3306
rect 12136 3320 12165 3336
rect 12179 3320 12208 3336
rect 12223 3326 12253 3342
rect 12281 3320 12287 3368
rect 12290 3362 12309 3368
rect 12324 3362 12354 3370
rect 12290 3354 12354 3362
rect 12290 3338 12370 3354
rect 12386 3347 12448 3378
rect 12464 3347 12526 3378
rect 12595 3376 12644 3401
rect 12659 3376 12689 3392
rect 12558 3362 12588 3370
rect 12595 3368 12705 3376
rect 12558 3354 12603 3362
rect 12290 3336 12309 3338
rect 12324 3336 12370 3338
rect 12290 3320 12370 3336
rect 12397 3334 12432 3347
rect 12473 3344 12510 3347
rect 12473 3342 12515 3344
rect 12402 3331 12432 3334
rect 12411 3327 12418 3331
rect 12418 3326 12419 3327
rect 12377 3320 12387 3326
rect 12136 3312 12171 3320
rect 12136 3286 12137 3312
rect 12144 3286 12171 3312
rect 12079 3268 12109 3282
rect 12136 3278 12171 3286
rect 12173 3312 12214 3320
rect 12173 3286 12188 3312
rect 12195 3286 12214 3312
rect 12278 3308 12309 3320
rect 12324 3308 12427 3320
rect 12439 3310 12465 3336
rect 12480 3331 12510 3342
rect 12542 3338 12604 3354
rect 12542 3336 12588 3338
rect 12542 3320 12604 3336
rect 12616 3320 12622 3368
rect 12625 3360 12705 3368
rect 12625 3358 12644 3360
rect 12659 3358 12693 3360
rect 12625 3342 12705 3358
rect 12625 3320 12644 3342
rect 12659 3326 12689 3342
rect 12717 3336 12723 3410
rect 12726 3336 12745 3480
rect 12760 3336 12766 3480
rect 12775 3410 12788 3480
rect 12840 3476 12862 3480
rect 12833 3454 12862 3468
rect 12915 3454 12931 3468
rect 12969 3464 12975 3466
rect 12982 3464 13090 3480
rect 13097 3464 13103 3466
rect 13111 3464 13126 3480
rect 13192 3474 13211 3477
rect 12833 3452 12931 3454
rect 12958 3452 13126 3464
rect 13141 3454 13157 3468
rect 13192 3455 13214 3474
rect 13224 3468 13240 3469
rect 13223 3466 13240 3468
rect 13224 3461 13240 3466
rect 13214 3454 13220 3455
rect 13223 3454 13252 3461
rect 13141 3453 13252 3454
rect 13141 3452 13258 3453
rect 12817 3444 12868 3452
rect 12915 3444 12949 3452
rect 12817 3432 12842 3444
rect 12849 3432 12868 3444
rect 12922 3442 12949 3444
rect 12958 3442 13179 3452
rect 13214 3449 13220 3452
rect 12922 3438 13179 3442
rect 12817 3424 12868 3432
rect 12915 3424 13179 3438
rect 13223 3444 13258 3452
rect 12769 3376 12788 3410
rect 12833 3416 12862 3424
rect 12833 3410 12850 3416
rect 12833 3408 12867 3410
rect 12915 3408 12931 3424
rect 12932 3414 13140 3424
rect 13141 3414 13157 3424
rect 13205 3420 13220 3435
rect 13223 3432 13224 3444
rect 13231 3432 13258 3444
rect 13223 3424 13258 3432
rect 13223 3423 13252 3424
rect 12943 3410 13157 3414
rect 12958 3408 13157 3410
rect 13192 3410 13205 3420
rect 13223 3410 13240 3423
rect 13192 3408 13240 3410
rect 12834 3404 12867 3408
rect 12830 3402 12867 3404
rect 12830 3401 12897 3402
rect 12830 3396 12861 3401
rect 12867 3396 12897 3401
rect 12830 3392 12897 3396
rect 12803 3389 12897 3392
rect 12803 3382 12852 3389
rect 12803 3376 12833 3382
rect 12852 3377 12857 3382
rect 12769 3360 12849 3376
rect 12861 3368 12897 3389
rect 12958 3384 13147 3408
rect 13192 3407 13239 3408
rect 13205 3402 13239 3407
rect 12973 3381 13147 3384
rect 12966 3378 13147 3381
rect 13175 3401 13239 3402
rect 12769 3358 12788 3360
rect 12803 3358 12837 3360
rect 12769 3342 12849 3358
rect 12769 3336 12788 3342
rect 12485 3310 12588 3320
rect 12439 3308 12588 3310
rect 12609 3308 12644 3320
rect 12278 3306 12440 3308
rect 12290 3286 12309 3306
rect 12324 3304 12354 3306
rect 12173 3278 12214 3286
rect 12296 3282 12309 3286
rect 12361 3290 12440 3306
rect 12472 3306 12644 3308
rect 12472 3290 12551 3306
rect 12558 3304 12588 3306
rect 12136 3268 12165 3278
rect 12179 3268 12208 3278
rect 12223 3268 12253 3282
rect 12296 3268 12339 3282
rect 12361 3278 12551 3290
rect 12616 3286 12622 3306
rect 12346 3268 12376 3278
rect 12377 3268 12535 3278
rect 12539 3268 12569 3278
rect 12573 3268 12603 3282
rect 12631 3268 12644 3306
rect 12716 3320 12745 3336
rect 12759 3320 12788 3336
rect 12803 3326 12833 3342
rect 12861 3320 12867 3368
rect 12870 3362 12889 3368
rect 12904 3362 12934 3370
rect 12870 3354 12934 3362
rect 12870 3338 12950 3354
rect 12966 3347 13028 3378
rect 13044 3347 13106 3378
rect 13175 3376 13224 3401
rect 13239 3376 13269 3392
rect 13138 3362 13168 3370
rect 13175 3368 13285 3376
rect 13138 3354 13183 3362
rect 12870 3336 12889 3338
rect 12904 3336 12950 3338
rect 12870 3320 12950 3336
rect 12977 3334 13012 3347
rect 13053 3344 13090 3347
rect 13053 3342 13095 3344
rect 12982 3331 13012 3334
rect 12991 3327 12998 3331
rect 12998 3326 12999 3327
rect 12957 3320 12967 3326
rect 12716 3312 12751 3320
rect 12716 3286 12717 3312
rect 12724 3286 12751 3312
rect 12659 3268 12689 3282
rect 12716 3278 12751 3286
rect 12753 3312 12794 3320
rect 12753 3286 12768 3312
rect 12775 3286 12794 3312
rect 12858 3308 12889 3320
rect 12904 3308 13007 3320
rect 13019 3310 13045 3336
rect 13060 3331 13090 3342
rect 13122 3338 13184 3354
rect 13122 3336 13168 3338
rect 13122 3320 13184 3336
rect 13196 3320 13202 3368
rect 13205 3360 13285 3368
rect 13205 3358 13224 3360
rect 13239 3358 13273 3360
rect 13205 3342 13285 3358
rect 13205 3320 13224 3342
rect 13239 3326 13269 3342
rect 13297 3336 13303 3410
rect 13306 3336 13325 3480
rect 13340 3336 13346 3480
rect 13355 3410 13368 3480
rect 13420 3476 13442 3480
rect 13413 3454 13442 3468
rect 13495 3454 13511 3468
rect 13549 3464 13555 3466
rect 13562 3464 13670 3480
rect 13677 3464 13683 3466
rect 13691 3464 13706 3480
rect 13772 3474 13791 3477
rect 13413 3452 13511 3454
rect 13538 3452 13706 3464
rect 13721 3454 13737 3468
rect 13772 3455 13794 3474
rect 13804 3468 13820 3469
rect 13803 3466 13820 3468
rect 13804 3461 13820 3466
rect 13794 3454 13800 3455
rect 13803 3454 13832 3461
rect 13721 3453 13832 3454
rect 13721 3452 13838 3453
rect 13397 3444 13448 3452
rect 13495 3444 13529 3452
rect 13397 3432 13422 3444
rect 13429 3432 13448 3444
rect 13502 3442 13529 3444
rect 13538 3442 13759 3452
rect 13794 3449 13800 3452
rect 13502 3438 13759 3442
rect 13397 3424 13448 3432
rect 13495 3424 13759 3438
rect 13803 3444 13838 3452
rect 13349 3376 13368 3410
rect 13413 3416 13442 3424
rect 13413 3410 13430 3416
rect 13413 3408 13447 3410
rect 13495 3408 13511 3424
rect 13512 3414 13720 3424
rect 13721 3414 13737 3424
rect 13785 3420 13800 3435
rect 13803 3432 13804 3444
rect 13811 3432 13838 3444
rect 13803 3424 13838 3432
rect 13803 3423 13832 3424
rect 13523 3410 13737 3414
rect 13538 3408 13737 3410
rect 13772 3410 13785 3420
rect 13803 3410 13820 3423
rect 13772 3408 13820 3410
rect 13414 3404 13447 3408
rect 13410 3402 13447 3404
rect 13410 3401 13477 3402
rect 13410 3396 13441 3401
rect 13447 3396 13477 3401
rect 13410 3392 13477 3396
rect 13383 3389 13477 3392
rect 13383 3382 13432 3389
rect 13383 3376 13413 3382
rect 13432 3377 13437 3382
rect 13349 3360 13429 3376
rect 13441 3368 13477 3389
rect 13538 3384 13727 3408
rect 13772 3407 13819 3408
rect 13785 3402 13819 3407
rect 13553 3381 13727 3384
rect 13546 3378 13727 3381
rect 13755 3401 13819 3402
rect 13349 3358 13368 3360
rect 13383 3358 13417 3360
rect 13349 3342 13429 3358
rect 13349 3336 13368 3342
rect 13065 3310 13168 3320
rect 13019 3308 13168 3310
rect 13189 3308 13224 3320
rect 12858 3306 13020 3308
rect 12870 3286 12889 3306
rect 12904 3304 12934 3306
rect 12753 3278 12794 3286
rect 12876 3282 12889 3286
rect 12941 3290 13020 3306
rect 13052 3306 13224 3308
rect 13052 3290 13131 3306
rect 13138 3304 13168 3306
rect 12716 3268 12745 3278
rect 12759 3268 12788 3278
rect 12803 3268 12833 3282
rect 12876 3268 12919 3282
rect 12941 3278 13131 3290
rect 13196 3286 13202 3306
rect 12926 3268 12956 3278
rect 12957 3268 13115 3278
rect 13119 3268 13149 3278
rect 13153 3268 13183 3282
rect 13211 3268 13224 3306
rect 13296 3320 13325 3336
rect 13339 3320 13368 3336
rect 13383 3326 13413 3342
rect 13441 3320 13447 3368
rect 13450 3362 13469 3368
rect 13484 3362 13514 3370
rect 13450 3354 13514 3362
rect 13450 3338 13530 3354
rect 13546 3347 13608 3378
rect 13624 3347 13686 3378
rect 13755 3376 13804 3401
rect 13819 3376 13849 3392
rect 13718 3362 13748 3370
rect 13755 3368 13865 3376
rect 13718 3354 13763 3362
rect 13450 3336 13469 3338
rect 13484 3336 13530 3338
rect 13450 3320 13530 3336
rect 13557 3334 13592 3347
rect 13633 3344 13670 3347
rect 13633 3342 13675 3344
rect 13562 3331 13592 3334
rect 13571 3327 13578 3331
rect 13578 3326 13579 3327
rect 13537 3320 13547 3326
rect 13296 3312 13331 3320
rect 13296 3286 13297 3312
rect 13304 3286 13331 3312
rect 13239 3268 13269 3282
rect 13296 3278 13331 3286
rect 13333 3312 13374 3320
rect 13333 3286 13348 3312
rect 13355 3286 13374 3312
rect 13438 3308 13469 3320
rect 13484 3308 13587 3320
rect 13599 3310 13625 3336
rect 13640 3331 13670 3342
rect 13702 3338 13764 3354
rect 13702 3336 13748 3338
rect 13702 3320 13764 3336
rect 13776 3320 13782 3368
rect 13785 3360 13865 3368
rect 13785 3358 13804 3360
rect 13819 3358 13853 3360
rect 13785 3342 13865 3358
rect 13785 3320 13804 3342
rect 13819 3326 13849 3342
rect 13877 3336 13883 3410
rect 13886 3336 13905 3480
rect 13920 3336 13926 3480
rect 13935 3410 13948 3480
rect 14000 3476 14022 3480
rect 13993 3454 14022 3468
rect 14075 3454 14091 3468
rect 14129 3464 14135 3466
rect 14142 3464 14250 3480
rect 14257 3464 14263 3466
rect 14271 3464 14286 3480
rect 14352 3474 14371 3477
rect 13993 3452 14091 3454
rect 14118 3452 14286 3464
rect 14301 3454 14317 3468
rect 14352 3455 14374 3474
rect 14384 3468 14400 3469
rect 14383 3466 14400 3468
rect 14384 3461 14400 3466
rect 14374 3454 14380 3455
rect 14383 3454 14412 3461
rect 14301 3453 14412 3454
rect 14301 3452 14418 3453
rect 13977 3444 14028 3452
rect 14075 3444 14109 3452
rect 13977 3432 14002 3444
rect 14009 3432 14028 3444
rect 14082 3442 14109 3444
rect 14118 3442 14339 3452
rect 14374 3449 14380 3452
rect 14082 3438 14339 3442
rect 13977 3424 14028 3432
rect 14075 3424 14339 3438
rect 14383 3444 14418 3452
rect 13929 3376 13948 3410
rect 13993 3416 14022 3424
rect 13993 3410 14010 3416
rect 13993 3408 14027 3410
rect 14075 3408 14091 3424
rect 14092 3414 14300 3424
rect 14301 3414 14317 3424
rect 14365 3420 14380 3435
rect 14383 3432 14384 3444
rect 14391 3432 14418 3444
rect 14383 3424 14418 3432
rect 14383 3423 14412 3424
rect 14103 3410 14317 3414
rect 14118 3408 14317 3410
rect 14352 3410 14365 3420
rect 14383 3410 14400 3423
rect 14352 3408 14400 3410
rect 13994 3404 14027 3408
rect 13990 3402 14027 3404
rect 13990 3401 14057 3402
rect 13990 3396 14021 3401
rect 14027 3396 14057 3401
rect 13990 3392 14057 3396
rect 13963 3389 14057 3392
rect 13963 3382 14012 3389
rect 13963 3376 13993 3382
rect 14012 3377 14017 3382
rect 13929 3360 14009 3376
rect 14021 3368 14057 3389
rect 14118 3384 14307 3408
rect 14352 3407 14399 3408
rect 14365 3402 14399 3407
rect 14133 3381 14307 3384
rect 14126 3378 14307 3381
rect 14335 3401 14399 3402
rect 13929 3358 13948 3360
rect 13963 3358 13997 3360
rect 13929 3342 14009 3358
rect 13929 3336 13948 3342
rect 13645 3310 13748 3320
rect 13599 3308 13748 3310
rect 13769 3308 13804 3320
rect 13438 3306 13600 3308
rect 13450 3286 13469 3306
rect 13484 3304 13514 3306
rect 13333 3278 13374 3286
rect 13456 3282 13469 3286
rect 13521 3290 13600 3306
rect 13632 3306 13804 3308
rect 13632 3290 13711 3306
rect 13718 3304 13748 3306
rect 13296 3268 13325 3278
rect 13339 3268 13368 3278
rect 13383 3268 13413 3282
rect 13456 3268 13499 3282
rect 13521 3278 13711 3290
rect 13776 3286 13782 3306
rect 13506 3268 13536 3278
rect 13537 3268 13695 3278
rect 13699 3268 13729 3278
rect 13733 3268 13763 3282
rect 13791 3268 13804 3306
rect 13876 3320 13905 3336
rect 13919 3320 13948 3336
rect 13963 3326 13993 3342
rect 14021 3320 14027 3368
rect 14030 3362 14049 3368
rect 14064 3362 14094 3370
rect 14030 3354 14094 3362
rect 14030 3338 14110 3354
rect 14126 3347 14188 3378
rect 14204 3347 14266 3378
rect 14335 3376 14384 3401
rect 14399 3376 14429 3392
rect 14298 3362 14328 3370
rect 14335 3368 14445 3376
rect 14298 3354 14343 3362
rect 14030 3336 14049 3338
rect 14064 3336 14110 3338
rect 14030 3320 14110 3336
rect 14137 3334 14172 3347
rect 14213 3344 14250 3347
rect 14213 3342 14255 3344
rect 14142 3331 14172 3334
rect 14151 3327 14158 3331
rect 14158 3326 14159 3327
rect 14117 3320 14127 3326
rect 13876 3312 13911 3320
rect 13876 3286 13877 3312
rect 13884 3286 13911 3312
rect 13819 3268 13849 3282
rect 13876 3278 13911 3286
rect 13913 3312 13954 3320
rect 13913 3286 13928 3312
rect 13935 3286 13954 3312
rect 14018 3308 14049 3320
rect 14064 3308 14167 3320
rect 14179 3310 14205 3336
rect 14220 3331 14250 3342
rect 14282 3338 14344 3354
rect 14282 3336 14328 3338
rect 14282 3320 14344 3336
rect 14356 3320 14362 3368
rect 14365 3360 14445 3368
rect 14365 3358 14384 3360
rect 14399 3358 14433 3360
rect 14365 3342 14445 3358
rect 14365 3320 14384 3342
rect 14399 3326 14429 3342
rect 14457 3336 14463 3410
rect 14466 3336 14485 3480
rect 14500 3336 14506 3480
rect 14515 3410 14528 3480
rect 14580 3476 14602 3480
rect 14573 3454 14602 3468
rect 14655 3454 14671 3468
rect 14709 3464 14715 3466
rect 14722 3464 14830 3480
rect 14837 3464 14843 3466
rect 14851 3464 14866 3480
rect 14932 3474 14951 3477
rect 14573 3452 14671 3454
rect 14698 3452 14866 3464
rect 14881 3454 14897 3468
rect 14932 3455 14954 3474
rect 14964 3468 14980 3469
rect 14963 3466 14980 3468
rect 14964 3461 14980 3466
rect 14954 3454 14960 3455
rect 14963 3454 14992 3461
rect 14881 3453 14992 3454
rect 14881 3452 14998 3453
rect 14557 3444 14608 3452
rect 14655 3444 14689 3452
rect 14557 3432 14582 3444
rect 14589 3432 14608 3444
rect 14662 3442 14689 3444
rect 14698 3442 14919 3452
rect 14954 3449 14960 3452
rect 14662 3438 14919 3442
rect 14557 3424 14608 3432
rect 14655 3424 14919 3438
rect 14963 3444 14998 3452
rect 14509 3376 14528 3410
rect 14573 3416 14602 3424
rect 14573 3410 14590 3416
rect 14573 3408 14607 3410
rect 14655 3408 14671 3424
rect 14672 3414 14880 3424
rect 14881 3414 14897 3424
rect 14945 3420 14960 3435
rect 14963 3432 14964 3444
rect 14971 3432 14998 3444
rect 14963 3424 14998 3432
rect 14963 3423 14992 3424
rect 14683 3410 14897 3414
rect 14698 3408 14897 3410
rect 14932 3410 14945 3420
rect 14963 3410 14980 3423
rect 14932 3408 14980 3410
rect 14574 3404 14607 3408
rect 14570 3402 14607 3404
rect 14570 3401 14637 3402
rect 14570 3396 14601 3401
rect 14607 3396 14637 3401
rect 14570 3392 14637 3396
rect 14543 3389 14637 3392
rect 14543 3382 14592 3389
rect 14543 3376 14573 3382
rect 14592 3377 14597 3382
rect 14509 3360 14589 3376
rect 14601 3368 14637 3389
rect 14698 3384 14887 3408
rect 14932 3407 14979 3408
rect 14945 3402 14979 3407
rect 14713 3381 14887 3384
rect 14706 3378 14887 3381
rect 14915 3401 14979 3402
rect 14509 3358 14528 3360
rect 14543 3358 14577 3360
rect 14509 3342 14589 3358
rect 14509 3336 14528 3342
rect 14225 3310 14328 3320
rect 14179 3308 14328 3310
rect 14349 3308 14384 3320
rect 14018 3306 14180 3308
rect 14030 3286 14049 3306
rect 14064 3304 14094 3306
rect 13913 3278 13954 3286
rect 14036 3282 14049 3286
rect 14101 3290 14180 3306
rect 14212 3306 14384 3308
rect 14212 3290 14291 3306
rect 14298 3304 14328 3306
rect 13876 3268 13905 3278
rect 13919 3268 13948 3278
rect 13963 3268 13993 3282
rect 14036 3268 14079 3282
rect 14101 3278 14291 3290
rect 14356 3286 14362 3306
rect 14086 3268 14116 3278
rect 14117 3268 14275 3278
rect 14279 3268 14309 3278
rect 14313 3268 14343 3282
rect 14371 3268 14384 3306
rect 14456 3320 14485 3336
rect 14499 3320 14528 3336
rect 14543 3326 14573 3342
rect 14601 3320 14607 3368
rect 14610 3362 14629 3368
rect 14644 3362 14674 3370
rect 14610 3354 14674 3362
rect 14610 3338 14690 3354
rect 14706 3347 14768 3378
rect 14784 3347 14846 3378
rect 14915 3376 14964 3401
rect 14979 3376 15009 3392
rect 14878 3362 14908 3370
rect 14915 3368 15025 3376
rect 14878 3354 14923 3362
rect 14610 3336 14629 3338
rect 14644 3336 14690 3338
rect 14610 3320 14690 3336
rect 14717 3334 14752 3347
rect 14793 3344 14830 3347
rect 14793 3342 14835 3344
rect 14722 3331 14752 3334
rect 14731 3327 14738 3331
rect 14738 3326 14739 3327
rect 14697 3320 14707 3326
rect 14456 3312 14491 3320
rect 14456 3286 14457 3312
rect 14464 3286 14491 3312
rect 14399 3268 14429 3282
rect 14456 3278 14491 3286
rect 14493 3312 14534 3320
rect 14493 3286 14508 3312
rect 14515 3286 14534 3312
rect 14598 3308 14629 3320
rect 14644 3308 14747 3320
rect 14759 3310 14785 3336
rect 14800 3331 14830 3342
rect 14862 3338 14924 3354
rect 14862 3336 14908 3338
rect 14862 3320 14924 3336
rect 14936 3320 14942 3368
rect 14945 3360 15025 3368
rect 14945 3358 14964 3360
rect 14979 3358 15013 3360
rect 14945 3342 15025 3358
rect 14945 3320 14964 3342
rect 14979 3326 15009 3342
rect 15037 3336 15043 3410
rect 15046 3336 15065 3480
rect 15080 3336 15086 3480
rect 15095 3410 15108 3480
rect 15160 3476 15182 3480
rect 15153 3454 15182 3468
rect 15235 3454 15251 3468
rect 15289 3464 15295 3466
rect 15302 3464 15410 3480
rect 15417 3464 15423 3466
rect 15431 3464 15446 3480
rect 15512 3474 15531 3477
rect 15153 3452 15251 3454
rect 15278 3452 15446 3464
rect 15461 3454 15477 3468
rect 15512 3455 15534 3474
rect 15544 3468 15560 3469
rect 15543 3466 15560 3468
rect 15544 3461 15560 3466
rect 15534 3454 15540 3455
rect 15543 3454 15572 3461
rect 15461 3453 15572 3454
rect 15461 3452 15578 3453
rect 15137 3444 15188 3452
rect 15235 3444 15269 3452
rect 15137 3432 15162 3444
rect 15169 3432 15188 3444
rect 15242 3442 15269 3444
rect 15278 3442 15499 3452
rect 15534 3449 15540 3452
rect 15242 3438 15499 3442
rect 15137 3424 15188 3432
rect 15235 3424 15499 3438
rect 15543 3444 15578 3452
rect 15089 3376 15108 3410
rect 15153 3416 15182 3424
rect 15153 3410 15170 3416
rect 15153 3408 15187 3410
rect 15235 3408 15251 3424
rect 15252 3414 15460 3424
rect 15461 3414 15477 3424
rect 15525 3420 15540 3435
rect 15543 3432 15544 3444
rect 15551 3432 15578 3444
rect 15543 3424 15578 3432
rect 15543 3423 15572 3424
rect 15263 3410 15477 3414
rect 15278 3408 15477 3410
rect 15512 3410 15525 3420
rect 15543 3410 15560 3423
rect 15512 3408 15560 3410
rect 15154 3404 15187 3408
rect 15150 3402 15187 3404
rect 15150 3401 15217 3402
rect 15150 3396 15181 3401
rect 15187 3396 15217 3401
rect 15150 3392 15217 3396
rect 15123 3389 15217 3392
rect 15123 3382 15172 3389
rect 15123 3376 15153 3382
rect 15172 3377 15177 3382
rect 15089 3360 15169 3376
rect 15181 3368 15217 3389
rect 15278 3384 15467 3408
rect 15512 3407 15559 3408
rect 15525 3402 15559 3407
rect 15293 3381 15467 3384
rect 15286 3378 15467 3381
rect 15495 3401 15559 3402
rect 15089 3358 15108 3360
rect 15123 3358 15157 3360
rect 15089 3342 15169 3358
rect 15089 3336 15108 3342
rect 14805 3310 14908 3320
rect 14759 3308 14908 3310
rect 14929 3308 14964 3320
rect 14598 3306 14760 3308
rect 14610 3286 14629 3306
rect 14644 3304 14674 3306
rect 14493 3278 14534 3286
rect 14616 3282 14629 3286
rect 14681 3290 14760 3306
rect 14792 3306 14964 3308
rect 14792 3290 14871 3306
rect 14878 3304 14908 3306
rect 14456 3268 14485 3278
rect 14499 3268 14528 3278
rect 14543 3268 14573 3282
rect 14616 3268 14659 3282
rect 14681 3278 14871 3290
rect 14936 3286 14942 3306
rect 14666 3268 14696 3278
rect 14697 3268 14855 3278
rect 14859 3268 14889 3278
rect 14893 3268 14923 3282
rect 14951 3268 14964 3306
rect 15036 3320 15065 3336
rect 15079 3320 15108 3336
rect 15123 3326 15153 3342
rect 15181 3320 15187 3368
rect 15190 3362 15209 3368
rect 15224 3362 15254 3370
rect 15190 3354 15254 3362
rect 15190 3338 15270 3354
rect 15286 3347 15348 3378
rect 15364 3347 15426 3378
rect 15495 3376 15544 3401
rect 15559 3376 15589 3392
rect 15458 3362 15488 3370
rect 15495 3368 15605 3376
rect 15458 3354 15503 3362
rect 15190 3336 15209 3338
rect 15224 3336 15270 3338
rect 15190 3320 15270 3336
rect 15297 3334 15332 3347
rect 15373 3344 15410 3347
rect 15373 3342 15415 3344
rect 15302 3331 15332 3334
rect 15311 3327 15318 3331
rect 15318 3326 15319 3327
rect 15277 3320 15287 3326
rect 15036 3312 15071 3320
rect 15036 3286 15037 3312
rect 15044 3286 15071 3312
rect 14979 3268 15009 3282
rect 15036 3278 15071 3286
rect 15073 3312 15114 3320
rect 15073 3286 15088 3312
rect 15095 3286 15114 3312
rect 15178 3308 15209 3320
rect 15224 3308 15327 3320
rect 15339 3310 15365 3336
rect 15380 3331 15410 3342
rect 15442 3338 15504 3354
rect 15442 3336 15488 3338
rect 15442 3320 15504 3336
rect 15516 3320 15522 3368
rect 15525 3360 15605 3368
rect 15525 3358 15544 3360
rect 15559 3358 15593 3360
rect 15525 3342 15605 3358
rect 15525 3320 15544 3342
rect 15559 3326 15589 3342
rect 15617 3336 15623 3410
rect 15626 3336 15645 3480
rect 15660 3336 15666 3480
rect 15675 3410 15688 3480
rect 15740 3476 15762 3480
rect 15733 3454 15762 3468
rect 15815 3454 15831 3468
rect 15869 3464 15875 3466
rect 15882 3464 15990 3480
rect 15997 3464 16003 3466
rect 16011 3464 16026 3480
rect 16092 3474 16111 3477
rect 15733 3452 15831 3454
rect 15858 3452 16026 3464
rect 16041 3454 16057 3468
rect 16092 3455 16114 3474
rect 16124 3468 16140 3469
rect 16123 3466 16140 3468
rect 16124 3461 16140 3466
rect 16114 3454 16120 3455
rect 16123 3454 16152 3461
rect 16041 3453 16152 3454
rect 16041 3452 16158 3453
rect 15717 3444 15768 3452
rect 15815 3444 15849 3452
rect 15717 3432 15742 3444
rect 15749 3432 15768 3444
rect 15822 3442 15849 3444
rect 15858 3442 16079 3452
rect 16114 3449 16120 3452
rect 15822 3438 16079 3442
rect 15717 3424 15768 3432
rect 15815 3424 16079 3438
rect 16123 3444 16158 3452
rect 15669 3376 15688 3410
rect 15733 3416 15762 3424
rect 15733 3410 15750 3416
rect 15733 3408 15767 3410
rect 15815 3408 15831 3424
rect 15832 3414 16040 3424
rect 16041 3414 16057 3424
rect 16105 3420 16120 3435
rect 16123 3432 16124 3444
rect 16131 3432 16158 3444
rect 16123 3424 16158 3432
rect 16123 3423 16152 3424
rect 15843 3410 16057 3414
rect 15858 3408 16057 3410
rect 16092 3410 16105 3420
rect 16123 3410 16140 3423
rect 16092 3408 16140 3410
rect 15734 3404 15767 3408
rect 15730 3402 15767 3404
rect 15730 3401 15797 3402
rect 15730 3396 15761 3401
rect 15767 3396 15797 3401
rect 15730 3392 15797 3396
rect 15703 3389 15797 3392
rect 15703 3382 15752 3389
rect 15703 3376 15733 3382
rect 15752 3377 15757 3382
rect 15669 3360 15749 3376
rect 15761 3368 15797 3389
rect 15858 3384 16047 3408
rect 16092 3407 16139 3408
rect 16105 3402 16139 3407
rect 15873 3381 16047 3384
rect 15866 3378 16047 3381
rect 16075 3401 16139 3402
rect 15669 3358 15688 3360
rect 15703 3358 15737 3360
rect 15669 3342 15749 3358
rect 15669 3336 15688 3342
rect 15385 3310 15488 3320
rect 15339 3308 15488 3310
rect 15509 3308 15544 3320
rect 15178 3306 15340 3308
rect 15190 3286 15209 3306
rect 15224 3304 15254 3306
rect 15073 3278 15114 3286
rect 15196 3282 15209 3286
rect 15261 3290 15340 3306
rect 15372 3306 15544 3308
rect 15372 3290 15451 3306
rect 15458 3304 15488 3306
rect 15036 3268 15065 3278
rect 15079 3268 15108 3278
rect 15123 3268 15153 3282
rect 15196 3268 15239 3282
rect 15261 3278 15451 3290
rect 15516 3286 15522 3306
rect 15246 3268 15276 3278
rect 15277 3268 15435 3278
rect 15439 3268 15469 3278
rect 15473 3268 15503 3282
rect 15531 3268 15544 3306
rect 15616 3320 15645 3336
rect 15659 3320 15688 3336
rect 15703 3326 15733 3342
rect 15761 3320 15767 3368
rect 15770 3362 15789 3368
rect 15804 3362 15834 3370
rect 15770 3354 15834 3362
rect 15770 3338 15850 3354
rect 15866 3347 15928 3378
rect 15944 3347 16006 3378
rect 16075 3376 16124 3401
rect 16139 3376 16169 3392
rect 16038 3362 16068 3370
rect 16075 3368 16185 3376
rect 16038 3354 16083 3362
rect 15770 3336 15789 3338
rect 15804 3336 15850 3338
rect 15770 3320 15850 3336
rect 15877 3334 15912 3347
rect 15953 3344 15990 3347
rect 15953 3342 15995 3344
rect 15882 3331 15912 3334
rect 15891 3327 15898 3331
rect 15898 3326 15899 3327
rect 15857 3320 15867 3326
rect 15616 3312 15651 3320
rect 15616 3286 15617 3312
rect 15624 3286 15651 3312
rect 15559 3268 15589 3282
rect 15616 3278 15651 3286
rect 15653 3312 15694 3320
rect 15653 3286 15668 3312
rect 15675 3286 15694 3312
rect 15758 3308 15789 3320
rect 15804 3308 15907 3320
rect 15919 3310 15945 3336
rect 15960 3331 15990 3342
rect 16022 3338 16084 3354
rect 16022 3336 16068 3338
rect 16022 3320 16084 3336
rect 16096 3320 16102 3368
rect 16105 3360 16185 3368
rect 16105 3358 16124 3360
rect 16139 3358 16173 3360
rect 16105 3342 16185 3358
rect 16105 3320 16124 3342
rect 16139 3326 16169 3342
rect 16197 3336 16203 3410
rect 16206 3336 16225 3480
rect 16240 3336 16246 3480
rect 16255 3410 16268 3480
rect 16320 3476 16342 3480
rect 16313 3454 16342 3468
rect 16395 3454 16411 3468
rect 16449 3464 16455 3466
rect 16462 3464 16570 3480
rect 16577 3464 16583 3466
rect 16591 3464 16606 3480
rect 16672 3474 16691 3477
rect 16313 3452 16411 3454
rect 16438 3452 16606 3464
rect 16621 3454 16637 3468
rect 16672 3455 16694 3474
rect 16704 3468 16720 3469
rect 16703 3466 16720 3468
rect 16704 3461 16720 3466
rect 16694 3454 16700 3455
rect 16703 3454 16732 3461
rect 16621 3453 16732 3454
rect 16621 3452 16738 3453
rect 16297 3444 16348 3452
rect 16395 3444 16429 3452
rect 16297 3432 16322 3444
rect 16329 3432 16348 3444
rect 16402 3442 16429 3444
rect 16438 3442 16659 3452
rect 16694 3449 16700 3452
rect 16402 3438 16659 3442
rect 16297 3424 16348 3432
rect 16395 3424 16659 3438
rect 16703 3444 16738 3452
rect 16249 3376 16268 3410
rect 16313 3416 16342 3424
rect 16313 3410 16330 3416
rect 16313 3408 16347 3410
rect 16395 3408 16411 3424
rect 16412 3414 16620 3424
rect 16621 3414 16637 3424
rect 16685 3420 16700 3435
rect 16703 3432 16704 3444
rect 16711 3432 16738 3444
rect 16703 3424 16738 3432
rect 16703 3423 16732 3424
rect 16423 3410 16637 3414
rect 16438 3408 16637 3410
rect 16672 3410 16685 3420
rect 16703 3410 16720 3423
rect 16672 3408 16720 3410
rect 16314 3404 16347 3408
rect 16310 3402 16347 3404
rect 16310 3401 16377 3402
rect 16310 3396 16341 3401
rect 16347 3396 16377 3401
rect 16310 3392 16377 3396
rect 16283 3389 16377 3392
rect 16283 3382 16332 3389
rect 16283 3376 16313 3382
rect 16332 3377 16337 3382
rect 16249 3360 16329 3376
rect 16341 3368 16377 3389
rect 16438 3384 16627 3408
rect 16672 3407 16719 3408
rect 16685 3402 16719 3407
rect 16453 3381 16627 3384
rect 16446 3378 16627 3381
rect 16655 3401 16719 3402
rect 16249 3358 16268 3360
rect 16283 3358 16317 3360
rect 16249 3342 16329 3358
rect 16249 3336 16268 3342
rect 15965 3310 16068 3320
rect 15919 3308 16068 3310
rect 16089 3308 16124 3320
rect 15758 3306 15920 3308
rect 15770 3286 15789 3306
rect 15804 3304 15834 3306
rect 15653 3278 15694 3286
rect 15776 3282 15789 3286
rect 15841 3290 15920 3306
rect 15952 3306 16124 3308
rect 15952 3290 16031 3306
rect 16038 3304 16068 3306
rect 15616 3268 15645 3278
rect 15659 3268 15688 3278
rect 15703 3268 15733 3282
rect 15776 3268 15819 3282
rect 15841 3278 16031 3290
rect 16096 3286 16102 3306
rect 15826 3268 15856 3278
rect 15857 3268 16015 3278
rect 16019 3268 16049 3278
rect 16053 3268 16083 3282
rect 16111 3268 16124 3306
rect 16196 3320 16225 3336
rect 16239 3320 16268 3336
rect 16283 3326 16313 3342
rect 16341 3320 16347 3368
rect 16350 3362 16369 3368
rect 16384 3362 16414 3370
rect 16350 3354 16414 3362
rect 16350 3338 16430 3354
rect 16446 3347 16508 3378
rect 16524 3347 16586 3378
rect 16655 3376 16704 3401
rect 16719 3376 16749 3392
rect 16618 3362 16648 3370
rect 16655 3368 16765 3376
rect 16618 3354 16663 3362
rect 16350 3336 16369 3338
rect 16384 3336 16430 3338
rect 16350 3320 16430 3336
rect 16457 3334 16492 3347
rect 16533 3344 16570 3347
rect 16533 3342 16575 3344
rect 16462 3331 16492 3334
rect 16471 3327 16478 3331
rect 16478 3326 16479 3327
rect 16437 3320 16447 3326
rect 16196 3312 16231 3320
rect 16196 3286 16197 3312
rect 16204 3286 16231 3312
rect 16139 3268 16169 3282
rect 16196 3278 16231 3286
rect 16233 3312 16274 3320
rect 16233 3286 16248 3312
rect 16255 3286 16274 3312
rect 16338 3308 16369 3320
rect 16384 3308 16487 3320
rect 16499 3310 16525 3336
rect 16540 3331 16570 3342
rect 16602 3338 16664 3354
rect 16602 3336 16648 3338
rect 16602 3320 16664 3336
rect 16676 3320 16682 3368
rect 16685 3360 16765 3368
rect 16685 3358 16704 3360
rect 16719 3358 16753 3360
rect 16685 3342 16765 3358
rect 16685 3320 16704 3342
rect 16719 3326 16749 3342
rect 16777 3336 16783 3410
rect 16786 3336 16805 3480
rect 16820 3336 16826 3480
rect 16835 3410 16848 3480
rect 16900 3476 16922 3480
rect 16893 3454 16922 3468
rect 16975 3454 16991 3468
rect 17029 3464 17035 3466
rect 17042 3464 17150 3480
rect 17157 3464 17163 3466
rect 17171 3464 17186 3480
rect 17252 3474 17271 3477
rect 16893 3452 16991 3454
rect 17018 3452 17186 3464
rect 17201 3454 17217 3468
rect 17252 3455 17274 3474
rect 17284 3468 17300 3469
rect 17283 3466 17300 3468
rect 17284 3461 17300 3466
rect 17274 3454 17280 3455
rect 17283 3454 17312 3461
rect 17201 3453 17312 3454
rect 17201 3452 17318 3453
rect 16877 3444 16928 3452
rect 16975 3444 17009 3452
rect 16877 3432 16902 3444
rect 16909 3432 16928 3444
rect 16982 3442 17009 3444
rect 17018 3442 17239 3452
rect 17274 3449 17280 3452
rect 16982 3438 17239 3442
rect 16877 3424 16928 3432
rect 16975 3424 17239 3438
rect 17283 3444 17318 3452
rect 16829 3376 16848 3410
rect 16893 3416 16922 3424
rect 16893 3410 16910 3416
rect 16893 3408 16927 3410
rect 16975 3408 16991 3424
rect 16992 3414 17200 3424
rect 17201 3414 17217 3424
rect 17265 3420 17280 3435
rect 17283 3432 17284 3444
rect 17291 3432 17318 3444
rect 17283 3424 17318 3432
rect 17283 3423 17312 3424
rect 17003 3410 17217 3414
rect 17018 3408 17217 3410
rect 17252 3410 17265 3420
rect 17283 3410 17300 3423
rect 17252 3408 17300 3410
rect 16894 3404 16927 3408
rect 16890 3402 16927 3404
rect 16890 3401 16957 3402
rect 16890 3396 16921 3401
rect 16927 3396 16957 3401
rect 16890 3392 16957 3396
rect 16863 3389 16957 3392
rect 16863 3382 16912 3389
rect 16863 3376 16893 3382
rect 16912 3377 16917 3382
rect 16829 3360 16909 3376
rect 16921 3368 16957 3389
rect 17018 3384 17207 3408
rect 17252 3407 17299 3408
rect 17265 3402 17299 3407
rect 17033 3381 17207 3384
rect 17026 3378 17207 3381
rect 17235 3401 17299 3402
rect 16829 3358 16848 3360
rect 16863 3358 16897 3360
rect 16829 3342 16909 3358
rect 16829 3336 16848 3342
rect 16545 3310 16648 3320
rect 16499 3308 16648 3310
rect 16669 3308 16704 3320
rect 16338 3306 16500 3308
rect 16350 3286 16369 3306
rect 16384 3304 16414 3306
rect 16233 3278 16274 3286
rect 16356 3282 16369 3286
rect 16421 3290 16500 3306
rect 16532 3306 16704 3308
rect 16532 3290 16611 3306
rect 16618 3304 16648 3306
rect 16196 3268 16225 3278
rect 16239 3268 16268 3278
rect 16283 3268 16313 3282
rect 16356 3268 16399 3282
rect 16421 3278 16611 3290
rect 16676 3286 16682 3306
rect 16406 3268 16436 3278
rect 16437 3268 16595 3278
rect 16599 3268 16629 3278
rect 16633 3268 16663 3282
rect 16691 3268 16704 3306
rect 16776 3320 16805 3336
rect 16819 3320 16848 3336
rect 16863 3326 16893 3342
rect 16921 3320 16927 3368
rect 16930 3362 16949 3368
rect 16964 3362 16994 3370
rect 16930 3354 16994 3362
rect 16930 3338 17010 3354
rect 17026 3347 17088 3378
rect 17104 3347 17166 3378
rect 17235 3376 17284 3401
rect 17299 3376 17329 3392
rect 17198 3362 17228 3370
rect 17235 3368 17345 3376
rect 17198 3354 17243 3362
rect 16930 3336 16949 3338
rect 16964 3336 17010 3338
rect 16930 3320 17010 3336
rect 17037 3334 17072 3347
rect 17113 3344 17150 3347
rect 17113 3342 17155 3344
rect 17042 3331 17072 3334
rect 17051 3327 17058 3331
rect 17058 3326 17059 3327
rect 17017 3320 17027 3326
rect 16776 3312 16811 3320
rect 16776 3286 16777 3312
rect 16784 3286 16811 3312
rect 16719 3268 16749 3282
rect 16776 3278 16811 3286
rect 16813 3312 16854 3320
rect 16813 3286 16828 3312
rect 16835 3286 16854 3312
rect 16918 3308 16949 3320
rect 16964 3308 17067 3320
rect 17079 3310 17105 3336
rect 17120 3331 17150 3342
rect 17182 3338 17244 3354
rect 17182 3336 17228 3338
rect 17182 3320 17244 3336
rect 17256 3320 17262 3368
rect 17265 3360 17345 3368
rect 17265 3358 17284 3360
rect 17299 3358 17333 3360
rect 17265 3342 17345 3358
rect 17265 3320 17284 3342
rect 17299 3326 17329 3342
rect 17357 3336 17363 3410
rect 17366 3336 17385 3480
rect 17400 3336 17406 3480
rect 17415 3410 17428 3480
rect 17480 3476 17502 3480
rect 17473 3454 17502 3468
rect 17555 3454 17571 3468
rect 17609 3464 17615 3466
rect 17622 3464 17730 3480
rect 17737 3464 17743 3466
rect 17751 3464 17766 3480
rect 17832 3474 17851 3477
rect 17473 3452 17571 3454
rect 17598 3452 17766 3464
rect 17781 3454 17797 3468
rect 17832 3455 17854 3474
rect 17864 3468 17880 3469
rect 17863 3466 17880 3468
rect 17864 3461 17880 3466
rect 17854 3454 17860 3455
rect 17863 3454 17892 3461
rect 17781 3453 17892 3454
rect 17781 3452 17898 3453
rect 17457 3444 17508 3452
rect 17555 3444 17589 3452
rect 17457 3432 17482 3444
rect 17489 3432 17508 3444
rect 17562 3442 17589 3444
rect 17598 3442 17819 3452
rect 17854 3449 17860 3452
rect 17562 3438 17819 3442
rect 17457 3424 17508 3432
rect 17555 3424 17819 3438
rect 17863 3444 17898 3452
rect 17409 3376 17428 3410
rect 17473 3416 17502 3424
rect 17473 3410 17490 3416
rect 17473 3408 17507 3410
rect 17555 3408 17571 3424
rect 17572 3414 17780 3424
rect 17781 3414 17797 3424
rect 17845 3420 17860 3435
rect 17863 3432 17864 3444
rect 17871 3432 17898 3444
rect 17863 3424 17898 3432
rect 17863 3423 17892 3424
rect 17583 3410 17797 3414
rect 17598 3408 17797 3410
rect 17832 3410 17845 3420
rect 17863 3410 17880 3423
rect 17832 3408 17880 3410
rect 17474 3404 17507 3408
rect 17470 3402 17507 3404
rect 17470 3401 17537 3402
rect 17470 3396 17501 3401
rect 17507 3396 17537 3401
rect 17470 3392 17537 3396
rect 17443 3389 17537 3392
rect 17443 3382 17492 3389
rect 17443 3376 17473 3382
rect 17492 3377 17497 3382
rect 17409 3360 17489 3376
rect 17501 3368 17537 3389
rect 17598 3384 17787 3408
rect 17832 3407 17879 3408
rect 17845 3402 17879 3407
rect 17613 3381 17787 3384
rect 17606 3378 17787 3381
rect 17815 3401 17879 3402
rect 17409 3358 17428 3360
rect 17443 3358 17477 3360
rect 17409 3342 17489 3358
rect 17409 3336 17428 3342
rect 17125 3310 17228 3320
rect 17079 3308 17228 3310
rect 17249 3308 17284 3320
rect 16918 3306 17080 3308
rect 16930 3286 16949 3306
rect 16964 3304 16994 3306
rect 16813 3278 16854 3286
rect 16936 3282 16949 3286
rect 17001 3290 17080 3306
rect 17112 3306 17284 3308
rect 17112 3290 17191 3306
rect 17198 3304 17228 3306
rect 16776 3268 16805 3278
rect 16819 3268 16848 3278
rect 16863 3268 16893 3282
rect 16936 3268 16979 3282
rect 17001 3278 17191 3290
rect 17256 3286 17262 3306
rect 16986 3268 17016 3278
rect 17017 3268 17175 3278
rect 17179 3268 17209 3278
rect 17213 3268 17243 3282
rect 17271 3268 17284 3306
rect 17356 3320 17385 3336
rect 17399 3320 17428 3336
rect 17443 3326 17473 3342
rect 17501 3320 17507 3368
rect 17510 3362 17529 3368
rect 17544 3362 17574 3370
rect 17510 3354 17574 3362
rect 17510 3338 17590 3354
rect 17606 3347 17668 3378
rect 17684 3347 17746 3378
rect 17815 3376 17864 3401
rect 17879 3376 17909 3392
rect 17778 3362 17808 3370
rect 17815 3368 17925 3376
rect 17778 3354 17823 3362
rect 17510 3336 17529 3338
rect 17544 3336 17590 3338
rect 17510 3320 17590 3336
rect 17617 3334 17652 3347
rect 17693 3344 17730 3347
rect 17693 3342 17735 3344
rect 17622 3331 17652 3334
rect 17631 3327 17638 3331
rect 17638 3326 17639 3327
rect 17597 3320 17607 3326
rect 17356 3312 17391 3320
rect 17356 3286 17357 3312
rect 17364 3286 17391 3312
rect 17299 3268 17329 3282
rect 17356 3278 17391 3286
rect 17393 3312 17434 3320
rect 17393 3286 17408 3312
rect 17415 3286 17434 3312
rect 17498 3308 17529 3320
rect 17544 3308 17647 3320
rect 17659 3310 17685 3336
rect 17700 3331 17730 3342
rect 17762 3338 17824 3354
rect 17762 3336 17808 3338
rect 17762 3320 17824 3336
rect 17836 3320 17842 3368
rect 17845 3360 17925 3368
rect 17845 3358 17864 3360
rect 17879 3358 17913 3360
rect 17845 3342 17925 3358
rect 17845 3320 17864 3342
rect 17879 3326 17909 3342
rect 17937 3336 17943 3410
rect 17946 3336 17965 3480
rect 17980 3336 17986 3480
rect 17995 3410 18008 3480
rect 18060 3476 18082 3480
rect 18053 3454 18082 3468
rect 18135 3454 18151 3468
rect 18189 3464 18195 3466
rect 18202 3464 18310 3480
rect 18317 3464 18323 3466
rect 18331 3464 18346 3480
rect 18412 3474 18431 3477
rect 18053 3452 18151 3454
rect 18178 3452 18346 3464
rect 18361 3454 18377 3468
rect 18412 3455 18434 3474
rect 18444 3468 18460 3469
rect 18443 3466 18460 3468
rect 18444 3461 18460 3466
rect 18434 3454 18440 3455
rect 18443 3454 18472 3461
rect 18361 3453 18472 3454
rect 18361 3452 18478 3453
rect 18037 3444 18088 3452
rect 18135 3444 18169 3452
rect 18037 3432 18062 3444
rect 18069 3432 18088 3444
rect 18142 3442 18169 3444
rect 18178 3442 18399 3452
rect 18434 3449 18440 3452
rect 18142 3438 18399 3442
rect 18037 3424 18088 3432
rect 18135 3424 18399 3438
rect 18443 3444 18478 3452
rect 17989 3376 18008 3410
rect 18053 3416 18082 3424
rect 18053 3410 18070 3416
rect 18053 3408 18087 3410
rect 18135 3408 18151 3424
rect 18152 3414 18360 3424
rect 18361 3414 18377 3424
rect 18425 3420 18440 3435
rect 18443 3432 18444 3444
rect 18451 3432 18478 3444
rect 18443 3424 18478 3432
rect 18443 3423 18472 3424
rect 18163 3410 18377 3414
rect 18178 3408 18377 3410
rect 18412 3410 18425 3420
rect 18443 3410 18460 3423
rect 18412 3408 18460 3410
rect 18054 3404 18087 3408
rect 18050 3402 18087 3404
rect 18050 3401 18117 3402
rect 18050 3396 18081 3401
rect 18087 3396 18117 3401
rect 18050 3392 18117 3396
rect 18023 3389 18117 3392
rect 18023 3382 18072 3389
rect 18023 3376 18053 3382
rect 18072 3377 18077 3382
rect 17989 3360 18069 3376
rect 18081 3368 18117 3389
rect 18178 3384 18367 3408
rect 18412 3407 18459 3408
rect 18425 3402 18459 3407
rect 18193 3381 18367 3384
rect 18186 3378 18367 3381
rect 18395 3401 18459 3402
rect 17989 3358 18008 3360
rect 18023 3358 18057 3360
rect 17989 3342 18069 3358
rect 17989 3336 18008 3342
rect 17705 3310 17808 3320
rect 17659 3308 17808 3310
rect 17829 3308 17864 3320
rect 17498 3306 17660 3308
rect 17510 3286 17529 3306
rect 17544 3304 17574 3306
rect 17393 3278 17434 3286
rect 17516 3282 17529 3286
rect 17581 3290 17660 3306
rect 17692 3306 17864 3308
rect 17692 3290 17771 3306
rect 17778 3304 17808 3306
rect 17356 3268 17385 3278
rect 17399 3268 17428 3278
rect 17443 3268 17473 3282
rect 17516 3268 17559 3282
rect 17581 3278 17771 3290
rect 17836 3286 17842 3306
rect 17566 3268 17596 3278
rect 17597 3268 17755 3278
rect 17759 3268 17789 3278
rect 17793 3268 17823 3282
rect 17851 3268 17864 3306
rect 17936 3320 17965 3336
rect 17979 3320 18008 3336
rect 18023 3326 18053 3342
rect 18081 3320 18087 3368
rect 18090 3362 18109 3368
rect 18124 3362 18154 3370
rect 18090 3354 18154 3362
rect 18090 3338 18170 3354
rect 18186 3347 18248 3378
rect 18264 3347 18326 3378
rect 18395 3376 18444 3401
rect 18459 3376 18489 3392
rect 18358 3362 18388 3370
rect 18395 3368 18505 3376
rect 18358 3354 18403 3362
rect 18090 3336 18109 3338
rect 18124 3336 18170 3338
rect 18090 3320 18170 3336
rect 18197 3334 18232 3347
rect 18273 3344 18310 3347
rect 18273 3342 18315 3344
rect 18202 3331 18232 3334
rect 18211 3327 18218 3331
rect 18218 3326 18219 3327
rect 18177 3320 18187 3326
rect 17936 3312 17971 3320
rect 17936 3286 17937 3312
rect 17944 3286 17971 3312
rect 17879 3268 17909 3282
rect 17936 3278 17971 3286
rect 17973 3312 18014 3320
rect 17973 3286 17988 3312
rect 17995 3286 18014 3312
rect 18078 3308 18109 3320
rect 18124 3308 18227 3320
rect 18239 3310 18265 3336
rect 18280 3331 18310 3342
rect 18342 3338 18404 3354
rect 18342 3336 18388 3338
rect 18342 3320 18404 3336
rect 18416 3320 18422 3368
rect 18425 3360 18505 3368
rect 18425 3358 18444 3360
rect 18459 3358 18493 3360
rect 18425 3342 18505 3358
rect 18425 3320 18444 3342
rect 18459 3326 18489 3342
rect 18517 3336 18523 3410
rect 18532 3336 18545 3480
rect 18285 3310 18388 3320
rect 18239 3308 18388 3310
rect 18409 3308 18444 3320
rect 18078 3306 18240 3308
rect 18090 3286 18109 3306
rect 18124 3304 18154 3306
rect 17973 3278 18014 3286
rect 18096 3282 18109 3286
rect 18161 3290 18240 3306
rect 18272 3306 18444 3308
rect 18272 3290 18351 3306
rect 18358 3304 18388 3306
rect 17936 3268 17965 3278
rect 17979 3268 18008 3278
rect 18023 3268 18053 3282
rect 18096 3268 18139 3282
rect 18161 3278 18351 3290
rect 18416 3286 18422 3306
rect 18146 3268 18176 3278
rect 18177 3268 18335 3278
rect 18339 3268 18369 3278
rect 18373 3268 18403 3282
rect 18431 3268 18444 3306
rect 18516 3320 18545 3336
rect 18516 3312 18551 3320
rect 18516 3286 18517 3312
rect 18524 3286 18551 3312
rect 18459 3268 18489 3282
rect 18516 3278 18551 3286
rect 18516 3268 18545 3278
rect -1 3262 18545 3268
rect 0 3254 18545 3262
rect 15 3224 28 3254
rect 43 3240 73 3254
rect 116 3240 159 3254
rect 166 3240 386 3254
rect 393 3240 423 3254
rect 83 3226 98 3238
rect 117 3226 130 3240
rect 198 3236 351 3240
rect 80 3224 102 3226
rect 180 3224 372 3236
rect 451 3224 464 3254
rect 479 3240 509 3254
rect 546 3224 565 3254
rect 580 3224 586 3254
rect 595 3224 608 3254
rect 623 3240 653 3254
rect 696 3240 739 3254
rect 746 3240 966 3254
rect 973 3240 1003 3254
rect 663 3226 678 3238
rect 697 3226 710 3240
rect 778 3236 931 3240
rect 660 3224 682 3226
rect 760 3224 952 3236
rect 1031 3224 1044 3254
rect 1059 3240 1089 3254
rect 1126 3224 1145 3254
rect 1160 3224 1166 3254
rect 1175 3224 1188 3254
rect 1203 3240 1233 3254
rect 1276 3240 1319 3254
rect 1326 3240 1546 3254
rect 1553 3240 1583 3254
rect 1243 3226 1258 3238
rect 1277 3226 1290 3240
rect 1358 3236 1511 3240
rect 1240 3224 1262 3226
rect 1340 3224 1532 3236
rect 1611 3224 1624 3254
rect 1639 3240 1669 3254
rect 1706 3224 1725 3254
rect 1740 3224 1746 3254
rect 1755 3224 1768 3254
rect 1783 3240 1813 3254
rect 1856 3240 1899 3254
rect 1906 3240 2126 3254
rect 2133 3240 2163 3254
rect 1823 3226 1838 3238
rect 1857 3226 1870 3240
rect 1938 3236 2091 3240
rect 1820 3224 1842 3226
rect 1920 3224 2112 3236
rect 2191 3224 2204 3254
rect 2219 3240 2249 3254
rect 2286 3224 2305 3254
rect 2320 3224 2326 3254
rect 2335 3224 2348 3254
rect 2363 3240 2393 3254
rect 2436 3240 2479 3254
rect 2486 3240 2706 3254
rect 2713 3240 2743 3254
rect 2403 3226 2418 3238
rect 2437 3226 2450 3240
rect 2518 3236 2671 3240
rect 2400 3224 2422 3226
rect 2500 3224 2692 3236
rect 2771 3224 2784 3254
rect 2799 3240 2829 3254
rect 2866 3224 2885 3254
rect 2900 3224 2906 3254
rect 2915 3224 2928 3254
rect 2943 3240 2973 3254
rect 3016 3240 3059 3254
rect 3066 3240 3286 3254
rect 3293 3240 3323 3254
rect 2983 3226 2998 3238
rect 3017 3226 3030 3240
rect 3098 3236 3251 3240
rect 2980 3224 3002 3226
rect 3080 3224 3272 3236
rect 3351 3224 3364 3254
rect 3379 3240 3409 3254
rect 3446 3224 3465 3254
rect 3480 3224 3486 3254
rect 3495 3224 3508 3254
rect 3523 3240 3553 3254
rect 3596 3240 3639 3254
rect 3646 3240 3866 3254
rect 3873 3240 3903 3254
rect 3563 3226 3578 3238
rect 3597 3226 3610 3240
rect 3678 3236 3831 3240
rect 3560 3224 3582 3226
rect 3660 3224 3852 3236
rect 3931 3224 3944 3254
rect 3959 3240 3989 3254
rect 4026 3224 4045 3254
rect 4060 3224 4066 3254
rect 4075 3224 4088 3254
rect 4103 3240 4133 3254
rect 4176 3240 4219 3254
rect 4226 3240 4446 3254
rect 4453 3240 4483 3254
rect 4143 3226 4158 3238
rect 4177 3226 4190 3240
rect 4258 3236 4411 3240
rect 4140 3224 4162 3226
rect 4240 3224 4432 3236
rect 4511 3224 4524 3254
rect 4539 3240 4569 3254
rect 4606 3224 4625 3254
rect 4640 3224 4646 3254
rect 4655 3224 4668 3254
rect 4683 3240 4713 3254
rect 4756 3240 4799 3254
rect 4806 3240 5026 3254
rect 5033 3240 5063 3254
rect 4723 3226 4738 3238
rect 4757 3226 4770 3240
rect 4838 3236 4991 3240
rect 4720 3224 4742 3226
rect 4820 3224 5012 3236
rect 5091 3224 5104 3254
rect 5119 3240 5149 3254
rect 5186 3224 5205 3254
rect 5220 3224 5226 3254
rect 5235 3224 5248 3254
rect 5263 3240 5293 3254
rect 5336 3240 5379 3254
rect 5386 3240 5606 3254
rect 5613 3240 5643 3254
rect 5303 3226 5318 3238
rect 5337 3226 5350 3240
rect 5418 3236 5571 3240
rect 5300 3224 5322 3226
rect 5400 3224 5592 3236
rect 5671 3224 5684 3254
rect 5699 3240 5729 3254
rect 5766 3224 5785 3254
rect 5800 3224 5806 3254
rect 5815 3224 5828 3254
rect 5843 3240 5873 3254
rect 5916 3240 5959 3254
rect 5966 3240 6186 3254
rect 6193 3240 6223 3254
rect 5883 3226 5898 3238
rect 5917 3226 5930 3240
rect 5998 3236 6151 3240
rect 5880 3224 5902 3226
rect 5980 3224 6172 3236
rect 6251 3224 6264 3254
rect 6279 3240 6309 3254
rect 6346 3224 6365 3254
rect 6380 3224 6386 3254
rect 6395 3224 6408 3254
rect 6423 3240 6453 3254
rect 6496 3240 6539 3254
rect 6546 3240 6766 3254
rect 6773 3240 6803 3254
rect 6463 3226 6478 3238
rect 6497 3226 6510 3240
rect 6578 3236 6731 3240
rect 6460 3224 6482 3226
rect 6560 3224 6752 3236
rect 6831 3224 6844 3254
rect 6859 3240 6889 3254
rect 6926 3224 6945 3254
rect 6960 3224 6966 3254
rect 6975 3224 6988 3254
rect 7003 3240 7033 3254
rect 7076 3240 7119 3254
rect 7126 3240 7346 3254
rect 7353 3240 7383 3254
rect 7043 3226 7058 3238
rect 7077 3226 7090 3240
rect 7158 3236 7311 3240
rect 7040 3224 7062 3226
rect 7140 3224 7332 3236
rect 7411 3224 7424 3254
rect 7439 3240 7469 3254
rect 7506 3224 7525 3254
rect 7540 3224 7546 3254
rect 7555 3224 7568 3254
rect 7583 3240 7613 3254
rect 7656 3240 7699 3254
rect 7706 3240 7926 3254
rect 7933 3240 7963 3254
rect 7623 3226 7638 3238
rect 7657 3226 7670 3240
rect 7738 3236 7891 3240
rect 7620 3224 7642 3226
rect 7720 3224 7912 3236
rect 7991 3224 8004 3254
rect 8019 3240 8049 3254
rect 8086 3224 8105 3254
rect 8120 3224 8126 3254
rect 8135 3224 8148 3254
rect 8163 3240 8193 3254
rect 8236 3240 8279 3254
rect 8286 3240 8506 3254
rect 8513 3240 8543 3254
rect 8203 3226 8218 3238
rect 8237 3226 8250 3240
rect 8318 3236 8471 3240
rect 8200 3224 8222 3226
rect 8300 3224 8492 3236
rect 8571 3224 8584 3254
rect 8599 3240 8629 3254
rect 8666 3224 8685 3254
rect 8700 3224 8706 3254
rect 8715 3224 8728 3254
rect 8743 3240 8773 3254
rect 8816 3240 8859 3254
rect 8866 3240 9086 3254
rect 9093 3240 9123 3254
rect 8783 3226 8798 3238
rect 8817 3226 8830 3240
rect 8898 3236 9051 3240
rect 8780 3224 8802 3226
rect 8880 3224 9072 3236
rect 9151 3224 9164 3254
rect 9179 3240 9209 3254
rect 9246 3224 9265 3254
rect 9280 3224 9286 3254
rect 9295 3224 9308 3254
rect 9323 3240 9353 3254
rect 9396 3240 9439 3254
rect 9446 3240 9666 3254
rect 9673 3240 9703 3254
rect 9363 3226 9378 3238
rect 9397 3226 9410 3240
rect 9478 3236 9631 3240
rect 9360 3224 9382 3226
rect 9460 3224 9652 3236
rect 9731 3224 9744 3254
rect 9759 3240 9789 3254
rect 9826 3224 9845 3254
rect 9860 3224 9866 3254
rect 9875 3224 9888 3254
rect 9903 3240 9933 3254
rect 9976 3240 10019 3254
rect 10026 3240 10246 3254
rect 10253 3240 10283 3254
rect 9943 3226 9958 3238
rect 9977 3226 9990 3240
rect 10058 3236 10211 3240
rect 9940 3224 9962 3226
rect 10040 3224 10232 3236
rect 10311 3224 10324 3254
rect 10339 3240 10369 3254
rect 10406 3224 10425 3254
rect 10440 3224 10446 3254
rect 10455 3224 10468 3254
rect 10483 3240 10513 3254
rect 10556 3240 10599 3254
rect 10606 3240 10826 3254
rect 10833 3240 10863 3254
rect 10523 3226 10538 3238
rect 10557 3226 10570 3240
rect 10638 3236 10791 3240
rect 10520 3224 10542 3226
rect 10620 3224 10812 3236
rect 10891 3224 10904 3254
rect 10919 3240 10949 3254
rect 10986 3224 11005 3254
rect 11020 3224 11026 3254
rect 11035 3224 11048 3254
rect 11063 3240 11093 3254
rect 11136 3240 11179 3254
rect 11186 3240 11406 3254
rect 11413 3240 11443 3254
rect 11103 3226 11118 3238
rect 11137 3226 11150 3240
rect 11218 3236 11371 3240
rect 11100 3224 11122 3226
rect 11200 3224 11392 3236
rect 11471 3224 11484 3254
rect 11499 3240 11529 3254
rect 11566 3224 11585 3254
rect 11600 3224 11606 3254
rect 11615 3224 11628 3254
rect 11643 3240 11673 3254
rect 11716 3240 11759 3254
rect 11766 3240 11986 3254
rect 11993 3240 12023 3254
rect 11683 3226 11698 3238
rect 11717 3226 11730 3240
rect 11798 3236 11951 3240
rect 11680 3224 11702 3226
rect 11780 3224 11972 3236
rect 12051 3224 12064 3254
rect 12079 3240 12109 3254
rect 12146 3224 12165 3254
rect 12180 3224 12186 3254
rect 12195 3224 12208 3254
rect 12223 3240 12253 3254
rect 12296 3240 12339 3254
rect 12346 3240 12566 3254
rect 12573 3240 12603 3254
rect 12263 3226 12278 3238
rect 12297 3226 12310 3240
rect 12378 3236 12531 3240
rect 12260 3224 12282 3226
rect 12360 3224 12552 3236
rect 12631 3224 12644 3254
rect 12659 3240 12689 3254
rect 12726 3224 12745 3254
rect 12760 3224 12766 3254
rect 12775 3224 12788 3254
rect 12803 3240 12833 3254
rect 12876 3240 12919 3254
rect 12926 3240 13146 3254
rect 13153 3240 13183 3254
rect 12843 3226 12858 3238
rect 12877 3226 12890 3240
rect 12958 3236 13111 3240
rect 12840 3224 12862 3226
rect 12940 3224 13132 3236
rect 13211 3224 13224 3254
rect 13239 3240 13269 3254
rect 13306 3224 13325 3254
rect 13340 3224 13346 3254
rect 13355 3224 13368 3254
rect 13383 3240 13413 3254
rect 13456 3240 13499 3254
rect 13506 3240 13726 3254
rect 13733 3240 13763 3254
rect 13423 3226 13438 3238
rect 13457 3226 13470 3240
rect 13538 3236 13691 3240
rect 13420 3224 13442 3226
rect 13520 3224 13712 3236
rect 13791 3224 13804 3254
rect 13819 3240 13849 3254
rect 13886 3224 13905 3254
rect 13920 3224 13926 3254
rect 13935 3224 13948 3254
rect 13963 3240 13993 3254
rect 14036 3240 14079 3254
rect 14086 3240 14306 3254
rect 14313 3240 14343 3254
rect 14003 3226 14018 3238
rect 14037 3226 14050 3240
rect 14118 3236 14271 3240
rect 14000 3224 14022 3226
rect 14100 3224 14292 3236
rect 14371 3224 14384 3254
rect 14399 3240 14429 3254
rect 14466 3224 14485 3254
rect 14500 3224 14506 3254
rect 14515 3224 14528 3254
rect 14543 3240 14573 3254
rect 14616 3240 14659 3254
rect 14666 3240 14886 3254
rect 14893 3240 14923 3254
rect 14583 3226 14598 3238
rect 14617 3226 14630 3240
rect 14698 3236 14851 3240
rect 14580 3224 14602 3226
rect 14680 3224 14872 3236
rect 14951 3224 14964 3254
rect 14979 3240 15009 3254
rect 15046 3224 15065 3254
rect 15080 3224 15086 3254
rect 15095 3224 15108 3254
rect 15123 3240 15153 3254
rect 15196 3240 15239 3254
rect 15246 3240 15466 3254
rect 15473 3240 15503 3254
rect 15163 3226 15178 3238
rect 15197 3226 15210 3240
rect 15278 3236 15431 3240
rect 15160 3224 15182 3226
rect 15260 3224 15452 3236
rect 15531 3224 15544 3254
rect 15559 3240 15589 3254
rect 15626 3224 15645 3254
rect 15660 3224 15666 3254
rect 15675 3224 15688 3254
rect 15703 3240 15733 3254
rect 15776 3240 15819 3254
rect 15826 3240 16046 3254
rect 16053 3240 16083 3254
rect 15743 3226 15758 3238
rect 15777 3226 15790 3240
rect 15858 3236 16011 3240
rect 15740 3224 15762 3226
rect 15840 3224 16032 3236
rect 16111 3224 16124 3254
rect 16139 3240 16169 3254
rect 16206 3224 16225 3254
rect 16240 3224 16246 3254
rect 16255 3224 16268 3254
rect 16283 3240 16313 3254
rect 16356 3240 16399 3254
rect 16406 3240 16626 3254
rect 16633 3240 16663 3254
rect 16323 3226 16338 3238
rect 16357 3226 16370 3240
rect 16438 3236 16591 3240
rect 16320 3224 16342 3226
rect 16420 3224 16612 3236
rect 16691 3224 16704 3254
rect 16719 3240 16749 3254
rect 16786 3224 16805 3254
rect 16820 3224 16826 3254
rect 16835 3224 16848 3254
rect 16863 3240 16893 3254
rect 16936 3240 16979 3254
rect 16986 3240 17206 3254
rect 17213 3240 17243 3254
rect 16903 3226 16918 3238
rect 16937 3226 16950 3240
rect 17018 3236 17171 3240
rect 16900 3224 16922 3226
rect 17000 3224 17192 3236
rect 17271 3224 17284 3254
rect 17299 3240 17329 3254
rect 17366 3224 17385 3254
rect 17400 3224 17406 3254
rect 17415 3224 17428 3254
rect 17443 3240 17473 3254
rect 17516 3240 17559 3254
rect 17566 3240 17786 3254
rect 17793 3240 17823 3254
rect 17483 3226 17498 3238
rect 17517 3226 17530 3240
rect 17598 3236 17751 3240
rect 17480 3224 17502 3226
rect 17580 3224 17772 3236
rect 17851 3224 17864 3254
rect 17879 3240 17909 3254
rect 17946 3224 17965 3254
rect 17980 3224 17986 3254
rect 17995 3224 18008 3254
rect 18023 3240 18053 3254
rect 18096 3240 18139 3254
rect 18146 3240 18366 3254
rect 18373 3240 18403 3254
rect 18063 3226 18078 3238
rect 18097 3226 18110 3240
rect 18178 3236 18331 3240
rect 18060 3224 18082 3226
rect 18160 3224 18352 3236
rect 18431 3224 18444 3254
rect 18459 3240 18489 3254
rect 18532 3224 18545 3254
rect 0 3210 18545 3224
rect 15 3140 28 3210
rect 80 3206 102 3210
rect 73 3184 102 3198
rect 155 3184 171 3198
rect 209 3194 215 3196
rect 222 3194 330 3210
rect 337 3194 343 3196
rect 351 3194 366 3210
rect 432 3204 451 3207
rect 73 3182 171 3184
rect 198 3182 366 3194
rect 381 3184 397 3198
rect 432 3185 454 3204
rect 464 3198 480 3199
rect 463 3196 480 3198
rect 464 3191 480 3196
rect 454 3184 460 3185
rect 463 3184 492 3191
rect 381 3183 492 3184
rect 381 3182 498 3183
rect 57 3174 108 3182
rect 155 3174 189 3182
rect 57 3162 82 3174
rect 89 3162 108 3174
rect 162 3172 189 3174
rect 198 3172 419 3182
rect 454 3179 460 3182
rect 162 3168 419 3172
rect 57 3154 108 3162
rect 155 3154 419 3168
rect 463 3174 498 3182
rect 9 3106 28 3140
rect 73 3146 102 3154
rect 73 3140 90 3146
rect 73 3138 107 3140
rect 155 3138 171 3154
rect 172 3144 380 3154
rect 381 3144 397 3154
rect 445 3150 460 3165
rect 463 3162 464 3174
rect 471 3162 498 3174
rect 463 3154 498 3162
rect 463 3153 492 3154
rect 183 3140 397 3144
rect 198 3138 397 3140
rect 432 3140 445 3150
rect 463 3140 480 3153
rect 432 3138 480 3140
rect 74 3134 107 3138
rect 70 3132 107 3134
rect 70 3131 137 3132
rect 70 3126 101 3131
rect 107 3126 137 3131
rect 70 3122 137 3126
rect 43 3119 137 3122
rect 43 3112 92 3119
rect 43 3106 73 3112
rect 92 3107 97 3112
rect 9 3090 89 3106
rect 101 3098 137 3119
rect 198 3114 387 3138
rect 432 3137 479 3138
rect 445 3132 479 3137
rect 213 3111 387 3114
rect 206 3108 387 3111
rect 415 3131 479 3132
rect 9 3088 28 3090
rect 43 3088 77 3090
rect 9 3072 89 3088
rect 9 3066 28 3072
rect -1 3050 28 3066
rect 43 3056 73 3072
rect 101 3050 107 3098
rect 110 3092 129 3098
rect 144 3092 174 3100
rect 110 3084 174 3092
rect 110 3068 190 3084
rect 206 3077 268 3108
rect 284 3077 346 3108
rect 415 3106 464 3131
rect 479 3106 509 3122
rect 378 3092 408 3100
rect 415 3098 525 3106
rect 378 3084 423 3092
rect 110 3066 129 3068
rect 144 3066 190 3068
rect 110 3050 190 3066
rect 217 3064 252 3077
rect 293 3074 330 3077
rect 293 3072 335 3074
rect 222 3061 252 3064
rect 231 3057 238 3061
rect 238 3056 239 3057
rect 197 3050 207 3056
rect -7 3042 34 3050
rect -7 3016 8 3042
rect 15 3016 34 3042
rect 98 3038 129 3050
rect 144 3038 247 3050
rect 259 3040 285 3066
rect 300 3061 330 3072
rect 362 3068 424 3084
rect 362 3066 408 3068
rect 362 3050 424 3066
rect 436 3050 442 3098
rect 445 3090 525 3098
rect 445 3088 464 3090
rect 479 3088 513 3090
rect 445 3072 525 3088
rect 445 3050 464 3072
rect 479 3056 509 3072
rect 537 3066 543 3140
rect 546 3066 565 3210
rect 580 3066 586 3210
rect 595 3140 608 3210
rect 660 3206 682 3210
rect 653 3184 682 3198
rect 735 3184 751 3198
rect 789 3194 795 3196
rect 802 3194 910 3210
rect 917 3194 923 3196
rect 931 3194 946 3210
rect 1012 3204 1031 3207
rect 653 3182 751 3184
rect 778 3182 946 3194
rect 961 3184 977 3198
rect 1012 3185 1034 3204
rect 1044 3198 1060 3199
rect 1043 3196 1060 3198
rect 1044 3191 1060 3196
rect 1034 3184 1040 3185
rect 1043 3184 1072 3191
rect 961 3183 1072 3184
rect 961 3182 1078 3183
rect 637 3174 688 3182
rect 735 3174 769 3182
rect 637 3162 662 3174
rect 669 3162 688 3174
rect 742 3172 769 3174
rect 778 3172 999 3182
rect 1034 3179 1040 3182
rect 742 3168 999 3172
rect 637 3154 688 3162
rect 735 3154 999 3168
rect 1043 3174 1078 3182
rect 589 3106 608 3140
rect 653 3146 682 3154
rect 653 3140 670 3146
rect 653 3138 687 3140
rect 735 3138 751 3154
rect 752 3144 960 3154
rect 961 3144 977 3154
rect 1025 3150 1040 3165
rect 1043 3162 1044 3174
rect 1051 3162 1078 3174
rect 1043 3154 1078 3162
rect 1043 3153 1072 3154
rect 763 3140 977 3144
rect 778 3138 977 3140
rect 1012 3140 1025 3150
rect 1043 3140 1060 3153
rect 1012 3138 1060 3140
rect 654 3134 687 3138
rect 650 3132 687 3134
rect 650 3131 717 3132
rect 650 3126 681 3131
rect 687 3126 717 3131
rect 650 3122 717 3126
rect 623 3119 717 3122
rect 623 3112 672 3119
rect 623 3106 653 3112
rect 672 3107 677 3112
rect 589 3090 669 3106
rect 681 3098 717 3119
rect 778 3114 967 3138
rect 1012 3137 1059 3138
rect 1025 3132 1059 3137
rect 793 3111 967 3114
rect 786 3108 967 3111
rect 995 3131 1059 3132
rect 589 3088 608 3090
rect 623 3088 657 3090
rect 589 3072 669 3088
rect 589 3066 608 3072
rect 305 3040 408 3050
rect 259 3038 408 3040
rect 429 3038 464 3050
rect 98 3036 260 3038
rect 110 3016 129 3036
rect 144 3034 174 3036
rect -7 3008 34 3016
rect 116 3012 129 3016
rect 181 3020 260 3036
rect 292 3036 464 3038
rect 292 3020 371 3036
rect 378 3034 408 3036
rect -1 2998 28 3008
rect 43 2998 73 3012
rect 116 2998 159 3012
rect 181 3008 371 3020
rect 436 3016 442 3036
rect 166 2998 196 3008
rect 197 2998 355 3008
rect 359 2998 389 3008
rect 393 2998 423 3012
rect 451 2998 464 3036
rect 536 3050 565 3066
rect 579 3050 608 3066
rect 623 3056 653 3072
rect 681 3050 687 3098
rect 690 3092 709 3098
rect 724 3092 754 3100
rect 690 3084 754 3092
rect 690 3068 770 3084
rect 786 3077 848 3108
rect 864 3077 926 3108
rect 995 3106 1044 3131
rect 1059 3106 1089 3122
rect 958 3092 988 3100
rect 995 3098 1105 3106
rect 958 3084 1003 3092
rect 690 3066 709 3068
rect 724 3066 770 3068
rect 690 3050 770 3066
rect 797 3064 832 3077
rect 873 3074 910 3077
rect 873 3072 915 3074
rect 802 3061 832 3064
rect 811 3057 818 3061
rect 818 3056 819 3057
rect 777 3050 787 3056
rect 536 3042 571 3050
rect 536 3016 537 3042
rect 544 3016 571 3042
rect 479 2998 509 3012
rect 536 3008 571 3016
rect 573 3042 614 3050
rect 573 3016 588 3042
rect 595 3016 614 3042
rect 678 3038 709 3050
rect 724 3038 827 3050
rect 839 3040 865 3066
rect 880 3061 910 3072
rect 942 3068 1004 3084
rect 942 3066 988 3068
rect 942 3050 1004 3066
rect 1016 3050 1022 3098
rect 1025 3090 1105 3098
rect 1025 3088 1044 3090
rect 1059 3088 1093 3090
rect 1025 3072 1105 3088
rect 1025 3050 1044 3072
rect 1059 3056 1089 3072
rect 1117 3066 1123 3140
rect 1126 3066 1145 3210
rect 1160 3066 1166 3210
rect 1175 3140 1188 3210
rect 1240 3206 1262 3210
rect 1233 3184 1262 3198
rect 1315 3184 1331 3198
rect 1369 3194 1375 3196
rect 1382 3194 1490 3210
rect 1497 3194 1503 3196
rect 1511 3194 1526 3210
rect 1592 3204 1611 3207
rect 1233 3182 1331 3184
rect 1358 3182 1526 3194
rect 1541 3184 1557 3198
rect 1592 3185 1614 3204
rect 1624 3198 1640 3199
rect 1623 3196 1640 3198
rect 1624 3191 1640 3196
rect 1614 3184 1620 3185
rect 1623 3184 1652 3191
rect 1541 3183 1652 3184
rect 1541 3182 1658 3183
rect 1217 3174 1268 3182
rect 1315 3174 1349 3182
rect 1217 3162 1242 3174
rect 1249 3162 1268 3174
rect 1322 3172 1349 3174
rect 1358 3172 1579 3182
rect 1614 3179 1620 3182
rect 1322 3168 1579 3172
rect 1217 3154 1268 3162
rect 1315 3154 1579 3168
rect 1623 3174 1658 3182
rect 1169 3106 1188 3140
rect 1233 3146 1262 3154
rect 1233 3140 1250 3146
rect 1233 3138 1267 3140
rect 1315 3138 1331 3154
rect 1332 3144 1540 3154
rect 1541 3144 1557 3154
rect 1605 3150 1620 3165
rect 1623 3162 1624 3174
rect 1631 3162 1658 3174
rect 1623 3154 1658 3162
rect 1623 3153 1652 3154
rect 1343 3140 1557 3144
rect 1358 3138 1557 3140
rect 1592 3140 1605 3150
rect 1623 3140 1640 3153
rect 1592 3138 1640 3140
rect 1234 3134 1267 3138
rect 1230 3132 1267 3134
rect 1230 3131 1297 3132
rect 1230 3126 1261 3131
rect 1267 3126 1297 3131
rect 1230 3122 1297 3126
rect 1203 3119 1297 3122
rect 1203 3112 1252 3119
rect 1203 3106 1233 3112
rect 1252 3107 1257 3112
rect 1169 3090 1249 3106
rect 1261 3098 1297 3119
rect 1358 3114 1547 3138
rect 1592 3137 1639 3138
rect 1605 3132 1639 3137
rect 1373 3111 1547 3114
rect 1366 3108 1547 3111
rect 1575 3131 1639 3132
rect 1169 3088 1188 3090
rect 1203 3088 1237 3090
rect 1169 3072 1249 3088
rect 1169 3066 1188 3072
rect 885 3040 988 3050
rect 839 3038 988 3040
rect 1009 3038 1044 3050
rect 678 3036 840 3038
rect 690 3016 709 3036
rect 724 3034 754 3036
rect 573 3008 614 3016
rect 696 3012 709 3016
rect 761 3020 840 3036
rect 872 3036 1044 3038
rect 872 3020 951 3036
rect 958 3034 988 3036
rect 536 2998 565 3008
rect 579 2998 608 3008
rect 623 2998 653 3012
rect 696 2998 739 3012
rect 761 3008 951 3020
rect 1016 3016 1022 3036
rect 746 2998 776 3008
rect 777 2998 935 3008
rect 939 2998 969 3008
rect 973 2998 1003 3012
rect 1031 2998 1044 3036
rect 1116 3050 1145 3066
rect 1159 3050 1188 3066
rect 1203 3056 1233 3072
rect 1261 3050 1267 3098
rect 1270 3092 1289 3098
rect 1304 3092 1334 3100
rect 1270 3084 1334 3092
rect 1270 3068 1350 3084
rect 1366 3077 1428 3108
rect 1444 3077 1506 3108
rect 1575 3106 1624 3131
rect 1639 3106 1669 3122
rect 1538 3092 1568 3100
rect 1575 3098 1685 3106
rect 1538 3084 1583 3092
rect 1270 3066 1289 3068
rect 1304 3066 1350 3068
rect 1270 3050 1350 3066
rect 1377 3064 1412 3077
rect 1453 3074 1490 3077
rect 1453 3072 1495 3074
rect 1382 3061 1412 3064
rect 1391 3057 1398 3061
rect 1398 3056 1399 3057
rect 1357 3050 1367 3056
rect 1116 3042 1151 3050
rect 1116 3016 1117 3042
rect 1124 3016 1151 3042
rect 1059 2998 1089 3012
rect 1116 3008 1151 3016
rect 1153 3042 1194 3050
rect 1153 3016 1168 3042
rect 1175 3016 1194 3042
rect 1258 3038 1289 3050
rect 1304 3038 1407 3050
rect 1419 3040 1445 3066
rect 1460 3061 1490 3072
rect 1522 3068 1584 3084
rect 1522 3066 1568 3068
rect 1522 3050 1584 3066
rect 1596 3050 1602 3098
rect 1605 3090 1685 3098
rect 1605 3088 1624 3090
rect 1639 3088 1673 3090
rect 1605 3072 1685 3088
rect 1605 3050 1624 3072
rect 1639 3056 1669 3072
rect 1697 3066 1703 3140
rect 1706 3066 1725 3210
rect 1740 3066 1746 3210
rect 1755 3140 1768 3210
rect 1820 3206 1842 3210
rect 1813 3184 1842 3198
rect 1895 3184 1911 3198
rect 1949 3194 1955 3196
rect 1962 3194 2070 3210
rect 2077 3194 2083 3196
rect 2091 3194 2106 3210
rect 2172 3204 2191 3207
rect 1813 3182 1911 3184
rect 1938 3182 2106 3194
rect 2121 3184 2137 3198
rect 2172 3185 2194 3204
rect 2204 3198 2220 3199
rect 2203 3196 2220 3198
rect 2204 3191 2220 3196
rect 2194 3184 2200 3185
rect 2203 3184 2232 3191
rect 2121 3183 2232 3184
rect 2121 3182 2238 3183
rect 1797 3174 1848 3182
rect 1895 3174 1929 3182
rect 1797 3162 1822 3174
rect 1829 3162 1848 3174
rect 1902 3172 1929 3174
rect 1938 3172 2159 3182
rect 2194 3179 2200 3182
rect 1902 3168 2159 3172
rect 1797 3154 1848 3162
rect 1895 3154 2159 3168
rect 2203 3174 2238 3182
rect 1749 3106 1768 3140
rect 1813 3146 1842 3154
rect 1813 3140 1830 3146
rect 1813 3138 1847 3140
rect 1895 3138 1911 3154
rect 1912 3144 2120 3154
rect 2121 3144 2137 3154
rect 2185 3150 2200 3165
rect 2203 3162 2204 3174
rect 2211 3162 2238 3174
rect 2203 3154 2238 3162
rect 2203 3153 2232 3154
rect 1923 3140 2137 3144
rect 1938 3138 2137 3140
rect 2172 3140 2185 3150
rect 2203 3140 2220 3153
rect 2172 3138 2220 3140
rect 1814 3134 1847 3138
rect 1810 3132 1847 3134
rect 1810 3131 1877 3132
rect 1810 3126 1841 3131
rect 1847 3126 1877 3131
rect 1810 3122 1877 3126
rect 1783 3119 1877 3122
rect 1783 3112 1832 3119
rect 1783 3106 1813 3112
rect 1832 3107 1837 3112
rect 1749 3090 1829 3106
rect 1841 3098 1877 3119
rect 1938 3114 2127 3138
rect 2172 3137 2219 3138
rect 2185 3132 2219 3137
rect 1953 3111 2127 3114
rect 1946 3108 2127 3111
rect 2155 3131 2219 3132
rect 1749 3088 1768 3090
rect 1783 3088 1817 3090
rect 1749 3072 1829 3088
rect 1749 3066 1768 3072
rect 1465 3040 1568 3050
rect 1419 3038 1568 3040
rect 1589 3038 1624 3050
rect 1258 3036 1420 3038
rect 1270 3016 1289 3036
rect 1304 3034 1334 3036
rect 1153 3008 1194 3016
rect 1276 3012 1289 3016
rect 1341 3020 1420 3036
rect 1452 3036 1624 3038
rect 1452 3020 1531 3036
rect 1538 3034 1568 3036
rect 1116 2998 1145 3008
rect 1159 2998 1188 3008
rect 1203 2998 1233 3012
rect 1276 2998 1319 3012
rect 1341 3008 1531 3020
rect 1596 3016 1602 3036
rect 1326 2998 1356 3008
rect 1357 2998 1515 3008
rect 1519 2998 1549 3008
rect 1553 2998 1583 3012
rect 1611 2998 1624 3036
rect 1696 3050 1725 3066
rect 1739 3050 1768 3066
rect 1783 3056 1813 3072
rect 1841 3050 1847 3098
rect 1850 3092 1869 3098
rect 1884 3092 1914 3100
rect 1850 3084 1914 3092
rect 1850 3068 1930 3084
rect 1946 3077 2008 3108
rect 2024 3077 2086 3108
rect 2155 3106 2204 3131
rect 2219 3106 2249 3122
rect 2118 3092 2148 3100
rect 2155 3098 2265 3106
rect 2118 3084 2163 3092
rect 1850 3066 1869 3068
rect 1884 3066 1930 3068
rect 1850 3050 1930 3066
rect 1957 3064 1992 3077
rect 2033 3074 2070 3077
rect 2033 3072 2075 3074
rect 1962 3061 1992 3064
rect 1971 3057 1978 3061
rect 1978 3056 1979 3057
rect 1937 3050 1947 3056
rect 1696 3042 1731 3050
rect 1696 3016 1697 3042
rect 1704 3016 1731 3042
rect 1639 2998 1669 3012
rect 1696 3008 1731 3016
rect 1733 3042 1774 3050
rect 1733 3016 1748 3042
rect 1755 3016 1774 3042
rect 1838 3038 1869 3050
rect 1884 3038 1987 3050
rect 1999 3040 2025 3066
rect 2040 3061 2070 3072
rect 2102 3068 2164 3084
rect 2102 3066 2148 3068
rect 2102 3050 2164 3066
rect 2176 3050 2182 3098
rect 2185 3090 2265 3098
rect 2185 3088 2204 3090
rect 2219 3088 2253 3090
rect 2185 3072 2265 3088
rect 2185 3050 2204 3072
rect 2219 3056 2249 3072
rect 2277 3066 2283 3140
rect 2286 3066 2305 3210
rect 2320 3066 2326 3210
rect 2335 3140 2348 3210
rect 2400 3206 2422 3210
rect 2393 3184 2422 3198
rect 2475 3184 2491 3198
rect 2529 3194 2535 3196
rect 2542 3194 2650 3210
rect 2657 3194 2663 3196
rect 2671 3194 2686 3210
rect 2752 3204 2771 3207
rect 2393 3182 2491 3184
rect 2518 3182 2686 3194
rect 2701 3184 2717 3198
rect 2752 3185 2774 3204
rect 2784 3198 2800 3199
rect 2783 3196 2800 3198
rect 2784 3191 2800 3196
rect 2774 3184 2780 3185
rect 2783 3184 2812 3191
rect 2701 3183 2812 3184
rect 2701 3182 2818 3183
rect 2377 3174 2428 3182
rect 2475 3174 2509 3182
rect 2377 3162 2402 3174
rect 2409 3162 2428 3174
rect 2482 3172 2509 3174
rect 2518 3172 2739 3182
rect 2774 3179 2780 3182
rect 2482 3168 2739 3172
rect 2377 3154 2428 3162
rect 2475 3154 2739 3168
rect 2783 3174 2818 3182
rect 2329 3106 2348 3140
rect 2393 3146 2422 3154
rect 2393 3140 2410 3146
rect 2393 3138 2427 3140
rect 2475 3138 2491 3154
rect 2492 3144 2700 3154
rect 2701 3144 2717 3154
rect 2765 3150 2780 3165
rect 2783 3162 2784 3174
rect 2791 3162 2818 3174
rect 2783 3154 2818 3162
rect 2783 3153 2812 3154
rect 2503 3140 2717 3144
rect 2518 3138 2717 3140
rect 2752 3140 2765 3150
rect 2783 3140 2800 3153
rect 2752 3138 2800 3140
rect 2394 3134 2427 3138
rect 2390 3132 2427 3134
rect 2390 3131 2457 3132
rect 2390 3126 2421 3131
rect 2427 3126 2457 3131
rect 2390 3122 2457 3126
rect 2363 3119 2457 3122
rect 2363 3112 2412 3119
rect 2363 3106 2393 3112
rect 2412 3107 2417 3112
rect 2329 3090 2409 3106
rect 2421 3098 2457 3119
rect 2518 3114 2707 3138
rect 2752 3137 2799 3138
rect 2765 3132 2799 3137
rect 2533 3111 2707 3114
rect 2526 3108 2707 3111
rect 2735 3131 2799 3132
rect 2329 3088 2348 3090
rect 2363 3088 2397 3090
rect 2329 3072 2409 3088
rect 2329 3066 2348 3072
rect 2045 3040 2148 3050
rect 1999 3038 2148 3040
rect 2169 3038 2204 3050
rect 1838 3036 2000 3038
rect 1850 3016 1869 3036
rect 1884 3034 1914 3036
rect 1733 3008 1774 3016
rect 1856 3012 1869 3016
rect 1921 3020 2000 3036
rect 2032 3036 2204 3038
rect 2032 3020 2111 3036
rect 2118 3034 2148 3036
rect 1696 2998 1725 3008
rect 1739 2998 1768 3008
rect 1783 2998 1813 3012
rect 1856 2998 1899 3012
rect 1921 3008 2111 3020
rect 2176 3016 2182 3036
rect 1906 2998 1936 3008
rect 1937 2998 2095 3008
rect 2099 2998 2129 3008
rect 2133 2998 2163 3012
rect 2191 2998 2204 3036
rect 2276 3050 2305 3066
rect 2319 3050 2348 3066
rect 2363 3056 2393 3072
rect 2421 3050 2427 3098
rect 2430 3092 2449 3098
rect 2464 3092 2494 3100
rect 2430 3084 2494 3092
rect 2430 3068 2510 3084
rect 2526 3077 2588 3108
rect 2604 3077 2666 3108
rect 2735 3106 2784 3131
rect 2799 3106 2829 3122
rect 2698 3092 2728 3100
rect 2735 3098 2845 3106
rect 2698 3084 2743 3092
rect 2430 3066 2449 3068
rect 2464 3066 2510 3068
rect 2430 3050 2510 3066
rect 2537 3064 2572 3077
rect 2613 3074 2650 3077
rect 2613 3072 2655 3074
rect 2542 3061 2572 3064
rect 2551 3057 2558 3061
rect 2558 3056 2559 3057
rect 2517 3050 2527 3056
rect 2276 3042 2311 3050
rect 2276 3016 2277 3042
rect 2284 3016 2311 3042
rect 2219 2998 2249 3012
rect 2276 3008 2311 3016
rect 2313 3042 2354 3050
rect 2313 3016 2328 3042
rect 2335 3016 2354 3042
rect 2418 3038 2449 3050
rect 2464 3038 2567 3050
rect 2579 3040 2605 3066
rect 2620 3061 2650 3072
rect 2682 3068 2744 3084
rect 2682 3066 2728 3068
rect 2682 3050 2744 3066
rect 2756 3050 2762 3098
rect 2765 3090 2845 3098
rect 2765 3088 2784 3090
rect 2799 3088 2833 3090
rect 2765 3072 2845 3088
rect 2765 3050 2784 3072
rect 2799 3056 2829 3072
rect 2857 3066 2863 3140
rect 2866 3066 2885 3210
rect 2900 3066 2906 3210
rect 2915 3140 2928 3210
rect 2980 3206 3002 3210
rect 2973 3184 3002 3198
rect 3055 3184 3071 3198
rect 3109 3194 3115 3196
rect 3122 3194 3230 3210
rect 3237 3194 3243 3196
rect 3251 3194 3266 3210
rect 3332 3204 3351 3207
rect 2973 3182 3071 3184
rect 3098 3182 3266 3194
rect 3281 3184 3297 3198
rect 3332 3185 3354 3204
rect 3364 3198 3380 3199
rect 3363 3196 3380 3198
rect 3364 3191 3380 3196
rect 3354 3184 3360 3185
rect 3363 3184 3392 3191
rect 3281 3183 3392 3184
rect 3281 3182 3398 3183
rect 2957 3174 3008 3182
rect 3055 3174 3089 3182
rect 2957 3162 2982 3174
rect 2989 3162 3008 3174
rect 3062 3172 3089 3174
rect 3098 3172 3319 3182
rect 3354 3179 3360 3182
rect 3062 3168 3319 3172
rect 2957 3154 3008 3162
rect 3055 3154 3319 3168
rect 3363 3174 3398 3182
rect 2909 3106 2928 3140
rect 2973 3146 3002 3154
rect 2973 3140 2990 3146
rect 2973 3138 3007 3140
rect 3055 3138 3071 3154
rect 3072 3144 3280 3154
rect 3281 3144 3297 3154
rect 3345 3150 3360 3165
rect 3363 3162 3364 3174
rect 3371 3162 3398 3174
rect 3363 3154 3398 3162
rect 3363 3153 3392 3154
rect 3083 3140 3297 3144
rect 3098 3138 3297 3140
rect 3332 3140 3345 3150
rect 3363 3140 3380 3153
rect 3332 3138 3380 3140
rect 2974 3134 3007 3138
rect 2970 3132 3007 3134
rect 2970 3131 3037 3132
rect 2970 3126 3001 3131
rect 3007 3126 3037 3131
rect 2970 3122 3037 3126
rect 2943 3119 3037 3122
rect 2943 3112 2992 3119
rect 2943 3106 2973 3112
rect 2992 3107 2997 3112
rect 2909 3090 2989 3106
rect 3001 3098 3037 3119
rect 3098 3114 3287 3138
rect 3332 3137 3379 3138
rect 3345 3132 3379 3137
rect 3113 3111 3287 3114
rect 3106 3108 3287 3111
rect 3315 3131 3379 3132
rect 2909 3088 2928 3090
rect 2943 3088 2977 3090
rect 2909 3072 2989 3088
rect 2909 3066 2928 3072
rect 2625 3040 2728 3050
rect 2579 3038 2728 3040
rect 2749 3038 2784 3050
rect 2418 3036 2580 3038
rect 2430 3016 2449 3036
rect 2464 3034 2494 3036
rect 2313 3008 2354 3016
rect 2436 3012 2449 3016
rect 2501 3020 2580 3036
rect 2612 3036 2784 3038
rect 2612 3020 2691 3036
rect 2698 3034 2728 3036
rect 2276 2998 2305 3008
rect 2319 2998 2348 3008
rect 2363 2998 2393 3012
rect 2436 2998 2479 3012
rect 2501 3008 2691 3020
rect 2756 3016 2762 3036
rect 2486 2998 2516 3008
rect 2517 2998 2675 3008
rect 2679 2998 2709 3008
rect 2713 2998 2743 3012
rect 2771 2998 2784 3036
rect 2856 3050 2885 3066
rect 2899 3050 2928 3066
rect 2943 3056 2973 3072
rect 3001 3050 3007 3098
rect 3010 3092 3029 3098
rect 3044 3092 3074 3100
rect 3010 3084 3074 3092
rect 3010 3068 3090 3084
rect 3106 3077 3168 3108
rect 3184 3077 3246 3108
rect 3315 3106 3364 3131
rect 3379 3106 3409 3122
rect 3278 3092 3308 3100
rect 3315 3098 3425 3106
rect 3278 3084 3323 3092
rect 3010 3066 3029 3068
rect 3044 3066 3090 3068
rect 3010 3050 3090 3066
rect 3117 3064 3152 3077
rect 3193 3074 3230 3077
rect 3193 3072 3235 3074
rect 3122 3061 3152 3064
rect 3131 3057 3138 3061
rect 3138 3056 3139 3057
rect 3097 3050 3107 3056
rect 2856 3042 2891 3050
rect 2856 3016 2857 3042
rect 2864 3016 2891 3042
rect 2799 2998 2829 3012
rect 2856 3008 2891 3016
rect 2893 3042 2934 3050
rect 2893 3016 2908 3042
rect 2915 3016 2934 3042
rect 2998 3038 3029 3050
rect 3044 3038 3147 3050
rect 3159 3040 3185 3066
rect 3200 3061 3230 3072
rect 3262 3068 3324 3084
rect 3262 3066 3308 3068
rect 3262 3050 3324 3066
rect 3336 3050 3342 3098
rect 3345 3090 3425 3098
rect 3345 3088 3364 3090
rect 3379 3088 3413 3090
rect 3345 3072 3425 3088
rect 3345 3050 3364 3072
rect 3379 3056 3409 3072
rect 3437 3066 3443 3140
rect 3446 3066 3465 3210
rect 3480 3066 3486 3210
rect 3495 3140 3508 3210
rect 3560 3206 3582 3210
rect 3553 3184 3582 3198
rect 3635 3184 3651 3198
rect 3689 3194 3695 3196
rect 3702 3194 3810 3210
rect 3817 3194 3823 3196
rect 3831 3194 3846 3210
rect 3912 3204 3931 3207
rect 3553 3182 3651 3184
rect 3678 3182 3846 3194
rect 3861 3184 3877 3198
rect 3912 3185 3934 3204
rect 3944 3198 3960 3199
rect 3943 3196 3960 3198
rect 3944 3191 3960 3196
rect 3934 3184 3940 3185
rect 3943 3184 3972 3191
rect 3861 3183 3972 3184
rect 3861 3182 3978 3183
rect 3537 3174 3588 3182
rect 3635 3174 3669 3182
rect 3537 3162 3562 3174
rect 3569 3162 3588 3174
rect 3642 3172 3669 3174
rect 3678 3172 3899 3182
rect 3934 3179 3940 3182
rect 3642 3168 3899 3172
rect 3537 3154 3588 3162
rect 3635 3154 3899 3168
rect 3943 3174 3978 3182
rect 3489 3106 3508 3140
rect 3553 3146 3582 3154
rect 3553 3140 3570 3146
rect 3553 3138 3587 3140
rect 3635 3138 3651 3154
rect 3652 3144 3860 3154
rect 3861 3144 3877 3154
rect 3925 3150 3940 3165
rect 3943 3162 3944 3174
rect 3951 3162 3978 3174
rect 3943 3154 3978 3162
rect 3943 3153 3972 3154
rect 3663 3140 3877 3144
rect 3678 3138 3877 3140
rect 3912 3140 3925 3150
rect 3943 3140 3960 3153
rect 3912 3138 3960 3140
rect 3554 3134 3587 3138
rect 3550 3132 3587 3134
rect 3550 3131 3617 3132
rect 3550 3126 3581 3131
rect 3587 3126 3617 3131
rect 3550 3122 3617 3126
rect 3523 3119 3617 3122
rect 3523 3112 3572 3119
rect 3523 3106 3553 3112
rect 3572 3107 3577 3112
rect 3489 3090 3569 3106
rect 3581 3098 3617 3119
rect 3678 3114 3867 3138
rect 3912 3137 3959 3138
rect 3925 3132 3959 3137
rect 3693 3111 3867 3114
rect 3686 3108 3867 3111
rect 3895 3131 3959 3132
rect 3489 3088 3508 3090
rect 3523 3088 3557 3090
rect 3489 3072 3569 3088
rect 3489 3066 3508 3072
rect 3205 3040 3308 3050
rect 3159 3038 3308 3040
rect 3329 3038 3364 3050
rect 2998 3036 3160 3038
rect 3010 3016 3029 3036
rect 3044 3034 3074 3036
rect 2893 3008 2934 3016
rect 3016 3012 3029 3016
rect 3081 3020 3160 3036
rect 3192 3036 3364 3038
rect 3192 3020 3271 3036
rect 3278 3034 3308 3036
rect 2856 2998 2885 3008
rect 2899 2998 2928 3008
rect 2943 2998 2973 3012
rect 3016 2998 3059 3012
rect 3081 3008 3271 3020
rect 3336 3016 3342 3036
rect 3066 2998 3096 3008
rect 3097 2998 3255 3008
rect 3259 2998 3289 3008
rect 3293 2998 3323 3012
rect 3351 2998 3364 3036
rect 3436 3050 3465 3066
rect 3479 3050 3508 3066
rect 3523 3056 3553 3072
rect 3581 3050 3587 3098
rect 3590 3092 3609 3098
rect 3624 3092 3654 3100
rect 3590 3084 3654 3092
rect 3590 3068 3670 3084
rect 3686 3077 3748 3108
rect 3764 3077 3826 3108
rect 3895 3106 3944 3131
rect 3959 3106 3989 3122
rect 3858 3092 3888 3100
rect 3895 3098 4005 3106
rect 3858 3084 3903 3092
rect 3590 3066 3609 3068
rect 3624 3066 3670 3068
rect 3590 3050 3670 3066
rect 3697 3064 3732 3077
rect 3773 3074 3810 3077
rect 3773 3072 3815 3074
rect 3702 3061 3732 3064
rect 3711 3057 3718 3061
rect 3718 3056 3719 3057
rect 3677 3050 3687 3056
rect 3436 3042 3471 3050
rect 3436 3016 3437 3042
rect 3444 3016 3471 3042
rect 3379 2998 3409 3012
rect 3436 3008 3471 3016
rect 3473 3042 3514 3050
rect 3473 3016 3488 3042
rect 3495 3016 3514 3042
rect 3578 3038 3609 3050
rect 3624 3038 3727 3050
rect 3739 3040 3765 3066
rect 3780 3061 3810 3072
rect 3842 3068 3904 3084
rect 3842 3066 3888 3068
rect 3842 3050 3904 3066
rect 3916 3050 3922 3098
rect 3925 3090 4005 3098
rect 3925 3088 3944 3090
rect 3959 3088 3993 3090
rect 3925 3072 4005 3088
rect 3925 3050 3944 3072
rect 3959 3056 3989 3072
rect 4017 3066 4023 3140
rect 4026 3066 4045 3210
rect 4060 3066 4066 3210
rect 4075 3140 4088 3210
rect 4140 3206 4162 3210
rect 4133 3184 4162 3198
rect 4215 3184 4231 3198
rect 4269 3194 4275 3196
rect 4282 3194 4390 3210
rect 4397 3194 4403 3196
rect 4411 3194 4426 3210
rect 4492 3204 4511 3207
rect 4133 3182 4231 3184
rect 4258 3182 4426 3194
rect 4441 3184 4457 3198
rect 4492 3185 4514 3204
rect 4524 3198 4540 3199
rect 4523 3196 4540 3198
rect 4524 3191 4540 3196
rect 4514 3184 4520 3185
rect 4523 3184 4552 3191
rect 4441 3183 4552 3184
rect 4441 3182 4558 3183
rect 4117 3174 4168 3182
rect 4215 3174 4249 3182
rect 4117 3162 4142 3174
rect 4149 3162 4168 3174
rect 4222 3172 4249 3174
rect 4258 3172 4479 3182
rect 4514 3179 4520 3182
rect 4222 3168 4479 3172
rect 4117 3154 4168 3162
rect 4215 3154 4479 3168
rect 4523 3174 4558 3182
rect 4069 3106 4088 3140
rect 4133 3146 4162 3154
rect 4133 3140 4150 3146
rect 4133 3138 4167 3140
rect 4215 3138 4231 3154
rect 4232 3144 4440 3154
rect 4441 3144 4457 3154
rect 4505 3150 4520 3165
rect 4523 3162 4524 3174
rect 4531 3162 4558 3174
rect 4523 3154 4558 3162
rect 4523 3153 4552 3154
rect 4243 3140 4457 3144
rect 4258 3138 4457 3140
rect 4492 3140 4505 3150
rect 4523 3140 4540 3153
rect 4492 3138 4540 3140
rect 4134 3134 4167 3138
rect 4130 3132 4167 3134
rect 4130 3131 4197 3132
rect 4130 3126 4161 3131
rect 4167 3126 4197 3131
rect 4130 3122 4197 3126
rect 4103 3119 4197 3122
rect 4103 3112 4152 3119
rect 4103 3106 4133 3112
rect 4152 3107 4157 3112
rect 4069 3090 4149 3106
rect 4161 3098 4197 3119
rect 4258 3114 4447 3138
rect 4492 3137 4539 3138
rect 4505 3132 4539 3137
rect 4273 3111 4447 3114
rect 4266 3108 4447 3111
rect 4475 3131 4539 3132
rect 4069 3088 4088 3090
rect 4103 3088 4137 3090
rect 4069 3072 4149 3088
rect 4069 3066 4088 3072
rect 3785 3040 3888 3050
rect 3739 3038 3888 3040
rect 3909 3038 3944 3050
rect 3578 3036 3740 3038
rect 3590 3016 3609 3036
rect 3624 3034 3654 3036
rect 3473 3008 3514 3016
rect 3596 3012 3609 3016
rect 3661 3020 3740 3036
rect 3772 3036 3944 3038
rect 3772 3020 3851 3036
rect 3858 3034 3888 3036
rect 3436 2998 3465 3008
rect 3479 2998 3508 3008
rect 3523 2998 3553 3012
rect 3596 2998 3639 3012
rect 3661 3008 3851 3020
rect 3916 3016 3922 3036
rect 3646 2998 3676 3008
rect 3677 2998 3835 3008
rect 3839 2998 3869 3008
rect 3873 2998 3903 3012
rect 3931 2998 3944 3036
rect 4016 3050 4045 3066
rect 4059 3050 4088 3066
rect 4103 3056 4133 3072
rect 4161 3050 4167 3098
rect 4170 3092 4189 3098
rect 4204 3092 4234 3100
rect 4170 3084 4234 3092
rect 4170 3068 4250 3084
rect 4266 3077 4328 3108
rect 4344 3077 4406 3108
rect 4475 3106 4524 3131
rect 4539 3106 4569 3122
rect 4438 3092 4468 3100
rect 4475 3098 4585 3106
rect 4438 3084 4483 3092
rect 4170 3066 4189 3068
rect 4204 3066 4250 3068
rect 4170 3050 4250 3066
rect 4277 3064 4312 3077
rect 4353 3074 4390 3077
rect 4353 3072 4395 3074
rect 4282 3061 4312 3064
rect 4291 3057 4298 3061
rect 4298 3056 4299 3057
rect 4257 3050 4267 3056
rect 4016 3042 4051 3050
rect 4016 3016 4017 3042
rect 4024 3016 4051 3042
rect 3959 2998 3989 3012
rect 4016 3008 4051 3016
rect 4053 3042 4094 3050
rect 4053 3016 4068 3042
rect 4075 3016 4094 3042
rect 4158 3038 4189 3050
rect 4204 3038 4307 3050
rect 4319 3040 4345 3066
rect 4360 3061 4390 3072
rect 4422 3068 4484 3084
rect 4422 3066 4468 3068
rect 4422 3050 4484 3066
rect 4496 3050 4502 3098
rect 4505 3090 4585 3098
rect 4505 3088 4524 3090
rect 4539 3088 4573 3090
rect 4505 3072 4585 3088
rect 4505 3050 4524 3072
rect 4539 3056 4569 3072
rect 4597 3066 4603 3140
rect 4606 3066 4625 3210
rect 4640 3066 4646 3210
rect 4655 3140 4668 3210
rect 4720 3206 4742 3210
rect 4713 3184 4742 3198
rect 4795 3184 4811 3198
rect 4849 3194 4855 3196
rect 4862 3194 4970 3210
rect 4977 3194 4983 3196
rect 4991 3194 5006 3210
rect 5072 3204 5091 3207
rect 4713 3182 4811 3184
rect 4838 3182 5006 3194
rect 5021 3184 5037 3198
rect 5072 3185 5094 3204
rect 5104 3198 5120 3199
rect 5103 3196 5120 3198
rect 5104 3191 5120 3196
rect 5094 3184 5100 3185
rect 5103 3184 5132 3191
rect 5021 3183 5132 3184
rect 5021 3182 5138 3183
rect 4697 3174 4748 3182
rect 4795 3174 4829 3182
rect 4697 3162 4722 3174
rect 4729 3162 4748 3174
rect 4802 3172 4829 3174
rect 4838 3172 5059 3182
rect 5094 3179 5100 3182
rect 4802 3168 5059 3172
rect 4697 3154 4748 3162
rect 4795 3154 5059 3168
rect 5103 3174 5138 3182
rect 4649 3106 4668 3140
rect 4713 3146 4742 3154
rect 4713 3140 4730 3146
rect 4713 3138 4747 3140
rect 4795 3138 4811 3154
rect 4812 3144 5020 3154
rect 5021 3144 5037 3154
rect 5085 3150 5100 3165
rect 5103 3162 5104 3174
rect 5111 3162 5138 3174
rect 5103 3154 5138 3162
rect 5103 3153 5132 3154
rect 4823 3140 5037 3144
rect 4838 3138 5037 3140
rect 5072 3140 5085 3150
rect 5103 3140 5120 3153
rect 5072 3138 5120 3140
rect 4714 3134 4747 3138
rect 4710 3132 4747 3134
rect 4710 3131 4777 3132
rect 4710 3126 4741 3131
rect 4747 3126 4777 3131
rect 4710 3122 4777 3126
rect 4683 3119 4777 3122
rect 4683 3112 4732 3119
rect 4683 3106 4713 3112
rect 4732 3107 4737 3112
rect 4649 3090 4729 3106
rect 4741 3098 4777 3119
rect 4838 3114 5027 3138
rect 5072 3137 5119 3138
rect 5085 3132 5119 3137
rect 4853 3111 5027 3114
rect 4846 3108 5027 3111
rect 5055 3131 5119 3132
rect 4649 3088 4668 3090
rect 4683 3088 4717 3090
rect 4649 3072 4729 3088
rect 4649 3066 4668 3072
rect 4365 3040 4468 3050
rect 4319 3038 4468 3040
rect 4489 3038 4524 3050
rect 4158 3036 4320 3038
rect 4170 3016 4189 3036
rect 4204 3034 4234 3036
rect 4053 3008 4094 3016
rect 4176 3012 4189 3016
rect 4241 3020 4320 3036
rect 4352 3036 4524 3038
rect 4352 3020 4431 3036
rect 4438 3034 4468 3036
rect 4016 2998 4045 3008
rect 4059 2998 4088 3008
rect 4103 2998 4133 3012
rect 4176 2998 4219 3012
rect 4241 3008 4431 3020
rect 4496 3016 4502 3036
rect 4226 2998 4256 3008
rect 4257 2998 4415 3008
rect 4419 2998 4449 3008
rect 4453 2998 4483 3012
rect 4511 2998 4524 3036
rect 4596 3050 4625 3066
rect 4639 3050 4668 3066
rect 4683 3056 4713 3072
rect 4741 3050 4747 3098
rect 4750 3092 4769 3098
rect 4784 3092 4814 3100
rect 4750 3084 4814 3092
rect 4750 3068 4830 3084
rect 4846 3077 4908 3108
rect 4924 3077 4986 3108
rect 5055 3106 5104 3131
rect 5119 3106 5149 3122
rect 5018 3092 5048 3100
rect 5055 3098 5165 3106
rect 5018 3084 5063 3092
rect 4750 3066 4769 3068
rect 4784 3066 4830 3068
rect 4750 3050 4830 3066
rect 4857 3064 4892 3077
rect 4933 3074 4970 3077
rect 4933 3072 4975 3074
rect 4862 3061 4892 3064
rect 4871 3057 4878 3061
rect 4878 3056 4879 3057
rect 4837 3050 4847 3056
rect 4596 3042 4631 3050
rect 4596 3016 4597 3042
rect 4604 3016 4631 3042
rect 4539 2998 4569 3012
rect 4596 3008 4631 3016
rect 4633 3042 4674 3050
rect 4633 3016 4648 3042
rect 4655 3016 4674 3042
rect 4738 3038 4769 3050
rect 4784 3038 4887 3050
rect 4899 3040 4925 3066
rect 4940 3061 4970 3072
rect 5002 3068 5064 3084
rect 5002 3066 5048 3068
rect 5002 3050 5064 3066
rect 5076 3050 5082 3098
rect 5085 3090 5165 3098
rect 5085 3088 5104 3090
rect 5119 3088 5153 3090
rect 5085 3072 5165 3088
rect 5085 3050 5104 3072
rect 5119 3056 5149 3072
rect 5177 3066 5183 3140
rect 5186 3066 5205 3210
rect 5220 3066 5226 3210
rect 5235 3140 5248 3210
rect 5300 3206 5322 3210
rect 5293 3184 5322 3198
rect 5375 3184 5391 3198
rect 5429 3194 5435 3196
rect 5442 3194 5550 3210
rect 5557 3194 5563 3196
rect 5571 3194 5586 3210
rect 5652 3204 5671 3207
rect 5293 3182 5391 3184
rect 5418 3182 5586 3194
rect 5601 3184 5617 3198
rect 5652 3185 5674 3204
rect 5684 3198 5700 3199
rect 5683 3196 5700 3198
rect 5684 3191 5700 3196
rect 5674 3184 5680 3185
rect 5683 3184 5712 3191
rect 5601 3183 5712 3184
rect 5601 3182 5718 3183
rect 5277 3174 5328 3182
rect 5375 3174 5409 3182
rect 5277 3162 5302 3174
rect 5309 3162 5328 3174
rect 5382 3172 5409 3174
rect 5418 3172 5639 3182
rect 5674 3179 5680 3182
rect 5382 3168 5639 3172
rect 5277 3154 5328 3162
rect 5375 3154 5639 3168
rect 5683 3174 5718 3182
rect 5229 3106 5248 3140
rect 5293 3146 5322 3154
rect 5293 3140 5310 3146
rect 5293 3138 5327 3140
rect 5375 3138 5391 3154
rect 5392 3144 5600 3154
rect 5601 3144 5617 3154
rect 5665 3150 5680 3165
rect 5683 3162 5684 3174
rect 5691 3162 5718 3174
rect 5683 3154 5718 3162
rect 5683 3153 5712 3154
rect 5403 3140 5617 3144
rect 5418 3138 5617 3140
rect 5652 3140 5665 3150
rect 5683 3140 5700 3153
rect 5652 3138 5700 3140
rect 5294 3134 5327 3138
rect 5290 3132 5327 3134
rect 5290 3131 5357 3132
rect 5290 3126 5321 3131
rect 5327 3126 5357 3131
rect 5290 3122 5357 3126
rect 5263 3119 5357 3122
rect 5263 3112 5312 3119
rect 5263 3106 5293 3112
rect 5312 3107 5317 3112
rect 5229 3090 5309 3106
rect 5321 3098 5357 3119
rect 5418 3114 5607 3138
rect 5652 3137 5699 3138
rect 5665 3132 5699 3137
rect 5433 3111 5607 3114
rect 5426 3108 5607 3111
rect 5635 3131 5699 3132
rect 5229 3088 5248 3090
rect 5263 3088 5297 3090
rect 5229 3072 5309 3088
rect 5229 3066 5248 3072
rect 4945 3040 5048 3050
rect 4899 3038 5048 3040
rect 5069 3038 5104 3050
rect 4738 3036 4900 3038
rect 4750 3016 4769 3036
rect 4784 3034 4814 3036
rect 4633 3008 4674 3016
rect 4756 3012 4769 3016
rect 4821 3020 4900 3036
rect 4932 3036 5104 3038
rect 4932 3020 5011 3036
rect 5018 3034 5048 3036
rect 4596 2998 4625 3008
rect 4639 2998 4668 3008
rect 4683 2998 4713 3012
rect 4756 2998 4799 3012
rect 4821 3008 5011 3020
rect 5076 3016 5082 3036
rect 4806 2998 4836 3008
rect 4837 2998 4995 3008
rect 4999 2998 5029 3008
rect 5033 2998 5063 3012
rect 5091 2998 5104 3036
rect 5176 3050 5205 3066
rect 5219 3050 5248 3066
rect 5263 3056 5293 3072
rect 5321 3050 5327 3098
rect 5330 3092 5349 3098
rect 5364 3092 5394 3100
rect 5330 3084 5394 3092
rect 5330 3068 5410 3084
rect 5426 3077 5488 3108
rect 5504 3077 5566 3108
rect 5635 3106 5684 3131
rect 5699 3106 5729 3122
rect 5598 3092 5628 3100
rect 5635 3098 5745 3106
rect 5598 3084 5643 3092
rect 5330 3066 5349 3068
rect 5364 3066 5410 3068
rect 5330 3050 5410 3066
rect 5437 3064 5472 3077
rect 5513 3074 5550 3077
rect 5513 3072 5555 3074
rect 5442 3061 5472 3064
rect 5451 3057 5458 3061
rect 5458 3056 5459 3057
rect 5417 3050 5427 3056
rect 5176 3042 5211 3050
rect 5176 3016 5177 3042
rect 5184 3016 5211 3042
rect 5119 2998 5149 3012
rect 5176 3008 5211 3016
rect 5213 3042 5254 3050
rect 5213 3016 5228 3042
rect 5235 3016 5254 3042
rect 5318 3038 5349 3050
rect 5364 3038 5467 3050
rect 5479 3040 5505 3066
rect 5520 3061 5550 3072
rect 5582 3068 5644 3084
rect 5582 3066 5628 3068
rect 5582 3050 5644 3066
rect 5656 3050 5662 3098
rect 5665 3090 5745 3098
rect 5665 3088 5684 3090
rect 5699 3088 5733 3090
rect 5665 3072 5745 3088
rect 5665 3050 5684 3072
rect 5699 3056 5729 3072
rect 5757 3066 5763 3140
rect 5766 3066 5785 3210
rect 5800 3066 5806 3210
rect 5815 3140 5828 3210
rect 5880 3206 5902 3210
rect 5873 3184 5902 3198
rect 5955 3184 5971 3198
rect 6009 3194 6015 3196
rect 6022 3194 6130 3210
rect 6137 3194 6143 3196
rect 6151 3194 6166 3210
rect 6232 3204 6251 3207
rect 5873 3182 5971 3184
rect 5998 3182 6166 3194
rect 6181 3184 6197 3198
rect 6232 3185 6254 3204
rect 6264 3198 6280 3199
rect 6263 3196 6280 3198
rect 6264 3191 6280 3196
rect 6254 3184 6260 3185
rect 6263 3184 6292 3191
rect 6181 3183 6292 3184
rect 6181 3182 6298 3183
rect 5857 3174 5908 3182
rect 5955 3174 5989 3182
rect 5857 3162 5882 3174
rect 5889 3162 5908 3174
rect 5962 3172 5989 3174
rect 5998 3172 6219 3182
rect 6254 3179 6260 3182
rect 5962 3168 6219 3172
rect 5857 3154 5908 3162
rect 5955 3154 6219 3168
rect 6263 3174 6298 3182
rect 5809 3106 5828 3140
rect 5873 3146 5902 3154
rect 5873 3140 5890 3146
rect 5873 3138 5907 3140
rect 5955 3138 5971 3154
rect 5972 3144 6180 3154
rect 6181 3144 6197 3154
rect 6245 3150 6260 3165
rect 6263 3162 6264 3174
rect 6271 3162 6298 3174
rect 6263 3154 6298 3162
rect 6263 3153 6292 3154
rect 5983 3140 6197 3144
rect 5998 3138 6197 3140
rect 6232 3140 6245 3150
rect 6263 3140 6280 3153
rect 6232 3138 6280 3140
rect 5874 3134 5907 3138
rect 5870 3132 5907 3134
rect 5870 3131 5937 3132
rect 5870 3126 5901 3131
rect 5907 3126 5937 3131
rect 5870 3122 5937 3126
rect 5843 3119 5937 3122
rect 5843 3112 5892 3119
rect 5843 3106 5873 3112
rect 5892 3107 5897 3112
rect 5809 3090 5889 3106
rect 5901 3098 5937 3119
rect 5998 3114 6187 3138
rect 6232 3137 6279 3138
rect 6245 3132 6279 3137
rect 6013 3111 6187 3114
rect 6006 3108 6187 3111
rect 6215 3131 6279 3132
rect 5809 3088 5828 3090
rect 5843 3088 5877 3090
rect 5809 3072 5889 3088
rect 5809 3066 5828 3072
rect 5525 3040 5628 3050
rect 5479 3038 5628 3040
rect 5649 3038 5684 3050
rect 5318 3036 5480 3038
rect 5330 3016 5349 3036
rect 5364 3034 5394 3036
rect 5213 3008 5254 3016
rect 5336 3012 5349 3016
rect 5401 3020 5480 3036
rect 5512 3036 5684 3038
rect 5512 3020 5591 3036
rect 5598 3034 5628 3036
rect 5176 2998 5205 3008
rect 5219 2998 5248 3008
rect 5263 2998 5293 3012
rect 5336 2998 5379 3012
rect 5401 3008 5591 3020
rect 5656 3016 5662 3036
rect 5386 2998 5416 3008
rect 5417 2998 5575 3008
rect 5579 2998 5609 3008
rect 5613 2998 5643 3012
rect 5671 2998 5684 3036
rect 5756 3050 5785 3066
rect 5799 3050 5828 3066
rect 5843 3056 5873 3072
rect 5901 3050 5907 3098
rect 5910 3092 5929 3098
rect 5944 3092 5974 3100
rect 5910 3084 5974 3092
rect 5910 3068 5990 3084
rect 6006 3077 6068 3108
rect 6084 3077 6146 3108
rect 6215 3106 6264 3131
rect 6279 3106 6309 3122
rect 6178 3092 6208 3100
rect 6215 3098 6325 3106
rect 6178 3084 6223 3092
rect 5910 3066 5929 3068
rect 5944 3066 5990 3068
rect 5910 3050 5990 3066
rect 6017 3064 6052 3077
rect 6093 3074 6130 3077
rect 6093 3072 6135 3074
rect 6022 3061 6052 3064
rect 6031 3057 6038 3061
rect 6038 3056 6039 3057
rect 5997 3050 6007 3056
rect 5756 3042 5791 3050
rect 5756 3016 5757 3042
rect 5764 3016 5791 3042
rect 5699 2998 5729 3012
rect 5756 3008 5791 3016
rect 5793 3042 5834 3050
rect 5793 3016 5808 3042
rect 5815 3016 5834 3042
rect 5898 3038 5929 3050
rect 5944 3038 6047 3050
rect 6059 3040 6085 3066
rect 6100 3061 6130 3072
rect 6162 3068 6224 3084
rect 6162 3066 6208 3068
rect 6162 3050 6224 3066
rect 6236 3050 6242 3098
rect 6245 3090 6325 3098
rect 6245 3088 6264 3090
rect 6279 3088 6313 3090
rect 6245 3072 6325 3088
rect 6245 3050 6264 3072
rect 6279 3056 6309 3072
rect 6337 3066 6343 3140
rect 6346 3066 6365 3210
rect 6380 3066 6386 3210
rect 6395 3140 6408 3210
rect 6460 3206 6482 3210
rect 6453 3184 6482 3198
rect 6535 3184 6551 3198
rect 6589 3194 6595 3196
rect 6602 3194 6710 3210
rect 6717 3194 6723 3196
rect 6731 3194 6746 3210
rect 6812 3204 6831 3207
rect 6453 3182 6551 3184
rect 6578 3182 6746 3194
rect 6761 3184 6777 3198
rect 6812 3185 6834 3204
rect 6844 3198 6860 3199
rect 6843 3196 6860 3198
rect 6844 3191 6860 3196
rect 6834 3184 6840 3185
rect 6843 3184 6872 3191
rect 6761 3183 6872 3184
rect 6761 3182 6878 3183
rect 6437 3174 6488 3182
rect 6535 3174 6569 3182
rect 6437 3162 6462 3174
rect 6469 3162 6488 3174
rect 6542 3172 6569 3174
rect 6578 3172 6799 3182
rect 6834 3179 6840 3182
rect 6542 3168 6799 3172
rect 6437 3154 6488 3162
rect 6535 3154 6799 3168
rect 6843 3174 6878 3182
rect 6389 3106 6408 3140
rect 6453 3146 6482 3154
rect 6453 3140 6470 3146
rect 6453 3138 6487 3140
rect 6535 3138 6551 3154
rect 6552 3144 6760 3154
rect 6761 3144 6777 3154
rect 6825 3150 6840 3165
rect 6843 3162 6844 3174
rect 6851 3162 6878 3174
rect 6843 3154 6878 3162
rect 6843 3153 6872 3154
rect 6563 3140 6777 3144
rect 6578 3138 6777 3140
rect 6812 3140 6825 3150
rect 6843 3140 6860 3153
rect 6812 3138 6860 3140
rect 6454 3134 6487 3138
rect 6450 3132 6487 3134
rect 6450 3131 6517 3132
rect 6450 3126 6481 3131
rect 6487 3126 6517 3131
rect 6450 3122 6517 3126
rect 6423 3119 6517 3122
rect 6423 3112 6472 3119
rect 6423 3106 6453 3112
rect 6472 3107 6477 3112
rect 6389 3090 6469 3106
rect 6481 3098 6517 3119
rect 6578 3114 6767 3138
rect 6812 3137 6859 3138
rect 6825 3132 6859 3137
rect 6593 3111 6767 3114
rect 6586 3108 6767 3111
rect 6795 3131 6859 3132
rect 6389 3088 6408 3090
rect 6423 3088 6457 3090
rect 6389 3072 6469 3088
rect 6389 3066 6408 3072
rect 6105 3040 6208 3050
rect 6059 3038 6208 3040
rect 6229 3038 6264 3050
rect 5898 3036 6060 3038
rect 5910 3016 5929 3036
rect 5944 3034 5974 3036
rect 5793 3008 5834 3016
rect 5916 3012 5929 3016
rect 5981 3020 6060 3036
rect 6092 3036 6264 3038
rect 6092 3020 6171 3036
rect 6178 3034 6208 3036
rect 5756 2998 5785 3008
rect 5799 2998 5828 3008
rect 5843 2998 5873 3012
rect 5916 2998 5959 3012
rect 5981 3008 6171 3020
rect 6236 3016 6242 3036
rect 5966 2998 5996 3008
rect 5997 2998 6155 3008
rect 6159 2998 6189 3008
rect 6193 2998 6223 3012
rect 6251 2998 6264 3036
rect 6336 3050 6365 3066
rect 6379 3050 6408 3066
rect 6423 3056 6453 3072
rect 6481 3050 6487 3098
rect 6490 3092 6509 3098
rect 6524 3092 6554 3100
rect 6490 3084 6554 3092
rect 6490 3068 6570 3084
rect 6586 3077 6648 3108
rect 6664 3077 6726 3108
rect 6795 3106 6844 3131
rect 6859 3106 6889 3122
rect 6758 3092 6788 3100
rect 6795 3098 6905 3106
rect 6758 3084 6803 3092
rect 6490 3066 6509 3068
rect 6524 3066 6570 3068
rect 6490 3050 6570 3066
rect 6597 3064 6632 3077
rect 6673 3074 6710 3077
rect 6673 3072 6715 3074
rect 6602 3061 6632 3064
rect 6611 3057 6618 3061
rect 6618 3056 6619 3057
rect 6577 3050 6587 3056
rect 6336 3042 6371 3050
rect 6336 3016 6337 3042
rect 6344 3016 6371 3042
rect 6279 2998 6309 3012
rect 6336 3008 6371 3016
rect 6373 3042 6414 3050
rect 6373 3016 6388 3042
rect 6395 3016 6414 3042
rect 6478 3038 6509 3050
rect 6524 3038 6627 3050
rect 6639 3040 6665 3066
rect 6680 3061 6710 3072
rect 6742 3068 6804 3084
rect 6742 3066 6788 3068
rect 6742 3050 6804 3066
rect 6816 3050 6822 3098
rect 6825 3090 6905 3098
rect 6825 3088 6844 3090
rect 6859 3088 6893 3090
rect 6825 3072 6905 3088
rect 6825 3050 6844 3072
rect 6859 3056 6889 3072
rect 6917 3066 6923 3140
rect 6926 3066 6945 3210
rect 6960 3066 6966 3210
rect 6975 3140 6988 3210
rect 7040 3206 7062 3210
rect 7033 3184 7062 3198
rect 7115 3184 7131 3198
rect 7169 3194 7175 3196
rect 7182 3194 7290 3210
rect 7297 3194 7303 3196
rect 7311 3194 7326 3210
rect 7392 3204 7411 3207
rect 7033 3182 7131 3184
rect 7158 3182 7326 3194
rect 7341 3184 7357 3198
rect 7392 3185 7414 3204
rect 7424 3198 7440 3199
rect 7423 3196 7440 3198
rect 7424 3191 7440 3196
rect 7414 3184 7420 3185
rect 7423 3184 7452 3191
rect 7341 3183 7452 3184
rect 7341 3182 7458 3183
rect 7017 3174 7068 3182
rect 7115 3174 7149 3182
rect 7017 3162 7042 3174
rect 7049 3162 7068 3174
rect 7122 3172 7149 3174
rect 7158 3172 7379 3182
rect 7414 3179 7420 3182
rect 7122 3168 7379 3172
rect 7017 3154 7068 3162
rect 7115 3154 7379 3168
rect 7423 3174 7458 3182
rect 6969 3106 6988 3140
rect 7033 3146 7062 3154
rect 7033 3140 7050 3146
rect 7033 3138 7067 3140
rect 7115 3138 7131 3154
rect 7132 3144 7340 3154
rect 7341 3144 7357 3154
rect 7405 3150 7420 3165
rect 7423 3162 7424 3174
rect 7431 3162 7458 3174
rect 7423 3154 7458 3162
rect 7423 3153 7452 3154
rect 7143 3140 7357 3144
rect 7158 3138 7357 3140
rect 7392 3140 7405 3150
rect 7423 3140 7440 3153
rect 7392 3138 7440 3140
rect 7034 3134 7067 3138
rect 7030 3132 7067 3134
rect 7030 3131 7097 3132
rect 7030 3126 7061 3131
rect 7067 3126 7097 3131
rect 7030 3122 7097 3126
rect 7003 3119 7097 3122
rect 7003 3112 7052 3119
rect 7003 3106 7033 3112
rect 7052 3107 7057 3112
rect 6969 3090 7049 3106
rect 7061 3098 7097 3119
rect 7158 3114 7347 3138
rect 7392 3137 7439 3138
rect 7405 3132 7439 3137
rect 7173 3111 7347 3114
rect 7166 3108 7347 3111
rect 7375 3131 7439 3132
rect 6969 3088 6988 3090
rect 7003 3088 7037 3090
rect 6969 3072 7049 3088
rect 6969 3066 6988 3072
rect 6685 3040 6788 3050
rect 6639 3038 6788 3040
rect 6809 3038 6844 3050
rect 6478 3036 6640 3038
rect 6490 3016 6509 3036
rect 6524 3034 6554 3036
rect 6373 3008 6414 3016
rect 6496 3012 6509 3016
rect 6561 3020 6640 3036
rect 6672 3036 6844 3038
rect 6672 3020 6751 3036
rect 6758 3034 6788 3036
rect 6336 2998 6365 3008
rect 6379 2998 6408 3008
rect 6423 2998 6453 3012
rect 6496 2998 6539 3012
rect 6561 3008 6751 3020
rect 6816 3016 6822 3036
rect 6546 2998 6576 3008
rect 6577 2998 6735 3008
rect 6739 2998 6769 3008
rect 6773 2998 6803 3012
rect 6831 2998 6844 3036
rect 6916 3050 6945 3066
rect 6959 3050 6988 3066
rect 7003 3056 7033 3072
rect 7061 3050 7067 3098
rect 7070 3092 7089 3098
rect 7104 3092 7134 3100
rect 7070 3084 7134 3092
rect 7070 3068 7150 3084
rect 7166 3077 7228 3108
rect 7244 3077 7306 3108
rect 7375 3106 7424 3131
rect 7439 3106 7469 3122
rect 7338 3092 7368 3100
rect 7375 3098 7485 3106
rect 7338 3084 7383 3092
rect 7070 3066 7089 3068
rect 7104 3066 7150 3068
rect 7070 3050 7150 3066
rect 7177 3064 7212 3077
rect 7253 3074 7290 3077
rect 7253 3072 7295 3074
rect 7182 3061 7212 3064
rect 7191 3057 7198 3061
rect 7198 3056 7199 3057
rect 7157 3050 7167 3056
rect 6916 3042 6951 3050
rect 6916 3016 6917 3042
rect 6924 3016 6951 3042
rect 6859 2998 6889 3012
rect 6916 3008 6951 3016
rect 6953 3042 6994 3050
rect 6953 3016 6968 3042
rect 6975 3016 6994 3042
rect 7058 3038 7089 3050
rect 7104 3038 7207 3050
rect 7219 3040 7245 3066
rect 7260 3061 7290 3072
rect 7322 3068 7384 3084
rect 7322 3066 7368 3068
rect 7322 3050 7384 3066
rect 7396 3050 7402 3098
rect 7405 3090 7485 3098
rect 7405 3088 7424 3090
rect 7439 3088 7473 3090
rect 7405 3072 7485 3088
rect 7405 3050 7424 3072
rect 7439 3056 7469 3072
rect 7497 3066 7503 3140
rect 7506 3066 7525 3210
rect 7540 3066 7546 3210
rect 7555 3140 7568 3210
rect 7620 3206 7642 3210
rect 7613 3184 7642 3198
rect 7695 3184 7711 3198
rect 7749 3194 7755 3196
rect 7762 3194 7870 3210
rect 7877 3194 7883 3196
rect 7891 3194 7906 3210
rect 7972 3204 7991 3207
rect 7613 3182 7711 3184
rect 7738 3182 7906 3194
rect 7921 3184 7937 3198
rect 7972 3185 7994 3204
rect 8004 3198 8020 3199
rect 8003 3196 8020 3198
rect 8004 3191 8020 3196
rect 7994 3184 8000 3185
rect 8003 3184 8032 3191
rect 7921 3183 8032 3184
rect 7921 3182 8038 3183
rect 7597 3174 7648 3182
rect 7695 3174 7729 3182
rect 7597 3162 7622 3174
rect 7629 3162 7648 3174
rect 7702 3172 7729 3174
rect 7738 3172 7959 3182
rect 7994 3179 8000 3182
rect 7702 3168 7959 3172
rect 7597 3154 7648 3162
rect 7695 3154 7959 3168
rect 8003 3174 8038 3182
rect 7549 3106 7568 3140
rect 7613 3146 7642 3154
rect 7613 3140 7630 3146
rect 7613 3138 7647 3140
rect 7695 3138 7711 3154
rect 7712 3144 7920 3154
rect 7921 3144 7937 3154
rect 7985 3150 8000 3165
rect 8003 3162 8004 3174
rect 8011 3162 8038 3174
rect 8003 3154 8038 3162
rect 8003 3153 8032 3154
rect 7723 3140 7937 3144
rect 7738 3138 7937 3140
rect 7972 3140 7985 3150
rect 8003 3140 8020 3153
rect 7972 3138 8020 3140
rect 7614 3134 7647 3138
rect 7610 3132 7647 3134
rect 7610 3131 7677 3132
rect 7610 3126 7641 3131
rect 7647 3126 7677 3131
rect 7610 3122 7677 3126
rect 7583 3119 7677 3122
rect 7583 3112 7632 3119
rect 7583 3106 7613 3112
rect 7632 3107 7637 3112
rect 7549 3090 7629 3106
rect 7641 3098 7677 3119
rect 7738 3114 7927 3138
rect 7972 3137 8019 3138
rect 7985 3132 8019 3137
rect 7753 3111 7927 3114
rect 7746 3108 7927 3111
rect 7955 3131 8019 3132
rect 7549 3088 7568 3090
rect 7583 3088 7617 3090
rect 7549 3072 7629 3088
rect 7549 3066 7568 3072
rect 7265 3040 7368 3050
rect 7219 3038 7368 3040
rect 7389 3038 7424 3050
rect 7058 3036 7220 3038
rect 7070 3016 7089 3036
rect 7104 3034 7134 3036
rect 6953 3008 6994 3016
rect 7076 3012 7089 3016
rect 7141 3020 7220 3036
rect 7252 3036 7424 3038
rect 7252 3020 7331 3036
rect 7338 3034 7368 3036
rect 6916 2998 6945 3008
rect 6959 2998 6988 3008
rect 7003 2998 7033 3012
rect 7076 2998 7119 3012
rect 7141 3008 7331 3020
rect 7396 3016 7402 3036
rect 7126 2998 7156 3008
rect 7157 2998 7315 3008
rect 7319 2998 7349 3008
rect 7353 2998 7383 3012
rect 7411 2998 7424 3036
rect 7496 3050 7525 3066
rect 7539 3050 7568 3066
rect 7583 3056 7613 3072
rect 7641 3050 7647 3098
rect 7650 3092 7669 3098
rect 7684 3092 7714 3100
rect 7650 3084 7714 3092
rect 7650 3068 7730 3084
rect 7746 3077 7808 3108
rect 7824 3077 7886 3108
rect 7955 3106 8004 3131
rect 8019 3106 8049 3122
rect 7918 3092 7948 3100
rect 7955 3098 8065 3106
rect 7918 3084 7963 3092
rect 7650 3066 7669 3068
rect 7684 3066 7730 3068
rect 7650 3050 7730 3066
rect 7757 3064 7792 3077
rect 7833 3074 7870 3077
rect 7833 3072 7875 3074
rect 7762 3061 7792 3064
rect 7771 3057 7778 3061
rect 7778 3056 7779 3057
rect 7737 3050 7747 3056
rect 7496 3042 7531 3050
rect 7496 3016 7497 3042
rect 7504 3016 7531 3042
rect 7439 2998 7469 3012
rect 7496 3008 7531 3016
rect 7533 3042 7574 3050
rect 7533 3016 7548 3042
rect 7555 3016 7574 3042
rect 7638 3038 7669 3050
rect 7684 3038 7787 3050
rect 7799 3040 7825 3066
rect 7840 3061 7870 3072
rect 7902 3068 7964 3084
rect 7902 3066 7948 3068
rect 7902 3050 7964 3066
rect 7976 3050 7982 3098
rect 7985 3090 8065 3098
rect 7985 3088 8004 3090
rect 8019 3088 8053 3090
rect 7985 3072 8065 3088
rect 7985 3050 8004 3072
rect 8019 3056 8049 3072
rect 8077 3066 8083 3140
rect 8086 3066 8105 3210
rect 8120 3066 8126 3210
rect 8135 3140 8148 3210
rect 8200 3206 8222 3210
rect 8193 3184 8222 3198
rect 8275 3184 8291 3198
rect 8329 3194 8335 3196
rect 8342 3194 8450 3210
rect 8457 3194 8463 3196
rect 8471 3194 8486 3210
rect 8552 3204 8571 3207
rect 8193 3182 8291 3184
rect 8318 3182 8486 3194
rect 8501 3184 8517 3198
rect 8552 3185 8574 3204
rect 8584 3198 8600 3199
rect 8583 3196 8600 3198
rect 8584 3191 8600 3196
rect 8574 3184 8580 3185
rect 8583 3184 8612 3191
rect 8501 3183 8612 3184
rect 8501 3182 8618 3183
rect 8177 3174 8228 3182
rect 8275 3174 8309 3182
rect 8177 3162 8202 3174
rect 8209 3162 8228 3174
rect 8282 3172 8309 3174
rect 8318 3172 8539 3182
rect 8574 3179 8580 3182
rect 8282 3168 8539 3172
rect 8177 3154 8228 3162
rect 8275 3154 8539 3168
rect 8583 3174 8618 3182
rect 8129 3106 8148 3140
rect 8193 3146 8222 3154
rect 8193 3140 8210 3146
rect 8193 3138 8227 3140
rect 8275 3138 8291 3154
rect 8292 3144 8500 3154
rect 8501 3144 8517 3154
rect 8565 3150 8580 3165
rect 8583 3162 8584 3174
rect 8591 3162 8618 3174
rect 8583 3154 8618 3162
rect 8583 3153 8612 3154
rect 8303 3140 8517 3144
rect 8318 3138 8517 3140
rect 8552 3140 8565 3150
rect 8583 3140 8600 3153
rect 8552 3138 8600 3140
rect 8194 3134 8227 3138
rect 8190 3132 8227 3134
rect 8190 3131 8257 3132
rect 8190 3126 8221 3131
rect 8227 3126 8257 3131
rect 8190 3122 8257 3126
rect 8163 3119 8257 3122
rect 8163 3112 8212 3119
rect 8163 3106 8193 3112
rect 8212 3107 8217 3112
rect 8129 3090 8209 3106
rect 8221 3098 8257 3119
rect 8318 3114 8507 3138
rect 8552 3137 8599 3138
rect 8565 3132 8599 3137
rect 8333 3111 8507 3114
rect 8326 3108 8507 3111
rect 8535 3131 8599 3132
rect 8129 3088 8148 3090
rect 8163 3088 8197 3090
rect 8129 3072 8209 3088
rect 8129 3066 8148 3072
rect 7845 3040 7948 3050
rect 7799 3038 7948 3040
rect 7969 3038 8004 3050
rect 7638 3036 7800 3038
rect 7650 3016 7669 3036
rect 7684 3034 7714 3036
rect 7533 3008 7574 3016
rect 7656 3012 7669 3016
rect 7721 3020 7800 3036
rect 7832 3036 8004 3038
rect 7832 3020 7911 3036
rect 7918 3034 7948 3036
rect 7496 2998 7525 3008
rect 7539 2998 7568 3008
rect 7583 2998 7613 3012
rect 7656 2998 7699 3012
rect 7721 3008 7911 3020
rect 7976 3016 7982 3036
rect 7706 2998 7736 3008
rect 7737 2998 7895 3008
rect 7899 2998 7929 3008
rect 7933 2998 7963 3012
rect 7991 2998 8004 3036
rect 8076 3050 8105 3066
rect 8119 3050 8148 3066
rect 8163 3056 8193 3072
rect 8221 3050 8227 3098
rect 8230 3092 8249 3098
rect 8264 3092 8294 3100
rect 8230 3084 8294 3092
rect 8230 3068 8310 3084
rect 8326 3077 8388 3108
rect 8404 3077 8466 3108
rect 8535 3106 8584 3131
rect 8599 3106 8629 3122
rect 8498 3092 8528 3100
rect 8535 3098 8645 3106
rect 8498 3084 8543 3092
rect 8230 3066 8249 3068
rect 8264 3066 8310 3068
rect 8230 3050 8310 3066
rect 8337 3064 8372 3077
rect 8413 3074 8450 3077
rect 8413 3072 8455 3074
rect 8342 3061 8372 3064
rect 8351 3057 8358 3061
rect 8358 3056 8359 3057
rect 8317 3050 8327 3056
rect 8076 3042 8111 3050
rect 8076 3016 8077 3042
rect 8084 3016 8111 3042
rect 8019 2998 8049 3012
rect 8076 3008 8111 3016
rect 8113 3042 8154 3050
rect 8113 3016 8128 3042
rect 8135 3016 8154 3042
rect 8218 3038 8249 3050
rect 8264 3038 8367 3050
rect 8379 3040 8405 3066
rect 8420 3061 8450 3072
rect 8482 3068 8544 3084
rect 8482 3066 8528 3068
rect 8482 3050 8544 3066
rect 8556 3050 8562 3098
rect 8565 3090 8645 3098
rect 8565 3088 8584 3090
rect 8599 3088 8633 3090
rect 8565 3072 8645 3088
rect 8565 3050 8584 3072
rect 8599 3056 8629 3072
rect 8657 3066 8663 3140
rect 8666 3066 8685 3210
rect 8700 3066 8706 3210
rect 8715 3140 8728 3210
rect 8780 3206 8802 3210
rect 8773 3184 8802 3198
rect 8855 3184 8871 3198
rect 8909 3194 8915 3196
rect 8922 3194 9030 3210
rect 9037 3194 9043 3196
rect 9051 3194 9066 3210
rect 9132 3204 9151 3207
rect 8773 3182 8871 3184
rect 8898 3182 9066 3194
rect 9081 3184 9097 3198
rect 9132 3185 9154 3204
rect 9164 3198 9180 3199
rect 9163 3196 9180 3198
rect 9164 3191 9180 3196
rect 9154 3184 9160 3185
rect 9163 3184 9192 3191
rect 9081 3183 9192 3184
rect 9081 3182 9198 3183
rect 8757 3174 8808 3182
rect 8855 3174 8889 3182
rect 8757 3162 8782 3174
rect 8789 3162 8808 3174
rect 8862 3172 8889 3174
rect 8898 3172 9119 3182
rect 9154 3179 9160 3182
rect 8862 3168 9119 3172
rect 8757 3154 8808 3162
rect 8855 3154 9119 3168
rect 9163 3174 9198 3182
rect 8709 3106 8728 3140
rect 8773 3146 8802 3154
rect 8773 3140 8790 3146
rect 8773 3138 8807 3140
rect 8855 3138 8871 3154
rect 8872 3144 9080 3154
rect 9081 3144 9097 3154
rect 9145 3150 9160 3165
rect 9163 3162 9164 3174
rect 9171 3162 9198 3174
rect 9163 3154 9198 3162
rect 9163 3153 9192 3154
rect 8883 3140 9097 3144
rect 8898 3138 9097 3140
rect 9132 3140 9145 3150
rect 9163 3140 9180 3153
rect 9132 3138 9180 3140
rect 8774 3134 8807 3138
rect 8770 3132 8807 3134
rect 8770 3131 8837 3132
rect 8770 3126 8801 3131
rect 8807 3126 8837 3131
rect 8770 3122 8837 3126
rect 8743 3119 8837 3122
rect 8743 3112 8792 3119
rect 8743 3106 8773 3112
rect 8792 3107 8797 3112
rect 8709 3090 8789 3106
rect 8801 3098 8837 3119
rect 8898 3114 9087 3138
rect 9132 3137 9179 3138
rect 9145 3132 9179 3137
rect 8913 3111 9087 3114
rect 8906 3108 9087 3111
rect 9115 3131 9179 3132
rect 8709 3088 8728 3090
rect 8743 3088 8777 3090
rect 8709 3072 8789 3088
rect 8709 3066 8728 3072
rect 8425 3040 8528 3050
rect 8379 3038 8528 3040
rect 8549 3038 8584 3050
rect 8218 3036 8380 3038
rect 8230 3016 8249 3036
rect 8264 3034 8294 3036
rect 8113 3008 8154 3016
rect 8236 3012 8249 3016
rect 8301 3020 8380 3036
rect 8412 3036 8584 3038
rect 8412 3020 8491 3036
rect 8498 3034 8528 3036
rect 8076 2998 8105 3008
rect 8119 2998 8148 3008
rect 8163 2998 8193 3012
rect 8236 2998 8279 3012
rect 8301 3008 8491 3020
rect 8556 3016 8562 3036
rect 8286 2998 8316 3008
rect 8317 2998 8475 3008
rect 8479 2998 8509 3008
rect 8513 2998 8543 3012
rect 8571 2998 8584 3036
rect 8656 3050 8685 3066
rect 8699 3050 8728 3066
rect 8743 3056 8773 3072
rect 8801 3050 8807 3098
rect 8810 3092 8829 3098
rect 8844 3092 8874 3100
rect 8810 3084 8874 3092
rect 8810 3068 8890 3084
rect 8906 3077 8968 3108
rect 8984 3077 9046 3108
rect 9115 3106 9164 3131
rect 9179 3106 9209 3122
rect 9078 3092 9108 3100
rect 9115 3098 9225 3106
rect 9078 3084 9123 3092
rect 8810 3066 8829 3068
rect 8844 3066 8890 3068
rect 8810 3050 8890 3066
rect 8917 3064 8952 3077
rect 8993 3074 9030 3077
rect 8993 3072 9035 3074
rect 8922 3061 8952 3064
rect 8931 3057 8938 3061
rect 8938 3056 8939 3057
rect 8897 3050 8907 3056
rect 8656 3042 8691 3050
rect 8656 3016 8657 3042
rect 8664 3016 8691 3042
rect 8599 2998 8629 3012
rect 8656 3008 8691 3016
rect 8693 3042 8734 3050
rect 8693 3016 8708 3042
rect 8715 3016 8734 3042
rect 8798 3038 8829 3050
rect 8844 3038 8947 3050
rect 8959 3040 8985 3066
rect 9000 3061 9030 3072
rect 9062 3068 9124 3084
rect 9062 3066 9108 3068
rect 9062 3050 9124 3066
rect 9136 3050 9142 3098
rect 9145 3090 9225 3098
rect 9145 3088 9164 3090
rect 9179 3088 9213 3090
rect 9145 3072 9225 3088
rect 9145 3050 9164 3072
rect 9179 3056 9209 3072
rect 9237 3066 9243 3140
rect 9246 3066 9265 3210
rect 9280 3066 9286 3210
rect 9295 3140 9308 3210
rect 9360 3206 9382 3210
rect 9353 3184 9382 3198
rect 9435 3184 9451 3198
rect 9489 3194 9495 3196
rect 9502 3194 9610 3210
rect 9617 3194 9623 3196
rect 9631 3194 9646 3210
rect 9712 3204 9731 3207
rect 9353 3182 9451 3184
rect 9478 3182 9646 3194
rect 9661 3184 9677 3198
rect 9712 3185 9734 3204
rect 9744 3198 9760 3199
rect 9743 3196 9760 3198
rect 9744 3191 9760 3196
rect 9734 3184 9740 3185
rect 9743 3184 9772 3191
rect 9661 3183 9772 3184
rect 9661 3182 9778 3183
rect 9337 3174 9388 3182
rect 9435 3174 9469 3182
rect 9337 3162 9362 3174
rect 9369 3162 9388 3174
rect 9442 3172 9469 3174
rect 9478 3172 9699 3182
rect 9734 3179 9740 3182
rect 9442 3168 9699 3172
rect 9337 3154 9388 3162
rect 9435 3154 9699 3168
rect 9743 3174 9778 3182
rect 9289 3106 9308 3140
rect 9353 3146 9382 3154
rect 9353 3140 9370 3146
rect 9353 3138 9387 3140
rect 9435 3138 9451 3154
rect 9452 3144 9660 3154
rect 9661 3144 9677 3154
rect 9725 3150 9740 3165
rect 9743 3162 9744 3174
rect 9751 3162 9778 3174
rect 9743 3154 9778 3162
rect 9743 3153 9772 3154
rect 9463 3140 9677 3144
rect 9478 3138 9677 3140
rect 9712 3140 9725 3150
rect 9743 3140 9760 3153
rect 9712 3138 9760 3140
rect 9354 3134 9387 3138
rect 9350 3132 9387 3134
rect 9350 3131 9417 3132
rect 9350 3126 9381 3131
rect 9387 3126 9417 3131
rect 9350 3122 9417 3126
rect 9323 3119 9417 3122
rect 9323 3112 9372 3119
rect 9323 3106 9353 3112
rect 9372 3107 9377 3112
rect 9289 3090 9369 3106
rect 9381 3098 9417 3119
rect 9478 3114 9667 3138
rect 9712 3137 9759 3138
rect 9725 3132 9759 3137
rect 9493 3111 9667 3114
rect 9486 3108 9667 3111
rect 9695 3131 9759 3132
rect 9289 3088 9308 3090
rect 9323 3088 9357 3090
rect 9289 3072 9369 3088
rect 9289 3066 9308 3072
rect 9005 3040 9108 3050
rect 8959 3038 9108 3040
rect 9129 3038 9164 3050
rect 8798 3036 8960 3038
rect 8810 3016 8829 3036
rect 8844 3034 8874 3036
rect 8693 3008 8734 3016
rect 8816 3012 8829 3016
rect 8881 3020 8960 3036
rect 8992 3036 9164 3038
rect 8992 3020 9071 3036
rect 9078 3034 9108 3036
rect 8656 2998 8685 3008
rect 8699 2998 8728 3008
rect 8743 2998 8773 3012
rect 8816 2998 8859 3012
rect 8881 3008 9071 3020
rect 9136 3016 9142 3036
rect 8866 2998 8896 3008
rect 8897 2998 9055 3008
rect 9059 2998 9089 3008
rect 9093 2998 9123 3012
rect 9151 2998 9164 3036
rect 9236 3050 9265 3066
rect 9279 3050 9308 3066
rect 9323 3056 9353 3072
rect 9381 3050 9387 3098
rect 9390 3092 9409 3098
rect 9424 3092 9454 3100
rect 9390 3084 9454 3092
rect 9390 3068 9470 3084
rect 9486 3077 9548 3108
rect 9564 3077 9626 3108
rect 9695 3106 9744 3131
rect 9759 3106 9789 3122
rect 9658 3092 9688 3100
rect 9695 3098 9805 3106
rect 9658 3084 9703 3092
rect 9390 3066 9409 3068
rect 9424 3066 9470 3068
rect 9390 3050 9470 3066
rect 9497 3064 9532 3077
rect 9573 3074 9610 3077
rect 9573 3072 9615 3074
rect 9502 3061 9532 3064
rect 9511 3057 9518 3061
rect 9518 3056 9519 3057
rect 9477 3050 9487 3056
rect 9236 3042 9271 3050
rect 9236 3016 9237 3042
rect 9244 3016 9271 3042
rect 9179 2998 9209 3012
rect 9236 3008 9271 3016
rect 9273 3042 9314 3050
rect 9273 3016 9288 3042
rect 9295 3016 9314 3042
rect 9378 3038 9409 3050
rect 9424 3038 9527 3050
rect 9539 3040 9565 3066
rect 9580 3061 9610 3072
rect 9642 3068 9704 3084
rect 9642 3066 9688 3068
rect 9642 3050 9704 3066
rect 9716 3050 9722 3098
rect 9725 3090 9805 3098
rect 9725 3088 9744 3090
rect 9759 3088 9793 3090
rect 9725 3072 9805 3088
rect 9725 3050 9744 3072
rect 9759 3056 9789 3072
rect 9817 3066 9823 3140
rect 9826 3066 9845 3210
rect 9860 3066 9866 3210
rect 9875 3140 9888 3210
rect 9940 3206 9962 3210
rect 9933 3184 9962 3198
rect 10015 3184 10031 3198
rect 10069 3194 10075 3196
rect 10082 3194 10190 3210
rect 10197 3194 10203 3196
rect 10211 3194 10226 3210
rect 10292 3204 10311 3207
rect 9933 3182 10031 3184
rect 10058 3182 10226 3194
rect 10241 3184 10257 3198
rect 10292 3185 10314 3204
rect 10324 3198 10340 3199
rect 10323 3196 10340 3198
rect 10324 3191 10340 3196
rect 10314 3184 10320 3185
rect 10323 3184 10352 3191
rect 10241 3183 10352 3184
rect 10241 3182 10358 3183
rect 9917 3174 9968 3182
rect 10015 3174 10049 3182
rect 9917 3162 9942 3174
rect 9949 3162 9968 3174
rect 10022 3172 10049 3174
rect 10058 3172 10279 3182
rect 10314 3179 10320 3182
rect 10022 3168 10279 3172
rect 9917 3154 9968 3162
rect 10015 3154 10279 3168
rect 10323 3174 10358 3182
rect 9869 3106 9888 3140
rect 9933 3146 9962 3154
rect 9933 3140 9950 3146
rect 9933 3138 9967 3140
rect 10015 3138 10031 3154
rect 10032 3144 10240 3154
rect 10241 3144 10257 3154
rect 10305 3150 10320 3165
rect 10323 3162 10324 3174
rect 10331 3162 10358 3174
rect 10323 3154 10358 3162
rect 10323 3153 10352 3154
rect 10043 3140 10257 3144
rect 10058 3138 10257 3140
rect 10292 3140 10305 3150
rect 10323 3140 10340 3153
rect 10292 3138 10340 3140
rect 9934 3134 9967 3138
rect 9930 3132 9967 3134
rect 9930 3131 9997 3132
rect 9930 3126 9961 3131
rect 9967 3126 9997 3131
rect 9930 3122 9997 3126
rect 9903 3119 9997 3122
rect 9903 3112 9952 3119
rect 9903 3106 9933 3112
rect 9952 3107 9957 3112
rect 9869 3090 9949 3106
rect 9961 3098 9997 3119
rect 10058 3114 10247 3138
rect 10292 3137 10339 3138
rect 10305 3132 10339 3137
rect 10073 3111 10247 3114
rect 10066 3108 10247 3111
rect 10275 3131 10339 3132
rect 9869 3088 9888 3090
rect 9903 3088 9937 3090
rect 9869 3072 9949 3088
rect 9869 3066 9888 3072
rect 9585 3040 9688 3050
rect 9539 3038 9688 3040
rect 9709 3038 9744 3050
rect 9378 3036 9540 3038
rect 9390 3016 9409 3036
rect 9424 3034 9454 3036
rect 9273 3008 9314 3016
rect 9396 3012 9409 3016
rect 9461 3020 9540 3036
rect 9572 3036 9744 3038
rect 9572 3020 9651 3036
rect 9658 3034 9688 3036
rect 9236 2998 9265 3008
rect 9279 2998 9308 3008
rect 9323 2998 9353 3012
rect 9396 2998 9439 3012
rect 9461 3008 9651 3020
rect 9716 3016 9722 3036
rect 9446 2998 9476 3008
rect 9477 2998 9635 3008
rect 9639 2998 9669 3008
rect 9673 2998 9703 3012
rect 9731 2998 9744 3036
rect 9816 3050 9845 3066
rect 9859 3050 9888 3066
rect 9903 3056 9933 3072
rect 9961 3050 9967 3098
rect 9970 3092 9989 3098
rect 10004 3092 10034 3100
rect 9970 3084 10034 3092
rect 9970 3068 10050 3084
rect 10066 3077 10128 3108
rect 10144 3077 10206 3108
rect 10275 3106 10324 3131
rect 10339 3106 10369 3122
rect 10238 3092 10268 3100
rect 10275 3098 10385 3106
rect 10238 3084 10283 3092
rect 9970 3066 9989 3068
rect 10004 3066 10050 3068
rect 9970 3050 10050 3066
rect 10077 3064 10112 3077
rect 10153 3074 10190 3077
rect 10153 3072 10195 3074
rect 10082 3061 10112 3064
rect 10091 3057 10098 3061
rect 10098 3056 10099 3057
rect 10057 3050 10067 3056
rect 9816 3042 9851 3050
rect 9816 3016 9817 3042
rect 9824 3016 9851 3042
rect 9759 2998 9789 3012
rect 9816 3008 9851 3016
rect 9853 3042 9894 3050
rect 9853 3016 9868 3042
rect 9875 3016 9894 3042
rect 9958 3038 9989 3050
rect 10004 3038 10107 3050
rect 10119 3040 10145 3066
rect 10160 3061 10190 3072
rect 10222 3068 10284 3084
rect 10222 3066 10268 3068
rect 10222 3050 10284 3066
rect 10296 3050 10302 3098
rect 10305 3090 10385 3098
rect 10305 3088 10324 3090
rect 10339 3088 10373 3090
rect 10305 3072 10385 3088
rect 10305 3050 10324 3072
rect 10339 3056 10369 3072
rect 10397 3066 10403 3140
rect 10406 3066 10425 3210
rect 10440 3066 10446 3210
rect 10455 3140 10468 3210
rect 10520 3206 10542 3210
rect 10513 3184 10542 3198
rect 10595 3184 10611 3198
rect 10649 3194 10655 3196
rect 10662 3194 10770 3210
rect 10777 3194 10783 3196
rect 10791 3194 10806 3210
rect 10872 3204 10891 3207
rect 10513 3182 10611 3184
rect 10638 3182 10806 3194
rect 10821 3184 10837 3198
rect 10872 3185 10894 3204
rect 10904 3198 10920 3199
rect 10903 3196 10920 3198
rect 10904 3191 10920 3196
rect 10894 3184 10900 3185
rect 10903 3184 10932 3191
rect 10821 3183 10932 3184
rect 10821 3182 10938 3183
rect 10497 3174 10548 3182
rect 10595 3174 10629 3182
rect 10497 3162 10522 3174
rect 10529 3162 10548 3174
rect 10602 3172 10629 3174
rect 10638 3172 10859 3182
rect 10894 3179 10900 3182
rect 10602 3168 10859 3172
rect 10497 3154 10548 3162
rect 10595 3154 10859 3168
rect 10903 3174 10938 3182
rect 10449 3106 10468 3140
rect 10513 3146 10542 3154
rect 10513 3140 10530 3146
rect 10513 3138 10547 3140
rect 10595 3138 10611 3154
rect 10612 3144 10820 3154
rect 10821 3144 10837 3154
rect 10885 3150 10900 3165
rect 10903 3162 10904 3174
rect 10911 3162 10938 3174
rect 10903 3154 10938 3162
rect 10903 3153 10932 3154
rect 10623 3140 10837 3144
rect 10638 3138 10837 3140
rect 10872 3140 10885 3150
rect 10903 3140 10920 3153
rect 10872 3138 10920 3140
rect 10514 3134 10547 3138
rect 10510 3132 10547 3134
rect 10510 3131 10577 3132
rect 10510 3126 10541 3131
rect 10547 3126 10577 3131
rect 10510 3122 10577 3126
rect 10483 3119 10577 3122
rect 10483 3112 10532 3119
rect 10483 3106 10513 3112
rect 10532 3107 10537 3112
rect 10449 3090 10529 3106
rect 10541 3098 10577 3119
rect 10638 3114 10827 3138
rect 10872 3137 10919 3138
rect 10885 3132 10919 3137
rect 10653 3111 10827 3114
rect 10646 3108 10827 3111
rect 10855 3131 10919 3132
rect 10449 3088 10468 3090
rect 10483 3088 10517 3090
rect 10449 3072 10529 3088
rect 10449 3066 10468 3072
rect 10165 3040 10268 3050
rect 10119 3038 10268 3040
rect 10289 3038 10324 3050
rect 9958 3036 10120 3038
rect 9970 3016 9989 3036
rect 10004 3034 10034 3036
rect 9853 3008 9894 3016
rect 9976 3012 9989 3016
rect 10041 3020 10120 3036
rect 10152 3036 10324 3038
rect 10152 3020 10231 3036
rect 10238 3034 10268 3036
rect 9816 2998 9845 3008
rect 9859 2998 9888 3008
rect 9903 2998 9933 3012
rect 9976 2998 10019 3012
rect 10041 3008 10231 3020
rect 10296 3016 10302 3036
rect 10026 2998 10056 3008
rect 10057 2998 10215 3008
rect 10219 2998 10249 3008
rect 10253 2998 10283 3012
rect 10311 2998 10324 3036
rect 10396 3050 10425 3066
rect 10439 3050 10468 3066
rect 10483 3056 10513 3072
rect 10541 3050 10547 3098
rect 10550 3092 10569 3098
rect 10584 3092 10614 3100
rect 10550 3084 10614 3092
rect 10550 3068 10630 3084
rect 10646 3077 10708 3108
rect 10724 3077 10786 3108
rect 10855 3106 10904 3131
rect 10919 3106 10949 3122
rect 10818 3092 10848 3100
rect 10855 3098 10965 3106
rect 10818 3084 10863 3092
rect 10550 3066 10569 3068
rect 10584 3066 10630 3068
rect 10550 3050 10630 3066
rect 10657 3064 10692 3077
rect 10733 3074 10770 3077
rect 10733 3072 10775 3074
rect 10662 3061 10692 3064
rect 10671 3057 10678 3061
rect 10678 3056 10679 3057
rect 10637 3050 10647 3056
rect 10396 3042 10431 3050
rect 10396 3016 10397 3042
rect 10404 3016 10431 3042
rect 10339 2998 10369 3012
rect 10396 3008 10431 3016
rect 10433 3042 10474 3050
rect 10433 3016 10448 3042
rect 10455 3016 10474 3042
rect 10538 3038 10569 3050
rect 10584 3038 10687 3050
rect 10699 3040 10725 3066
rect 10740 3061 10770 3072
rect 10802 3068 10864 3084
rect 10802 3066 10848 3068
rect 10802 3050 10864 3066
rect 10876 3050 10882 3098
rect 10885 3090 10965 3098
rect 10885 3088 10904 3090
rect 10919 3088 10953 3090
rect 10885 3072 10965 3088
rect 10885 3050 10904 3072
rect 10919 3056 10949 3072
rect 10977 3066 10983 3140
rect 10986 3066 11005 3210
rect 11020 3066 11026 3210
rect 11035 3140 11048 3210
rect 11100 3206 11122 3210
rect 11093 3184 11122 3198
rect 11175 3184 11191 3198
rect 11229 3194 11235 3196
rect 11242 3194 11350 3210
rect 11357 3194 11363 3196
rect 11371 3194 11386 3210
rect 11452 3204 11471 3207
rect 11093 3182 11191 3184
rect 11218 3182 11386 3194
rect 11401 3184 11417 3198
rect 11452 3185 11474 3204
rect 11484 3198 11500 3199
rect 11483 3196 11500 3198
rect 11484 3191 11500 3196
rect 11474 3184 11480 3185
rect 11483 3184 11512 3191
rect 11401 3183 11512 3184
rect 11401 3182 11518 3183
rect 11077 3174 11128 3182
rect 11175 3174 11209 3182
rect 11077 3162 11102 3174
rect 11109 3162 11128 3174
rect 11182 3172 11209 3174
rect 11218 3172 11439 3182
rect 11474 3179 11480 3182
rect 11182 3168 11439 3172
rect 11077 3154 11128 3162
rect 11175 3154 11439 3168
rect 11483 3174 11518 3182
rect 11029 3106 11048 3140
rect 11093 3146 11122 3154
rect 11093 3140 11110 3146
rect 11093 3138 11127 3140
rect 11175 3138 11191 3154
rect 11192 3144 11400 3154
rect 11401 3144 11417 3154
rect 11465 3150 11480 3165
rect 11483 3162 11484 3174
rect 11491 3162 11518 3174
rect 11483 3154 11518 3162
rect 11483 3153 11512 3154
rect 11203 3140 11417 3144
rect 11218 3138 11417 3140
rect 11452 3140 11465 3150
rect 11483 3140 11500 3153
rect 11452 3138 11500 3140
rect 11094 3134 11127 3138
rect 11090 3132 11127 3134
rect 11090 3131 11157 3132
rect 11090 3126 11121 3131
rect 11127 3126 11157 3131
rect 11090 3122 11157 3126
rect 11063 3119 11157 3122
rect 11063 3112 11112 3119
rect 11063 3106 11093 3112
rect 11112 3107 11117 3112
rect 11029 3090 11109 3106
rect 11121 3098 11157 3119
rect 11218 3114 11407 3138
rect 11452 3137 11499 3138
rect 11465 3132 11499 3137
rect 11233 3111 11407 3114
rect 11226 3108 11407 3111
rect 11435 3131 11499 3132
rect 11029 3088 11048 3090
rect 11063 3088 11097 3090
rect 11029 3072 11109 3088
rect 11029 3066 11048 3072
rect 10745 3040 10848 3050
rect 10699 3038 10848 3040
rect 10869 3038 10904 3050
rect 10538 3036 10700 3038
rect 10550 3016 10569 3036
rect 10584 3034 10614 3036
rect 10433 3008 10474 3016
rect 10556 3012 10569 3016
rect 10621 3020 10700 3036
rect 10732 3036 10904 3038
rect 10732 3020 10811 3036
rect 10818 3034 10848 3036
rect 10396 2998 10425 3008
rect 10439 2998 10468 3008
rect 10483 2998 10513 3012
rect 10556 2998 10599 3012
rect 10621 3008 10811 3020
rect 10876 3016 10882 3036
rect 10606 2998 10636 3008
rect 10637 2998 10795 3008
rect 10799 2998 10829 3008
rect 10833 2998 10863 3012
rect 10891 2998 10904 3036
rect 10976 3050 11005 3066
rect 11019 3050 11048 3066
rect 11063 3056 11093 3072
rect 11121 3050 11127 3098
rect 11130 3092 11149 3098
rect 11164 3092 11194 3100
rect 11130 3084 11194 3092
rect 11130 3068 11210 3084
rect 11226 3077 11288 3108
rect 11304 3077 11366 3108
rect 11435 3106 11484 3131
rect 11499 3106 11529 3122
rect 11398 3092 11428 3100
rect 11435 3098 11545 3106
rect 11398 3084 11443 3092
rect 11130 3066 11149 3068
rect 11164 3066 11210 3068
rect 11130 3050 11210 3066
rect 11237 3064 11272 3077
rect 11313 3074 11350 3077
rect 11313 3072 11355 3074
rect 11242 3061 11272 3064
rect 11251 3057 11258 3061
rect 11258 3056 11259 3057
rect 11217 3050 11227 3056
rect 10976 3042 11011 3050
rect 10976 3016 10977 3042
rect 10984 3016 11011 3042
rect 10919 2998 10949 3012
rect 10976 3008 11011 3016
rect 11013 3042 11054 3050
rect 11013 3016 11028 3042
rect 11035 3016 11054 3042
rect 11118 3038 11149 3050
rect 11164 3038 11267 3050
rect 11279 3040 11305 3066
rect 11320 3061 11350 3072
rect 11382 3068 11444 3084
rect 11382 3066 11428 3068
rect 11382 3050 11444 3066
rect 11456 3050 11462 3098
rect 11465 3090 11545 3098
rect 11465 3088 11484 3090
rect 11499 3088 11533 3090
rect 11465 3072 11545 3088
rect 11465 3050 11484 3072
rect 11499 3056 11529 3072
rect 11557 3066 11563 3140
rect 11566 3066 11585 3210
rect 11600 3066 11606 3210
rect 11615 3140 11628 3210
rect 11680 3206 11702 3210
rect 11673 3184 11702 3198
rect 11755 3184 11771 3198
rect 11809 3194 11815 3196
rect 11822 3194 11930 3210
rect 11937 3194 11943 3196
rect 11951 3194 11966 3210
rect 12032 3204 12051 3207
rect 11673 3182 11771 3184
rect 11798 3182 11966 3194
rect 11981 3184 11997 3198
rect 12032 3185 12054 3204
rect 12064 3198 12080 3199
rect 12063 3196 12080 3198
rect 12064 3191 12080 3196
rect 12054 3184 12060 3185
rect 12063 3184 12092 3191
rect 11981 3183 12092 3184
rect 11981 3182 12098 3183
rect 11657 3174 11708 3182
rect 11755 3174 11789 3182
rect 11657 3162 11682 3174
rect 11689 3162 11708 3174
rect 11762 3172 11789 3174
rect 11798 3172 12019 3182
rect 12054 3179 12060 3182
rect 11762 3168 12019 3172
rect 11657 3154 11708 3162
rect 11755 3154 12019 3168
rect 12063 3174 12098 3182
rect 11609 3106 11628 3140
rect 11673 3146 11702 3154
rect 11673 3140 11690 3146
rect 11673 3138 11707 3140
rect 11755 3138 11771 3154
rect 11772 3144 11980 3154
rect 11981 3144 11997 3154
rect 12045 3150 12060 3165
rect 12063 3162 12064 3174
rect 12071 3162 12098 3174
rect 12063 3154 12098 3162
rect 12063 3153 12092 3154
rect 11783 3140 11997 3144
rect 11798 3138 11997 3140
rect 12032 3140 12045 3150
rect 12063 3140 12080 3153
rect 12032 3138 12080 3140
rect 11674 3134 11707 3138
rect 11670 3132 11707 3134
rect 11670 3131 11737 3132
rect 11670 3126 11701 3131
rect 11707 3126 11737 3131
rect 11670 3122 11737 3126
rect 11643 3119 11737 3122
rect 11643 3112 11692 3119
rect 11643 3106 11673 3112
rect 11692 3107 11697 3112
rect 11609 3090 11689 3106
rect 11701 3098 11737 3119
rect 11798 3114 11987 3138
rect 12032 3137 12079 3138
rect 12045 3132 12079 3137
rect 11813 3111 11987 3114
rect 11806 3108 11987 3111
rect 12015 3131 12079 3132
rect 11609 3088 11628 3090
rect 11643 3088 11677 3090
rect 11609 3072 11689 3088
rect 11609 3066 11628 3072
rect 11325 3040 11428 3050
rect 11279 3038 11428 3040
rect 11449 3038 11484 3050
rect 11118 3036 11280 3038
rect 11130 3016 11149 3036
rect 11164 3034 11194 3036
rect 11013 3008 11054 3016
rect 11136 3012 11149 3016
rect 11201 3020 11280 3036
rect 11312 3036 11484 3038
rect 11312 3020 11391 3036
rect 11398 3034 11428 3036
rect 10976 2998 11005 3008
rect 11019 2998 11048 3008
rect 11063 2998 11093 3012
rect 11136 2998 11179 3012
rect 11201 3008 11391 3020
rect 11456 3016 11462 3036
rect 11186 2998 11216 3008
rect 11217 2998 11375 3008
rect 11379 2998 11409 3008
rect 11413 2998 11443 3012
rect 11471 2998 11484 3036
rect 11556 3050 11585 3066
rect 11599 3050 11628 3066
rect 11643 3056 11673 3072
rect 11701 3050 11707 3098
rect 11710 3092 11729 3098
rect 11744 3092 11774 3100
rect 11710 3084 11774 3092
rect 11710 3068 11790 3084
rect 11806 3077 11868 3108
rect 11884 3077 11946 3108
rect 12015 3106 12064 3131
rect 12079 3106 12109 3122
rect 11978 3092 12008 3100
rect 12015 3098 12125 3106
rect 11978 3084 12023 3092
rect 11710 3066 11729 3068
rect 11744 3066 11790 3068
rect 11710 3050 11790 3066
rect 11817 3064 11852 3077
rect 11893 3074 11930 3077
rect 11893 3072 11935 3074
rect 11822 3061 11852 3064
rect 11831 3057 11838 3061
rect 11838 3056 11839 3057
rect 11797 3050 11807 3056
rect 11556 3042 11591 3050
rect 11556 3016 11557 3042
rect 11564 3016 11591 3042
rect 11499 2998 11529 3012
rect 11556 3008 11591 3016
rect 11593 3042 11634 3050
rect 11593 3016 11608 3042
rect 11615 3016 11634 3042
rect 11698 3038 11729 3050
rect 11744 3038 11847 3050
rect 11859 3040 11885 3066
rect 11900 3061 11930 3072
rect 11962 3068 12024 3084
rect 11962 3066 12008 3068
rect 11962 3050 12024 3066
rect 12036 3050 12042 3098
rect 12045 3090 12125 3098
rect 12045 3088 12064 3090
rect 12079 3088 12113 3090
rect 12045 3072 12125 3088
rect 12045 3050 12064 3072
rect 12079 3056 12109 3072
rect 12137 3066 12143 3140
rect 12146 3066 12165 3210
rect 12180 3066 12186 3210
rect 12195 3140 12208 3210
rect 12260 3206 12282 3210
rect 12253 3184 12282 3198
rect 12335 3184 12351 3198
rect 12389 3194 12395 3196
rect 12402 3194 12510 3210
rect 12517 3194 12523 3196
rect 12531 3194 12546 3210
rect 12612 3204 12631 3207
rect 12253 3182 12351 3184
rect 12378 3182 12546 3194
rect 12561 3184 12577 3198
rect 12612 3185 12634 3204
rect 12644 3198 12660 3199
rect 12643 3196 12660 3198
rect 12644 3191 12660 3196
rect 12634 3184 12640 3185
rect 12643 3184 12672 3191
rect 12561 3183 12672 3184
rect 12561 3182 12678 3183
rect 12237 3174 12288 3182
rect 12335 3174 12369 3182
rect 12237 3162 12262 3174
rect 12269 3162 12288 3174
rect 12342 3172 12369 3174
rect 12378 3172 12599 3182
rect 12634 3179 12640 3182
rect 12342 3168 12599 3172
rect 12237 3154 12288 3162
rect 12335 3154 12599 3168
rect 12643 3174 12678 3182
rect 12189 3106 12208 3140
rect 12253 3146 12282 3154
rect 12253 3140 12270 3146
rect 12253 3138 12287 3140
rect 12335 3138 12351 3154
rect 12352 3144 12560 3154
rect 12561 3144 12577 3154
rect 12625 3150 12640 3165
rect 12643 3162 12644 3174
rect 12651 3162 12678 3174
rect 12643 3154 12678 3162
rect 12643 3153 12672 3154
rect 12363 3140 12577 3144
rect 12378 3138 12577 3140
rect 12612 3140 12625 3150
rect 12643 3140 12660 3153
rect 12612 3138 12660 3140
rect 12254 3134 12287 3138
rect 12250 3132 12287 3134
rect 12250 3131 12317 3132
rect 12250 3126 12281 3131
rect 12287 3126 12317 3131
rect 12250 3122 12317 3126
rect 12223 3119 12317 3122
rect 12223 3112 12272 3119
rect 12223 3106 12253 3112
rect 12272 3107 12277 3112
rect 12189 3090 12269 3106
rect 12281 3098 12317 3119
rect 12378 3114 12567 3138
rect 12612 3137 12659 3138
rect 12625 3132 12659 3137
rect 12393 3111 12567 3114
rect 12386 3108 12567 3111
rect 12595 3131 12659 3132
rect 12189 3088 12208 3090
rect 12223 3088 12257 3090
rect 12189 3072 12269 3088
rect 12189 3066 12208 3072
rect 11905 3040 12008 3050
rect 11859 3038 12008 3040
rect 12029 3038 12064 3050
rect 11698 3036 11860 3038
rect 11710 3016 11729 3036
rect 11744 3034 11774 3036
rect 11593 3008 11634 3016
rect 11716 3012 11729 3016
rect 11781 3020 11860 3036
rect 11892 3036 12064 3038
rect 11892 3020 11971 3036
rect 11978 3034 12008 3036
rect 11556 2998 11585 3008
rect 11599 2998 11628 3008
rect 11643 2998 11673 3012
rect 11716 2998 11759 3012
rect 11781 3008 11971 3020
rect 12036 3016 12042 3036
rect 11766 2998 11796 3008
rect 11797 2998 11955 3008
rect 11959 2998 11989 3008
rect 11993 2998 12023 3012
rect 12051 2998 12064 3036
rect 12136 3050 12165 3066
rect 12179 3050 12208 3066
rect 12223 3056 12253 3072
rect 12281 3050 12287 3098
rect 12290 3092 12309 3098
rect 12324 3092 12354 3100
rect 12290 3084 12354 3092
rect 12290 3068 12370 3084
rect 12386 3077 12448 3108
rect 12464 3077 12526 3108
rect 12595 3106 12644 3131
rect 12659 3106 12689 3122
rect 12558 3092 12588 3100
rect 12595 3098 12705 3106
rect 12558 3084 12603 3092
rect 12290 3066 12309 3068
rect 12324 3066 12370 3068
rect 12290 3050 12370 3066
rect 12397 3064 12432 3077
rect 12473 3074 12510 3077
rect 12473 3072 12515 3074
rect 12402 3061 12432 3064
rect 12411 3057 12418 3061
rect 12418 3056 12419 3057
rect 12377 3050 12387 3056
rect 12136 3042 12171 3050
rect 12136 3016 12137 3042
rect 12144 3016 12171 3042
rect 12079 2998 12109 3012
rect 12136 3008 12171 3016
rect 12173 3042 12214 3050
rect 12173 3016 12188 3042
rect 12195 3016 12214 3042
rect 12278 3038 12309 3050
rect 12324 3038 12427 3050
rect 12439 3040 12465 3066
rect 12480 3061 12510 3072
rect 12542 3068 12604 3084
rect 12542 3066 12588 3068
rect 12542 3050 12604 3066
rect 12616 3050 12622 3098
rect 12625 3090 12705 3098
rect 12625 3088 12644 3090
rect 12659 3088 12693 3090
rect 12625 3072 12705 3088
rect 12625 3050 12644 3072
rect 12659 3056 12689 3072
rect 12717 3066 12723 3140
rect 12726 3066 12745 3210
rect 12760 3066 12766 3210
rect 12775 3140 12788 3210
rect 12840 3206 12862 3210
rect 12833 3184 12862 3198
rect 12915 3184 12931 3198
rect 12969 3194 12975 3196
rect 12982 3194 13090 3210
rect 13097 3194 13103 3196
rect 13111 3194 13126 3210
rect 13192 3204 13211 3207
rect 12833 3182 12931 3184
rect 12958 3182 13126 3194
rect 13141 3184 13157 3198
rect 13192 3185 13214 3204
rect 13224 3198 13240 3199
rect 13223 3196 13240 3198
rect 13224 3191 13240 3196
rect 13214 3184 13220 3185
rect 13223 3184 13252 3191
rect 13141 3183 13252 3184
rect 13141 3182 13258 3183
rect 12817 3174 12868 3182
rect 12915 3174 12949 3182
rect 12817 3162 12842 3174
rect 12849 3162 12868 3174
rect 12922 3172 12949 3174
rect 12958 3172 13179 3182
rect 13214 3179 13220 3182
rect 12922 3168 13179 3172
rect 12817 3154 12868 3162
rect 12915 3154 13179 3168
rect 13223 3174 13258 3182
rect 12769 3106 12788 3140
rect 12833 3146 12862 3154
rect 12833 3140 12850 3146
rect 12833 3138 12867 3140
rect 12915 3138 12931 3154
rect 12932 3144 13140 3154
rect 13141 3144 13157 3154
rect 13205 3150 13220 3165
rect 13223 3162 13224 3174
rect 13231 3162 13258 3174
rect 13223 3154 13258 3162
rect 13223 3153 13252 3154
rect 12943 3140 13157 3144
rect 12958 3138 13157 3140
rect 13192 3140 13205 3150
rect 13223 3140 13240 3153
rect 13192 3138 13240 3140
rect 12834 3134 12867 3138
rect 12830 3132 12867 3134
rect 12830 3131 12897 3132
rect 12830 3126 12861 3131
rect 12867 3126 12897 3131
rect 12830 3122 12897 3126
rect 12803 3119 12897 3122
rect 12803 3112 12852 3119
rect 12803 3106 12833 3112
rect 12852 3107 12857 3112
rect 12769 3090 12849 3106
rect 12861 3098 12897 3119
rect 12958 3114 13147 3138
rect 13192 3137 13239 3138
rect 13205 3132 13239 3137
rect 12973 3111 13147 3114
rect 12966 3108 13147 3111
rect 13175 3131 13239 3132
rect 12769 3088 12788 3090
rect 12803 3088 12837 3090
rect 12769 3072 12849 3088
rect 12769 3066 12788 3072
rect 12485 3040 12588 3050
rect 12439 3038 12588 3040
rect 12609 3038 12644 3050
rect 12278 3036 12440 3038
rect 12290 3016 12309 3036
rect 12324 3034 12354 3036
rect 12173 3008 12214 3016
rect 12296 3012 12309 3016
rect 12361 3020 12440 3036
rect 12472 3036 12644 3038
rect 12472 3020 12551 3036
rect 12558 3034 12588 3036
rect 12136 2998 12165 3008
rect 12179 2998 12208 3008
rect 12223 2998 12253 3012
rect 12296 2998 12339 3012
rect 12361 3008 12551 3020
rect 12616 3016 12622 3036
rect 12346 2998 12376 3008
rect 12377 2998 12535 3008
rect 12539 2998 12569 3008
rect 12573 2998 12603 3012
rect 12631 2998 12644 3036
rect 12716 3050 12745 3066
rect 12759 3050 12788 3066
rect 12803 3056 12833 3072
rect 12861 3050 12867 3098
rect 12870 3092 12889 3098
rect 12904 3092 12934 3100
rect 12870 3084 12934 3092
rect 12870 3068 12950 3084
rect 12966 3077 13028 3108
rect 13044 3077 13106 3108
rect 13175 3106 13224 3131
rect 13239 3106 13269 3122
rect 13138 3092 13168 3100
rect 13175 3098 13285 3106
rect 13138 3084 13183 3092
rect 12870 3066 12889 3068
rect 12904 3066 12950 3068
rect 12870 3050 12950 3066
rect 12977 3064 13012 3077
rect 13053 3074 13090 3077
rect 13053 3072 13095 3074
rect 12982 3061 13012 3064
rect 12991 3057 12998 3061
rect 12998 3056 12999 3057
rect 12957 3050 12967 3056
rect 12716 3042 12751 3050
rect 12716 3016 12717 3042
rect 12724 3016 12751 3042
rect 12659 2998 12689 3012
rect 12716 3008 12751 3016
rect 12753 3042 12794 3050
rect 12753 3016 12768 3042
rect 12775 3016 12794 3042
rect 12858 3038 12889 3050
rect 12904 3038 13007 3050
rect 13019 3040 13045 3066
rect 13060 3061 13090 3072
rect 13122 3068 13184 3084
rect 13122 3066 13168 3068
rect 13122 3050 13184 3066
rect 13196 3050 13202 3098
rect 13205 3090 13285 3098
rect 13205 3088 13224 3090
rect 13239 3088 13273 3090
rect 13205 3072 13285 3088
rect 13205 3050 13224 3072
rect 13239 3056 13269 3072
rect 13297 3066 13303 3140
rect 13306 3066 13325 3210
rect 13340 3066 13346 3210
rect 13355 3140 13368 3210
rect 13420 3206 13442 3210
rect 13413 3184 13442 3198
rect 13495 3184 13511 3198
rect 13549 3194 13555 3196
rect 13562 3194 13670 3210
rect 13677 3194 13683 3196
rect 13691 3194 13706 3210
rect 13772 3204 13791 3207
rect 13413 3182 13511 3184
rect 13538 3182 13706 3194
rect 13721 3184 13737 3198
rect 13772 3185 13794 3204
rect 13804 3198 13820 3199
rect 13803 3196 13820 3198
rect 13804 3191 13820 3196
rect 13794 3184 13800 3185
rect 13803 3184 13832 3191
rect 13721 3183 13832 3184
rect 13721 3182 13838 3183
rect 13397 3174 13448 3182
rect 13495 3174 13529 3182
rect 13397 3162 13422 3174
rect 13429 3162 13448 3174
rect 13502 3172 13529 3174
rect 13538 3172 13759 3182
rect 13794 3179 13800 3182
rect 13502 3168 13759 3172
rect 13397 3154 13448 3162
rect 13495 3154 13759 3168
rect 13803 3174 13838 3182
rect 13349 3106 13368 3140
rect 13413 3146 13442 3154
rect 13413 3140 13430 3146
rect 13413 3138 13447 3140
rect 13495 3138 13511 3154
rect 13512 3144 13720 3154
rect 13721 3144 13737 3154
rect 13785 3150 13800 3165
rect 13803 3162 13804 3174
rect 13811 3162 13838 3174
rect 13803 3154 13838 3162
rect 13803 3153 13832 3154
rect 13523 3140 13737 3144
rect 13538 3138 13737 3140
rect 13772 3140 13785 3150
rect 13803 3140 13820 3153
rect 13772 3138 13820 3140
rect 13414 3134 13447 3138
rect 13410 3132 13447 3134
rect 13410 3131 13477 3132
rect 13410 3126 13441 3131
rect 13447 3126 13477 3131
rect 13410 3122 13477 3126
rect 13383 3119 13477 3122
rect 13383 3112 13432 3119
rect 13383 3106 13413 3112
rect 13432 3107 13437 3112
rect 13349 3090 13429 3106
rect 13441 3098 13477 3119
rect 13538 3114 13727 3138
rect 13772 3137 13819 3138
rect 13785 3132 13819 3137
rect 13553 3111 13727 3114
rect 13546 3108 13727 3111
rect 13755 3131 13819 3132
rect 13349 3088 13368 3090
rect 13383 3088 13417 3090
rect 13349 3072 13429 3088
rect 13349 3066 13368 3072
rect 13065 3040 13168 3050
rect 13019 3038 13168 3040
rect 13189 3038 13224 3050
rect 12858 3036 13020 3038
rect 12870 3016 12889 3036
rect 12904 3034 12934 3036
rect 12753 3008 12794 3016
rect 12876 3012 12889 3016
rect 12941 3020 13020 3036
rect 13052 3036 13224 3038
rect 13052 3020 13131 3036
rect 13138 3034 13168 3036
rect 12716 2998 12745 3008
rect 12759 2998 12788 3008
rect 12803 2998 12833 3012
rect 12876 2998 12919 3012
rect 12941 3008 13131 3020
rect 13196 3016 13202 3036
rect 12926 2998 12956 3008
rect 12957 2998 13115 3008
rect 13119 2998 13149 3008
rect 13153 2998 13183 3012
rect 13211 2998 13224 3036
rect 13296 3050 13325 3066
rect 13339 3050 13368 3066
rect 13383 3056 13413 3072
rect 13441 3050 13447 3098
rect 13450 3092 13469 3098
rect 13484 3092 13514 3100
rect 13450 3084 13514 3092
rect 13450 3068 13530 3084
rect 13546 3077 13608 3108
rect 13624 3077 13686 3108
rect 13755 3106 13804 3131
rect 13819 3106 13849 3122
rect 13718 3092 13748 3100
rect 13755 3098 13865 3106
rect 13718 3084 13763 3092
rect 13450 3066 13469 3068
rect 13484 3066 13530 3068
rect 13450 3050 13530 3066
rect 13557 3064 13592 3077
rect 13633 3074 13670 3077
rect 13633 3072 13675 3074
rect 13562 3061 13592 3064
rect 13571 3057 13578 3061
rect 13578 3056 13579 3057
rect 13537 3050 13547 3056
rect 13296 3042 13331 3050
rect 13296 3016 13297 3042
rect 13304 3016 13331 3042
rect 13239 2998 13269 3012
rect 13296 3008 13331 3016
rect 13333 3042 13374 3050
rect 13333 3016 13348 3042
rect 13355 3016 13374 3042
rect 13438 3038 13469 3050
rect 13484 3038 13587 3050
rect 13599 3040 13625 3066
rect 13640 3061 13670 3072
rect 13702 3068 13764 3084
rect 13702 3066 13748 3068
rect 13702 3050 13764 3066
rect 13776 3050 13782 3098
rect 13785 3090 13865 3098
rect 13785 3088 13804 3090
rect 13819 3088 13853 3090
rect 13785 3072 13865 3088
rect 13785 3050 13804 3072
rect 13819 3056 13849 3072
rect 13877 3066 13883 3140
rect 13886 3066 13905 3210
rect 13920 3066 13926 3210
rect 13935 3140 13948 3210
rect 14000 3206 14022 3210
rect 13993 3184 14022 3198
rect 14075 3184 14091 3198
rect 14129 3194 14135 3196
rect 14142 3194 14250 3210
rect 14257 3194 14263 3196
rect 14271 3194 14286 3210
rect 14352 3204 14371 3207
rect 13993 3182 14091 3184
rect 14118 3182 14286 3194
rect 14301 3184 14317 3198
rect 14352 3185 14374 3204
rect 14384 3198 14400 3199
rect 14383 3196 14400 3198
rect 14384 3191 14400 3196
rect 14374 3184 14380 3185
rect 14383 3184 14412 3191
rect 14301 3183 14412 3184
rect 14301 3182 14418 3183
rect 13977 3174 14028 3182
rect 14075 3174 14109 3182
rect 13977 3162 14002 3174
rect 14009 3162 14028 3174
rect 14082 3172 14109 3174
rect 14118 3172 14339 3182
rect 14374 3179 14380 3182
rect 14082 3168 14339 3172
rect 13977 3154 14028 3162
rect 14075 3154 14339 3168
rect 14383 3174 14418 3182
rect 13929 3106 13948 3140
rect 13993 3146 14022 3154
rect 13993 3140 14010 3146
rect 13993 3138 14027 3140
rect 14075 3138 14091 3154
rect 14092 3144 14300 3154
rect 14301 3144 14317 3154
rect 14365 3150 14380 3165
rect 14383 3162 14384 3174
rect 14391 3162 14418 3174
rect 14383 3154 14418 3162
rect 14383 3153 14412 3154
rect 14103 3140 14317 3144
rect 14118 3138 14317 3140
rect 14352 3140 14365 3150
rect 14383 3140 14400 3153
rect 14352 3138 14400 3140
rect 13994 3134 14027 3138
rect 13990 3132 14027 3134
rect 13990 3131 14057 3132
rect 13990 3126 14021 3131
rect 14027 3126 14057 3131
rect 13990 3122 14057 3126
rect 13963 3119 14057 3122
rect 13963 3112 14012 3119
rect 13963 3106 13993 3112
rect 14012 3107 14017 3112
rect 13929 3090 14009 3106
rect 14021 3098 14057 3119
rect 14118 3114 14307 3138
rect 14352 3137 14399 3138
rect 14365 3132 14399 3137
rect 14133 3111 14307 3114
rect 14126 3108 14307 3111
rect 14335 3131 14399 3132
rect 13929 3088 13948 3090
rect 13963 3088 13997 3090
rect 13929 3072 14009 3088
rect 13929 3066 13948 3072
rect 13645 3040 13748 3050
rect 13599 3038 13748 3040
rect 13769 3038 13804 3050
rect 13438 3036 13600 3038
rect 13450 3016 13469 3036
rect 13484 3034 13514 3036
rect 13333 3008 13374 3016
rect 13456 3012 13469 3016
rect 13521 3020 13600 3036
rect 13632 3036 13804 3038
rect 13632 3020 13711 3036
rect 13718 3034 13748 3036
rect 13296 2998 13325 3008
rect 13339 2998 13368 3008
rect 13383 2998 13413 3012
rect 13456 2998 13499 3012
rect 13521 3008 13711 3020
rect 13776 3016 13782 3036
rect 13506 2998 13536 3008
rect 13537 2998 13695 3008
rect 13699 2998 13729 3008
rect 13733 2998 13763 3012
rect 13791 2998 13804 3036
rect 13876 3050 13905 3066
rect 13919 3050 13948 3066
rect 13963 3056 13993 3072
rect 14021 3050 14027 3098
rect 14030 3092 14049 3098
rect 14064 3092 14094 3100
rect 14030 3084 14094 3092
rect 14030 3068 14110 3084
rect 14126 3077 14188 3108
rect 14204 3077 14266 3108
rect 14335 3106 14384 3131
rect 14399 3106 14429 3122
rect 14298 3092 14328 3100
rect 14335 3098 14445 3106
rect 14298 3084 14343 3092
rect 14030 3066 14049 3068
rect 14064 3066 14110 3068
rect 14030 3050 14110 3066
rect 14137 3064 14172 3077
rect 14213 3074 14250 3077
rect 14213 3072 14255 3074
rect 14142 3061 14172 3064
rect 14151 3057 14158 3061
rect 14158 3056 14159 3057
rect 14117 3050 14127 3056
rect 13876 3042 13911 3050
rect 13876 3016 13877 3042
rect 13884 3016 13911 3042
rect 13819 2998 13849 3012
rect 13876 3008 13911 3016
rect 13913 3042 13954 3050
rect 13913 3016 13928 3042
rect 13935 3016 13954 3042
rect 14018 3038 14049 3050
rect 14064 3038 14167 3050
rect 14179 3040 14205 3066
rect 14220 3061 14250 3072
rect 14282 3068 14344 3084
rect 14282 3066 14328 3068
rect 14282 3050 14344 3066
rect 14356 3050 14362 3098
rect 14365 3090 14445 3098
rect 14365 3088 14384 3090
rect 14399 3088 14433 3090
rect 14365 3072 14445 3088
rect 14365 3050 14384 3072
rect 14399 3056 14429 3072
rect 14457 3066 14463 3140
rect 14466 3066 14485 3210
rect 14500 3066 14506 3210
rect 14515 3140 14528 3210
rect 14580 3206 14602 3210
rect 14573 3184 14602 3198
rect 14655 3184 14671 3198
rect 14709 3194 14715 3196
rect 14722 3194 14830 3210
rect 14837 3194 14843 3196
rect 14851 3194 14866 3210
rect 14932 3204 14951 3207
rect 14573 3182 14671 3184
rect 14698 3182 14866 3194
rect 14881 3184 14897 3198
rect 14932 3185 14954 3204
rect 14964 3198 14980 3199
rect 14963 3196 14980 3198
rect 14964 3191 14980 3196
rect 14954 3184 14960 3185
rect 14963 3184 14992 3191
rect 14881 3183 14992 3184
rect 14881 3182 14998 3183
rect 14557 3174 14608 3182
rect 14655 3174 14689 3182
rect 14557 3162 14582 3174
rect 14589 3162 14608 3174
rect 14662 3172 14689 3174
rect 14698 3172 14919 3182
rect 14954 3179 14960 3182
rect 14662 3168 14919 3172
rect 14557 3154 14608 3162
rect 14655 3154 14919 3168
rect 14963 3174 14998 3182
rect 14509 3106 14528 3140
rect 14573 3146 14602 3154
rect 14573 3140 14590 3146
rect 14573 3138 14607 3140
rect 14655 3138 14671 3154
rect 14672 3144 14880 3154
rect 14881 3144 14897 3154
rect 14945 3150 14960 3165
rect 14963 3162 14964 3174
rect 14971 3162 14998 3174
rect 14963 3154 14998 3162
rect 14963 3153 14992 3154
rect 14683 3140 14897 3144
rect 14698 3138 14897 3140
rect 14932 3140 14945 3150
rect 14963 3140 14980 3153
rect 14932 3138 14980 3140
rect 14574 3134 14607 3138
rect 14570 3132 14607 3134
rect 14570 3131 14637 3132
rect 14570 3126 14601 3131
rect 14607 3126 14637 3131
rect 14570 3122 14637 3126
rect 14543 3119 14637 3122
rect 14543 3112 14592 3119
rect 14543 3106 14573 3112
rect 14592 3107 14597 3112
rect 14509 3090 14589 3106
rect 14601 3098 14637 3119
rect 14698 3114 14887 3138
rect 14932 3137 14979 3138
rect 14945 3132 14979 3137
rect 14713 3111 14887 3114
rect 14706 3108 14887 3111
rect 14915 3131 14979 3132
rect 14509 3088 14528 3090
rect 14543 3088 14577 3090
rect 14509 3072 14589 3088
rect 14509 3066 14528 3072
rect 14225 3040 14328 3050
rect 14179 3038 14328 3040
rect 14349 3038 14384 3050
rect 14018 3036 14180 3038
rect 14030 3016 14049 3036
rect 14064 3034 14094 3036
rect 13913 3008 13954 3016
rect 14036 3012 14049 3016
rect 14101 3020 14180 3036
rect 14212 3036 14384 3038
rect 14212 3020 14291 3036
rect 14298 3034 14328 3036
rect 13876 2998 13905 3008
rect 13919 2998 13948 3008
rect 13963 2998 13993 3012
rect 14036 2998 14079 3012
rect 14101 3008 14291 3020
rect 14356 3016 14362 3036
rect 14086 2998 14116 3008
rect 14117 2998 14275 3008
rect 14279 2998 14309 3008
rect 14313 2998 14343 3012
rect 14371 2998 14384 3036
rect 14456 3050 14485 3066
rect 14499 3050 14528 3066
rect 14543 3056 14573 3072
rect 14601 3050 14607 3098
rect 14610 3092 14629 3098
rect 14644 3092 14674 3100
rect 14610 3084 14674 3092
rect 14610 3068 14690 3084
rect 14706 3077 14768 3108
rect 14784 3077 14846 3108
rect 14915 3106 14964 3131
rect 14979 3106 15009 3122
rect 14878 3092 14908 3100
rect 14915 3098 15025 3106
rect 14878 3084 14923 3092
rect 14610 3066 14629 3068
rect 14644 3066 14690 3068
rect 14610 3050 14690 3066
rect 14717 3064 14752 3077
rect 14793 3074 14830 3077
rect 14793 3072 14835 3074
rect 14722 3061 14752 3064
rect 14731 3057 14738 3061
rect 14738 3056 14739 3057
rect 14697 3050 14707 3056
rect 14456 3042 14491 3050
rect 14456 3016 14457 3042
rect 14464 3016 14491 3042
rect 14399 2998 14429 3012
rect 14456 3008 14491 3016
rect 14493 3042 14534 3050
rect 14493 3016 14508 3042
rect 14515 3016 14534 3042
rect 14598 3038 14629 3050
rect 14644 3038 14747 3050
rect 14759 3040 14785 3066
rect 14800 3061 14830 3072
rect 14862 3068 14924 3084
rect 14862 3066 14908 3068
rect 14862 3050 14924 3066
rect 14936 3050 14942 3098
rect 14945 3090 15025 3098
rect 14945 3088 14964 3090
rect 14979 3088 15013 3090
rect 14945 3072 15025 3088
rect 14945 3050 14964 3072
rect 14979 3056 15009 3072
rect 15037 3066 15043 3140
rect 15046 3066 15065 3210
rect 15080 3066 15086 3210
rect 15095 3140 15108 3210
rect 15160 3206 15182 3210
rect 15153 3184 15182 3198
rect 15235 3184 15251 3198
rect 15289 3194 15295 3196
rect 15302 3194 15410 3210
rect 15417 3194 15423 3196
rect 15431 3194 15446 3210
rect 15512 3204 15531 3207
rect 15153 3182 15251 3184
rect 15278 3182 15446 3194
rect 15461 3184 15477 3198
rect 15512 3185 15534 3204
rect 15544 3198 15560 3199
rect 15543 3196 15560 3198
rect 15544 3191 15560 3196
rect 15534 3184 15540 3185
rect 15543 3184 15572 3191
rect 15461 3183 15572 3184
rect 15461 3182 15578 3183
rect 15137 3174 15188 3182
rect 15235 3174 15269 3182
rect 15137 3162 15162 3174
rect 15169 3162 15188 3174
rect 15242 3172 15269 3174
rect 15278 3172 15499 3182
rect 15534 3179 15540 3182
rect 15242 3168 15499 3172
rect 15137 3154 15188 3162
rect 15235 3154 15499 3168
rect 15543 3174 15578 3182
rect 15089 3106 15108 3140
rect 15153 3146 15182 3154
rect 15153 3140 15170 3146
rect 15153 3138 15187 3140
rect 15235 3138 15251 3154
rect 15252 3144 15460 3154
rect 15461 3144 15477 3154
rect 15525 3150 15540 3165
rect 15543 3162 15544 3174
rect 15551 3162 15578 3174
rect 15543 3154 15578 3162
rect 15543 3153 15572 3154
rect 15263 3140 15477 3144
rect 15278 3138 15477 3140
rect 15512 3140 15525 3150
rect 15543 3140 15560 3153
rect 15512 3138 15560 3140
rect 15154 3134 15187 3138
rect 15150 3132 15187 3134
rect 15150 3131 15217 3132
rect 15150 3126 15181 3131
rect 15187 3126 15217 3131
rect 15150 3122 15217 3126
rect 15123 3119 15217 3122
rect 15123 3112 15172 3119
rect 15123 3106 15153 3112
rect 15172 3107 15177 3112
rect 15089 3090 15169 3106
rect 15181 3098 15217 3119
rect 15278 3114 15467 3138
rect 15512 3137 15559 3138
rect 15525 3132 15559 3137
rect 15293 3111 15467 3114
rect 15286 3108 15467 3111
rect 15495 3131 15559 3132
rect 15089 3088 15108 3090
rect 15123 3088 15157 3090
rect 15089 3072 15169 3088
rect 15089 3066 15108 3072
rect 14805 3040 14908 3050
rect 14759 3038 14908 3040
rect 14929 3038 14964 3050
rect 14598 3036 14760 3038
rect 14610 3016 14629 3036
rect 14644 3034 14674 3036
rect 14493 3008 14534 3016
rect 14616 3012 14629 3016
rect 14681 3020 14760 3036
rect 14792 3036 14964 3038
rect 14792 3020 14871 3036
rect 14878 3034 14908 3036
rect 14456 2998 14485 3008
rect 14499 2998 14528 3008
rect 14543 2998 14573 3012
rect 14616 2998 14659 3012
rect 14681 3008 14871 3020
rect 14936 3016 14942 3036
rect 14666 2998 14696 3008
rect 14697 2998 14855 3008
rect 14859 2998 14889 3008
rect 14893 2998 14923 3012
rect 14951 2998 14964 3036
rect 15036 3050 15065 3066
rect 15079 3050 15108 3066
rect 15123 3056 15153 3072
rect 15181 3050 15187 3098
rect 15190 3092 15209 3098
rect 15224 3092 15254 3100
rect 15190 3084 15254 3092
rect 15190 3068 15270 3084
rect 15286 3077 15348 3108
rect 15364 3077 15426 3108
rect 15495 3106 15544 3131
rect 15559 3106 15589 3122
rect 15458 3092 15488 3100
rect 15495 3098 15605 3106
rect 15458 3084 15503 3092
rect 15190 3066 15209 3068
rect 15224 3066 15270 3068
rect 15190 3050 15270 3066
rect 15297 3064 15332 3077
rect 15373 3074 15410 3077
rect 15373 3072 15415 3074
rect 15302 3061 15332 3064
rect 15311 3057 15318 3061
rect 15318 3056 15319 3057
rect 15277 3050 15287 3056
rect 15036 3042 15071 3050
rect 15036 3016 15037 3042
rect 15044 3016 15071 3042
rect 14979 2998 15009 3012
rect 15036 3008 15071 3016
rect 15073 3042 15114 3050
rect 15073 3016 15088 3042
rect 15095 3016 15114 3042
rect 15178 3038 15209 3050
rect 15224 3038 15327 3050
rect 15339 3040 15365 3066
rect 15380 3061 15410 3072
rect 15442 3068 15504 3084
rect 15442 3066 15488 3068
rect 15442 3050 15504 3066
rect 15516 3050 15522 3098
rect 15525 3090 15605 3098
rect 15525 3088 15544 3090
rect 15559 3088 15593 3090
rect 15525 3072 15605 3088
rect 15525 3050 15544 3072
rect 15559 3056 15589 3072
rect 15617 3066 15623 3140
rect 15626 3066 15645 3210
rect 15660 3066 15666 3210
rect 15675 3140 15688 3210
rect 15740 3206 15762 3210
rect 15733 3184 15762 3198
rect 15815 3184 15831 3198
rect 15869 3194 15875 3196
rect 15882 3194 15990 3210
rect 15997 3194 16003 3196
rect 16011 3194 16026 3210
rect 16092 3204 16111 3207
rect 15733 3182 15831 3184
rect 15858 3182 16026 3194
rect 16041 3184 16057 3198
rect 16092 3185 16114 3204
rect 16124 3198 16140 3199
rect 16123 3196 16140 3198
rect 16124 3191 16140 3196
rect 16114 3184 16120 3185
rect 16123 3184 16152 3191
rect 16041 3183 16152 3184
rect 16041 3182 16158 3183
rect 15717 3174 15768 3182
rect 15815 3174 15849 3182
rect 15717 3162 15742 3174
rect 15749 3162 15768 3174
rect 15822 3172 15849 3174
rect 15858 3172 16079 3182
rect 16114 3179 16120 3182
rect 15822 3168 16079 3172
rect 15717 3154 15768 3162
rect 15815 3154 16079 3168
rect 16123 3174 16158 3182
rect 15669 3106 15688 3140
rect 15733 3146 15762 3154
rect 15733 3140 15750 3146
rect 15733 3138 15767 3140
rect 15815 3138 15831 3154
rect 15832 3144 16040 3154
rect 16041 3144 16057 3154
rect 16105 3150 16120 3165
rect 16123 3162 16124 3174
rect 16131 3162 16158 3174
rect 16123 3154 16158 3162
rect 16123 3153 16152 3154
rect 15843 3140 16057 3144
rect 15858 3138 16057 3140
rect 16092 3140 16105 3150
rect 16123 3140 16140 3153
rect 16092 3138 16140 3140
rect 15734 3134 15767 3138
rect 15730 3132 15767 3134
rect 15730 3131 15797 3132
rect 15730 3126 15761 3131
rect 15767 3126 15797 3131
rect 15730 3122 15797 3126
rect 15703 3119 15797 3122
rect 15703 3112 15752 3119
rect 15703 3106 15733 3112
rect 15752 3107 15757 3112
rect 15669 3090 15749 3106
rect 15761 3098 15797 3119
rect 15858 3114 16047 3138
rect 16092 3137 16139 3138
rect 16105 3132 16139 3137
rect 15873 3111 16047 3114
rect 15866 3108 16047 3111
rect 16075 3131 16139 3132
rect 15669 3088 15688 3090
rect 15703 3088 15737 3090
rect 15669 3072 15749 3088
rect 15669 3066 15688 3072
rect 15385 3040 15488 3050
rect 15339 3038 15488 3040
rect 15509 3038 15544 3050
rect 15178 3036 15340 3038
rect 15190 3016 15209 3036
rect 15224 3034 15254 3036
rect 15073 3008 15114 3016
rect 15196 3012 15209 3016
rect 15261 3020 15340 3036
rect 15372 3036 15544 3038
rect 15372 3020 15451 3036
rect 15458 3034 15488 3036
rect 15036 2998 15065 3008
rect 15079 2998 15108 3008
rect 15123 2998 15153 3012
rect 15196 2998 15239 3012
rect 15261 3008 15451 3020
rect 15516 3016 15522 3036
rect 15246 2998 15276 3008
rect 15277 2998 15435 3008
rect 15439 2998 15469 3008
rect 15473 2998 15503 3012
rect 15531 2998 15544 3036
rect 15616 3050 15645 3066
rect 15659 3050 15688 3066
rect 15703 3056 15733 3072
rect 15761 3050 15767 3098
rect 15770 3092 15789 3098
rect 15804 3092 15834 3100
rect 15770 3084 15834 3092
rect 15770 3068 15850 3084
rect 15866 3077 15928 3108
rect 15944 3077 16006 3108
rect 16075 3106 16124 3131
rect 16139 3106 16169 3122
rect 16038 3092 16068 3100
rect 16075 3098 16185 3106
rect 16038 3084 16083 3092
rect 15770 3066 15789 3068
rect 15804 3066 15850 3068
rect 15770 3050 15850 3066
rect 15877 3064 15912 3077
rect 15953 3074 15990 3077
rect 15953 3072 15995 3074
rect 15882 3061 15912 3064
rect 15891 3057 15898 3061
rect 15898 3056 15899 3057
rect 15857 3050 15867 3056
rect 15616 3042 15651 3050
rect 15616 3016 15617 3042
rect 15624 3016 15651 3042
rect 15559 2998 15589 3012
rect 15616 3008 15651 3016
rect 15653 3042 15694 3050
rect 15653 3016 15668 3042
rect 15675 3016 15694 3042
rect 15758 3038 15789 3050
rect 15804 3038 15907 3050
rect 15919 3040 15945 3066
rect 15960 3061 15990 3072
rect 16022 3068 16084 3084
rect 16022 3066 16068 3068
rect 16022 3050 16084 3066
rect 16096 3050 16102 3098
rect 16105 3090 16185 3098
rect 16105 3088 16124 3090
rect 16139 3088 16173 3090
rect 16105 3072 16185 3088
rect 16105 3050 16124 3072
rect 16139 3056 16169 3072
rect 16197 3066 16203 3140
rect 16206 3066 16225 3210
rect 16240 3066 16246 3210
rect 16255 3140 16268 3210
rect 16320 3206 16342 3210
rect 16313 3184 16342 3198
rect 16395 3184 16411 3198
rect 16449 3194 16455 3196
rect 16462 3194 16570 3210
rect 16577 3194 16583 3196
rect 16591 3194 16606 3210
rect 16672 3204 16691 3207
rect 16313 3182 16411 3184
rect 16438 3182 16606 3194
rect 16621 3184 16637 3198
rect 16672 3185 16694 3204
rect 16704 3198 16720 3199
rect 16703 3196 16720 3198
rect 16704 3191 16720 3196
rect 16694 3184 16700 3185
rect 16703 3184 16732 3191
rect 16621 3183 16732 3184
rect 16621 3182 16738 3183
rect 16297 3174 16348 3182
rect 16395 3174 16429 3182
rect 16297 3162 16322 3174
rect 16329 3162 16348 3174
rect 16402 3172 16429 3174
rect 16438 3172 16659 3182
rect 16694 3179 16700 3182
rect 16402 3168 16659 3172
rect 16297 3154 16348 3162
rect 16395 3154 16659 3168
rect 16703 3174 16738 3182
rect 16249 3106 16268 3140
rect 16313 3146 16342 3154
rect 16313 3140 16330 3146
rect 16313 3138 16347 3140
rect 16395 3138 16411 3154
rect 16412 3144 16620 3154
rect 16621 3144 16637 3154
rect 16685 3150 16700 3165
rect 16703 3162 16704 3174
rect 16711 3162 16738 3174
rect 16703 3154 16738 3162
rect 16703 3153 16732 3154
rect 16423 3140 16637 3144
rect 16438 3138 16637 3140
rect 16672 3140 16685 3150
rect 16703 3140 16720 3153
rect 16672 3138 16720 3140
rect 16314 3134 16347 3138
rect 16310 3132 16347 3134
rect 16310 3131 16377 3132
rect 16310 3126 16341 3131
rect 16347 3126 16377 3131
rect 16310 3122 16377 3126
rect 16283 3119 16377 3122
rect 16283 3112 16332 3119
rect 16283 3106 16313 3112
rect 16332 3107 16337 3112
rect 16249 3090 16329 3106
rect 16341 3098 16377 3119
rect 16438 3114 16627 3138
rect 16672 3137 16719 3138
rect 16685 3132 16719 3137
rect 16453 3111 16627 3114
rect 16446 3108 16627 3111
rect 16655 3131 16719 3132
rect 16249 3088 16268 3090
rect 16283 3088 16317 3090
rect 16249 3072 16329 3088
rect 16249 3066 16268 3072
rect 15965 3040 16068 3050
rect 15919 3038 16068 3040
rect 16089 3038 16124 3050
rect 15758 3036 15920 3038
rect 15770 3016 15789 3036
rect 15804 3034 15834 3036
rect 15653 3008 15694 3016
rect 15776 3012 15789 3016
rect 15841 3020 15920 3036
rect 15952 3036 16124 3038
rect 15952 3020 16031 3036
rect 16038 3034 16068 3036
rect 15616 2998 15645 3008
rect 15659 2998 15688 3008
rect 15703 2998 15733 3012
rect 15776 2998 15819 3012
rect 15841 3008 16031 3020
rect 16096 3016 16102 3036
rect 15826 2998 15856 3008
rect 15857 2998 16015 3008
rect 16019 2998 16049 3008
rect 16053 2998 16083 3012
rect 16111 2998 16124 3036
rect 16196 3050 16225 3066
rect 16239 3050 16268 3066
rect 16283 3056 16313 3072
rect 16341 3050 16347 3098
rect 16350 3092 16369 3098
rect 16384 3092 16414 3100
rect 16350 3084 16414 3092
rect 16350 3068 16430 3084
rect 16446 3077 16508 3108
rect 16524 3077 16586 3108
rect 16655 3106 16704 3131
rect 16719 3106 16749 3122
rect 16618 3092 16648 3100
rect 16655 3098 16765 3106
rect 16618 3084 16663 3092
rect 16350 3066 16369 3068
rect 16384 3066 16430 3068
rect 16350 3050 16430 3066
rect 16457 3064 16492 3077
rect 16533 3074 16570 3077
rect 16533 3072 16575 3074
rect 16462 3061 16492 3064
rect 16471 3057 16478 3061
rect 16478 3056 16479 3057
rect 16437 3050 16447 3056
rect 16196 3042 16231 3050
rect 16196 3016 16197 3042
rect 16204 3016 16231 3042
rect 16139 2998 16169 3012
rect 16196 3008 16231 3016
rect 16233 3042 16274 3050
rect 16233 3016 16248 3042
rect 16255 3016 16274 3042
rect 16338 3038 16369 3050
rect 16384 3038 16487 3050
rect 16499 3040 16525 3066
rect 16540 3061 16570 3072
rect 16602 3068 16664 3084
rect 16602 3066 16648 3068
rect 16602 3050 16664 3066
rect 16676 3050 16682 3098
rect 16685 3090 16765 3098
rect 16685 3088 16704 3090
rect 16719 3088 16753 3090
rect 16685 3072 16765 3088
rect 16685 3050 16704 3072
rect 16719 3056 16749 3072
rect 16777 3066 16783 3140
rect 16786 3066 16805 3210
rect 16820 3066 16826 3210
rect 16835 3140 16848 3210
rect 16900 3206 16922 3210
rect 16893 3184 16922 3198
rect 16975 3184 16991 3198
rect 17029 3194 17035 3196
rect 17042 3194 17150 3210
rect 17157 3194 17163 3196
rect 17171 3194 17186 3210
rect 17252 3204 17271 3207
rect 16893 3182 16991 3184
rect 17018 3182 17186 3194
rect 17201 3184 17217 3198
rect 17252 3185 17274 3204
rect 17284 3198 17300 3199
rect 17283 3196 17300 3198
rect 17284 3191 17300 3196
rect 17274 3184 17280 3185
rect 17283 3184 17312 3191
rect 17201 3183 17312 3184
rect 17201 3182 17318 3183
rect 16877 3174 16928 3182
rect 16975 3174 17009 3182
rect 16877 3162 16902 3174
rect 16909 3162 16928 3174
rect 16982 3172 17009 3174
rect 17018 3172 17239 3182
rect 17274 3179 17280 3182
rect 16982 3168 17239 3172
rect 16877 3154 16928 3162
rect 16975 3154 17239 3168
rect 17283 3174 17318 3182
rect 16829 3106 16848 3140
rect 16893 3146 16922 3154
rect 16893 3140 16910 3146
rect 16893 3138 16927 3140
rect 16975 3138 16991 3154
rect 16992 3144 17200 3154
rect 17201 3144 17217 3154
rect 17265 3150 17280 3165
rect 17283 3162 17284 3174
rect 17291 3162 17318 3174
rect 17283 3154 17318 3162
rect 17283 3153 17312 3154
rect 17003 3140 17217 3144
rect 17018 3138 17217 3140
rect 17252 3140 17265 3150
rect 17283 3140 17300 3153
rect 17252 3138 17300 3140
rect 16894 3134 16927 3138
rect 16890 3132 16927 3134
rect 16890 3131 16957 3132
rect 16890 3126 16921 3131
rect 16927 3126 16957 3131
rect 16890 3122 16957 3126
rect 16863 3119 16957 3122
rect 16863 3112 16912 3119
rect 16863 3106 16893 3112
rect 16912 3107 16917 3112
rect 16829 3090 16909 3106
rect 16921 3098 16957 3119
rect 17018 3114 17207 3138
rect 17252 3137 17299 3138
rect 17265 3132 17299 3137
rect 17033 3111 17207 3114
rect 17026 3108 17207 3111
rect 17235 3131 17299 3132
rect 16829 3088 16848 3090
rect 16863 3088 16897 3090
rect 16829 3072 16909 3088
rect 16829 3066 16848 3072
rect 16545 3040 16648 3050
rect 16499 3038 16648 3040
rect 16669 3038 16704 3050
rect 16338 3036 16500 3038
rect 16350 3016 16369 3036
rect 16384 3034 16414 3036
rect 16233 3008 16274 3016
rect 16356 3012 16369 3016
rect 16421 3020 16500 3036
rect 16532 3036 16704 3038
rect 16532 3020 16611 3036
rect 16618 3034 16648 3036
rect 16196 2998 16225 3008
rect 16239 2998 16268 3008
rect 16283 2998 16313 3012
rect 16356 2998 16399 3012
rect 16421 3008 16611 3020
rect 16676 3016 16682 3036
rect 16406 2998 16436 3008
rect 16437 2998 16595 3008
rect 16599 2998 16629 3008
rect 16633 2998 16663 3012
rect 16691 2998 16704 3036
rect 16776 3050 16805 3066
rect 16819 3050 16848 3066
rect 16863 3056 16893 3072
rect 16921 3050 16927 3098
rect 16930 3092 16949 3098
rect 16964 3092 16994 3100
rect 16930 3084 16994 3092
rect 16930 3068 17010 3084
rect 17026 3077 17088 3108
rect 17104 3077 17166 3108
rect 17235 3106 17284 3131
rect 17299 3106 17329 3122
rect 17198 3092 17228 3100
rect 17235 3098 17345 3106
rect 17198 3084 17243 3092
rect 16930 3066 16949 3068
rect 16964 3066 17010 3068
rect 16930 3050 17010 3066
rect 17037 3064 17072 3077
rect 17113 3074 17150 3077
rect 17113 3072 17155 3074
rect 17042 3061 17072 3064
rect 17051 3057 17058 3061
rect 17058 3056 17059 3057
rect 17017 3050 17027 3056
rect 16776 3042 16811 3050
rect 16776 3016 16777 3042
rect 16784 3016 16811 3042
rect 16719 2998 16749 3012
rect 16776 3008 16811 3016
rect 16813 3042 16854 3050
rect 16813 3016 16828 3042
rect 16835 3016 16854 3042
rect 16918 3038 16949 3050
rect 16964 3038 17067 3050
rect 17079 3040 17105 3066
rect 17120 3061 17150 3072
rect 17182 3068 17244 3084
rect 17182 3066 17228 3068
rect 17182 3050 17244 3066
rect 17256 3050 17262 3098
rect 17265 3090 17345 3098
rect 17265 3088 17284 3090
rect 17299 3088 17333 3090
rect 17265 3072 17345 3088
rect 17265 3050 17284 3072
rect 17299 3056 17329 3072
rect 17357 3066 17363 3140
rect 17366 3066 17385 3210
rect 17400 3066 17406 3210
rect 17415 3140 17428 3210
rect 17480 3206 17502 3210
rect 17473 3184 17502 3198
rect 17555 3184 17571 3198
rect 17609 3194 17615 3196
rect 17622 3194 17730 3210
rect 17737 3194 17743 3196
rect 17751 3194 17766 3210
rect 17832 3204 17851 3207
rect 17473 3182 17571 3184
rect 17598 3182 17766 3194
rect 17781 3184 17797 3198
rect 17832 3185 17854 3204
rect 17864 3198 17880 3199
rect 17863 3196 17880 3198
rect 17864 3191 17880 3196
rect 17854 3184 17860 3185
rect 17863 3184 17892 3191
rect 17781 3183 17892 3184
rect 17781 3182 17898 3183
rect 17457 3174 17508 3182
rect 17555 3174 17589 3182
rect 17457 3162 17482 3174
rect 17489 3162 17508 3174
rect 17562 3172 17589 3174
rect 17598 3172 17819 3182
rect 17854 3179 17860 3182
rect 17562 3168 17819 3172
rect 17457 3154 17508 3162
rect 17555 3154 17819 3168
rect 17863 3174 17898 3182
rect 17409 3106 17428 3140
rect 17473 3146 17502 3154
rect 17473 3140 17490 3146
rect 17473 3138 17507 3140
rect 17555 3138 17571 3154
rect 17572 3144 17780 3154
rect 17781 3144 17797 3154
rect 17845 3150 17860 3165
rect 17863 3162 17864 3174
rect 17871 3162 17898 3174
rect 17863 3154 17898 3162
rect 17863 3153 17892 3154
rect 17583 3140 17797 3144
rect 17598 3138 17797 3140
rect 17832 3140 17845 3150
rect 17863 3140 17880 3153
rect 17832 3138 17880 3140
rect 17474 3134 17507 3138
rect 17470 3132 17507 3134
rect 17470 3131 17537 3132
rect 17470 3126 17501 3131
rect 17507 3126 17537 3131
rect 17470 3122 17537 3126
rect 17443 3119 17537 3122
rect 17443 3112 17492 3119
rect 17443 3106 17473 3112
rect 17492 3107 17497 3112
rect 17409 3090 17489 3106
rect 17501 3098 17537 3119
rect 17598 3114 17787 3138
rect 17832 3137 17879 3138
rect 17845 3132 17879 3137
rect 17613 3111 17787 3114
rect 17606 3108 17787 3111
rect 17815 3131 17879 3132
rect 17409 3088 17428 3090
rect 17443 3088 17477 3090
rect 17409 3072 17489 3088
rect 17409 3066 17428 3072
rect 17125 3040 17228 3050
rect 17079 3038 17228 3040
rect 17249 3038 17284 3050
rect 16918 3036 17080 3038
rect 16930 3016 16949 3036
rect 16964 3034 16994 3036
rect 16813 3008 16854 3016
rect 16936 3012 16949 3016
rect 17001 3020 17080 3036
rect 17112 3036 17284 3038
rect 17112 3020 17191 3036
rect 17198 3034 17228 3036
rect 16776 2998 16805 3008
rect 16819 2998 16848 3008
rect 16863 2998 16893 3012
rect 16936 2998 16979 3012
rect 17001 3008 17191 3020
rect 17256 3016 17262 3036
rect 16986 2998 17016 3008
rect 17017 2998 17175 3008
rect 17179 2998 17209 3008
rect 17213 2998 17243 3012
rect 17271 2998 17284 3036
rect 17356 3050 17385 3066
rect 17399 3050 17428 3066
rect 17443 3056 17473 3072
rect 17501 3050 17507 3098
rect 17510 3092 17529 3098
rect 17544 3092 17574 3100
rect 17510 3084 17574 3092
rect 17510 3068 17590 3084
rect 17606 3077 17668 3108
rect 17684 3077 17746 3108
rect 17815 3106 17864 3131
rect 17879 3106 17909 3122
rect 17778 3092 17808 3100
rect 17815 3098 17925 3106
rect 17778 3084 17823 3092
rect 17510 3066 17529 3068
rect 17544 3066 17590 3068
rect 17510 3050 17590 3066
rect 17617 3064 17652 3077
rect 17693 3074 17730 3077
rect 17693 3072 17735 3074
rect 17622 3061 17652 3064
rect 17631 3057 17638 3061
rect 17638 3056 17639 3057
rect 17597 3050 17607 3056
rect 17356 3042 17391 3050
rect 17356 3016 17357 3042
rect 17364 3016 17391 3042
rect 17299 2998 17329 3012
rect 17356 3008 17391 3016
rect 17393 3042 17434 3050
rect 17393 3016 17408 3042
rect 17415 3016 17434 3042
rect 17498 3038 17529 3050
rect 17544 3038 17647 3050
rect 17659 3040 17685 3066
rect 17700 3061 17730 3072
rect 17762 3068 17824 3084
rect 17762 3066 17808 3068
rect 17762 3050 17824 3066
rect 17836 3050 17842 3098
rect 17845 3090 17925 3098
rect 17845 3088 17864 3090
rect 17879 3088 17913 3090
rect 17845 3072 17925 3088
rect 17845 3050 17864 3072
rect 17879 3056 17909 3072
rect 17937 3066 17943 3140
rect 17946 3066 17965 3210
rect 17980 3066 17986 3210
rect 17995 3140 18008 3210
rect 18060 3206 18082 3210
rect 18053 3184 18082 3198
rect 18135 3184 18151 3198
rect 18189 3194 18195 3196
rect 18202 3194 18310 3210
rect 18317 3194 18323 3196
rect 18331 3194 18346 3210
rect 18412 3204 18431 3207
rect 18053 3182 18151 3184
rect 18178 3182 18346 3194
rect 18361 3184 18377 3198
rect 18412 3185 18434 3204
rect 18444 3198 18460 3199
rect 18443 3196 18460 3198
rect 18444 3191 18460 3196
rect 18434 3184 18440 3185
rect 18443 3184 18472 3191
rect 18361 3183 18472 3184
rect 18361 3182 18478 3183
rect 18037 3174 18088 3182
rect 18135 3174 18169 3182
rect 18037 3162 18062 3174
rect 18069 3162 18088 3174
rect 18142 3172 18169 3174
rect 18178 3172 18399 3182
rect 18434 3179 18440 3182
rect 18142 3168 18399 3172
rect 18037 3154 18088 3162
rect 18135 3154 18399 3168
rect 18443 3174 18478 3182
rect 17989 3106 18008 3140
rect 18053 3146 18082 3154
rect 18053 3140 18070 3146
rect 18053 3138 18087 3140
rect 18135 3138 18151 3154
rect 18152 3144 18360 3154
rect 18361 3144 18377 3154
rect 18425 3150 18440 3165
rect 18443 3162 18444 3174
rect 18451 3162 18478 3174
rect 18443 3154 18478 3162
rect 18443 3153 18472 3154
rect 18163 3140 18377 3144
rect 18178 3138 18377 3140
rect 18412 3140 18425 3150
rect 18443 3140 18460 3153
rect 18412 3138 18460 3140
rect 18054 3134 18087 3138
rect 18050 3132 18087 3134
rect 18050 3131 18117 3132
rect 18050 3126 18081 3131
rect 18087 3126 18117 3131
rect 18050 3122 18117 3126
rect 18023 3119 18117 3122
rect 18023 3112 18072 3119
rect 18023 3106 18053 3112
rect 18072 3107 18077 3112
rect 17989 3090 18069 3106
rect 18081 3098 18117 3119
rect 18178 3114 18367 3138
rect 18412 3137 18459 3138
rect 18425 3132 18459 3137
rect 18193 3111 18367 3114
rect 18186 3108 18367 3111
rect 18395 3131 18459 3132
rect 17989 3088 18008 3090
rect 18023 3088 18057 3090
rect 17989 3072 18069 3088
rect 17989 3066 18008 3072
rect 17705 3040 17808 3050
rect 17659 3038 17808 3040
rect 17829 3038 17864 3050
rect 17498 3036 17660 3038
rect 17510 3016 17529 3036
rect 17544 3034 17574 3036
rect 17393 3008 17434 3016
rect 17516 3012 17529 3016
rect 17581 3020 17660 3036
rect 17692 3036 17864 3038
rect 17692 3020 17771 3036
rect 17778 3034 17808 3036
rect 17356 2998 17385 3008
rect 17399 2998 17428 3008
rect 17443 2998 17473 3012
rect 17516 2998 17559 3012
rect 17581 3008 17771 3020
rect 17836 3016 17842 3036
rect 17566 2998 17596 3008
rect 17597 2998 17755 3008
rect 17759 2998 17789 3008
rect 17793 2998 17823 3012
rect 17851 2998 17864 3036
rect 17936 3050 17965 3066
rect 17979 3050 18008 3066
rect 18023 3056 18053 3072
rect 18081 3050 18087 3098
rect 18090 3092 18109 3098
rect 18124 3092 18154 3100
rect 18090 3084 18154 3092
rect 18090 3068 18170 3084
rect 18186 3077 18248 3108
rect 18264 3077 18326 3108
rect 18395 3106 18444 3131
rect 18459 3106 18489 3122
rect 18358 3092 18388 3100
rect 18395 3098 18505 3106
rect 18358 3084 18403 3092
rect 18090 3066 18109 3068
rect 18124 3066 18170 3068
rect 18090 3050 18170 3066
rect 18197 3064 18232 3077
rect 18273 3074 18310 3077
rect 18273 3072 18315 3074
rect 18202 3061 18232 3064
rect 18211 3057 18218 3061
rect 18218 3056 18219 3057
rect 18177 3050 18187 3056
rect 17936 3042 17971 3050
rect 17936 3016 17937 3042
rect 17944 3016 17971 3042
rect 17879 2998 17909 3012
rect 17936 3008 17971 3016
rect 17973 3042 18014 3050
rect 17973 3016 17988 3042
rect 17995 3016 18014 3042
rect 18078 3038 18109 3050
rect 18124 3038 18227 3050
rect 18239 3040 18265 3066
rect 18280 3061 18310 3072
rect 18342 3068 18404 3084
rect 18342 3066 18388 3068
rect 18342 3050 18404 3066
rect 18416 3050 18422 3098
rect 18425 3090 18505 3098
rect 18425 3088 18444 3090
rect 18459 3088 18493 3090
rect 18425 3072 18505 3088
rect 18425 3050 18444 3072
rect 18459 3056 18489 3072
rect 18517 3066 18523 3140
rect 18532 3066 18545 3210
rect 18285 3040 18388 3050
rect 18239 3038 18388 3040
rect 18409 3038 18444 3050
rect 18078 3036 18240 3038
rect 18090 3016 18109 3036
rect 18124 3034 18154 3036
rect 17973 3008 18014 3016
rect 18096 3012 18109 3016
rect 18161 3020 18240 3036
rect 18272 3036 18444 3038
rect 18272 3020 18351 3036
rect 18358 3034 18388 3036
rect 17936 2998 17965 3008
rect 17979 2998 18008 3008
rect 18023 2998 18053 3012
rect 18096 2998 18139 3012
rect 18161 3008 18351 3020
rect 18416 3016 18422 3036
rect 18146 2998 18176 3008
rect 18177 2998 18335 3008
rect 18339 2998 18369 3008
rect 18373 2998 18403 3012
rect 18431 2998 18444 3036
rect 18516 3050 18545 3066
rect 18516 3042 18551 3050
rect 18516 3016 18517 3042
rect 18524 3016 18551 3042
rect 18459 2998 18489 3012
rect 18516 3008 18551 3016
rect 18516 2998 18545 3008
rect -1 2992 18545 2998
rect 0 2984 18545 2992
rect 15 2954 28 2984
rect 43 2970 73 2984
rect 116 2970 159 2984
rect 166 2970 386 2984
rect 393 2970 423 2984
rect 83 2956 98 2968
rect 117 2956 130 2970
rect 198 2966 351 2970
rect 80 2954 102 2956
rect 180 2954 372 2966
rect 451 2954 464 2984
rect 479 2970 509 2984
rect 546 2954 565 2984
rect 580 2954 586 2984
rect 595 2954 608 2984
rect 623 2970 653 2984
rect 696 2970 739 2984
rect 746 2970 966 2984
rect 973 2970 1003 2984
rect 663 2956 678 2968
rect 697 2956 710 2970
rect 778 2966 931 2970
rect 660 2954 682 2956
rect 760 2954 952 2966
rect 1031 2954 1044 2984
rect 1059 2970 1089 2984
rect 1126 2954 1145 2984
rect 1160 2954 1166 2984
rect 1175 2954 1188 2984
rect 1203 2970 1233 2984
rect 1276 2970 1319 2984
rect 1326 2970 1546 2984
rect 1553 2970 1583 2984
rect 1243 2956 1258 2968
rect 1277 2956 1290 2970
rect 1358 2966 1511 2970
rect 1240 2954 1262 2956
rect 1340 2954 1532 2966
rect 1611 2954 1624 2984
rect 1639 2970 1669 2984
rect 1706 2954 1725 2984
rect 1740 2954 1746 2984
rect 1755 2954 1768 2984
rect 1783 2970 1813 2984
rect 1856 2970 1899 2984
rect 1906 2970 2126 2984
rect 2133 2970 2163 2984
rect 1823 2956 1838 2968
rect 1857 2956 1870 2970
rect 1938 2966 2091 2970
rect 1820 2954 1842 2956
rect 1920 2954 2112 2966
rect 2191 2954 2204 2984
rect 2219 2970 2249 2984
rect 2286 2954 2305 2984
rect 2320 2954 2326 2984
rect 2335 2954 2348 2984
rect 2363 2970 2393 2984
rect 2436 2970 2479 2984
rect 2486 2970 2706 2984
rect 2713 2970 2743 2984
rect 2403 2956 2418 2968
rect 2437 2956 2450 2970
rect 2518 2966 2671 2970
rect 2400 2954 2422 2956
rect 2500 2954 2692 2966
rect 2771 2954 2784 2984
rect 2799 2970 2829 2984
rect 2866 2954 2885 2984
rect 2900 2954 2906 2984
rect 2915 2954 2928 2984
rect 2943 2970 2973 2984
rect 3016 2970 3059 2984
rect 3066 2970 3286 2984
rect 3293 2970 3323 2984
rect 2983 2956 2998 2968
rect 3017 2956 3030 2970
rect 3098 2966 3251 2970
rect 2980 2954 3002 2956
rect 3080 2954 3272 2966
rect 3351 2954 3364 2984
rect 3379 2970 3409 2984
rect 3446 2954 3465 2984
rect 3480 2954 3486 2984
rect 3495 2954 3508 2984
rect 3523 2970 3553 2984
rect 3596 2970 3639 2984
rect 3646 2970 3866 2984
rect 3873 2970 3903 2984
rect 3563 2956 3578 2968
rect 3597 2956 3610 2970
rect 3678 2966 3831 2970
rect 3560 2954 3582 2956
rect 3660 2954 3852 2966
rect 3931 2954 3944 2984
rect 3959 2970 3989 2984
rect 4026 2954 4045 2984
rect 4060 2954 4066 2984
rect 4075 2954 4088 2984
rect 4103 2970 4133 2984
rect 4176 2970 4219 2984
rect 4226 2970 4446 2984
rect 4453 2970 4483 2984
rect 4143 2956 4158 2968
rect 4177 2956 4190 2970
rect 4258 2966 4411 2970
rect 4140 2954 4162 2956
rect 4240 2954 4432 2966
rect 4511 2954 4524 2984
rect 4539 2970 4569 2984
rect 4606 2954 4625 2984
rect 4640 2954 4646 2984
rect 4655 2954 4668 2984
rect 4683 2970 4713 2984
rect 4756 2970 4799 2984
rect 4806 2970 5026 2984
rect 5033 2970 5063 2984
rect 4723 2956 4738 2968
rect 4757 2956 4770 2970
rect 4838 2966 4991 2970
rect 4720 2954 4742 2956
rect 4820 2954 5012 2966
rect 5091 2954 5104 2984
rect 5119 2970 5149 2984
rect 5186 2954 5205 2984
rect 5220 2954 5226 2984
rect 5235 2954 5248 2984
rect 5263 2970 5293 2984
rect 5336 2970 5379 2984
rect 5386 2970 5606 2984
rect 5613 2970 5643 2984
rect 5303 2956 5318 2968
rect 5337 2956 5350 2970
rect 5418 2966 5571 2970
rect 5300 2954 5322 2956
rect 5400 2954 5592 2966
rect 5671 2954 5684 2984
rect 5699 2970 5729 2984
rect 5766 2954 5785 2984
rect 5800 2954 5806 2984
rect 5815 2954 5828 2984
rect 5843 2970 5873 2984
rect 5916 2970 5959 2984
rect 5966 2970 6186 2984
rect 6193 2970 6223 2984
rect 5883 2956 5898 2968
rect 5917 2956 5930 2970
rect 5998 2966 6151 2970
rect 5880 2954 5902 2956
rect 5980 2954 6172 2966
rect 6251 2954 6264 2984
rect 6279 2970 6309 2984
rect 6346 2954 6365 2984
rect 6380 2954 6386 2984
rect 6395 2954 6408 2984
rect 6423 2970 6453 2984
rect 6496 2970 6539 2984
rect 6546 2970 6766 2984
rect 6773 2970 6803 2984
rect 6463 2956 6478 2968
rect 6497 2956 6510 2970
rect 6578 2966 6731 2970
rect 6460 2954 6482 2956
rect 6560 2954 6752 2966
rect 6831 2954 6844 2984
rect 6859 2970 6889 2984
rect 6926 2954 6945 2984
rect 6960 2954 6966 2984
rect 6975 2954 6988 2984
rect 7003 2970 7033 2984
rect 7076 2970 7119 2984
rect 7126 2970 7346 2984
rect 7353 2970 7383 2984
rect 7043 2956 7058 2968
rect 7077 2956 7090 2970
rect 7158 2966 7311 2970
rect 7040 2954 7062 2956
rect 7140 2954 7332 2966
rect 7411 2954 7424 2984
rect 7439 2970 7469 2984
rect 7506 2954 7525 2984
rect 7540 2954 7546 2984
rect 7555 2954 7568 2984
rect 7583 2970 7613 2984
rect 7656 2970 7699 2984
rect 7706 2970 7926 2984
rect 7933 2970 7963 2984
rect 7623 2956 7638 2968
rect 7657 2956 7670 2970
rect 7738 2966 7891 2970
rect 7620 2954 7642 2956
rect 7720 2954 7912 2966
rect 7991 2954 8004 2984
rect 8019 2970 8049 2984
rect 8086 2954 8105 2984
rect 8120 2954 8126 2984
rect 8135 2954 8148 2984
rect 8163 2970 8193 2984
rect 8236 2970 8279 2984
rect 8286 2970 8506 2984
rect 8513 2970 8543 2984
rect 8203 2956 8218 2968
rect 8237 2956 8250 2970
rect 8318 2966 8471 2970
rect 8200 2954 8222 2956
rect 8300 2954 8492 2966
rect 8571 2954 8584 2984
rect 8599 2970 8629 2984
rect 8666 2954 8685 2984
rect 8700 2954 8706 2984
rect 8715 2954 8728 2984
rect 8743 2970 8773 2984
rect 8816 2970 8859 2984
rect 8866 2970 9086 2984
rect 9093 2970 9123 2984
rect 8783 2956 8798 2968
rect 8817 2956 8830 2970
rect 8898 2966 9051 2970
rect 8780 2954 8802 2956
rect 8880 2954 9072 2966
rect 9151 2954 9164 2984
rect 9179 2970 9209 2984
rect 9246 2954 9265 2984
rect 9280 2954 9286 2984
rect 9295 2954 9308 2984
rect 9323 2970 9353 2984
rect 9396 2970 9439 2984
rect 9446 2970 9666 2984
rect 9673 2970 9703 2984
rect 9363 2956 9378 2968
rect 9397 2956 9410 2970
rect 9478 2966 9631 2970
rect 9360 2954 9382 2956
rect 9460 2954 9652 2966
rect 9731 2954 9744 2984
rect 9759 2970 9789 2984
rect 9826 2954 9845 2984
rect 9860 2954 9866 2984
rect 9875 2954 9888 2984
rect 9903 2970 9933 2984
rect 9976 2970 10019 2984
rect 10026 2970 10246 2984
rect 10253 2970 10283 2984
rect 9943 2956 9958 2968
rect 9977 2956 9990 2970
rect 10058 2966 10211 2970
rect 9940 2954 9962 2956
rect 10040 2954 10232 2966
rect 10311 2954 10324 2984
rect 10339 2970 10369 2984
rect 10406 2954 10425 2984
rect 10440 2954 10446 2984
rect 10455 2954 10468 2984
rect 10483 2970 10513 2984
rect 10556 2970 10599 2984
rect 10606 2970 10826 2984
rect 10833 2970 10863 2984
rect 10523 2956 10538 2968
rect 10557 2956 10570 2970
rect 10638 2966 10791 2970
rect 10520 2954 10542 2956
rect 10620 2954 10812 2966
rect 10891 2954 10904 2984
rect 10919 2970 10949 2984
rect 10986 2954 11005 2984
rect 11020 2954 11026 2984
rect 11035 2954 11048 2984
rect 11063 2970 11093 2984
rect 11136 2970 11179 2984
rect 11186 2970 11406 2984
rect 11413 2970 11443 2984
rect 11103 2956 11118 2968
rect 11137 2956 11150 2970
rect 11218 2966 11371 2970
rect 11100 2954 11122 2956
rect 11200 2954 11392 2966
rect 11471 2954 11484 2984
rect 11499 2970 11529 2984
rect 11566 2954 11585 2984
rect 11600 2954 11606 2984
rect 11615 2954 11628 2984
rect 11643 2970 11673 2984
rect 11716 2970 11759 2984
rect 11766 2970 11986 2984
rect 11993 2970 12023 2984
rect 11683 2956 11698 2968
rect 11717 2956 11730 2970
rect 11798 2966 11951 2970
rect 11680 2954 11702 2956
rect 11780 2954 11972 2966
rect 12051 2954 12064 2984
rect 12079 2970 12109 2984
rect 12146 2954 12165 2984
rect 12180 2954 12186 2984
rect 12195 2954 12208 2984
rect 12223 2970 12253 2984
rect 12296 2970 12339 2984
rect 12346 2970 12566 2984
rect 12573 2970 12603 2984
rect 12263 2956 12278 2968
rect 12297 2956 12310 2970
rect 12378 2966 12531 2970
rect 12260 2954 12282 2956
rect 12360 2954 12552 2966
rect 12631 2954 12644 2984
rect 12659 2970 12689 2984
rect 12726 2954 12745 2984
rect 12760 2954 12766 2984
rect 12775 2954 12788 2984
rect 12803 2970 12833 2984
rect 12876 2970 12919 2984
rect 12926 2970 13146 2984
rect 13153 2970 13183 2984
rect 12843 2956 12858 2968
rect 12877 2956 12890 2970
rect 12958 2966 13111 2970
rect 12840 2954 12862 2956
rect 12940 2954 13132 2966
rect 13211 2954 13224 2984
rect 13239 2970 13269 2984
rect 13306 2954 13325 2984
rect 13340 2954 13346 2984
rect 13355 2954 13368 2984
rect 13383 2970 13413 2984
rect 13456 2970 13499 2984
rect 13506 2970 13726 2984
rect 13733 2970 13763 2984
rect 13423 2956 13438 2968
rect 13457 2956 13470 2970
rect 13538 2966 13691 2970
rect 13420 2954 13442 2956
rect 13520 2954 13712 2966
rect 13791 2954 13804 2984
rect 13819 2970 13849 2984
rect 13886 2954 13905 2984
rect 13920 2954 13926 2984
rect 13935 2954 13948 2984
rect 13963 2970 13993 2984
rect 14036 2970 14079 2984
rect 14086 2970 14306 2984
rect 14313 2970 14343 2984
rect 14003 2956 14018 2968
rect 14037 2956 14050 2970
rect 14118 2966 14271 2970
rect 14000 2954 14022 2956
rect 14100 2954 14292 2966
rect 14371 2954 14384 2984
rect 14399 2970 14429 2984
rect 14466 2954 14485 2984
rect 14500 2954 14506 2984
rect 14515 2954 14528 2984
rect 14543 2970 14573 2984
rect 14616 2970 14659 2984
rect 14666 2970 14886 2984
rect 14893 2970 14923 2984
rect 14583 2956 14598 2968
rect 14617 2956 14630 2970
rect 14698 2966 14851 2970
rect 14580 2954 14602 2956
rect 14680 2954 14872 2966
rect 14951 2954 14964 2984
rect 14979 2970 15009 2984
rect 15046 2954 15065 2984
rect 15080 2954 15086 2984
rect 15095 2954 15108 2984
rect 15123 2970 15153 2984
rect 15196 2970 15239 2984
rect 15246 2970 15466 2984
rect 15473 2970 15503 2984
rect 15163 2956 15178 2968
rect 15197 2956 15210 2970
rect 15278 2966 15431 2970
rect 15160 2954 15182 2956
rect 15260 2954 15452 2966
rect 15531 2954 15544 2984
rect 15559 2970 15589 2984
rect 15626 2954 15645 2984
rect 15660 2954 15666 2984
rect 15675 2954 15688 2984
rect 15703 2970 15733 2984
rect 15776 2970 15819 2984
rect 15826 2970 16046 2984
rect 16053 2970 16083 2984
rect 15743 2956 15758 2968
rect 15777 2956 15790 2970
rect 15858 2966 16011 2970
rect 15740 2954 15762 2956
rect 15840 2954 16032 2966
rect 16111 2954 16124 2984
rect 16139 2970 16169 2984
rect 16206 2954 16225 2984
rect 16240 2954 16246 2984
rect 16255 2954 16268 2984
rect 16283 2970 16313 2984
rect 16356 2970 16399 2984
rect 16406 2970 16626 2984
rect 16633 2970 16663 2984
rect 16323 2956 16338 2968
rect 16357 2956 16370 2970
rect 16438 2966 16591 2970
rect 16320 2954 16342 2956
rect 16420 2954 16612 2966
rect 16691 2954 16704 2984
rect 16719 2970 16749 2984
rect 16786 2954 16805 2984
rect 16820 2954 16826 2984
rect 16835 2954 16848 2984
rect 16863 2970 16893 2984
rect 16936 2970 16979 2984
rect 16986 2970 17206 2984
rect 17213 2970 17243 2984
rect 16903 2956 16918 2968
rect 16937 2956 16950 2970
rect 17018 2966 17171 2970
rect 16900 2954 16922 2956
rect 17000 2954 17192 2966
rect 17271 2954 17284 2984
rect 17299 2970 17329 2984
rect 17366 2954 17385 2984
rect 17400 2954 17406 2984
rect 17415 2954 17428 2984
rect 17443 2970 17473 2984
rect 17516 2970 17559 2984
rect 17566 2970 17786 2984
rect 17793 2970 17823 2984
rect 17483 2956 17498 2968
rect 17517 2956 17530 2970
rect 17598 2966 17751 2970
rect 17480 2954 17502 2956
rect 17580 2954 17772 2966
rect 17851 2954 17864 2984
rect 17879 2970 17909 2984
rect 17946 2954 17965 2984
rect 17980 2954 17986 2984
rect 17995 2954 18008 2984
rect 18023 2970 18053 2984
rect 18096 2970 18139 2984
rect 18146 2970 18366 2984
rect 18373 2970 18403 2984
rect 18063 2956 18078 2968
rect 18097 2956 18110 2970
rect 18178 2966 18331 2970
rect 18060 2954 18082 2956
rect 18160 2954 18352 2966
rect 18431 2954 18444 2984
rect 18459 2970 18489 2984
rect 18532 2954 18545 2984
rect 0 2940 18545 2954
rect 15 2870 28 2940
rect 80 2936 102 2940
rect 73 2914 102 2928
rect 155 2914 171 2928
rect 209 2924 215 2926
rect 222 2924 330 2940
rect 337 2924 343 2926
rect 351 2924 366 2940
rect 432 2934 451 2937
rect 73 2912 171 2914
rect 198 2912 366 2924
rect 381 2914 397 2928
rect 432 2915 454 2934
rect 464 2928 480 2929
rect 463 2926 480 2928
rect 464 2921 480 2926
rect 454 2914 460 2915
rect 463 2914 492 2921
rect 381 2913 492 2914
rect 381 2912 498 2913
rect 57 2904 108 2912
rect 155 2904 189 2912
rect 57 2892 82 2904
rect 89 2892 108 2904
rect 162 2902 189 2904
rect 198 2902 419 2912
rect 454 2909 460 2912
rect 162 2898 419 2902
rect 57 2884 108 2892
rect 155 2884 419 2898
rect 463 2904 498 2912
rect 9 2836 28 2870
rect 73 2876 102 2884
rect 73 2870 90 2876
rect 73 2868 107 2870
rect 155 2868 171 2884
rect 172 2874 380 2884
rect 381 2874 397 2884
rect 445 2880 460 2895
rect 463 2892 464 2904
rect 471 2892 498 2904
rect 463 2884 498 2892
rect 463 2883 492 2884
rect 183 2870 397 2874
rect 198 2868 397 2870
rect 432 2870 445 2880
rect 463 2870 480 2883
rect 432 2868 480 2870
rect 74 2864 107 2868
rect 70 2862 107 2864
rect 70 2861 137 2862
rect 70 2856 101 2861
rect 107 2856 137 2861
rect 70 2852 137 2856
rect 43 2849 137 2852
rect 43 2842 92 2849
rect 43 2836 73 2842
rect 92 2837 97 2842
rect 9 2820 89 2836
rect 101 2828 137 2849
rect 198 2844 387 2868
rect 432 2867 479 2868
rect 445 2862 479 2867
rect 213 2841 387 2844
rect 206 2838 387 2841
rect 415 2861 479 2862
rect 9 2818 28 2820
rect 43 2818 77 2820
rect 9 2802 89 2818
rect 9 2796 28 2802
rect -1 2780 28 2796
rect 43 2786 73 2802
rect 101 2780 107 2828
rect 110 2822 129 2828
rect 144 2822 174 2830
rect 110 2814 174 2822
rect 110 2798 190 2814
rect 206 2807 268 2838
rect 284 2807 346 2838
rect 415 2836 464 2861
rect 479 2836 509 2852
rect 378 2822 408 2830
rect 415 2828 525 2836
rect 378 2814 423 2822
rect 110 2796 129 2798
rect 144 2796 190 2798
rect 110 2780 190 2796
rect 217 2794 252 2807
rect 293 2804 330 2807
rect 293 2802 335 2804
rect 222 2791 252 2794
rect 231 2787 238 2791
rect 238 2786 239 2787
rect 197 2780 207 2786
rect -7 2772 34 2780
rect -7 2746 8 2772
rect 15 2746 34 2772
rect 98 2768 129 2780
rect 144 2768 247 2780
rect 259 2770 285 2796
rect 300 2791 330 2802
rect 362 2798 424 2814
rect 362 2796 408 2798
rect 362 2780 424 2796
rect 436 2780 442 2828
rect 445 2820 525 2828
rect 445 2818 464 2820
rect 479 2818 513 2820
rect 445 2802 525 2818
rect 445 2780 464 2802
rect 479 2786 509 2802
rect 537 2796 543 2870
rect 546 2796 565 2940
rect 580 2796 586 2940
rect 595 2870 608 2940
rect 660 2936 682 2940
rect 653 2914 682 2928
rect 735 2914 751 2928
rect 789 2924 795 2926
rect 802 2924 910 2940
rect 917 2924 923 2926
rect 931 2924 946 2940
rect 1012 2934 1031 2937
rect 653 2912 751 2914
rect 778 2912 946 2924
rect 961 2914 977 2928
rect 1012 2915 1034 2934
rect 1044 2928 1060 2929
rect 1043 2926 1060 2928
rect 1044 2921 1060 2926
rect 1034 2914 1040 2915
rect 1043 2914 1072 2921
rect 961 2913 1072 2914
rect 961 2912 1078 2913
rect 637 2904 688 2912
rect 735 2904 769 2912
rect 637 2892 662 2904
rect 669 2892 688 2904
rect 742 2902 769 2904
rect 778 2902 999 2912
rect 1034 2909 1040 2912
rect 742 2898 999 2902
rect 637 2884 688 2892
rect 735 2884 999 2898
rect 1043 2904 1078 2912
rect 589 2836 608 2870
rect 653 2876 682 2884
rect 653 2870 670 2876
rect 653 2868 687 2870
rect 735 2868 751 2884
rect 752 2874 960 2884
rect 961 2874 977 2884
rect 1025 2880 1040 2895
rect 1043 2892 1044 2904
rect 1051 2892 1078 2904
rect 1043 2884 1078 2892
rect 1043 2883 1072 2884
rect 763 2870 977 2874
rect 778 2868 977 2870
rect 1012 2870 1025 2880
rect 1043 2870 1060 2883
rect 1012 2868 1060 2870
rect 654 2864 687 2868
rect 650 2862 687 2864
rect 650 2861 717 2862
rect 650 2856 681 2861
rect 687 2856 717 2861
rect 650 2852 717 2856
rect 623 2849 717 2852
rect 623 2842 672 2849
rect 623 2836 653 2842
rect 672 2837 677 2842
rect 589 2820 669 2836
rect 681 2828 717 2849
rect 778 2844 967 2868
rect 1012 2867 1059 2868
rect 1025 2862 1059 2867
rect 793 2841 967 2844
rect 786 2838 967 2841
rect 995 2861 1059 2862
rect 589 2818 608 2820
rect 623 2818 657 2820
rect 589 2802 669 2818
rect 589 2796 608 2802
rect 305 2770 408 2780
rect 259 2768 408 2770
rect 429 2768 464 2780
rect 98 2766 260 2768
rect 110 2746 129 2766
rect 144 2764 174 2766
rect -7 2738 34 2746
rect 116 2742 129 2746
rect 181 2750 260 2766
rect 292 2766 464 2768
rect 292 2750 371 2766
rect 378 2764 408 2766
rect -1 2728 28 2738
rect 43 2728 73 2742
rect 116 2728 159 2742
rect 181 2738 371 2750
rect 436 2746 442 2766
rect 166 2728 196 2738
rect 197 2728 355 2738
rect 359 2728 389 2738
rect 393 2728 423 2742
rect 451 2728 464 2766
rect 536 2780 565 2796
rect 579 2780 608 2796
rect 623 2786 653 2802
rect 681 2780 687 2828
rect 690 2822 709 2828
rect 724 2822 754 2830
rect 690 2814 754 2822
rect 690 2798 770 2814
rect 786 2807 848 2838
rect 864 2807 926 2838
rect 995 2836 1044 2861
rect 1059 2836 1089 2852
rect 958 2822 988 2830
rect 995 2828 1105 2836
rect 958 2814 1003 2822
rect 690 2796 709 2798
rect 724 2796 770 2798
rect 690 2780 770 2796
rect 797 2794 832 2807
rect 873 2804 910 2807
rect 873 2802 915 2804
rect 802 2791 832 2794
rect 811 2787 818 2791
rect 818 2786 819 2787
rect 777 2780 787 2786
rect 536 2772 571 2780
rect 536 2746 537 2772
rect 544 2746 571 2772
rect 479 2728 509 2742
rect 536 2738 571 2746
rect 573 2772 614 2780
rect 573 2746 588 2772
rect 595 2746 614 2772
rect 678 2768 709 2780
rect 724 2768 827 2780
rect 839 2770 865 2796
rect 880 2791 910 2802
rect 942 2798 1004 2814
rect 942 2796 988 2798
rect 942 2780 1004 2796
rect 1016 2780 1022 2828
rect 1025 2820 1105 2828
rect 1025 2818 1044 2820
rect 1059 2818 1093 2820
rect 1025 2802 1105 2818
rect 1025 2780 1044 2802
rect 1059 2786 1089 2802
rect 1117 2796 1123 2870
rect 1126 2796 1145 2940
rect 1160 2796 1166 2940
rect 1175 2870 1188 2940
rect 1240 2936 1262 2940
rect 1233 2914 1262 2928
rect 1315 2914 1331 2928
rect 1369 2924 1375 2926
rect 1382 2924 1490 2940
rect 1497 2924 1503 2926
rect 1511 2924 1526 2940
rect 1592 2934 1611 2937
rect 1233 2912 1331 2914
rect 1358 2912 1526 2924
rect 1541 2914 1557 2928
rect 1592 2915 1614 2934
rect 1624 2928 1640 2929
rect 1623 2926 1640 2928
rect 1624 2921 1640 2926
rect 1614 2914 1620 2915
rect 1623 2914 1652 2921
rect 1541 2913 1652 2914
rect 1541 2912 1658 2913
rect 1217 2904 1268 2912
rect 1315 2904 1349 2912
rect 1217 2892 1242 2904
rect 1249 2892 1268 2904
rect 1322 2902 1349 2904
rect 1358 2902 1579 2912
rect 1614 2909 1620 2912
rect 1322 2898 1579 2902
rect 1217 2884 1268 2892
rect 1315 2884 1579 2898
rect 1623 2904 1658 2912
rect 1169 2836 1188 2870
rect 1233 2876 1262 2884
rect 1233 2870 1250 2876
rect 1233 2868 1267 2870
rect 1315 2868 1331 2884
rect 1332 2874 1540 2884
rect 1541 2874 1557 2884
rect 1605 2880 1620 2895
rect 1623 2892 1624 2904
rect 1631 2892 1658 2904
rect 1623 2884 1658 2892
rect 1623 2883 1652 2884
rect 1343 2870 1557 2874
rect 1358 2868 1557 2870
rect 1592 2870 1605 2880
rect 1623 2870 1640 2883
rect 1592 2868 1640 2870
rect 1234 2864 1267 2868
rect 1230 2862 1267 2864
rect 1230 2861 1297 2862
rect 1230 2856 1261 2861
rect 1267 2856 1297 2861
rect 1230 2852 1297 2856
rect 1203 2849 1297 2852
rect 1203 2842 1252 2849
rect 1203 2836 1233 2842
rect 1252 2837 1257 2842
rect 1169 2820 1249 2836
rect 1261 2828 1297 2849
rect 1358 2844 1547 2868
rect 1592 2867 1639 2868
rect 1605 2862 1639 2867
rect 1373 2841 1547 2844
rect 1366 2838 1547 2841
rect 1575 2861 1639 2862
rect 1169 2818 1188 2820
rect 1203 2818 1237 2820
rect 1169 2802 1249 2818
rect 1169 2796 1188 2802
rect 885 2770 988 2780
rect 839 2768 988 2770
rect 1009 2768 1044 2780
rect 678 2766 840 2768
rect 690 2746 709 2766
rect 724 2764 754 2766
rect 573 2738 614 2746
rect 696 2742 709 2746
rect 761 2750 840 2766
rect 872 2766 1044 2768
rect 872 2750 951 2766
rect 958 2764 988 2766
rect 536 2728 565 2738
rect 579 2728 608 2738
rect 623 2728 653 2742
rect 696 2728 739 2742
rect 761 2738 951 2750
rect 1016 2746 1022 2766
rect 746 2728 776 2738
rect 777 2728 935 2738
rect 939 2728 969 2738
rect 973 2728 1003 2742
rect 1031 2728 1044 2766
rect 1116 2780 1145 2796
rect 1159 2780 1188 2796
rect 1203 2786 1233 2802
rect 1261 2780 1267 2828
rect 1270 2822 1289 2828
rect 1304 2822 1334 2830
rect 1270 2814 1334 2822
rect 1270 2798 1350 2814
rect 1366 2807 1428 2838
rect 1444 2807 1506 2838
rect 1575 2836 1624 2861
rect 1639 2836 1669 2852
rect 1538 2822 1568 2830
rect 1575 2828 1685 2836
rect 1538 2814 1583 2822
rect 1270 2796 1289 2798
rect 1304 2796 1350 2798
rect 1270 2780 1350 2796
rect 1377 2794 1412 2807
rect 1453 2804 1490 2807
rect 1453 2802 1495 2804
rect 1382 2791 1412 2794
rect 1391 2787 1398 2791
rect 1398 2786 1399 2787
rect 1357 2780 1367 2786
rect 1116 2772 1151 2780
rect 1116 2746 1117 2772
rect 1124 2746 1151 2772
rect 1059 2728 1089 2742
rect 1116 2738 1151 2746
rect 1153 2772 1194 2780
rect 1153 2746 1168 2772
rect 1175 2746 1194 2772
rect 1258 2768 1289 2780
rect 1304 2768 1407 2780
rect 1419 2770 1445 2796
rect 1460 2791 1490 2802
rect 1522 2798 1584 2814
rect 1522 2796 1568 2798
rect 1522 2780 1584 2796
rect 1596 2780 1602 2828
rect 1605 2820 1685 2828
rect 1605 2818 1624 2820
rect 1639 2818 1673 2820
rect 1605 2802 1685 2818
rect 1605 2780 1624 2802
rect 1639 2786 1669 2802
rect 1697 2796 1703 2870
rect 1706 2796 1725 2940
rect 1740 2796 1746 2940
rect 1755 2870 1768 2940
rect 1820 2936 1842 2940
rect 1813 2914 1842 2928
rect 1895 2914 1911 2928
rect 1949 2924 1955 2926
rect 1962 2924 2070 2940
rect 2077 2924 2083 2926
rect 2091 2924 2106 2940
rect 2172 2934 2191 2937
rect 1813 2912 1911 2914
rect 1938 2912 2106 2924
rect 2121 2914 2137 2928
rect 2172 2915 2194 2934
rect 2204 2928 2220 2929
rect 2203 2926 2220 2928
rect 2204 2921 2220 2926
rect 2194 2914 2200 2915
rect 2203 2914 2232 2921
rect 2121 2913 2232 2914
rect 2121 2912 2238 2913
rect 1797 2904 1848 2912
rect 1895 2904 1929 2912
rect 1797 2892 1822 2904
rect 1829 2892 1848 2904
rect 1902 2902 1929 2904
rect 1938 2902 2159 2912
rect 2194 2909 2200 2912
rect 1902 2898 2159 2902
rect 1797 2884 1848 2892
rect 1895 2884 2159 2898
rect 2203 2904 2238 2912
rect 1749 2836 1768 2870
rect 1813 2876 1842 2884
rect 1813 2870 1830 2876
rect 1813 2868 1847 2870
rect 1895 2868 1911 2884
rect 1912 2874 2120 2884
rect 2121 2874 2137 2884
rect 2185 2880 2200 2895
rect 2203 2892 2204 2904
rect 2211 2892 2238 2904
rect 2203 2884 2238 2892
rect 2203 2883 2232 2884
rect 1923 2870 2137 2874
rect 1938 2868 2137 2870
rect 2172 2870 2185 2880
rect 2203 2870 2220 2883
rect 2172 2868 2220 2870
rect 1814 2864 1847 2868
rect 1810 2862 1847 2864
rect 1810 2861 1877 2862
rect 1810 2856 1841 2861
rect 1847 2856 1877 2861
rect 1810 2852 1877 2856
rect 1783 2849 1877 2852
rect 1783 2842 1832 2849
rect 1783 2836 1813 2842
rect 1832 2837 1837 2842
rect 1749 2820 1829 2836
rect 1841 2828 1877 2849
rect 1938 2844 2127 2868
rect 2172 2867 2219 2868
rect 2185 2862 2219 2867
rect 1953 2841 2127 2844
rect 1946 2838 2127 2841
rect 2155 2861 2219 2862
rect 1749 2818 1768 2820
rect 1783 2818 1817 2820
rect 1749 2802 1829 2818
rect 1749 2796 1768 2802
rect 1465 2770 1568 2780
rect 1419 2768 1568 2770
rect 1589 2768 1624 2780
rect 1258 2766 1420 2768
rect 1270 2746 1289 2766
rect 1304 2764 1334 2766
rect 1153 2738 1194 2746
rect 1276 2742 1289 2746
rect 1341 2750 1420 2766
rect 1452 2766 1624 2768
rect 1452 2750 1531 2766
rect 1538 2764 1568 2766
rect 1116 2728 1145 2738
rect 1159 2728 1188 2738
rect 1203 2728 1233 2742
rect 1276 2728 1319 2742
rect 1341 2738 1531 2750
rect 1596 2746 1602 2766
rect 1326 2728 1356 2738
rect 1357 2728 1515 2738
rect 1519 2728 1549 2738
rect 1553 2728 1583 2742
rect 1611 2728 1624 2766
rect 1696 2780 1725 2796
rect 1739 2780 1768 2796
rect 1783 2786 1813 2802
rect 1841 2780 1847 2828
rect 1850 2822 1869 2828
rect 1884 2822 1914 2830
rect 1850 2814 1914 2822
rect 1850 2798 1930 2814
rect 1946 2807 2008 2838
rect 2024 2807 2086 2838
rect 2155 2836 2204 2861
rect 2219 2836 2249 2852
rect 2118 2822 2148 2830
rect 2155 2828 2265 2836
rect 2118 2814 2163 2822
rect 1850 2796 1869 2798
rect 1884 2796 1930 2798
rect 1850 2780 1930 2796
rect 1957 2794 1992 2807
rect 2033 2804 2070 2807
rect 2033 2802 2075 2804
rect 1962 2791 1992 2794
rect 1971 2787 1978 2791
rect 1978 2786 1979 2787
rect 1937 2780 1947 2786
rect 1696 2772 1731 2780
rect 1696 2746 1697 2772
rect 1704 2746 1731 2772
rect 1639 2728 1669 2742
rect 1696 2738 1731 2746
rect 1733 2772 1774 2780
rect 1733 2746 1748 2772
rect 1755 2746 1774 2772
rect 1838 2768 1869 2780
rect 1884 2768 1987 2780
rect 1999 2770 2025 2796
rect 2040 2791 2070 2802
rect 2102 2798 2164 2814
rect 2102 2796 2148 2798
rect 2102 2780 2164 2796
rect 2176 2780 2182 2828
rect 2185 2820 2265 2828
rect 2185 2818 2204 2820
rect 2219 2818 2253 2820
rect 2185 2802 2265 2818
rect 2185 2780 2204 2802
rect 2219 2786 2249 2802
rect 2277 2796 2283 2870
rect 2286 2796 2305 2940
rect 2320 2796 2326 2940
rect 2335 2870 2348 2940
rect 2400 2936 2422 2940
rect 2393 2914 2422 2928
rect 2475 2914 2491 2928
rect 2529 2924 2535 2926
rect 2542 2924 2650 2940
rect 2657 2924 2663 2926
rect 2671 2924 2686 2940
rect 2752 2934 2771 2937
rect 2393 2912 2491 2914
rect 2518 2912 2686 2924
rect 2701 2914 2717 2928
rect 2752 2915 2774 2934
rect 2784 2928 2800 2929
rect 2783 2926 2800 2928
rect 2784 2921 2800 2926
rect 2774 2914 2780 2915
rect 2783 2914 2812 2921
rect 2701 2913 2812 2914
rect 2701 2912 2818 2913
rect 2377 2904 2428 2912
rect 2475 2904 2509 2912
rect 2377 2892 2402 2904
rect 2409 2892 2428 2904
rect 2482 2902 2509 2904
rect 2518 2902 2739 2912
rect 2774 2909 2780 2912
rect 2482 2898 2739 2902
rect 2377 2884 2428 2892
rect 2475 2884 2739 2898
rect 2783 2904 2818 2912
rect 2329 2836 2348 2870
rect 2393 2876 2422 2884
rect 2393 2870 2410 2876
rect 2393 2868 2427 2870
rect 2475 2868 2491 2884
rect 2492 2874 2700 2884
rect 2701 2874 2717 2884
rect 2765 2880 2780 2895
rect 2783 2892 2784 2904
rect 2791 2892 2818 2904
rect 2783 2884 2818 2892
rect 2783 2883 2812 2884
rect 2503 2870 2717 2874
rect 2518 2868 2717 2870
rect 2752 2870 2765 2880
rect 2783 2870 2800 2883
rect 2752 2868 2800 2870
rect 2394 2864 2427 2868
rect 2390 2862 2427 2864
rect 2390 2861 2457 2862
rect 2390 2856 2421 2861
rect 2427 2856 2457 2861
rect 2390 2852 2457 2856
rect 2363 2849 2457 2852
rect 2363 2842 2412 2849
rect 2363 2836 2393 2842
rect 2412 2837 2417 2842
rect 2329 2820 2409 2836
rect 2421 2828 2457 2849
rect 2518 2844 2707 2868
rect 2752 2867 2799 2868
rect 2765 2862 2799 2867
rect 2533 2841 2707 2844
rect 2526 2838 2707 2841
rect 2735 2861 2799 2862
rect 2329 2818 2348 2820
rect 2363 2818 2397 2820
rect 2329 2802 2409 2818
rect 2329 2796 2348 2802
rect 2045 2770 2148 2780
rect 1999 2768 2148 2770
rect 2169 2768 2204 2780
rect 1838 2766 2000 2768
rect 1850 2746 1869 2766
rect 1884 2764 1914 2766
rect 1733 2738 1774 2746
rect 1856 2742 1869 2746
rect 1921 2750 2000 2766
rect 2032 2766 2204 2768
rect 2032 2750 2111 2766
rect 2118 2764 2148 2766
rect 1696 2728 1725 2738
rect 1739 2728 1768 2738
rect 1783 2728 1813 2742
rect 1856 2728 1899 2742
rect 1921 2738 2111 2750
rect 2176 2746 2182 2766
rect 1906 2728 1936 2738
rect 1937 2728 2095 2738
rect 2099 2728 2129 2738
rect 2133 2728 2163 2742
rect 2191 2728 2204 2766
rect 2276 2780 2305 2796
rect 2319 2780 2348 2796
rect 2363 2786 2393 2802
rect 2421 2780 2427 2828
rect 2430 2822 2449 2828
rect 2464 2822 2494 2830
rect 2430 2814 2494 2822
rect 2430 2798 2510 2814
rect 2526 2807 2588 2838
rect 2604 2807 2666 2838
rect 2735 2836 2784 2861
rect 2799 2836 2829 2852
rect 2698 2822 2728 2830
rect 2735 2828 2845 2836
rect 2698 2814 2743 2822
rect 2430 2796 2449 2798
rect 2464 2796 2510 2798
rect 2430 2780 2510 2796
rect 2537 2794 2572 2807
rect 2613 2804 2650 2807
rect 2613 2802 2655 2804
rect 2542 2791 2572 2794
rect 2551 2787 2558 2791
rect 2558 2786 2559 2787
rect 2517 2780 2527 2786
rect 2276 2772 2311 2780
rect 2276 2746 2277 2772
rect 2284 2746 2311 2772
rect 2219 2728 2249 2742
rect 2276 2738 2311 2746
rect 2313 2772 2354 2780
rect 2313 2746 2328 2772
rect 2335 2746 2354 2772
rect 2418 2768 2449 2780
rect 2464 2768 2567 2780
rect 2579 2770 2605 2796
rect 2620 2791 2650 2802
rect 2682 2798 2744 2814
rect 2682 2796 2728 2798
rect 2682 2780 2744 2796
rect 2756 2780 2762 2828
rect 2765 2820 2845 2828
rect 2765 2818 2784 2820
rect 2799 2818 2833 2820
rect 2765 2802 2845 2818
rect 2765 2780 2784 2802
rect 2799 2786 2829 2802
rect 2857 2796 2863 2870
rect 2866 2796 2885 2940
rect 2900 2796 2906 2940
rect 2915 2870 2928 2940
rect 2980 2936 3002 2940
rect 2973 2914 3002 2928
rect 3055 2914 3071 2928
rect 3109 2924 3115 2926
rect 3122 2924 3230 2940
rect 3237 2924 3243 2926
rect 3251 2924 3266 2940
rect 3332 2934 3351 2937
rect 2973 2912 3071 2914
rect 3098 2912 3266 2924
rect 3281 2914 3297 2928
rect 3332 2915 3354 2934
rect 3364 2928 3380 2929
rect 3363 2926 3380 2928
rect 3364 2921 3380 2926
rect 3354 2914 3360 2915
rect 3363 2914 3392 2921
rect 3281 2913 3392 2914
rect 3281 2912 3398 2913
rect 2957 2904 3008 2912
rect 3055 2904 3089 2912
rect 2957 2892 2982 2904
rect 2989 2892 3008 2904
rect 3062 2902 3089 2904
rect 3098 2902 3319 2912
rect 3354 2909 3360 2912
rect 3062 2898 3319 2902
rect 2957 2884 3008 2892
rect 3055 2884 3319 2898
rect 3363 2904 3398 2912
rect 2909 2836 2928 2870
rect 2973 2876 3002 2884
rect 2973 2870 2990 2876
rect 2973 2868 3007 2870
rect 3055 2868 3071 2884
rect 3072 2874 3280 2884
rect 3281 2874 3297 2884
rect 3345 2880 3360 2895
rect 3363 2892 3364 2904
rect 3371 2892 3398 2904
rect 3363 2884 3398 2892
rect 3363 2883 3392 2884
rect 3083 2870 3297 2874
rect 3098 2868 3297 2870
rect 3332 2870 3345 2880
rect 3363 2870 3380 2883
rect 3332 2868 3380 2870
rect 2974 2864 3007 2868
rect 2970 2862 3007 2864
rect 2970 2861 3037 2862
rect 2970 2856 3001 2861
rect 3007 2856 3037 2861
rect 2970 2852 3037 2856
rect 2943 2849 3037 2852
rect 2943 2842 2992 2849
rect 2943 2836 2973 2842
rect 2992 2837 2997 2842
rect 2909 2820 2989 2836
rect 3001 2828 3037 2849
rect 3098 2844 3287 2868
rect 3332 2867 3379 2868
rect 3345 2862 3379 2867
rect 3113 2841 3287 2844
rect 3106 2838 3287 2841
rect 3315 2861 3379 2862
rect 2909 2818 2928 2820
rect 2943 2818 2977 2820
rect 2909 2802 2989 2818
rect 2909 2796 2928 2802
rect 2625 2770 2728 2780
rect 2579 2768 2728 2770
rect 2749 2768 2784 2780
rect 2418 2766 2580 2768
rect 2430 2746 2449 2766
rect 2464 2764 2494 2766
rect 2313 2738 2354 2746
rect 2436 2742 2449 2746
rect 2501 2750 2580 2766
rect 2612 2766 2784 2768
rect 2612 2750 2691 2766
rect 2698 2764 2728 2766
rect 2276 2728 2305 2738
rect 2319 2728 2348 2738
rect 2363 2728 2393 2742
rect 2436 2728 2479 2742
rect 2501 2738 2691 2750
rect 2756 2746 2762 2766
rect 2486 2728 2516 2738
rect 2517 2728 2675 2738
rect 2679 2728 2709 2738
rect 2713 2728 2743 2742
rect 2771 2728 2784 2766
rect 2856 2780 2885 2796
rect 2899 2780 2928 2796
rect 2943 2786 2973 2802
rect 3001 2780 3007 2828
rect 3010 2822 3029 2828
rect 3044 2822 3074 2830
rect 3010 2814 3074 2822
rect 3010 2798 3090 2814
rect 3106 2807 3168 2838
rect 3184 2807 3246 2838
rect 3315 2836 3364 2861
rect 3379 2836 3409 2852
rect 3278 2822 3308 2830
rect 3315 2828 3425 2836
rect 3278 2814 3323 2822
rect 3010 2796 3029 2798
rect 3044 2796 3090 2798
rect 3010 2780 3090 2796
rect 3117 2794 3152 2807
rect 3193 2804 3230 2807
rect 3193 2802 3235 2804
rect 3122 2791 3152 2794
rect 3131 2787 3138 2791
rect 3138 2786 3139 2787
rect 3097 2780 3107 2786
rect 2856 2772 2891 2780
rect 2856 2746 2857 2772
rect 2864 2746 2891 2772
rect 2799 2728 2829 2742
rect 2856 2738 2891 2746
rect 2893 2772 2934 2780
rect 2893 2746 2908 2772
rect 2915 2746 2934 2772
rect 2998 2768 3029 2780
rect 3044 2768 3147 2780
rect 3159 2770 3185 2796
rect 3200 2791 3230 2802
rect 3262 2798 3324 2814
rect 3262 2796 3308 2798
rect 3262 2780 3324 2796
rect 3336 2780 3342 2828
rect 3345 2820 3425 2828
rect 3345 2818 3364 2820
rect 3379 2818 3413 2820
rect 3345 2802 3425 2818
rect 3345 2780 3364 2802
rect 3379 2786 3409 2802
rect 3437 2796 3443 2870
rect 3446 2796 3465 2940
rect 3480 2796 3486 2940
rect 3495 2870 3508 2940
rect 3560 2936 3582 2940
rect 3553 2914 3582 2928
rect 3635 2914 3651 2928
rect 3689 2924 3695 2926
rect 3702 2924 3810 2940
rect 3817 2924 3823 2926
rect 3831 2924 3846 2940
rect 3912 2934 3931 2937
rect 3553 2912 3651 2914
rect 3678 2912 3846 2924
rect 3861 2914 3877 2928
rect 3912 2915 3934 2934
rect 3944 2928 3960 2929
rect 3943 2926 3960 2928
rect 3944 2921 3960 2926
rect 3934 2914 3940 2915
rect 3943 2914 3972 2921
rect 3861 2913 3972 2914
rect 3861 2912 3978 2913
rect 3537 2904 3588 2912
rect 3635 2904 3669 2912
rect 3537 2892 3562 2904
rect 3569 2892 3588 2904
rect 3642 2902 3669 2904
rect 3678 2902 3899 2912
rect 3934 2909 3940 2912
rect 3642 2898 3899 2902
rect 3537 2884 3588 2892
rect 3635 2884 3899 2898
rect 3943 2904 3978 2912
rect 3489 2836 3508 2870
rect 3553 2876 3582 2884
rect 3553 2870 3570 2876
rect 3553 2868 3587 2870
rect 3635 2868 3651 2884
rect 3652 2874 3860 2884
rect 3861 2874 3877 2884
rect 3925 2880 3940 2895
rect 3943 2892 3944 2904
rect 3951 2892 3978 2904
rect 3943 2884 3978 2892
rect 3943 2883 3972 2884
rect 3663 2870 3877 2874
rect 3678 2868 3877 2870
rect 3912 2870 3925 2880
rect 3943 2870 3960 2883
rect 3912 2868 3960 2870
rect 3554 2864 3587 2868
rect 3550 2862 3587 2864
rect 3550 2861 3617 2862
rect 3550 2856 3581 2861
rect 3587 2856 3617 2861
rect 3550 2852 3617 2856
rect 3523 2849 3617 2852
rect 3523 2842 3572 2849
rect 3523 2836 3553 2842
rect 3572 2837 3577 2842
rect 3489 2820 3569 2836
rect 3581 2828 3617 2849
rect 3678 2844 3867 2868
rect 3912 2867 3959 2868
rect 3925 2862 3959 2867
rect 3693 2841 3867 2844
rect 3686 2838 3867 2841
rect 3895 2861 3959 2862
rect 3489 2818 3508 2820
rect 3523 2818 3557 2820
rect 3489 2802 3569 2818
rect 3489 2796 3508 2802
rect 3205 2770 3308 2780
rect 3159 2768 3308 2770
rect 3329 2768 3364 2780
rect 2998 2766 3160 2768
rect 3010 2746 3029 2766
rect 3044 2764 3074 2766
rect 2893 2738 2934 2746
rect 3016 2742 3029 2746
rect 3081 2750 3160 2766
rect 3192 2766 3364 2768
rect 3192 2750 3271 2766
rect 3278 2764 3308 2766
rect 2856 2728 2885 2738
rect 2899 2728 2928 2738
rect 2943 2728 2973 2742
rect 3016 2728 3059 2742
rect 3081 2738 3271 2750
rect 3336 2746 3342 2766
rect 3066 2728 3096 2738
rect 3097 2728 3255 2738
rect 3259 2728 3289 2738
rect 3293 2728 3323 2742
rect 3351 2728 3364 2766
rect 3436 2780 3465 2796
rect 3479 2780 3508 2796
rect 3523 2786 3553 2802
rect 3581 2780 3587 2828
rect 3590 2822 3609 2828
rect 3624 2822 3654 2830
rect 3590 2814 3654 2822
rect 3590 2798 3670 2814
rect 3686 2807 3748 2838
rect 3764 2807 3826 2838
rect 3895 2836 3944 2861
rect 3959 2836 3989 2852
rect 3858 2822 3888 2830
rect 3895 2828 4005 2836
rect 3858 2814 3903 2822
rect 3590 2796 3609 2798
rect 3624 2796 3670 2798
rect 3590 2780 3670 2796
rect 3697 2794 3732 2807
rect 3773 2804 3810 2807
rect 3773 2802 3815 2804
rect 3702 2791 3732 2794
rect 3711 2787 3718 2791
rect 3718 2786 3719 2787
rect 3677 2780 3687 2786
rect 3436 2772 3471 2780
rect 3436 2746 3437 2772
rect 3444 2746 3471 2772
rect 3379 2728 3409 2742
rect 3436 2738 3471 2746
rect 3473 2772 3514 2780
rect 3473 2746 3488 2772
rect 3495 2746 3514 2772
rect 3578 2768 3609 2780
rect 3624 2768 3727 2780
rect 3739 2770 3765 2796
rect 3780 2791 3810 2802
rect 3842 2798 3904 2814
rect 3842 2796 3888 2798
rect 3842 2780 3904 2796
rect 3916 2780 3922 2828
rect 3925 2820 4005 2828
rect 3925 2818 3944 2820
rect 3959 2818 3993 2820
rect 3925 2802 4005 2818
rect 3925 2780 3944 2802
rect 3959 2786 3989 2802
rect 4017 2796 4023 2870
rect 4026 2796 4045 2940
rect 4060 2796 4066 2940
rect 4075 2870 4088 2940
rect 4140 2936 4162 2940
rect 4133 2914 4162 2928
rect 4215 2914 4231 2928
rect 4269 2924 4275 2926
rect 4282 2924 4390 2940
rect 4397 2924 4403 2926
rect 4411 2924 4426 2940
rect 4492 2934 4511 2937
rect 4133 2912 4231 2914
rect 4258 2912 4426 2924
rect 4441 2914 4457 2928
rect 4492 2915 4514 2934
rect 4524 2928 4540 2929
rect 4523 2926 4540 2928
rect 4524 2921 4540 2926
rect 4514 2914 4520 2915
rect 4523 2914 4552 2921
rect 4441 2913 4552 2914
rect 4441 2912 4558 2913
rect 4117 2904 4168 2912
rect 4215 2904 4249 2912
rect 4117 2892 4142 2904
rect 4149 2892 4168 2904
rect 4222 2902 4249 2904
rect 4258 2902 4479 2912
rect 4514 2909 4520 2912
rect 4222 2898 4479 2902
rect 4117 2884 4168 2892
rect 4215 2884 4479 2898
rect 4523 2904 4558 2912
rect 4069 2836 4088 2870
rect 4133 2876 4162 2884
rect 4133 2870 4150 2876
rect 4133 2868 4167 2870
rect 4215 2868 4231 2884
rect 4232 2874 4440 2884
rect 4441 2874 4457 2884
rect 4505 2880 4520 2895
rect 4523 2892 4524 2904
rect 4531 2892 4558 2904
rect 4523 2884 4558 2892
rect 4523 2883 4552 2884
rect 4243 2870 4457 2874
rect 4258 2868 4457 2870
rect 4492 2870 4505 2880
rect 4523 2870 4540 2883
rect 4492 2868 4540 2870
rect 4134 2864 4167 2868
rect 4130 2862 4167 2864
rect 4130 2861 4197 2862
rect 4130 2856 4161 2861
rect 4167 2856 4197 2861
rect 4130 2852 4197 2856
rect 4103 2849 4197 2852
rect 4103 2842 4152 2849
rect 4103 2836 4133 2842
rect 4152 2837 4157 2842
rect 4069 2820 4149 2836
rect 4161 2828 4197 2849
rect 4258 2844 4447 2868
rect 4492 2867 4539 2868
rect 4505 2862 4539 2867
rect 4273 2841 4447 2844
rect 4266 2838 4447 2841
rect 4475 2861 4539 2862
rect 4069 2818 4088 2820
rect 4103 2818 4137 2820
rect 4069 2802 4149 2818
rect 4069 2796 4088 2802
rect 3785 2770 3888 2780
rect 3739 2768 3888 2770
rect 3909 2768 3944 2780
rect 3578 2766 3740 2768
rect 3590 2746 3609 2766
rect 3624 2764 3654 2766
rect 3473 2738 3514 2746
rect 3596 2742 3609 2746
rect 3661 2750 3740 2766
rect 3772 2766 3944 2768
rect 3772 2750 3851 2766
rect 3858 2764 3888 2766
rect 3436 2728 3465 2738
rect 3479 2728 3508 2738
rect 3523 2728 3553 2742
rect 3596 2728 3639 2742
rect 3661 2738 3851 2750
rect 3916 2746 3922 2766
rect 3646 2728 3676 2738
rect 3677 2728 3835 2738
rect 3839 2728 3869 2738
rect 3873 2728 3903 2742
rect 3931 2728 3944 2766
rect 4016 2780 4045 2796
rect 4059 2780 4088 2796
rect 4103 2786 4133 2802
rect 4161 2780 4167 2828
rect 4170 2822 4189 2828
rect 4204 2822 4234 2830
rect 4170 2814 4234 2822
rect 4170 2798 4250 2814
rect 4266 2807 4328 2838
rect 4344 2807 4406 2838
rect 4475 2836 4524 2861
rect 4539 2836 4569 2852
rect 4438 2822 4468 2830
rect 4475 2828 4585 2836
rect 4438 2814 4483 2822
rect 4170 2796 4189 2798
rect 4204 2796 4250 2798
rect 4170 2780 4250 2796
rect 4277 2794 4312 2807
rect 4353 2804 4390 2807
rect 4353 2802 4395 2804
rect 4282 2791 4312 2794
rect 4291 2787 4298 2791
rect 4298 2786 4299 2787
rect 4257 2780 4267 2786
rect 4016 2772 4051 2780
rect 4016 2746 4017 2772
rect 4024 2746 4051 2772
rect 3959 2728 3989 2742
rect 4016 2738 4051 2746
rect 4053 2772 4094 2780
rect 4053 2746 4068 2772
rect 4075 2746 4094 2772
rect 4158 2768 4189 2780
rect 4204 2768 4307 2780
rect 4319 2770 4345 2796
rect 4360 2791 4390 2802
rect 4422 2798 4484 2814
rect 4422 2796 4468 2798
rect 4422 2780 4484 2796
rect 4496 2780 4502 2828
rect 4505 2820 4585 2828
rect 4505 2818 4524 2820
rect 4539 2818 4573 2820
rect 4505 2802 4585 2818
rect 4505 2780 4524 2802
rect 4539 2786 4569 2802
rect 4597 2796 4603 2870
rect 4606 2796 4625 2940
rect 4640 2796 4646 2940
rect 4655 2870 4668 2940
rect 4720 2936 4742 2940
rect 4713 2914 4742 2928
rect 4795 2914 4811 2928
rect 4849 2924 4855 2926
rect 4862 2924 4970 2940
rect 4977 2924 4983 2926
rect 4991 2924 5006 2940
rect 5072 2934 5091 2937
rect 4713 2912 4811 2914
rect 4838 2912 5006 2924
rect 5021 2914 5037 2928
rect 5072 2915 5094 2934
rect 5104 2928 5120 2929
rect 5103 2926 5120 2928
rect 5104 2921 5120 2926
rect 5094 2914 5100 2915
rect 5103 2914 5132 2921
rect 5021 2913 5132 2914
rect 5021 2912 5138 2913
rect 4697 2904 4748 2912
rect 4795 2904 4829 2912
rect 4697 2892 4722 2904
rect 4729 2892 4748 2904
rect 4802 2902 4829 2904
rect 4838 2902 5059 2912
rect 5094 2909 5100 2912
rect 4802 2898 5059 2902
rect 4697 2884 4748 2892
rect 4795 2884 5059 2898
rect 5103 2904 5138 2912
rect 4649 2836 4668 2870
rect 4713 2876 4742 2884
rect 4713 2870 4730 2876
rect 4713 2868 4747 2870
rect 4795 2868 4811 2884
rect 4812 2874 5020 2884
rect 5021 2874 5037 2884
rect 5085 2880 5100 2895
rect 5103 2892 5104 2904
rect 5111 2892 5138 2904
rect 5103 2884 5138 2892
rect 5103 2883 5132 2884
rect 4823 2870 5037 2874
rect 4838 2868 5037 2870
rect 5072 2870 5085 2880
rect 5103 2870 5120 2883
rect 5072 2868 5120 2870
rect 4714 2864 4747 2868
rect 4710 2862 4747 2864
rect 4710 2861 4777 2862
rect 4710 2856 4741 2861
rect 4747 2856 4777 2861
rect 4710 2852 4777 2856
rect 4683 2849 4777 2852
rect 4683 2842 4732 2849
rect 4683 2836 4713 2842
rect 4732 2837 4737 2842
rect 4649 2820 4729 2836
rect 4741 2828 4777 2849
rect 4838 2844 5027 2868
rect 5072 2867 5119 2868
rect 5085 2862 5119 2867
rect 4853 2841 5027 2844
rect 4846 2838 5027 2841
rect 5055 2861 5119 2862
rect 4649 2818 4668 2820
rect 4683 2818 4717 2820
rect 4649 2802 4729 2818
rect 4649 2796 4668 2802
rect 4365 2770 4468 2780
rect 4319 2768 4468 2770
rect 4489 2768 4524 2780
rect 4158 2766 4320 2768
rect 4170 2746 4189 2766
rect 4204 2764 4234 2766
rect 4053 2738 4094 2746
rect 4176 2742 4189 2746
rect 4241 2750 4320 2766
rect 4352 2766 4524 2768
rect 4352 2750 4431 2766
rect 4438 2764 4468 2766
rect 4016 2728 4045 2738
rect 4059 2728 4088 2738
rect 4103 2728 4133 2742
rect 4176 2728 4219 2742
rect 4241 2738 4431 2750
rect 4496 2746 4502 2766
rect 4226 2728 4256 2738
rect 4257 2728 4415 2738
rect 4419 2728 4449 2738
rect 4453 2728 4483 2742
rect 4511 2728 4524 2766
rect 4596 2780 4625 2796
rect 4639 2780 4668 2796
rect 4683 2786 4713 2802
rect 4741 2780 4747 2828
rect 4750 2822 4769 2828
rect 4784 2822 4814 2830
rect 4750 2814 4814 2822
rect 4750 2798 4830 2814
rect 4846 2807 4908 2838
rect 4924 2807 4986 2838
rect 5055 2836 5104 2861
rect 5119 2836 5149 2852
rect 5018 2822 5048 2830
rect 5055 2828 5165 2836
rect 5018 2814 5063 2822
rect 4750 2796 4769 2798
rect 4784 2796 4830 2798
rect 4750 2780 4830 2796
rect 4857 2794 4892 2807
rect 4933 2804 4970 2807
rect 4933 2802 4975 2804
rect 4862 2791 4892 2794
rect 4871 2787 4878 2791
rect 4878 2786 4879 2787
rect 4837 2780 4847 2786
rect 4596 2772 4631 2780
rect 4596 2746 4597 2772
rect 4604 2746 4631 2772
rect 4539 2728 4569 2742
rect 4596 2738 4631 2746
rect 4633 2772 4674 2780
rect 4633 2746 4648 2772
rect 4655 2746 4674 2772
rect 4738 2768 4769 2780
rect 4784 2768 4887 2780
rect 4899 2770 4925 2796
rect 4940 2791 4970 2802
rect 5002 2798 5064 2814
rect 5002 2796 5048 2798
rect 5002 2780 5064 2796
rect 5076 2780 5082 2828
rect 5085 2820 5165 2828
rect 5085 2818 5104 2820
rect 5119 2818 5153 2820
rect 5085 2802 5165 2818
rect 5085 2780 5104 2802
rect 5119 2786 5149 2802
rect 5177 2796 5183 2870
rect 5186 2796 5205 2940
rect 5220 2796 5226 2940
rect 5235 2870 5248 2940
rect 5300 2936 5322 2940
rect 5293 2914 5322 2928
rect 5375 2914 5391 2928
rect 5429 2924 5435 2926
rect 5442 2924 5550 2940
rect 5557 2924 5563 2926
rect 5571 2924 5586 2940
rect 5652 2934 5671 2937
rect 5293 2912 5391 2914
rect 5418 2912 5586 2924
rect 5601 2914 5617 2928
rect 5652 2915 5674 2934
rect 5684 2928 5700 2929
rect 5683 2926 5700 2928
rect 5684 2921 5700 2926
rect 5674 2914 5680 2915
rect 5683 2914 5712 2921
rect 5601 2913 5712 2914
rect 5601 2912 5718 2913
rect 5277 2904 5328 2912
rect 5375 2904 5409 2912
rect 5277 2892 5302 2904
rect 5309 2892 5328 2904
rect 5382 2902 5409 2904
rect 5418 2902 5639 2912
rect 5674 2909 5680 2912
rect 5382 2898 5639 2902
rect 5277 2884 5328 2892
rect 5375 2884 5639 2898
rect 5683 2904 5718 2912
rect 5229 2836 5248 2870
rect 5293 2876 5322 2884
rect 5293 2870 5310 2876
rect 5293 2868 5327 2870
rect 5375 2868 5391 2884
rect 5392 2874 5600 2884
rect 5601 2874 5617 2884
rect 5665 2880 5680 2895
rect 5683 2892 5684 2904
rect 5691 2892 5718 2904
rect 5683 2884 5718 2892
rect 5683 2883 5712 2884
rect 5403 2870 5617 2874
rect 5418 2868 5617 2870
rect 5652 2870 5665 2880
rect 5683 2870 5700 2883
rect 5652 2868 5700 2870
rect 5294 2864 5327 2868
rect 5290 2862 5327 2864
rect 5290 2861 5357 2862
rect 5290 2856 5321 2861
rect 5327 2856 5357 2861
rect 5290 2852 5357 2856
rect 5263 2849 5357 2852
rect 5263 2842 5312 2849
rect 5263 2836 5293 2842
rect 5312 2837 5317 2842
rect 5229 2820 5309 2836
rect 5321 2828 5357 2849
rect 5418 2844 5607 2868
rect 5652 2867 5699 2868
rect 5665 2862 5699 2867
rect 5433 2841 5607 2844
rect 5426 2838 5607 2841
rect 5635 2861 5699 2862
rect 5229 2818 5248 2820
rect 5263 2818 5297 2820
rect 5229 2802 5309 2818
rect 5229 2796 5248 2802
rect 4945 2770 5048 2780
rect 4899 2768 5048 2770
rect 5069 2768 5104 2780
rect 4738 2766 4900 2768
rect 4750 2746 4769 2766
rect 4784 2764 4814 2766
rect 4633 2738 4674 2746
rect 4756 2742 4769 2746
rect 4821 2750 4900 2766
rect 4932 2766 5104 2768
rect 4932 2750 5011 2766
rect 5018 2764 5048 2766
rect 4596 2728 4625 2738
rect 4639 2728 4668 2738
rect 4683 2728 4713 2742
rect 4756 2728 4799 2742
rect 4821 2738 5011 2750
rect 5076 2746 5082 2766
rect 4806 2728 4836 2738
rect 4837 2728 4995 2738
rect 4999 2728 5029 2738
rect 5033 2728 5063 2742
rect 5091 2728 5104 2766
rect 5176 2780 5205 2796
rect 5219 2780 5248 2796
rect 5263 2786 5293 2802
rect 5321 2780 5327 2828
rect 5330 2822 5349 2828
rect 5364 2822 5394 2830
rect 5330 2814 5394 2822
rect 5330 2798 5410 2814
rect 5426 2807 5488 2838
rect 5504 2807 5566 2838
rect 5635 2836 5684 2861
rect 5699 2836 5729 2852
rect 5598 2822 5628 2830
rect 5635 2828 5745 2836
rect 5598 2814 5643 2822
rect 5330 2796 5349 2798
rect 5364 2796 5410 2798
rect 5330 2780 5410 2796
rect 5437 2794 5472 2807
rect 5513 2804 5550 2807
rect 5513 2802 5555 2804
rect 5442 2791 5472 2794
rect 5451 2787 5458 2791
rect 5458 2786 5459 2787
rect 5417 2780 5427 2786
rect 5176 2772 5211 2780
rect 5176 2746 5177 2772
rect 5184 2746 5211 2772
rect 5119 2728 5149 2742
rect 5176 2738 5211 2746
rect 5213 2772 5254 2780
rect 5213 2746 5228 2772
rect 5235 2746 5254 2772
rect 5318 2768 5349 2780
rect 5364 2768 5467 2780
rect 5479 2770 5505 2796
rect 5520 2791 5550 2802
rect 5582 2798 5644 2814
rect 5582 2796 5628 2798
rect 5582 2780 5644 2796
rect 5656 2780 5662 2828
rect 5665 2820 5745 2828
rect 5665 2818 5684 2820
rect 5699 2818 5733 2820
rect 5665 2802 5745 2818
rect 5665 2780 5684 2802
rect 5699 2786 5729 2802
rect 5757 2796 5763 2870
rect 5766 2796 5785 2940
rect 5800 2796 5806 2940
rect 5815 2870 5828 2940
rect 5880 2936 5902 2940
rect 5873 2914 5902 2928
rect 5955 2914 5971 2928
rect 6009 2924 6015 2926
rect 6022 2924 6130 2940
rect 6137 2924 6143 2926
rect 6151 2924 6166 2940
rect 6232 2934 6251 2937
rect 5873 2912 5971 2914
rect 5998 2912 6166 2924
rect 6181 2914 6197 2928
rect 6232 2915 6254 2934
rect 6264 2928 6280 2929
rect 6263 2926 6280 2928
rect 6264 2921 6280 2926
rect 6254 2914 6260 2915
rect 6263 2914 6292 2921
rect 6181 2913 6292 2914
rect 6181 2912 6298 2913
rect 5857 2904 5908 2912
rect 5955 2904 5989 2912
rect 5857 2892 5882 2904
rect 5889 2892 5908 2904
rect 5962 2902 5989 2904
rect 5998 2902 6219 2912
rect 6254 2909 6260 2912
rect 5962 2898 6219 2902
rect 5857 2884 5908 2892
rect 5955 2884 6219 2898
rect 6263 2904 6298 2912
rect 5809 2836 5828 2870
rect 5873 2876 5902 2884
rect 5873 2870 5890 2876
rect 5873 2868 5907 2870
rect 5955 2868 5971 2884
rect 5972 2874 6180 2884
rect 6181 2874 6197 2884
rect 6245 2880 6260 2895
rect 6263 2892 6264 2904
rect 6271 2892 6298 2904
rect 6263 2884 6298 2892
rect 6263 2883 6292 2884
rect 5983 2870 6197 2874
rect 5998 2868 6197 2870
rect 6232 2870 6245 2880
rect 6263 2870 6280 2883
rect 6232 2868 6280 2870
rect 5874 2864 5907 2868
rect 5870 2862 5907 2864
rect 5870 2861 5937 2862
rect 5870 2856 5901 2861
rect 5907 2856 5937 2861
rect 5870 2852 5937 2856
rect 5843 2849 5937 2852
rect 5843 2842 5892 2849
rect 5843 2836 5873 2842
rect 5892 2837 5897 2842
rect 5809 2820 5889 2836
rect 5901 2828 5937 2849
rect 5998 2844 6187 2868
rect 6232 2867 6279 2868
rect 6245 2862 6279 2867
rect 6013 2841 6187 2844
rect 6006 2838 6187 2841
rect 6215 2861 6279 2862
rect 5809 2818 5828 2820
rect 5843 2818 5877 2820
rect 5809 2802 5889 2818
rect 5809 2796 5828 2802
rect 5525 2770 5628 2780
rect 5479 2768 5628 2770
rect 5649 2768 5684 2780
rect 5318 2766 5480 2768
rect 5330 2746 5349 2766
rect 5364 2764 5394 2766
rect 5213 2738 5254 2746
rect 5336 2742 5349 2746
rect 5401 2750 5480 2766
rect 5512 2766 5684 2768
rect 5512 2750 5591 2766
rect 5598 2764 5628 2766
rect 5176 2728 5205 2738
rect 5219 2728 5248 2738
rect 5263 2728 5293 2742
rect 5336 2728 5379 2742
rect 5401 2738 5591 2750
rect 5656 2746 5662 2766
rect 5386 2728 5416 2738
rect 5417 2728 5575 2738
rect 5579 2728 5609 2738
rect 5613 2728 5643 2742
rect 5671 2728 5684 2766
rect 5756 2780 5785 2796
rect 5799 2780 5828 2796
rect 5843 2786 5873 2802
rect 5901 2780 5907 2828
rect 5910 2822 5929 2828
rect 5944 2822 5974 2830
rect 5910 2814 5974 2822
rect 5910 2798 5990 2814
rect 6006 2807 6068 2838
rect 6084 2807 6146 2838
rect 6215 2836 6264 2861
rect 6279 2836 6309 2852
rect 6178 2822 6208 2830
rect 6215 2828 6325 2836
rect 6178 2814 6223 2822
rect 5910 2796 5929 2798
rect 5944 2796 5990 2798
rect 5910 2780 5990 2796
rect 6017 2794 6052 2807
rect 6093 2804 6130 2807
rect 6093 2802 6135 2804
rect 6022 2791 6052 2794
rect 6031 2787 6038 2791
rect 6038 2786 6039 2787
rect 5997 2780 6007 2786
rect 5756 2772 5791 2780
rect 5756 2746 5757 2772
rect 5764 2746 5791 2772
rect 5699 2728 5729 2742
rect 5756 2738 5791 2746
rect 5793 2772 5834 2780
rect 5793 2746 5808 2772
rect 5815 2746 5834 2772
rect 5898 2768 5929 2780
rect 5944 2768 6047 2780
rect 6059 2770 6085 2796
rect 6100 2791 6130 2802
rect 6162 2798 6224 2814
rect 6162 2796 6208 2798
rect 6162 2780 6224 2796
rect 6236 2780 6242 2828
rect 6245 2820 6325 2828
rect 6245 2818 6264 2820
rect 6279 2818 6313 2820
rect 6245 2802 6325 2818
rect 6245 2780 6264 2802
rect 6279 2786 6309 2802
rect 6337 2796 6343 2870
rect 6346 2796 6365 2940
rect 6380 2796 6386 2940
rect 6395 2870 6408 2940
rect 6460 2936 6482 2940
rect 6453 2914 6482 2928
rect 6535 2914 6551 2928
rect 6589 2924 6595 2926
rect 6602 2924 6710 2940
rect 6717 2924 6723 2926
rect 6731 2924 6746 2940
rect 6812 2934 6831 2937
rect 6453 2912 6551 2914
rect 6578 2912 6746 2924
rect 6761 2914 6777 2928
rect 6812 2915 6834 2934
rect 6844 2928 6860 2929
rect 6843 2926 6860 2928
rect 6844 2921 6860 2926
rect 6834 2914 6840 2915
rect 6843 2914 6872 2921
rect 6761 2913 6872 2914
rect 6761 2912 6878 2913
rect 6437 2904 6488 2912
rect 6535 2904 6569 2912
rect 6437 2892 6462 2904
rect 6469 2892 6488 2904
rect 6542 2902 6569 2904
rect 6578 2902 6799 2912
rect 6834 2909 6840 2912
rect 6542 2898 6799 2902
rect 6437 2884 6488 2892
rect 6535 2884 6799 2898
rect 6843 2904 6878 2912
rect 6389 2836 6408 2870
rect 6453 2876 6482 2884
rect 6453 2870 6470 2876
rect 6453 2868 6487 2870
rect 6535 2868 6551 2884
rect 6552 2874 6760 2884
rect 6761 2874 6777 2884
rect 6825 2880 6840 2895
rect 6843 2892 6844 2904
rect 6851 2892 6878 2904
rect 6843 2884 6878 2892
rect 6843 2883 6872 2884
rect 6563 2870 6777 2874
rect 6578 2868 6777 2870
rect 6812 2870 6825 2880
rect 6843 2870 6860 2883
rect 6812 2868 6860 2870
rect 6454 2864 6487 2868
rect 6450 2862 6487 2864
rect 6450 2861 6517 2862
rect 6450 2856 6481 2861
rect 6487 2856 6517 2861
rect 6450 2852 6517 2856
rect 6423 2849 6517 2852
rect 6423 2842 6472 2849
rect 6423 2836 6453 2842
rect 6472 2837 6477 2842
rect 6389 2820 6469 2836
rect 6481 2828 6517 2849
rect 6578 2844 6767 2868
rect 6812 2867 6859 2868
rect 6825 2862 6859 2867
rect 6593 2841 6767 2844
rect 6586 2838 6767 2841
rect 6795 2861 6859 2862
rect 6389 2818 6408 2820
rect 6423 2818 6457 2820
rect 6389 2802 6469 2818
rect 6389 2796 6408 2802
rect 6105 2770 6208 2780
rect 6059 2768 6208 2770
rect 6229 2768 6264 2780
rect 5898 2766 6060 2768
rect 5910 2746 5929 2766
rect 5944 2764 5974 2766
rect 5793 2738 5834 2746
rect 5916 2742 5929 2746
rect 5981 2750 6060 2766
rect 6092 2766 6264 2768
rect 6092 2750 6171 2766
rect 6178 2764 6208 2766
rect 5756 2728 5785 2738
rect 5799 2728 5828 2738
rect 5843 2728 5873 2742
rect 5916 2728 5959 2742
rect 5981 2738 6171 2750
rect 6236 2746 6242 2766
rect 5966 2728 5996 2738
rect 5997 2728 6155 2738
rect 6159 2728 6189 2738
rect 6193 2728 6223 2742
rect 6251 2728 6264 2766
rect 6336 2780 6365 2796
rect 6379 2780 6408 2796
rect 6423 2786 6453 2802
rect 6481 2780 6487 2828
rect 6490 2822 6509 2828
rect 6524 2822 6554 2830
rect 6490 2814 6554 2822
rect 6490 2798 6570 2814
rect 6586 2807 6648 2838
rect 6664 2807 6726 2838
rect 6795 2836 6844 2861
rect 6859 2836 6889 2852
rect 6758 2822 6788 2830
rect 6795 2828 6905 2836
rect 6758 2814 6803 2822
rect 6490 2796 6509 2798
rect 6524 2796 6570 2798
rect 6490 2780 6570 2796
rect 6597 2794 6632 2807
rect 6673 2804 6710 2807
rect 6673 2802 6715 2804
rect 6602 2791 6632 2794
rect 6611 2787 6618 2791
rect 6618 2786 6619 2787
rect 6577 2780 6587 2786
rect 6336 2772 6371 2780
rect 6336 2746 6337 2772
rect 6344 2746 6371 2772
rect 6279 2728 6309 2742
rect 6336 2738 6371 2746
rect 6373 2772 6414 2780
rect 6373 2746 6388 2772
rect 6395 2746 6414 2772
rect 6478 2768 6509 2780
rect 6524 2768 6627 2780
rect 6639 2770 6665 2796
rect 6680 2791 6710 2802
rect 6742 2798 6804 2814
rect 6742 2796 6788 2798
rect 6742 2780 6804 2796
rect 6816 2780 6822 2828
rect 6825 2820 6905 2828
rect 6825 2818 6844 2820
rect 6859 2818 6893 2820
rect 6825 2802 6905 2818
rect 6825 2780 6844 2802
rect 6859 2786 6889 2802
rect 6917 2796 6923 2870
rect 6926 2796 6945 2940
rect 6960 2796 6966 2940
rect 6975 2870 6988 2940
rect 7040 2936 7062 2940
rect 7033 2914 7062 2928
rect 7115 2914 7131 2928
rect 7169 2924 7175 2926
rect 7182 2924 7290 2940
rect 7297 2924 7303 2926
rect 7311 2924 7326 2940
rect 7392 2934 7411 2937
rect 7033 2912 7131 2914
rect 7158 2912 7326 2924
rect 7341 2914 7357 2928
rect 7392 2915 7414 2934
rect 7424 2928 7440 2929
rect 7423 2926 7440 2928
rect 7424 2921 7440 2926
rect 7414 2914 7420 2915
rect 7423 2914 7452 2921
rect 7341 2913 7452 2914
rect 7341 2912 7458 2913
rect 7017 2904 7068 2912
rect 7115 2904 7149 2912
rect 7017 2892 7042 2904
rect 7049 2892 7068 2904
rect 7122 2902 7149 2904
rect 7158 2902 7379 2912
rect 7414 2909 7420 2912
rect 7122 2898 7379 2902
rect 7017 2884 7068 2892
rect 7115 2884 7379 2898
rect 7423 2904 7458 2912
rect 6969 2836 6988 2870
rect 7033 2876 7062 2884
rect 7033 2870 7050 2876
rect 7033 2868 7067 2870
rect 7115 2868 7131 2884
rect 7132 2874 7340 2884
rect 7341 2874 7357 2884
rect 7405 2880 7420 2895
rect 7423 2892 7424 2904
rect 7431 2892 7458 2904
rect 7423 2884 7458 2892
rect 7423 2883 7452 2884
rect 7151 2870 7357 2874
rect 7158 2868 7357 2870
rect 7392 2870 7405 2880
rect 7423 2870 7440 2883
rect 7392 2868 7440 2870
rect 7034 2864 7067 2868
rect 7030 2862 7067 2864
rect 7030 2861 7097 2862
rect 7030 2856 7061 2861
rect 7067 2856 7097 2861
rect 7030 2852 7097 2856
rect 7003 2849 7097 2852
rect 7003 2842 7052 2849
rect 7003 2836 7033 2842
rect 7052 2837 7057 2842
rect 6969 2820 7049 2836
rect 7061 2828 7097 2849
rect 7158 2844 7347 2868
rect 7392 2867 7439 2868
rect 7405 2862 7439 2867
rect 7173 2841 7347 2844
rect 7166 2838 7347 2841
rect 7375 2861 7439 2862
rect 6969 2818 6988 2820
rect 7003 2818 7037 2820
rect 6969 2802 7049 2818
rect 6969 2796 6988 2802
rect 6685 2770 6788 2780
rect 6639 2768 6788 2770
rect 6809 2768 6844 2780
rect 6478 2766 6640 2768
rect 6490 2746 6509 2766
rect 6524 2764 6554 2766
rect 6373 2738 6414 2746
rect 6496 2742 6509 2746
rect 6561 2750 6640 2766
rect 6672 2766 6844 2768
rect 6672 2750 6751 2766
rect 6758 2764 6788 2766
rect 6336 2728 6365 2738
rect 6379 2728 6408 2738
rect 6423 2728 6453 2742
rect 6496 2728 6539 2742
rect 6561 2738 6751 2750
rect 6816 2746 6822 2766
rect 6546 2728 6576 2738
rect 6577 2728 6735 2738
rect 6739 2728 6769 2738
rect 6773 2728 6803 2742
rect 6831 2728 6844 2766
rect 6916 2780 6945 2796
rect 6959 2780 6988 2796
rect 7003 2786 7033 2802
rect 7061 2780 7067 2828
rect 7070 2822 7089 2828
rect 7104 2822 7134 2830
rect 7070 2814 7134 2822
rect 7070 2798 7150 2814
rect 7166 2807 7228 2838
rect 7244 2807 7306 2838
rect 7375 2836 7424 2861
rect 7439 2836 7469 2852
rect 7338 2822 7368 2830
rect 7375 2828 7485 2836
rect 7338 2814 7383 2822
rect 7070 2796 7089 2798
rect 7104 2796 7150 2798
rect 7070 2780 7150 2796
rect 7177 2794 7212 2807
rect 7253 2804 7290 2807
rect 7253 2802 7295 2804
rect 7182 2791 7212 2794
rect 7191 2787 7198 2791
rect 7198 2786 7199 2787
rect 7157 2780 7167 2786
rect 6916 2772 6951 2780
rect 6916 2746 6917 2772
rect 6924 2746 6951 2772
rect 6859 2728 6889 2742
rect 6916 2738 6951 2746
rect 6953 2772 6994 2780
rect 6953 2746 6968 2772
rect 6975 2746 6994 2772
rect 7058 2768 7089 2780
rect 7104 2768 7207 2780
rect 7219 2770 7245 2796
rect 7260 2791 7290 2802
rect 7322 2798 7384 2814
rect 7322 2796 7368 2798
rect 7322 2780 7384 2796
rect 7396 2780 7402 2828
rect 7405 2820 7485 2828
rect 7405 2818 7424 2820
rect 7439 2818 7473 2820
rect 7405 2802 7485 2818
rect 7405 2780 7424 2802
rect 7439 2786 7469 2802
rect 7497 2796 7503 2870
rect 7506 2796 7525 2940
rect 7540 2796 7546 2940
rect 7555 2870 7568 2940
rect 7620 2936 7642 2940
rect 7613 2914 7642 2928
rect 7695 2914 7711 2928
rect 7749 2924 7755 2926
rect 7762 2924 7870 2940
rect 7877 2924 7883 2926
rect 7891 2924 7906 2940
rect 7972 2934 7991 2937
rect 7613 2912 7711 2914
rect 7738 2912 7906 2924
rect 7921 2914 7937 2928
rect 7972 2915 7994 2934
rect 8004 2928 8020 2929
rect 8003 2926 8020 2928
rect 8004 2921 8020 2926
rect 7994 2914 8000 2915
rect 8003 2914 8032 2921
rect 7921 2913 8032 2914
rect 7921 2912 8038 2913
rect 7597 2904 7648 2912
rect 7695 2904 7729 2912
rect 7597 2892 7622 2904
rect 7629 2892 7648 2904
rect 7702 2902 7729 2904
rect 7738 2902 7959 2912
rect 7994 2909 8000 2912
rect 7702 2898 7959 2902
rect 7597 2884 7648 2892
rect 7695 2884 7959 2898
rect 8003 2904 8038 2912
rect 7549 2836 7568 2870
rect 7613 2876 7642 2884
rect 7613 2870 7630 2876
rect 7613 2868 7647 2870
rect 7695 2868 7711 2884
rect 7712 2874 7920 2884
rect 7921 2874 7937 2884
rect 7985 2880 8000 2895
rect 8003 2892 8004 2904
rect 8011 2892 8038 2904
rect 8003 2884 8038 2892
rect 8003 2883 8032 2884
rect 7723 2870 7937 2874
rect 7738 2868 7937 2870
rect 7972 2870 7985 2880
rect 8003 2870 8020 2883
rect 7972 2868 8020 2870
rect 7614 2864 7647 2868
rect 7610 2862 7647 2864
rect 7610 2861 7677 2862
rect 7610 2856 7641 2861
rect 7647 2856 7677 2861
rect 7610 2852 7677 2856
rect 7583 2849 7677 2852
rect 7583 2842 7632 2849
rect 7583 2836 7613 2842
rect 7632 2837 7637 2842
rect 7549 2820 7629 2836
rect 7641 2828 7677 2849
rect 7738 2844 7927 2868
rect 7972 2867 8019 2868
rect 7985 2862 8019 2867
rect 7753 2841 7927 2844
rect 7746 2838 7927 2841
rect 7955 2861 8019 2862
rect 7549 2818 7568 2820
rect 7583 2818 7617 2820
rect 7549 2802 7629 2818
rect 7549 2796 7568 2802
rect 7265 2770 7368 2780
rect 7219 2768 7368 2770
rect 7389 2768 7424 2780
rect 7058 2766 7220 2768
rect 7070 2746 7089 2766
rect 7104 2764 7134 2766
rect 6953 2738 6994 2746
rect 7076 2742 7089 2746
rect 7141 2750 7220 2766
rect 7252 2766 7424 2768
rect 7252 2750 7331 2766
rect 7338 2764 7368 2766
rect 6916 2728 6945 2738
rect 6959 2728 6988 2738
rect 7003 2728 7033 2742
rect 7076 2728 7119 2742
rect 7141 2738 7331 2750
rect 7396 2746 7402 2766
rect 7126 2728 7156 2738
rect 7157 2728 7315 2738
rect 7319 2728 7349 2738
rect 7353 2728 7383 2742
rect 7411 2728 7424 2766
rect 7496 2780 7525 2796
rect 7539 2780 7568 2796
rect 7583 2786 7613 2802
rect 7641 2780 7647 2828
rect 7650 2822 7669 2828
rect 7684 2822 7714 2830
rect 7650 2814 7714 2822
rect 7650 2798 7730 2814
rect 7746 2807 7808 2838
rect 7824 2807 7886 2838
rect 7955 2836 8004 2861
rect 8019 2836 8049 2852
rect 7918 2822 7948 2830
rect 7955 2828 8065 2836
rect 7918 2814 7963 2822
rect 7650 2796 7669 2798
rect 7684 2796 7730 2798
rect 7650 2780 7730 2796
rect 7757 2794 7792 2807
rect 7833 2804 7870 2807
rect 7833 2802 7875 2804
rect 7762 2791 7792 2794
rect 7771 2787 7778 2791
rect 7778 2786 7779 2787
rect 7737 2780 7747 2786
rect 7496 2772 7531 2780
rect 7496 2746 7497 2772
rect 7504 2746 7531 2772
rect 7439 2728 7469 2742
rect 7496 2738 7531 2746
rect 7533 2772 7574 2780
rect 7533 2746 7548 2772
rect 7555 2746 7574 2772
rect 7638 2768 7669 2780
rect 7684 2768 7787 2780
rect 7799 2770 7825 2796
rect 7840 2791 7870 2802
rect 7902 2798 7964 2814
rect 7902 2796 7948 2798
rect 7902 2780 7964 2796
rect 7976 2780 7982 2828
rect 7985 2820 8065 2828
rect 7985 2818 8004 2820
rect 8019 2818 8053 2820
rect 7985 2802 8065 2818
rect 7985 2780 8004 2802
rect 8019 2786 8049 2802
rect 8077 2796 8083 2870
rect 8086 2796 8105 2940
rect 8120 2796 8126 2940
rect 8135 2870 8148 2940
rect 8200 2936 8222 2940
rect 8193 2914 8222 2928
rect 8275 2914 8291 2928
rect 8329 2924 8335 2926
rect 8342 2924 8450 2940
rect 8457 2924 8463 2926
rect 8471 2924 8486 2940
rect 8552 2934 8571 2937
rect 8193 2912 8291 2914
rect 8318 2912 8486 2924
rect 8501 2914 8517 2928
rect 8552 2915 8574 2934
rect 8584 2928 8600 2929
rect 8583 2926 8600 2928
rect 8584 2921 8600 2926
rect 8574 2914 8580 2915
rect 8583 2914 8612 2921
rect 8501 2913 8612 2914
rect 8501 2912 8618 2913
rect 8177 2904 8228 2912
rect 8275 2904 8309 2912
rect 8177 2892 8202 2904
rect 8209 2892 8228 2904
rect 8282 2902 8309 2904
rect 8318 2902 8539 2912
rect 8574 2909 8580 2912
rect 8282 2898 8539 2902
rect 8177 2884 8228 2892
rect 8275 2884 8539 2898
rect 8583 2904 8618 2912
rect 8129 2836 8148 2870
rect 8193 2876 8222 2884
rect 8193 2870 8210 2876
rect 8193 2868 8227 2870
rect 8275 2868 8291 2884
rect 8292 2874 8500 2884
rect 8501 2874 8517 2884
rect 8565 2880 8580 2895
rect 8583 2892 8584 2904
rect 8591 2892 8618 2904
rect 8583 2884 8618 2892
rect 8583 2883 8612 2884
rect 8303 2870 8517 2874
rect 8318 2868 8517 2870
rect 8552 2870 8565 2880
rect 8583 2870 8600 2883
rect 8552 2868 8600 2870
rect 8194 2864 8227 2868
rect 8190 2862 8227 2864
rect 8190 2861 8257 2862
rect 8190 2856 8221 2861
rect 8227 2856 8257 2861
rect 8190 2852 8257 2856
rect 8163 2849 8257 2852
rect 8163 2842 8212 2849
rect 8163 2836 8193 2842
rect 8212 2837 8217 2842
rect 8129 2820 8209 2836
rect 8221 2828 8257 2849
rect 8318 2844 8507 2868
rect 8552 2867 8599 2868
rect 8565 2862 8599 2867
rect 8333 2841 8507 2844
rect 8326 2838 8507 2841
rect 8535 2861 8599 2862
rect 8129 2818 8148 2820
rect 8163 2818 8197 2820
rect 8129 2802 8209 2818
rect 8129 2796 8148 2802
rect 7845 2770 7948 2780
rect 7799 2768 7948 2770
rect 7969 2768 8004 2780
rect 7638 2766 7800 2768
rect 7650 2746 7669 2766
rect 7684 2764 7714 2766
rect 7533 2738 7574 2746
rect 7656 2742 7669 2746
rect 7721 2750 7800 2766
rect 7832 2766 8004 2768
rect 7832 2750 7911 2766
rect 7918 2764 7948 2766
rect 7496 2728 7525 2738
rect 7539 2728 7568 2738
rect 7583 2728 7613 2742
rect 7656 2728 7699 2742
rect 7721 2738 7911 2750
rect 7976 2746 7982 2766
rect 7706 2728 7736 2738
rect 7737 2728 7895 2738
rect 7899 2728 7929 2738
rect 7933 2728 7963 2742
rect 7991 2728 8004 2766
rect 8076 2780 8105 2796
rect 8119 2780 8148 2796
rect 8163 2786 8193 2802
rect 8221 2780 8227 2828
rect 8230 2822 8249 2828
rect 8264 2822 8294 2830
rect 8230 2814 8294 2822
rect 8230 2798 8310 2814
rect 8326 2807 8388 2838
rect 8404 2807 8466 2838
rect 8535 2836 8584 2861
rect 8599 2836 8629 2852
rect 8498 2822 8528 2830
rect 8535 2828 8645 2836
rect 8498 2814 8543 2822
rect 8230 2796 8249 2798
rect 8264 2796 8310 2798
rect 8230 2780 8310 2796
rect 8337 2794 8372 2807
rect 8413 2804 8450 2807
rect 8413 2802 8455 2804
rect 8342 2791 8372 2794
rect 8351 2787 8358 2791
rect 8358 2786 8359 2787
rect 8317 2780 8327 2786
rect 8076 2772 8111 2780
rect 8076 2746 8077 2772
rect 8084 2746 8111 2772
rect 8019 2728 8049 2742
rect 8076 2738 8111 2746
rect 8113 2772 8154 2780
rect 8113 2746 8128 2772
rect 8135 2746 8154 2772
rect 8218 2768 8249 2780
rect 8264 2768 8367 2780
rect 8379 2770 8405 2796
rect 8420 2791 8450 2802
rect 8482 2798 8544 2814
rect 8482 2796 8528 2798
rect 8482 2780 8544 2796
rect 8556 2780 8562 2828
rect 8565 2820 8645 2828
rect 8565 2818 8584 2820
rect 8599 2818 8633 2820
rect 8565 2802 8645 2818
rect 8565 2780 8584 2802
rect 8599 2786 8629 2802
rect 8657 2796 8663 2870
rect 8666 2796 8685 2940
rect 8700 2796 8706 2940
rect 8715 2870 8728 2940
rect 8780 2936 8802 2940
rect 8773 2914 8802 2928
rect 8855 2914 8871 2928
rect 8909 2924 8915 2926
rect 8922 2924 9030 2940
rect 9037 2924 9043 2926
rect 9051 2924 9066 2940
rect 9132 2934 9151 2937
rect 8773 2912 8871 2914
rect 8898 2912 9066 2924
rect 9081 2914 9097 2928
rect 9132 2915 9154 2934
rect 9164 2928 9180 2929
rect 9163 2926 9180 2928
rect 9164 2921 9180 2926
rect 9154 2914 9160 2915
rect 9163 2914 9192 2921
rect 9081 2913 9192 2914
rect 9081 2912 9198 2913
rect 8757 2904 8808 2912
rect 8855 2904 8889 2912
rect 8757 2892 8782 2904
rect 8789 2892 8808 2904
rect 8862 2902 8889 2904
rect 8898 2902 9119 2912
rect 9154 2909 9160 2912
rect 8862 2898 9119 2902
rect 8757 2884 8808 2892
rect 8855 2884 9119 2898
rect 9163 2904 9198 2912
rect 8709 2836 8728 2870
rect 8773 2876 8802 2884
rect 8773 2870 8790 2876
rect 8773 2868 8807 2870
rect 8855 2868 8871 2884
rect 8872 2874 9080 2884
rect 9081 2874 9097 2884
rect 9145 2880 9160 2895
rect 9163 2892 9164 2904
rect 9171 2892 9198 2904
rect 9163 2884 9198 2892
rect 9163 2883 9192 2884
rect 8883 2870 9097 2874
rect 8898 2868 9097 2870
rect 9132 2870 9145 2880
rect 9163 2870 9180 2883
rect 9132 2868 9180 2870
rect 8774 2864 8807 2868
rect 8770 2862 8807 2864
rect 8770 2861 8837 2862
rect 8770 2856 8801 2861
rect 8807 2856 8837 2861
rect 8770 2852 8837 2856
rect 8743 2849 8837 2852
rect 8743 2842 8792 2849
rect 8743 2836 8773 2842
rect 8792 2837 8797 2842
rect 8709 2820 8789 2836
rect 8801 2828 8837 2849
rect 8898 2844 9087 2868
rect 9132 2867 9179 2868
rect 9145 2862 9179 2867
rect 8913 2841 9087 2844
rect 8906 2838 9087 2841
rect 9115 2861 9179 2862
rect 8709 2818 8728 2820
rect 8743 2818 8777 2820
rect 8709 2802 8789 2818
rect 8709 2796 8728 2802
rect 8425 2770 8528 2780
rect 8379 2768 8528 2770
rect 8549 2768 8584 2780
rect 8218 2766 8380 2768
rect 8230 2746 8249 2766
rect 8264 2764 8294 2766
rect 8113 2738 8154 2746
rect 8236 2742 8249 2746
rect 8301 2750 8380 2766
rect 8412 2766 8584 2768
rect 8412 2750 8491 2766
rect 8498 2764 8528 2766
rect 8076 2728 8105 2738
rect 8119 2728 8148 2738
rect 8163 2728 8193 2742
rect 8236 2728 8279 2742
rect 8301 2738 8491 2750
rect 8556 2746 8562 2766
rect 8286 2728 8316 2738
rect 8317 2728 8475 2738
rect 8479 2728 8509 2738
rect 8513 2728 8543 2742
rect 8571 2728 8584 2766
rect 8656 2780 8685 2796
rect 8699 2780 8728 2796
rect 8743 2786 8773 2802
rect 8801 2780 8807 2828
rect 8810 2822 8829 2828
rect 8844 2822 8874 2830
rect 8810 2814 8874 2822
rect 8810 2798 8890 2814
rect 8906 2807 8968 2838
rect 8984 2807 9046 2838
rect 9115 2836 9164 2861
rect 9179 2836 9209 2852
rect 9078 2822 9108 2830
rect 9115 2828 9225 2836
rect 9078 2814 9123 2822
rect 8810 2796 8829 2798
rect 8844 2796 8890 2798
rect 8810 2780 8890 2796
rect 8917 2794 8952 2807
rect 8993 2804 9030 2807
rect 8993 2802 9035 2804
rect 8922 2791 8952 2794
rect 8931 2787 8938 2791
rect 8938 2786 8939 2787
rect 8897 2780 8907 2786
rect 8656 2772 8691 2780
rect 8656 2746 8657 2772
rect 8664 2746 8691 2772
rect 8599 2728 8629 2742
rect 8656 2738 8691 2746
rect 8693 2772 8734 2780
rect 8693 2746 8708 2772
rect 8715 2746 8734 2772
rect 8798 2768 8829 2780
rect 8844 2768 8947 2780
rect 8959 2770 8985 2796
rect 9000 2791 9030 2802
rect 9062 2798 9124 2814
rect 9062 2796 9108 2798
rect 9062 2780 9124 2796
rect 9136 2780 9142 2828
rect 9145 2820 9225 2828
rect 9145 2818 9164 2820
rect 9179 2818 9213 2820
rect 9145 2802 9225 2818
rect 9145 2780 9164 2802
rect 9179 2786 9209 2802
rect 9237 2796 9243 2870
rect 9246 2796 9265 2940
rect 9280 2796 9286 2940
rect 9295 2870 9308 2940
rect 9360 2936 9382 2940
rect 9353 2914 9382 2928
rect 9435 2914 9451 2928
rect 9489 2924 9495 2926
rect 9502 2924 9610 2940
rect 9617 2924 9623 2926
rect 9631 2924 9646 2940
rect 9712 2934 9731 2937
rect 9353 2912 9451 2914
rect 9478 2912 9646 2924
rect 9661 2914 9677 2928
rect 9712 2915 9734 2934
rect 9744 2928 9760 2929
rect 9743 2926 9760 2928
rect 9744 2921 9760 2926
rect 9734 2914 9740 2915
rect 9743 2914 9772 2921
rect 9661 2913 9772 2914
rect 9661 2912 9778 2913
rect 9337 2904 9388 2912
rect 9435 2904 9469 2912
rect 9337 2892 9362 2904
rect 9369 2892 9388 2904
rect 9442 2902 9469 2904
rect 9478 2902 9699 2912
rect 9734 2909 9740 2912
rect 9442 2898 9699 2902
rect 9337 2884 9388 2892
rect 9435 2884 9699 2898
rect 9743 2904 9778 2912
rect 9289 2836 9308 2870
rect 9353 2876 9382 2884
rect 9353 2870 9370 2876
rect 9353 2868 9387 2870
rect 9435 2868 9451 2884
rect 9452 2874 9660 2884
rect 9661 2874 9677 2884
rect 9725 2880 9740 2895
rect 9743 2892 9744 2904
rect 9751 2892 9778 2904
rect 9743 2884 9778 2892
rect 9743 2883 9772 2884
rect 9463 2870 9677 2874
rect 9478 2868 9677 2870
rect 9712 2870 9725 2880
rect 9743 2870 9760 2883
rect 9712 2868 9760 2870
rect 9354 2864 9387 2868
rect 9350 2862 9387 2864
rect 9350 2861 9417 2862
rect 9350 2856 9381 2861
rect 9387 2856 9417 2861
rect 9350 2852 9417 2856
rect 9323 2849 9417 2852
rect 9323 2842 9372 2849
rect 9323 2836 9353 2842
rect 9372 2837 9377 2842
rect 9289 2820 9369 2836
rect 9381 2828 9417 2849
rect 9478 2844 9667 2868
rect 9712 2867 9759 2868
rect 9725 2862 9759 2867
rect 9493 2841 9667 2844
rect 9486 2838 9667 2841
rect 9695 2861 9759 2862
rect 9289 2818 9308 2820
rect 9323 2818 9357 2820
rect 9289 2802 9369 2818
rect 9289 2796 9308 2802
rect 9005 2770 9108 2780
rect 8959 2768 9108 2770
rect 9129 2768 9164 2780
rect 8798 2766 8960 2768
rect 8810 2746 8829 2766
rect 8844 2764 8874 2766
rect 8693 2738 8734 2746
rect 8816 2742 8829 2746
rect 8881 2750 8960 2766
rect 8992 2766 9164 2768
rect 8992 2750 9071 2766
rect 9078 2764 9108 2766
rect 8656 2728 8685 2738
rect 8699 2728 8728 2738
rect 8743 2728 8773 2742
rect 8816 2728 8859 2742
rect 8881 2738 9071 2750
rect 9136 2746 9142 2766
rect 8866 2728 8896 2738
rect 8897 2728 9055 2738
rect 9059 2728 9089 2738
rect 9093 2728 9123 2742
rect 9151 2728 9164 2766
rect 9236 2780 9265 2796
rect 9279 2780 9308 2796
rect 9323 2786 9353 2802
rect 9381 2780 9387 2828
rect 9390 2822 9409 2828
rect 9424 2822 9454 2830
rect 9390 2814 9454 2822
rect 9390 2798 9470 2814
rect 9486 2807 9548 2838
rect 9564 2807 9626 2838
rect 9695 2836 9744 2861
rect 9759 2836 9789 2852
rect 9658 2822 9688 2830
rect 9695 2828 9805 2836
rect 9658 2814 9703 2822
rect 9390 2796 9409 2798
rect 9424 2796 9470 2798
rect 9390 2780 9470 2796
rect 9497 2794 9532 2807
rect 9573 2804 9610 2807
rect 9573 2802 9615 2804
rect 9502 2791 9532 2794
rect 9511 2787 9518 2791
rect 9518 2786 9519 2787
rect 9477 2780 9487 2786
rect 9236 2772 9271 2780
rect 9236 2746 9237 2772
rect 9244 2746 9271 2772
rect 9179 2728 9209 2742
rect 9236 2738 9271 2746
rect 9273 2772 9314 2780
rect 9273 2746 9288 2772
rect 9295 2746 9314 2772
rect 9378 2768 9409 2780
rect 9424 2768 9527 2780
rect 9539 2770 9565 2796
rect 9580 2791 9610 2802
rect 9642 2798 9704 2814
rect 9642 2796 9688 2798
rect 9642 2780 9704 2796
rect 9716 2780 9722 2828
rect 9725 2820 9805 2828
rect 9725 2818 9744 2820
rect 9759 2818 9793 2820
rect 9725 2802 9805 2818
rect 9725 2780 9744 2802
rect 9759 2786 9789 2802
rect 9817 2796 9823 2870
rect 9826 2796 9845 2940
rect 9860 2796 9866 2940
rect 9875 2870 9888 2940
rect 9940 2936 9962 2940
rect 9933 2914 9962 2928
rect 10015 2914 10031 2928
rect 10069 2924 10075 2926
rect 10082 2924 10190 2940
rect 10197 2924 10203 2926
rect 10211 2924 10226 2940
rect 10292 2934 10311 2937
rect 9933 2912 10031 2914
rect 10058 2912 10226 2924
rect 10241 2914 10257 2928
rect 10292 2915 10314 2934
rect 10324 2928 10340 2929
rect 10323 2926 10340 2928
rect 10324 2921 10340 2926
rect 10314 2914 10320 2915
rect 10323 2914 10352 2921
rect 10241 2913 10352 2914
rect 10241 2912 10358 2913
rect 9917 2904 9968 2912
rect 10015 2904 10049 2912
rect 9917 2892 9942 2904
rect 9949 2892 9968 2904
rect 10022 2902 10049 2904
rect 10058 2902 10279 2912
rect 10314 2909 10320 2912
rect 10022 2898 10279 2902
rect 9917 2884 9968 2892
rect 10015 2884 10279 2898
rect 10323 2904 10358 2912
rect 9869 2836 9888 2870
rect 9933 2876 9962 2884
rect 9933 2870 9950 2876
rect 9933 2868 9967 2870
rect 10015 2868 10031 2884
rect 10032 2874 10240 2884
rect 10241 2874 10257 2884
rect 10305 2880 10320 2895
rect 10323 2892 10324 2904
rect 10331 2892 10358 2904
rect 10323 2884 10358 2892
rect 10323 2883 10352 2884
rect 10043 2870 10257 2874
rect 10058 2868 10257 2870
rect 10292 2870 10305 2880
rect 10323 2870 10340 2883
rect 10292 2868 10340 2870
rect 9934 2864 9967 2868
rect 9930 2862 9967 2864
rect 9930 2861 9997 2862
rect 9930 2856 9961 2861
rect 9967 2856 9997 2861
rect 9930 2852 9997 2856
rect 9903 2849 9997 2852
rect 9903 2842 9952 2849
rect 9903 2836 9933 2842
rect 9952 2837 9957 2842
rect 9869 2820 9949 2836
rect 9961 2828 9997 2849
rect 10058 2844 10247 2868
rect 10292 2867 10339 2868
rect 10305 2862 10339 2867
rect 10073 2841 10247 2844
rect 10066 2838 10247 2841
rect 10275 2861 10339 2862
rect 9869 2818 9888 2820
rect 9903 2818 9937 2820
rect 9869 2802 9949 2818
rect 9869 2796 9888 2802
rect 9585 2770 9688 2780
rect 9539 2768 9688 2770
rect 9709 2768 9744 2780
rect 9378 2766 9540 2768
rect 9390 2746 9409 2766
rect 9424 2764 9454 2766
rect 9273 2738 9314 2746
rect 9396 2742 9409 2746
rect 9461 2750 9540 2766
rect 9572 2766 9744 2768
rect 9572 2750 9651 2766
rect 9658 2764 9688 2766
rect 9236 2728 9265 2738
rect 9279 2728 9308 2738
rect 9323 2728 9353 2742
rect 9396 2728 9439 2742
rect 9461 2738 9651 2750
rect 9716 2746 9722 2766
rect 9446 2728 9476 2738
rect 9477 2728 9635 2738
rect 9639 2728 9669 2738
rect 9673 2728 9703 2742
rect 9731 2728 9744 2766
rect 9816 2780 9845 2796
rect 9859 2780 9888 2796
rect 9903 2786 9933 2802
rect 9961 2780 9967 2828
rect 9970 2822 9989 2828
rect 10004 2822 10034 2830
rect 9970 2814 10034 2822
rect 9970 2798 10050 2814
rect 10066 2807 10128 2838
rect 10144 2807 10206 2838
rect 10275 2836 10324 2861
rect 10339 2836 10369 2852
rect 10238 2822 10268 2830
rect 10275 2828 10385 2836
rect 10238 2814 10283 2822
rect 9970 2796 9989 2798
rect 10004 2796 10050 2798
rect 9970 2780 10050 2796
rect 10077 2794 10112 2807
rect 10153 2804 10190 2807
rect 10153 2802 10195 2804
rect 10082 2791 10112 2794
rect 10091 2787 10098 2791
rect 10098 2786 10099 2787
rect 10057 2780 10067 2786
rect 9816 2772 9851 2780
rect 9816 2746 9817 2772
rect 9824 2746 9851 2772
rect 9759 2728 9789 2742
rect 9816 2738 9851 2746
rect 9853 2772 9894 2780
rect 9853 2746 9868 2772
rect 9875 2746 9894 2772
rect 9958 2768 9989 2780
rect 10004 2768 10107 2780
rect 10119 2770 10145 2796
rect 10160 2791 10190 2802
rect 10222 2798 10284 2814
rect 10222 2796 10268 2798
rect 10222 2780 10284 2796
rect 10296 2780 10302 2828
rect 10305 2820 10385 2828
rect 10305 2818 10324 2820
rect 10339 2818 10373 2820
rect 10305 2802 10385 2818
rect 10305 2780 10324 2802
rect 10339 2786 10369 2802
rect 10397 2796 10403 2870
rect 10406 2796 10425 2940
rect 10440 2796 10446 2940
rect 10455 2870 10468 2940
rect 10520 2936 10542 2940
rect 10513 2914 10542 2928
rect 10595 2914 10611 2928
rect 10649 2924 10655 2926
rect 10662 2924 10770 2940
rect 10777 2924 10783 2926
rect 10791 2924 10806 2940
rect 10872 2934 10891 2937
rect 10513 2912 10611 2914
rect 10638 2912 10806 2924
rect 10821 2914 10837 2928
rect 10872 2915 10894 2934
rect 10904 2928 10920 2929
rect 10903 2926 10920 2928
rect 10904 2921 10920 2926
rect 10894 2914 10900 2915
rect 10903 2914 10932 2921
rect 10821 2913 10932 2914
rect 10821 2912 10938 2913
rect 10497 2904 10548 2912
rect 10595 2904 10629 2912
rect 10497 2892 10522 2904
rect 10529 2892 10548 2904
rect 10602 2902 10629 2904
rect 10638 2902 10859 2912
rect 10894 2909 10900 2912
rect 10602 2898 10859 2902
rect 10497 2884 10548 2892
rect 10595 2884 10859 2898
rect 10903 2904 10938 2912
rect 10449 2836 10468 2870
rect 10513 2876 10542 2884
rect 10513 2870 10530 2876
rect 10513 2868 10547 2870
rect 10595 2868 10611 2884
rect 10612 2874 10820 2884
rect 10821 2874 10837 2884
rect 10885 2880 10900 2895
rect 10903 2892 10904 2904
rect 10911 2892 10938 2904
rect 10903 2884 10938 2892
rect 10903 2883 10932 2884
rect 10623 2870 10837 2874
rect 10638 2868 10837 2870
rect 10872 2870 10885 2880
rect 10903 2870 10920 2883
rect 10872 2868 10920 2870
rect 10514 2864 10547 2868
rect 10510 2862 10547 2864
rect 10510 2861 10577 2862
rect 10510 2856 10541 2861
rect 10547 2856 10577 2861
rect 10510 2852 10577 2856
rect 10483 2849 10577 2852
rect 10483 2842 10532 2849
rect 10483 2836 10513 2842
rect 10532 2837 10537 2842
rect 10449 2820 10529 2836
rect 10541 2828 10577 2849
rect 10638 2844 10827 2868
rect 10872 2867 10919 2868
rect 10885 2862 10919 2867
rect 10653 2841 10827 2844
rect 10646 2838 10827 2841
rect 10855 2861 10919 2862
rect 10449 2818 10468 2820
rect 10483 2818 10517 2820
rect 10449 2802 10529 2818
rect 10449 2796 10468 2802
rect 10165 2770 10268 2780
rect 10119 2768 10268 2770
rect 10289 2768 10324 2780
rect 9958 2766 10120 2768
rect 9970 2746 9989 2766
rect 10004 2764 10034 2766
rect 9853 2738 9894 2746
rect 9976 2742 9989 2746
rect 10041 2750 10120 2766
rect 10152 2766 10324 2768
rect 10152 2750 10231 2766
rect 10238 2764 10268 2766
rect 9816 2728 9845 2738
rect 9859 2728 9888 2738
rect 9903 2728 9933 2742
rect 9976 2728 10019 2742
rect 10041 2738 10231 2750
rect 10296 2746 10302 2766
rect 10026 2728 10056 2738
rect 10057 2728 10215 2738
rect 10219 2728 10249 2738
rect 10253 2728 10283 2742
rect 10311 2728 10324 2766
rect 10396 2780 10425 2796
rect 10439 2780 10468 2796
rect 10483 2786 10513 2802
rect 10541 2780 10547 2828
rect 10550 2822 10569 2828
rect 10584 2822 10614 2830
rect 10550 2814 10614 2822
rect 10550 2798 10630 2814
rect 10646 2807 10708 2838
rect 10724 2807 10786 2838
rect 10855 2836 10904 2861
rect 10919 2836 10949 2852
rect 10818 2822 10848 2830
rect 10855 2828 10965 2836
rect 10818 2814 10863 2822
rect 10550 2796 10569 2798
rect 10584 2796 10630 2798
rect 10550 2780 10630 2796
rect 10657 2794 10692 2807
rect 10733 2804 10770 2807
rect 10733 2802 10775 2804
rect 10662 2791 10692 2794
rect 10671 2787 10678 2791
rect 10678 2786 10679 2787
rect 10637 2780 10647 2786
rect 10396 2772 10431 2780
rect 10396 2746 10397 2772
rect 10404 2746 10431 2772
rect 10339 2728 10369 2742
rect 10396 2738 10431 2746
rect 10433 2772 10474 2780
rect 10433 2746 10448 2772
rect 10455 2746 10474 2772
rect 10538 2768 10569 2780
rect 10584 2768 10687 2780
rect 10699 2770 10725 2796
rect 10740 2791 10770 2802
rect 10802 2798 10864 2814
rect 10802 2796 10848 2798
rect 10802 2780 10864 2796
rect 10876 2780 10882 2828
rect 10885 2820 10965 2828
rect 10885 2818 10904 2820
rect 10919 2818 10953 2820
rect 10885 2802 10965 2818
rect 10885 2780 10904 2802
rect 10919 2786 10949 2802
rect 10977 2796 10983 2870
rect 10986 2796 11005 2940
rect 11020 2796 11026 2940
rect 11035 2870 11048 2940
rect 11100 2936 11122 2940
rect 11093 2914 11122 2928
rect 11175 2914 11191 2928
rect 11229 2924 11235 2926
rect 11242 2924 11350 2940
rect 11357 2924 11363 2926
rect 11371 2924 11386 2940
rect 11452 2934 11471 2937
rect 11093 2912 11191 2914
rect 11218 2912 11386 2924
rect 11401 2914 11417 2928
rect 11452 2915 11474 2934
rect 11484 2928 11500 2929
rect 11483 2926 11500 2928
rect 11484 2921 11500 2926
rect 11474 2914 11480 2915
rect 11483 2914 11512 2921
rect 11401 2913 11512 2914
rect 11401 2912 11518 2913
rect 11077 2904 11128 2912
rect 11175 2904 11209 2912
rect 11077 2892 11102 2904
rect 11109 2892 11128 2904
rect 11182 2902 11209 2904
rect 11218 2902 11439 2912
rect 11474 2909 11480 2912
rect 11182 2898 11439 2902
rect 11077 2884 11128 2892
rect 11175 2884 11439 2898
rect 11483 2904 11518 2912
rect 11029 2836 11048 2870
rect 11093 2876 11122 2884
rect 11093 2870 11110 2876
rect 11093 2868 11127 2870
rect 11175 2868 11191 2884
rect 11192 2874 11400 2884
rect 11401 2874 11417 2884
rect 11465 2880 11480 2895
rect 11483 2892 11484 2904
rect 11491 2892 11518 2904
rect 11483 2884 11518 2892
rect 11483 2883 11512 2884
rect 11203 2870 11417 2874
rect 11218 2868 11417 2870
rect 11452 2870 11465 2880
rect 11483 2870 11500 2883
rect 11452 2868 11500 2870
rect 11094 2864 11127 2868
rect 11090 2862 11127 2864
rect 11090 2861 11157 2862
rect 11090 2856 11121 2861
rect 11127 2856 11157 2861
rect 11090 2852 11157 2856
rect 11063 2849 11157 2852
rect 11063 2842 11112 2849
rect 11063 2836 11093 2842
rect 11112 2837 11117 2842
rect 11029 2820 11109 2836
rect 11121 2828 11157 2849
rect 11218 2844 11407 2868
rect 11452 2867 11499 2868
rect 11465 2862 11499 2867
rect 11233 2841 11407 2844
rect 11226 2838 11407 2841
rect 11435 2861 11499 2862
rect 11029 2818 11048 2820
rect 11063 2818 11097 2820
rect 11029 2802 11109 2818
rect 11029 2796 11048 2802
rect 10745 2770 10848 2780
rect 10699 2768 10848 2770
rect 10869 2768 10904 2780
rect 10538 2766 10700 2768
rect 10550 2746 10569 2766
rect 10584 2764 10614 2766
rect 10433 2738 10474 2746
rect 10556 2742 10569 2746
rect 10621 2750 10700 2766
rect 10732 2766 10904 2768
rect 10732 2750 10811 2766
rect 10818 2764 10848 2766
rect 10396 2728 10425 2738
rect 10439 2728 10468 2738
rect 10483 2728 10513 2742
rect 10556 2728 10599 2742
rect 10621 2738 10811 2750
rect 10876 2746 10882 2766
rect 10606 2728 10636 2738
rect 10637 2728 10795 2738
rect 10799 2728 10829 2738
rect 10833 2728 10863 2742
rect 10891 2728 10904 2766
rect 10976 2780 11005 2796
rect 11019 2780 11048 2796
rect 11063 2786 11093 2802
rect 11121 2780 11127 2828
rect 11130 2822 11149 2828
rect 11164 2822 11194 2830
rect 11130 2814 11194 2822
rect 11130 2798 11210 2814
rect 11226 2807 11288 2838
rect 11304 2807 11366 2838
rect 11435 2836 11484 2861
rect 11499 2836 11529 2852
rect 11398 2822 11428 2830
rect 11435 2828 11545 2836
rect 11398 2814 11443 2822
rect 11130 2796 11149 2798
rect 11164 2796 11210 2798
rect 11130 2780 11210 2796
rect 11237 2794 11272 2807
rect 11313 2804 11350 2807
rect 11313 2802 11355 2804
rect 11242 2791 11272 2794
rect 11251 2787 11258 2791
rect 11258 2786 11259 2787
rect 11217 2780 11227 2786
rect 10976 2772 11011 2780
rect 10976 2746 10977 2772
rect 10984 2746 11011 2772
rect 10919 2728 10949 2742
rect 10976 2738 11011 2746
rect 11013 2772 11054 2780
rect 11013 2746 11028 2772
rect 11035 2746 11054 2772
rect 11118 2768 11149 2780
rect 11164 2768 11267 2780
rect 11279 2770 11305 2796
rect 11320 2791 11350 2802
rect 11382 2798 11444 2814
rect 11382 2796 11428 2798
rect 11382 2780 11444 2796
rect 11456 2780 11462 2828
rect 11465 2820 11545 2828
rect 11465 2818 11484 2820
rect 11499 2818 11533 2820
rect 11465 2802 11545 2818
rect 11465 2780 11484 2802
rect 11499 2786 11529 2802
rect 11557 2796 11563 2870
rect 11566 2796 11585 2940
rect 11600 2796 11606 2940
rect 11615 2870 11628 2940
rect 11680 2936 11702 2940
rect 11673 2914 11702 2928
rect 11755 2914 11771 2928
rect 11809 2924 11815 2926
rect 11822 2924 11930 2940
rect 11937 2924 11943 2926
rect 11951 2924 11966 2940
rect 12032 2934 12051 2937
rect 11673 2912 11771 2914
rect 11798 2912 11966 2924
rect 11981 2914 11997 2928
rect 12032 2915 12054 2934
rect 12064 2928 12080 2929
rect 12063 2926 12080 2928
rect 12064 2921 12080 2926
rect 12054 2914 12060 2915
rect 12063 2914 12092 2921
rect 11981 2913 12092 2914
rect 11981 2912 12098 2913
rect 11657 2904 11708 2912
rect 11755 2904 11789 2912
rect 11657 2892 11682 2904
rect 11689 2892 11708 2904
rect 11762 2902 11789 2904
rect 11798 2902 12019 2912
rect 12054 2909 12060 2912
rect 11762 2898 12019 2902
rect 11657 2884 11708 2892
rect 11755 2884 12019 2898
rect 12063 2904 12098 2912
rect 11609 2836 11628 2870
rect 11673 2876 11702 2884
rect 11673 2870 11690 2876
rect 11673 2868 11707 2870
rect 11755 2868 11771 2884
rect 11772 2874 11980 2884
rect 11981 2874 11997 2884
rect 12045 2880 12060 2895
rect 12063 2892 12064 2904
rect 12071 2892 12098 2904
rect 12063 2884 12098 2892
rect 12063 2883 12092 2884
rect 11783 2870 11997 2874
rect 11798 2868 11997 2870
rect 12032 2870 12045 2880
rect 12063 2870 12080 2883
rect 12032 2868 12080 2870
rect 11674 2864 11707 2868
rect 11670 2862 11707 2864
rect 11670 2861 11737 2862
rect 11670 2856 11701 2861
rect 11707 2856 11737 2861
rect 11670 2852 11737 2856
rect 11643 2849 11737 2852
rect 11643 2842 11692 2849
rect 11643 2836 11673 2842
rect 11692 2837 11697 2842
rect 11609 2820 11689 2836
rect 11701 2828 11737 2849
rect 11798 2844 11987 2868
rect 12032 2867 12079 2868
rect 12045 2862 12079 2867
rect 11813 2841 11987 2844
rect 11806 2838 11987 2841
rect 12015 2861 12079 2862
rect 11609 2818 11628 2820
rect 11643 2818 11677 2820
rect 11609 2802 11689 2818
rect 11609 2796 11628 2802
rect 11325 2770 11428 2780
rect 11279 2768 11428 2770
rect 11449 2768 11484 2780
rect 11118 2766 11280 2768
rect 11130 2746 11149 2766
rect 11164 2764 11194 2766
rect 11013 2738 11054 2746
rect 11136 2742 11149 2746
rect 11201 2750 11280 2766
rect 11312 2766 11484 2768
rect 11312 2750 11391 2766
rect 11398 2764 11428 2766
rect 10976 2728 11005 2738
rect 11019 2728 11048 2738
rect 11063 2728 11093 2742
rect 11136 2728 11179 2742
rect 11201 2738 11391 2750
rect 11456 2746 11462 2766
rect 11186 2728 11216 2738
rect 11217 2728 11375 2738
rect 11379 2728 11409 2738
rect 11413 2728 11443 2742
rect 11471 2728 11484 2766
rect 11556 2780 11585 2796
rect 11599 2780 11628 2796
rect 11643 2786 11673 2802
rect 11701 2780 11707 2828
rect 11710 2822 11729 2828
rect 11744 2822 11774 2830
rect 11710 2814 11774 2822
rect 11710 2798 11790 2814
rect 11806 2807 11868 2838
rect 11884 2807 11946 2838
rect 12015 2836 12064 2861
rect 12079 2836 12109 2852
rect 11978 2822 12008 2830
rect 12015 2828 12125 2836
rect 11978 2814 12023 2822
rect 11710 2796 11729 2798
rect 11744 2796 11790 2798
rect 11710 2780 11790 2796
rect 11817 2794 11852 2807
rect 11893 2804 11930 2807
rect 11893 2802 11935 2804
rect 11822 2791 11852 2794
rect 11831 2787 11838 2791
rect 11838 2786 11839 2787
rect 11797 2780 11807 2786
rect 11556 2772 11591 2780
rect 11556 2746 11557 2772
rect 11564 2746 11591 2772
rect 11499 2728 11529 2742
rect 11556 2738 11591 2746
rect 11593 2772 11634 2780
rect 11593 2746 11608 2772
rect 11615 2746 11634 2772
rect 11698 2768 11729 2780
rect 11744 2768 11847 2780
rect 11859 2770 11885 2796
rect 11900 2791 11930 2802
rect 11962 2798 12024 2814
rect 11962 2796 12008 2798
rect 11962 2780 12024 2796
rect 12036 2780 12042 2828
rect 12045 2820 12125 2828
rect 12045 2818 12064 2820
rect 12079 2818 12113 2820
rect 12045 2802 12125 2818
rect 12045 2780 12064 2802
rect 12079 2786 12109 2802
rect 12137 2796 12143 2870
rect 12146 2796 12165 2940
rect 12180 2796 12186 2940
rect 12195 2870 12208 2940
rect 12260 2936 12282 2940
rect 12253 2914 12282 2928
rect 12335 2914 12351 2928
rect 12389 2924 12395 2926
rect 12402 2924 12510 2940
rect 12517 2924 12523 2926
rect 12531 2924 12546 2940
rect 12612 2934 12631 2937
rect 12253 2912 12351 2914
rect 12378 2912 12546 2924
rect 12561 2914 12577 2928
rect 12612 2915 12634 2934
rect 12644 2928 12660 2929
rect 12643 2926 12660 2928
rect 12644 2921 12660 2926
rect 12634 2914 12640 2915
rect 12643 2914 12672 2921
rect 12561 2913 12672 2914
rect 12561 2912 12678 2913
rect 12237 2904 12288 2912
rect 12335 2904 12369 2912
rect 12237 2892 12262 2904
rect 12269 2892 12288 2904
rect 12342 2902 12369 2904
rect 12378 2902 12599 2912
rect 12634 2909 12640 2912
rect 12342 2898 12599 2902
rect 12237 2884 12288 2892
rect 12335 2884 12599 2898
rect 12643 2904 12678 2912
rect 12189 2836 12208 2870
rect 12253 2876 12282 2884
rect 12253 2870 12270 2876
rect 12253 2868 12287 2870
rect 12335 2868 12351 2884
rect 12352 2874 12560 2884
rect 12561 2874 12577 2884
rect 12625 2880 12640 2895
rect 12643 2892 12644 2904
rect 12651 2892 12678 2904
rect 12643 2884 12678 2892
rect 12643 2883 12672 2884
rect 12363 2870 12577 2874
rect 12378 2868 12577 2870
rect 12612 2870 12625 2880
rect 12643 2870 12660 2883
rect 12612 2868 12660 2870
rect 12254 2864 12287 2868
rect 12250 2862 12287 2864
rect 12250 2861 12317 2862
rect 12250 2856 12281 2861
rect 12287 2856 12317 2861
rect 12250 2852 12317 2856
rect 12223 2849 12317 2852
rect 12223 2842 12272 2849
rect 12223 2836 12253 2842
rect 12272 2837 12277 2842
rect 12189 2820 12269 2836
rect 12281 2828 12317 2849
rect 12378 2844 12567 2868
rect 12612 2867 12659 2868
rect 12625 2862 12659 2867
rect 12393 2841 12567 2844
rect 12386 2838 12567 2841
rect 12595 2861 12659 2862
rect 12189 2818 12208 2820
rect 12223 2818 12257 2820
rect 12189 2802 12269 2818
rect 12189 2796 12208 2802
rect 11905 2770 12008 2780
rect 11859 2768 12008 2770
rect 12029 2768 12064 2780
rect 11698 2766 11860 2768
rect 11710 2746 11729 2766
rect 11744 2764 11774 2766
rect 11593 2738 11634 2746
rect 11716 2742 11729 2746
rect 11781 2750 11860 2766
rect 11892 2766 12064 2768
rect 11892 2750 11971 2766
rect 11978 2764 12008 2766
rect 11556 2728 11585 2738
rect 11599 2728 11628 2738
rect 11643 2728 11673 2742
rect 11716 2728 11759 2742
rect 11781 2738 11971 2750
rect 12036 2746 12042 2766
rect 11766 2728 11796 2738
rect 11797 2728 11955 2738
rect 11959 2728 11989 2738
rect 11993 2728 12023 2742
rect 12051 2728 12064 2766
rect 12136 2780 12165 2796
rect 12179 2780 12208 2796
rect 12223 2786 12253 2802
rect 12281 2780 12287 2828
rect 12290 2822 12309 2828
rect 12324 2822 12354 2830
rect 12290 2814 12354 2822
rect 12290 2798 12370 2814
rect 12386 2807 12448 2838
rect 12464 2807 12526 2838
rect 12595 2836 12644 2861
rect 12659 2836 12689 2852
rect 12558 2822 12588 2830
rect 12595 2828 12705 2836
rect 12558 2814 12603 2822
rect 12290 2796 12309 2798
rect 12324 2796 12370 2798
rect 12290 2780 12370 2796
rect 12397 2794 12432 2807
rect 12473 2804 12510 2807
rect 12473 2802 12515 2804
rect 12402 2791 12432 2794
rect 12411 2787 12418 2791
rect 12418 2786 12419 2787
rect 12377 2780 12387 2786
rect 12136 2772 12171 2780
rect 12136 2746 12137 2772
rect 12144 2746 12171 2772
rect 12079 2728 12109 2742
rect 12136 2738 12171 2746
rect 12173 2772 12214 2780
rect 12173 2746 12188 2772
rect 12195 2746 12214 2772
rect 12278 2768 12309 2780
rect 12324 2768 12427 2780
rect 12439 2770 12465 2796
rect 12480 2791 12510 2802
rect 12542 2798 12604 2814
rect 12542 2796 12588 2798
rect 12542 2780 12604 2796
rect 12616 2780 12622 2828
rect 12625 2820 12705 2828
rect 12625 2818 12644 2820
rect 12659 2818 12693 2820
rect 12625 2802 12705 2818
rect 12625 2780 12644 2802
rect 12659 2786 12689 2802
rect 12717 2796 12723 2870
rect 12726 2796 12745 2940
rect 12760 2796 12766 2940
rect 12775 2870 12788 2940
rect 12840 2936 12862 2940
rect 12833 2914 12862 2928
rect 12915 2914 12931 2928
rect 12969 2924 12975 2926
rect 12982 2924 13090 2940
rect 13097 2924 13103 2926
rect 13111 2924 13126 2940
rect 13192 2934 13211 2937
rect 12833 2912 12931 2914
rect 12958 2912 13126 2924
rect 13141 2914 13157 2928
rect 13192 2915 13214 2934
rect 13224 2928 13240 2929
rect 13223 2926 13240 2928
rect 13224 2921 13240 2926
rect 13214 2914 13220 2915
rect 13223 2914 13252 2921
rect 13141 2913 13252 2914
rect 13141 2912 13258 2913
rect 12817 2904 12868 2912
rect 12915 2904 12949 2912
rect 12817 2892 12842 2904
rect 12849 2892 12868 2904
rect 12922 2902 12949 2904
rect 12958 2902 13179 2912
rect 13214 2909 13220 2912
rect 12922 2898 13179 2902
rect 12817 2884 12868 2892
rect 12915 2884 13179 2898
rect 13223 2904 13258 2912
rect 12769 2836 12788 2870
rect 12833 2876 12862 2884
rect 12833 2870 12850 2876
rect 12833 2868 12867 2870
rect 12915 2868 12931 2884
rect 12932 2874 13140 2884
rect 13141 2874 13157 2884
rect 13205 2880 13220 2895
rect 13223 2892 13224 2904
rect 13231 2892 13258 2904
rect 13223 2884 13258 2892
rect 13223 2883 13252 2884
rect 12943 2870 13157 2874
rect 12958 2868 13157 2870
rect 13192 2870 13205 2880
rect 13223 2870 13240 2883
rect 13192 2868 13240 2870
rect 12834 2864 12867 2868
rect 12830 2862 12867 2864
rect 12830 2861 12897 2862
rect 12830 2856 12861 2861
rect 12867 2856 12897 2861
rect 12830 2852 12897 2856
rect 12803 2849 12897 2852
rect 12803 2842 12852 2849
rect 12803 2836 12833 2842
rect 12852 2837 12857 2842
rect 12769 2820 12849 2836
rect 12861 2828 12897 2849
rect 12958 2844 13147 2868
rect 13192 2867 13239 2868
rect 13205 2862 13239 2867
rect 12973 2841 13147 2844
rect 12966 2838 13147 2841
rect 13175 2861 13239 2862
rect 12769 2818 12788 2820
rect 12803 2818 12837 2820
rect 12769 2802 12849 2818
rect 12769 2796 12788 2802
rect 12485 2770 12588 2780
rect 12439 2768 12588 2770
rect 12609 2768 12644 2780
rect 12278 2766 12440 2768
rect 12290 2746 12309 2766
rect 12324 2764 12354 2766
rect 12173 2738 12214 2746
rect 12296 2742 12309 2746
rect 12361 2750 12440 2766
rect 12472 2766 12644 2768
rect 12472 2750 12551 2766
rect 12558 2764 12588 2766
rect 12136 2728 12165 2738
rect 12179 2728 12208 2738
rect 12223 2728 12253 2742
rect 12296 2728 12339 2742
rect 12361 2738 12551 2750
rect 12616 2746 12622 2766
rect 12346 2728 12376 2738
rect 12377 2728 12535 2738
rect 12539 2728 12569 2738
rect 12573 2728 12603 2742
rect 12631 2728 12644 2766
rect 12716 2780 12745 2796
rect 12759 2780 12788 2796
rect 12803 2786 12833 2802
rect 12861 2780 12867 2828
rect 12870 2822 12889 2828
rect 12904 2822 12934 2830
rect 12870 2814 12934 2822
rect 12870 2798 12950 2814
rect 12966 2807 13028 2838
rect 13044 2807 13106 2838
rect 13175 2836 13224 2861
rect 13239 2836 13269 2852
rect 13138 2822 13168 2830
rect 13175 2828 13285 2836
rect 13138 2814 13183 2822
rect 12870 2796 12889 2798
rect 12904 2796 12950 2798
rect 12870 2780 12950 2796
rect 12977 2794 13012 2807
rect 13053 2804 13090 2807
rect 13053 2802 13095 2804
rect 12982 2791 13012 2794
rect 12991 2787 12998 2791
rect 12998 2786 12999 2787
rect 12957 2780 12967 2786
rect 12716 2772 12751 2780
rect 12716 2746 12717 2772
rect 12724 2746 12751 2772
rect 12659 2728 12689 2742
rect 12716 2738 12751 2746
rect 12753 2772 12794 2780
rect 12753 2746 12768 2772
rect 12775 2746 12794 2772
rect 12858 2768 12889 2780
rect 12904 2768 13007 2780
rect 13019 2770 13045 2796
rect 13060 2791 13090 2802
rect 13122 2798 13184 2814
rect 13122 2796 13168 2798
rect 13122 2780 13184 2796
rect 13196 2780 13202 2828
rect 13205 2820 13285 2828
rect 13205 2818 13224 2820
rect 13239 2818 13273 2820
rect 13205 2802 13285 2818
rect 13205 2780 13224 2802
rect 13239 2786 13269 2802
rect 13297 2796 13303 2870
rect 13306 2796 13325 2940
rect 13340 2796 13346 2940
rect 13355 2870 13368 2940
rect 13420 2936 13442 2940
rect 13413 2914 13442 2928
rect 13495 2914 13511 2928
rect 13549 2924 13555 2926
rect 13562 2924 13670 2940
rect 13677 2924 13683 2926
rect 13691 2924 13706 2940
rect 13772 2934 13791 2937
rect 13413 2912 13511 2914
rect 13538 2912 13706 2924
rect 13721 2914 13737 2928
rect 13772 2915 13794 2934
rect 13804 2928 13820 2929
rect 13803 2926 13820 2928
rect 13804 2921 13820 2926
rect 13794 2914 13800 2915
rect 13803 2914 13832 2921
rect 13721 2913 13832 2914
rect 13721 2912 13838 2913
rect 13397 2904 13448 2912
rect 13495 2904 13529 2912
rect 13397 2892 13422 2904
rect 13429 2892 13448 2904
rect 13502 2902 13529 2904
rect 13538 2902 13759 2912
rect 13794 2909 13800 2912
rect 13502 2898 13759 2902
rect 13397 2884 13448 2892
rect 13495 2884 13759 2898
rect 13803 2904 13838 2912
rect 13349 2836 13368 2870
rect 13413 2876 13442 2884
rect 13413 2870 13430 2876
rect 13413 2868 13447 2870
rect 13495 2868 13511 2884
rect 13512 2874 13720 2884
rect 13721 2874 13737 2884
rect 13785 2880 13800 2895
rect 13803 2892 13804 2904
rect 13811 2892 13838 2904
rect 13803 2884 13838 2892
rect 13803 2883 13832 2884
rect 13523 2870 13737 2874
rect 13538 2868 13737 2870
rect 13772 2870 13785 2880
rect 13803 2870 13820 2883
rect 13772 2868 13820 2870
rect 13414 2864 13447 2868
rect 13410 2862 13447 2864
rect 13410 2861 13477 2862
rect 13410 2856 13441 2861
rect 13447 2856 13477 2861
rect 13410 2852 13477 2856
rect 13383 2849 13477 2852
rect 13383 2842 13432 2849
rect 13383 2836 13413 2842
rect 13432 2837 13437 2842
rect 13349 2820 13429 2836
rect 13441 2828 13477 2849
rect 13538 2844 13727 2868
rect 13772 2867 13819 2868
rect 13785 2862 13819 2867
rect 13553 2841 13727 2844
rect 13546 2838 13727 2841
rect 13755 2861 13819 2862
rect 13349 2818 13368 2820
rect 13383 2818 13417 2820
rect 13349 2802 13429 2818
rect 13349 2796 13368 2802
rect 13065 2770 13168 2780
rect 13019 2768 13168 2770
rect 13189 2768 13224 2780
rect 12858 2766 13020 2768
rect 12870 2746 12889 2766
rect 12904 2764 12934 2766
rect 12753 2738 12794 2746
rect 12876 2742 12889 2746
rect 12941 2750 13020 2766
rect 13052 2766 13224 2768
rect 13052 2750 13131 2766
rect 13138 2764 13168 2766
rect 12716 2728 12745 2738
rect 12759 2728 12788 2738
rect 12803 2728 12833 2742
rect 12876 2728 12919 2742
rect 12941 2738 13131 2750
rect 13196 2746 13202 2766
rect 12926 2728 12956 2738
rect 12957 2728 13115 2738
rect 13119 2728 13149 2738
rect 13153 2728 13183 2742
rect 13211 2728 13224 2766
rect 13296 2780 13325 2796
rect 13339 2780 13368 2796
rect 13383 2786 13413 2802
rect 13441 2780 13447 2828
rect 13450 2822 13469 2828
rect 13484 2822 13514 2830
rect 13450 2814 13514 2822
rect 13450 2798 13530 2814
rect 13546 2807 13608 2838
rect 13624 2807 13686 2838
rect 13755 2836 13804 2861
rect 13819 2836 13849 2852
rect 13718 2822 13748 2830
rect 13755 2828 13865 2836
rect 13718 2814 13763 2822
rect 13450 2796 13469 2798
rect 13484 2796 13530 2798
rect 13450 2780 13530 2796
rect 13557 2794 13592 2807
rect 13633 2804 13670 2807
rect 13633 2802 13675 2804
rect 13562 2791 13592 2794
rect 13571 2787 13578 2791
rect 13578 2786 13579 2787
rect 13537 2780 13547 2786
rect 13296 2772 13331 2780
rect 13296 2746 13297 2772
rect 13304 2746 13331 2772
rect 13239 2728 13269 2742
rect 13296 2738 13331 2746
rect 13333 2772 13374 2780
rect 13333 2746 13348 2772
rect 13355 2746 13374 2772
rect 13438 2768 13469 2780
rect 13484 2768 13587 2780
rect 13599 2770 13625 2796
rect 13640 2791 13670 2802
rect 13702 2798 13764 2814
rect 13702 2796 13748 2798
rect 13702 2780 13764 2796
rect 13776 2780 13782 2828
rect 13785 2820 13865 2828
rect 13785 2818 13804 2820
rect 13819 2818 13853 2820
rect 13785 2802 13865 2818
rect 13785 2780 13804 2802
rect 13819 2786 13849 2802
rect 13877 2796 13883 2870
rect 13886 2796 13905 2940
rect 13920 2796 13926 2940
rect 13935 2870 13948 2940
rect 14000 2936 14022 2940
rect 13993 2914 14022 2928
rect 14075 2914 14091 2928
rect 14129 2924 14135 2926
rect 14142 2924 14250 2940
rect 14257 2924 14263 2926
rect 14271 2924 14286 2940
rect 14352 2934 14371 2937
rect 13993 2912 14091 2914
rect 14118 2912 14286 2924
rect 14301 2914 14317 2928
rect 14352 2915 14374 2934
rect 14384 2928 14400 2929
rect 14383 2926 14400 2928
rect 14384 2921 14400 2926
rect 14374 2914 14380 2915
rect 14383 2914 14412 2921
rect 14301 2913 14412 2914
rect 14301 2912 14418 2913
rect 13977 2904 14028 2912
rect 14075 2904 14109 2912
rect 13977 2892 14002 2904
rect 14009 2892 14028 2904
rect 14082 2902 14109 2904
rect 14118 2902 14339 2912
rect 14374 2909 14380 2912
rect 14082 2898 14339 2902
rect 13977 2884 14028 2892
rect 14075 2884 14339 2898
rect 14383 2904 14418 2912
rect 13929 2836 13948 2870
rect 13993 2876 14022 2884
rect 13993 2870 14010 2876
rect 13993 2868 14027 2870
rect 14075 2868 14091 2884
rect 14092 2874 14300 2884
rect 14301 2874 14317 2884
rect 14365 2880 14380 2895
rect 14383 2892 14384 2904
rect 14391 2892 14418 2904
rect 14383 2884 14418 2892
rect 14383 2883 14412 2884
rect 14103 2870 14317 2874
rect 14118 2868 14317 2870
rect 14352 2870 14365 2880
rect 14383 2870 14400 2883
rect 14352 2868 14400 2870
rect 13994 2864 14027 2868
rect 13990 2862 14027 2864
rect 13990 2861 14057 2862
rect 13990 2856 14021 2861
rect 14027 2856 14057 2861
rect 13990 2852 14057 2856
rect 13963 2849 14057 2852
rect 13963 2842 14012 2849
rect 13963 2836 13993 2842
rect 14012 2837 14017 2842
rect 13929 2820 14009 2836
rect 14021 2828 14057 2849
rect 14118 2844 14307 2868
rect 14352 2867 14399 2868
rect 14365 2862 14399 2867
rect 14133 2841 14307 2844
rect 14126 2838 14307 2841
rect 14335 2861 14399 2862
rect 13929 2818 13948 2820
rect 13963 2818 13997 2820
rect 13929 2802 14009 2818
rect 13929 2796 13948 2802
rect 13645 2770 13748 2780
rect 13599 2768 13748 2770
rect 13769 2768 13804 2780
rect 13438 2766 13600 2768
rect 13450 2746 13469 2766
rect 13484 2764 13514 2766
rect 13333 2738 13374 2746
rect 13456 2742 13469 2746
rect 13521 2750 13600 2766
rect 13632 2766 13804 2768
rect 13632 2750 13711 2766
rect 13718 2764 13748 2766
rect 13296 2728 13325 2738
rect 13339 2728 13368 2738
rect 13383 2728 13413 2742
rect 13456 2728 13499 2742
rect 13521 2738 13711 2750
rect 13776 2746 13782 2766
rect 13506 2728 13536 2738
rect 13537 2728 13695 2738
rect 13699 2728 13729 2738
rect 13733 2728 13763 2742
rect 13791 2728 13804 2766
rect 13876 2780 13905 2796
rect 13919 2780 13948 2796
rect 13963 2786 13993 2802
rect 14021 2780 14027 2828
rect 14030 2822 14049 2828
rect 14064 2822 14094 2830
rect 14030 2814 14094 2822
rect 14030 2798 14110 2814
rect 14126 2807 14188 2838
rect 14204 2807 14266 2838
rect 14335 2836 14384 2861
rect 14399 2836 14429 2852
rect 14298 2822 14328 2830
rect 14335 2828 14445 2836
rect 14298 2814 14343 2822
rect 14030 2796 14049 2798
rect 14064 2796 14110 2798
rect 14030 2780 14110 2796
rect 14137 2794 14172 2807
rect 14213 2804 14250 2807
rect 14213 2802 14255 2804
rect 14142 2791 14172 2794
rect 14151 2787 14158 2791
rect 14158 2786 14159 2787
rect 14117 2780 14127 2786
rect 13876 2772 13911 2780
rect 13876 2746 13877 2772
rect 13884 2746 13911 2772
rect 13819 2728 13849 2742
rect 13876 2738 13911 2746
rect 13913 2772 13954 2780
rect 13913 2746 13928 2772
rect 13935 2746 13954 2772
rect 14018 2768 14049 2780
rect 14064 2768 14167 2780
rect 14179 2770 14205 2796
rect 14220 2791 14250 2802
rect 14282 2798 14344 2814
rect 14282 2796 14328 2798
rect 14282 2780 14344 2796
rect 14356 2780 14362 2828
rect 14365 2820 14445 2828
rect 14365 2818 14384 2820
rect 14399 2818 14433 2820
rect 14365 2802 14445 2818
rect 14365 2780 14384 2802
rect 14399 2786 14429 2802
rect 14457 2796 14463 2870
rect 14466 2796 14485 2940
rect 14500 2796 14506 2940
rect 14515 2870 14528 2940
rect 14580 2936 14602 2940
rect 14573 2914 14602 2928
rect 14655 2914 14671 2928
rect 14709 2924 14715 2926
rect 14722 2924 14830 2940
rect 14837 2924 14843 2926
rect 14851 2924 14866 2940
rect 14932 2934 14951 2937
rect 14573 2912 14671 2914
rect 14698 2912 14866 2924
rect 14881 2914 14897 2928
rect 14932 2915 14954 2934
rect 14964 2928 14980 2929
rect 14963 2926 14980 2928
rect 14964 2921 14980 2926
rect 14954 2914 14960 2915
rect 14963 2914 14992 2921
rect 14881 2913 14992 2914
rect 14881 2912 14998 2913
rect 14557 2904 14608 2912
rect 14655 2904 14689 2912
rect 14557 2892 14582 2904
rect 14589 2892 14608 2904
rect 14662 2902 14689 2904
rect 14698 2902 14919 2912
rect 14954 2909 14960 2912
rect 14662 2898 14919 2902
rect 14557 2884 14608 2892
rect 14655 2884 14919 2898
rect 14963 2904 14998 2912
rect 14509 2836 14528 2870
rect 14573 2876 14602 2884
rect 14573 2870 14590 2876
rect 14573 2868 14607 2870
rect 14655 2868 14671 2884
rect 14672 2874 14880 2884
rect 14881 2874 14897 2884
rect 14945 2880 14960 2895
rect 14963 2892 14964 2904
rect 14971 2892 14998 2904
rect 14963 2884 14998 2892
rect 14963 2883 14992 2884
rect 14683 2870 14897 2874
rect 14698 2868 14897 2870
rect 14932 2870 14945 2880
rect 14963 2870 14980 2883
rect 14932 2868 14980 2870
rect 14574 2864 14607 2868
rect 14570 2862 14607 2864
rect 14570 2861 14637 2862
rect 14570 2856 14601 2861
rect 14607 2856 14637 2861
rect 14570 2852 14637 2856
rect 14543 2849 14637 2852
rect 14543 2842 14592 2849
rect 14543 2836 14573 2842
rect 14592 2837 14597 2842
rect 14509 2820 14589 2836
rect 14601 2828 14637 2849
rect 14698 2844 14887 2868
rect 14932 2867 14979 2868
rect 14945 2862 14979 2867
rect 14713 2841 14887 2844
rect 14706 2838 14887 2841
rect 14915 2861 14979 2862
rect 14509 2818 14528 2820
rect 14543 2818 14577 2820
rect 14509 2802 14589 2818
rect 14509 2796 14528 2802
rect 14225 2770 14328 2780
rect 14179 2768 14328 2770
rect 14349 2768 14384 2780
rect 14018 2766 14180 2768
rect 14030 2746 14049 2766
rect 14064 2764 14094 2766
rect 13913 2738 13954 2746
rect 14036 2742 14049 2746
rect 14101 2750 14180 2766
rect 14212 2766 14384 2768
rect 14212 2750 14291 2766
rect 14298 2764 14328 2766
rect 13876 2728 13905 2738
rect 13919 2728 13948 2738
rect 13963 2728 13993 2742
rect 14036 2728 14079 2742
rect 14101 2738 14291 2750
rect 14356 2746 14362 2766
rect 14086 2728 14116 2738
rect 14117 2728 14275 2738
rect 14279 2728 14309 2738
rect 14313 2728 14343 2742
rect 14371 2728 14384 2766
rect 14456 2780 14485 2796
rect 14499 2780 14528 2796
rect 14543 2786 14573 2802
rect 14601 2780 14607 2828
rect 14610 2822 14629 2828
rect 14644 2822 14674 2830
rect 14610 2814 14674 2822
rect 14610 2798 14690 2814
rect 14706 2807 14768 2838
rect 14784 2807 14846 2838
rect 14915 2836 14964 2861
rect 14979 2836 15009 2852
rect 14878 2822 14908 2830
rect 14915 2828 15025 2836
rect 14878 2814 14923 2822
rect 14610 2796 14629 2798
rect 14644 2796 14690 2798
rect 14610 2780 14690 2796
rect 14717 2794 14752 2807
rect 14793 2804 14830 2807
rect 14793 2802 14835 2804
rect 14722 2791 14752 2794
rect 14731 2787 14738 2791
rect 14738 2786 14739 2787
rect 14697 2780 14707 2786
rect 14456 2772 14491 2780
rect 14456 2746 14457 2772
rect 14464 2746 14491 2772
rect 14399 2728 14429 2742
rect 14456 2738 14491 2746
rect 14493 2772 14534 2780
rect 14493 2746 14508 2772
rect 14515 2746 14534 2772
rect 14598 2768 14629 2780
rect 14644 2768 14747 2780
rect 14759 2770 14785 2796
rect 14800 2791 14830 2802
rect 14862 2798 14924 2814
rect 14862 2796 14908 2798
rect 14862 2780 14924 2796
rect 14936 2780 14942 2828
rect 14945 2820 15025 2828
rect 14945 2818 14964 2820
rect 14979 2818 15013 2820
rect 14945 2802 15025 2818
rect 14945 2780 14964 2802
rect 14979 2786 15009 2802
rect 15037 2796 15043 2870
rect 15046 2796 15065 2940
rect 15080 2796 15086 2940
rect 15095 2870 15108 2940
rect 15160 2936 15182 2940
rect 15153 2914 15182 2928
rect 15235 2914 15251 2928
rect 15289 2924 15295 2926
rect 15302 2924 15410 2940
rect 15417 2924 15423 2926
rect 15431 2924 15446 2940
rect 15512 2934 15531 2937
rect 15153 2912 15251 2914
rect 15278 2912 15446 2924
rect 15461 2914 15477 2928
rect 15512 2915 15534 2934
rect 15544 2928 15560 2929
rect 15543 2926 15560 2928
rect 15544 2921 15560 2926
rect 15534 2914 15540 2915
rect 15543 2914 15572 2921
rect 15461 2913 15572 2914
rect 15461 2912 15578 2913
rect 15137 2904 15188 2912
rect 15235 2904 15269 2912
rect 15137 2892 15162 2904
rect 15169 2892 15188 2904
rect 15242 2902 15269 2904
rect 15278 2902 15499 2912
rect 15534 2909 15540 2912
rect 15242 2898 15499 2902
rect 15137 2884 15188 2892
rect 15235 2884 15499 2898
rect 15543 2904 15578 2912
rect 15089 2836 15108 2870
rect 15153 2876 15182 2884
rect 15153 2870 15170 2876
rect 15153 2868 15187 2870
rect 15235 2868 15251 2884
rect 15252 2874 15460 2884
rect 15461 2874 15477 2884
rect 15525 2880 15540 2895
rect 15543 2892 15544 2904
rect 15551 2892 15578 2904
rect 15543 2884 15578 2892
rect 15543 2883 15572 2884
rect 15263 2870 15477 2874
rect 15278 2868 15477 2870
rect 15512 2870 15525 2880
rect 15543 2870 15560 2883
rect 15512 2868 15560 2870
rect 15154 2864 15187 2868
rect 15150 2862 15187 2864
rect 15150 2861 15217 2862
rect 15150 2856 15181 2861
rect 15187 2856 15217 2861
rect 15150 2852 15217 2856
rect 15123 2849 15217 2852
rect 15123 2842 15172 2849
rect 15123 2836 15153 2842
rect 15172 2837 15177 2842
rect 15089 2820 15169 2836
rect 15181 2828 15217 2849
rect 15278 2844 15467 2868
rect 15512 2867 15559 2868
rect 15525 2862 15559 2867
rect 15293 2841 15467 2844
rect 15286 2838 15467 2841
rect 15495 2861 15559 2862
rect 15089 2818 15108 2820
rect 15123 2818 15157 2820
rect 15089 2802 15169 2818
rect 15089 2796 15108 2802
rect 14805 2770 14908 2780
rect 14759 2768 14908 2770
rect 14929 2768 14964 2780
rect 14598 2766 14760 2768
rect 14610 2746 14629 2766
rect 14644 2764 14674 2766
rect 14493 2738 14534 2746
rect 14616 2742 14629 2746
rect 14681 2750 14760 2766
rect 14792 2766 14964 2768
rect 14792 2750 14871 2766
rect 14878 2764 14908 2766
rect 14456 2728 14485 2738
rect 14499 2728 14528 2738
rect 14543 2728 14573 2742
rect 14616 2728 14659 2742
rect 14681 2738 14871 2750
rect 14936 2746 14942 2766
rect 14666 2728 14696 2738
rect 14697 2728 14855 2738
rect 14859 2728 14889 2738
rect 14893 2728 14923 2742
rect 14951 2728 14964 2766
rect 15036 2780 15065 2796
rect 15079 2780 15108 2796
rect 15123 2786 15153 2802
rect 15181 2780 15187 2828
rect 15190 2822 15209 2828
rect 15224 2822 15254 2830
rect 15190 2814 15254 2822
rect 15190 2798 15270 2814
rect 15286 2807 15348 2838
rect 15364 2807 15426 2838
rect 15495 2836 15544 2861
rect 15559 2836 15589 2852
rect 15458 2822 15488 2830
rect 15495 2828 15605 2836
rect 15458 2814 15503 2822
rect 15190 2796 15209 2798
rect 15224 2796 15270 2798
rect 15190 2780 15270 2796
rect 15297 2794 15332 2807
rect 15373 2804 15410 2807
rect 15373 2802 15415 2804
rect 15302 2791 15332 2794
rect 15311 2787 15318 2791
rect 15318 2786 15319 2787
rect 15277 2780 15287 2786
rect 15036 2772 15071 2780
rect 15036 2746 15037 2772
rect 15044 2746 15071 2772
rect 14979 2728 15009 2742
rect 15036 2738 15071 2746
rect 15073 2772 15114 2780
rect 15073 2746 15088 2772
rect 15095 2746 15114 2772
rect 15178 2768 15209 2780
rect 15224 2768 15327 2780
rect 15339 2770 15365 2796
rect 15380 2791 15410 2802
rect 15442 2798 15504 2814
rect 15442 2796 15488 2798
rect 15442 2780 15504 2796
rect 15516 2780 15522 2828
rect 15525 2820 15605 2828
rect 15525 2818 15544 2820
rect 15559 2818 15593 2820
rect 15525 2802 15605 2818
rect 15525 2780 15544 2802
rect 15559 2786 15589 2802
rect 15617 2796 15623 2870
rect 15626 2796 15645 2940
rect 15660 2796 15666 2940
rect 15675 2870 15688 2940
rect 15740 2936 15762 2940
rect 15733 2914 15762 2928
rect 15815 2914 15831 2928
rect 15869 2924 15875 2926
rect 15882 2924 15990 2940
rect 15997 2924 16003 2926
rect 16011 2924 16026 2940
rect 16092 2934 16111 2937
rect 15733 2912 15831 2914
rect 15858 2912 16026 2924
rect 16041 2914 16057 2928
rect 16092 2915 16114 2934
rect 16124 2928 16140 2929
rect 16123 2926 16140 2928
rect 16124 2921 16140 2926
rect 16114 2914 16120 2915
rect 16123 2914 16152 2921
rect 16041 2913 16152 2914
rect 16041 2912 16158 2913
rect 15717 2904 15768 2912
rect 15815 2904 15849 2912
rect 15717 2892 15742 2904
rect 15749 2892 15768 2904
rect 15822 2902 15849 2904
rect 15858 2902 16079 2912
rect 16114 2909 16120 2912
rect 15822 2898 16079 2902
rect 15717 2884 15768 2892
rect 15815 2884 16079 2898
rect 16123 2904 16158 2912
rect 15669 2836 15688 2870
rect 15733 2876 15762 2884
rect 15733 2870 15750 2876
rect 15733 2868 15767 2870
rect 15815 2868 15831 2884
rect 15832 2874 16040 2884
rect 16041 2874 16057 2884
rect 16105 2880 16120 2895
rect 16123 2892 16124 2904
rect 16131 2892 16158 2904
rect 16123 2884 16158 2892
rect 16123 2883 16152 2884
rect 15843 2870 16057 2874
rect 15858 2868 16057 2870
rect 16092 2870 16105 2880
rect 16123 2870 16140 2883
rect 16092 2868 16140 2870
rect 15734 2864 15767 2868
rect 15730 2862 15767 2864
rect 15730 2861 15797 2862
rect 15730 2856 15761 2861
rect 15767 2856 15797 2861
rect 15730 2852 15797 2856
rect 15703 2849 15797 2852
rect 15703 2842 15752 2849
rect 15703 2836 15733 2842
rect 15752 2837 15757 2842
rect 15669 2820 15749 2836
rect 15761 2828 15797 2849
rect 15858 2844 16047 2868
rect 16092 2867 16139 2868
rect 16105 2862 16139 2867
rect 15873 2841 16047 2844
rect 15866 2838 16047 2841
rect 16075 2861 16139 2862
rect 15669 2818 15688 2820
rect 15703 2818 15737 2820
rect 15669 2802 15749 2818
rect 15669 2796 15688 2802
rect 15385 2770 15488 2780
rect 15339 2768 15488 2770
rect 15509 2768 15544 2780
rect 15178 2766 15340 2768
rect 15190 2746 15209 2766
rect 15224 2764 15254 2766
rect 15073 2738 15114 2746
rect 15196 2742 15209 2746
rect 15261 2750 15340 2766
rect 15372 2766 15544 2768
rect 15372 2750 15451 2766
rect 15458 2764 15488 2766
rect 15036 2728 15065 2738
rect 15079 2728 15108 2738
rect 15123 2728 15153 2742
rect 15196 2728 15239 2742
rect 15261 2738 15451 2750
rect 15516 2746 15522 2766
rect 15246 2728 15276 2738
rect 15277 2728 15435 2738
rect 15439 2728 15469 2738
rect 15473 2728 15503 2742
rect 15531 2728 15544 2766
rect 15616 2780 15645 2796
rect 15659 2780 15688 2796
rect 15703 2786 15733 2802
rect 15761 2780 15767 2828
rect 15770 2822 15789 2828
rect 15804 2822 15834 2830
rect 15770 2814 15834 2822
rect 15770 2798 15850 2814
rect 15866 2807 15928 2838
rect 15944 2807 16006 2838
rect 16075 2836 16124 2861
rect 16139 2836 16169 2852
rect 16038 2822 16068 2830
rect 16075 2828 16185 2836
rect 16038 2814 16083 2822
rect 15770 2796 15789 2798
rect 15804 2796 15850 2798
rect 15770 2780 15850 2796
rect 15877 2794 15912 2807
rect 15953 2804 15990 2807
rect 15953 2802 15995 2804
rect 15882 2791 15912 2794
rect 15891 2787 15898 2791
rect 15898 2786 15899 2787
rect 15857 2780 15867 2786
rect 15616 2772 15651 2780
rect 15616 2746 15617 2772
rect 15624 2746 15651 2772
rect 15559 2728 15589 2742
rect 15616 2738 15651 2746
rect 15653 2772 15694 2780
rect 15653 2746 15668 2772
rect 15675 2746 15694 2772
rect 15758 2768 15789 2780
rect 15804 2768 15907 2780
rect 15919 2770 15945 2796
rect 15960 2791 15990 2802
rect 16022 2798 16084 2814
rect 16022 2796 16068 2798
rect 16022 2780 16084 2796
rect 16096 2780 16102 2828
rect 16105 2820 16185 2828
rect 16105 2818 16124 2820
rect 16139 2818 16173 2820
rect 16105 2802 16185 2818
rect 16105 2780 16124 2802
rect 16139 2786 16169 2802
rect 16197 2796 16203 2870
rect 16206 2796 16225 2940
rect 16240 2796 16246 2940
rect 16255 2870 16268 2940
rect 16320 2936 16342 2940
rect 16313 2914 16342 2928
rect 16395 2914 16411 2928
rect 16449 2924 16455 2926
rect 16462 2924 16570 2940
rect 16577 2924 16583 2926
rect 16591 2924 16606 2940
rect 16672 2934 16691 2937
rect 16313 2912 16411 2914
rect 16438 2912 16606 2924
rect 16621 2914 16637 2928
rect 16672 2915 16694 2934
rect 16704 2928 16720 2929
rect 16703 2926 16720 2928
rect 16704 2921 16720 2926
rect 16694 2914 16700 2915
rect 16703 2914 16732 2921
rect 16621 2913 16732 2914
rect 16621 2912 16738 2913
rect 16297 2904 16348 2912
rect 16395 2904 16429 2912
rect 16297 2892 16322 2904
rect 16329 2892 16348 2904
rect 16402 2902 16429 2904
rect 16438 2902 16659 2912
rect 16694 2909 16700 2912
rect 16402 2898 16659 2902
rect 16297 2884 16348 2892
rect 16395 2884 16659 2898
rect 16703 2904 16738 2912
rect 16249 2836 16268 2870
rect 16313 2876 16342 2884
rect 16313 2870 16330 2876
rect 16313 2868 16347 2870
rect 16395 2868 16411 2884
rect 16412 2874 16620 2884
rect 16621 2874 16637 2884
rect 16685 2880 16700 2895
rect 16703 2892 16704 2904
rect 16711 2892 16738 2904
rect 16703 2884 16738 2892
rect 16703 2883 16732 2884
rect 16423 2870 16637 2874
rect 16438 2868 16637 2870
rect 16672 2870 16685 2880
rect 16703 2870 16720 2883
rect 16672 2868 16720 2870
rect 16314 2864 16347 2868
rect 16310 2862 16347 2864
rect 16310 2861 16377 2862
rect 16310 2856 16341 2861
rect 16347 2856 16377 2861
rect 16310 2852 16377 2856
rect 16283 2849 16377 2852
rect 16283 2842 16332 2849
rect 16283 2836 16313 2842
rect 16332 2837 16337 2842
rect 16249 2820 16329 2836
rect 16341 2828 16377 2849
rect 16438 2844 16627 2868
rect 16672 2867 16719 2868
rect 16685 2862 16719 2867
rect 16453 2841 16627 2844
rect 16446 2838 16627 2841
rect 16655 2861 16719 2862
rect 16249 2818 16268 2820
rect 16283 2818 16317 2820
rect 16249 2802 16329 2818
rect 16249 2796 16268 2802
rect 15965 2770 16068 2780
rect 15919 2768 16068 2770
rect 16089 2768 16124 2780
rect 15758 2766 15920 2768
rect 15770 2746 15789 2766
rect 15804 2764 15834 2766
rect 15653 2738 15694 2746
rect 15776 2742 15789 2746
rect 15841 2750 15920 2766
rect 15952 2766 16124 2768
rect 15952 2750 16031 2766
rect 16038 2764 16068 2766
rect 15616 2728 15645 2738
rect 15659 2728 15688 2738
rect 15703 2728 15733 2742
rect 15776 2728 15819 2742
rect 15841 2738 16031 2750
rect 16096 2746 16102 2766
rect 15826 2728 15856 2738
rect 15857 2728 16015 2738
rect 16019 2728 16049 2738
rect 16053 2728 16083 2742
rect 16111 2728 16124 2766
rect 16196 2780 16225 2796
rect 16239 2780 16268 2796
rect 16283 2786 16313 2802
rect 16341 2780 16347 2828
rect 16350 2822 16369 2828
rect 16384 2822 16414 2830
rect 16350 2814 16414 2822
rect 16350 2798 16430 2814
rect 16446 2807 16508 2838
rect 16524 2807 16586 2838
rect 16655 2836 16704 2861
rect 16719 2836 16749 2852
rect 16618 2822 16648 2830
rect 16655 2828 16765 2836
rect 16618 2814 16663 2822
rect 16350 2796 16369 2798
rect 16384 2796 16430 2798
rect 16350 2780 16430 2796
rect 16457 2794 16492 2807
rect 16533 2804 16570 2807
rect 16533 2802 16575 2804
rect 16462 2791 16492 2794
rect 16471 2787 16478 2791
rect 16478 2786 16479 2787
rect 16437 2780 16447 2786
rect 16196 2772 16231 2780
rect 16196 2746 16197 2772
rect 16204 2746 16231 2772
rect 16139 2728 16169 2742
rect 16196 2738 16231 2746
rect 16233 2772 16274 2780
rect 16233 2746 16248 2772
rect 16255 2746 16274 2772
rect 16338 2768 16369 2780
rect 16384 2768 16487 2780
rect 16499 2770 16525 2796
rect 16540 2791 16570 2802
rect 16602 2798 16664 2814
rect 16602 2796 16648 2798
rect 16602 2780 16664 2796
rect 16676 2780 16682 2828
rect 16685 2820 16765 2828
rect 16685 2818 16704 2820
rect 16719 2818 16753 2820
rect 16685 2802 16765 2818
rect 16685 2780 16704 2802
rect 16719 2786 16749 2802
rect 16777 2796 16783 2870
rect 16786 2796 16805 2940
rect 16820 2796 16826 2940
rect 16835 2870 16848 2940
rect 16900 2936 16922 2940
rect 16893 2914 16922 2928
rect 16975 2914 16991 2928
rect 17029 2924 17035 2926
rect 17042 2924 17150 2940
rect 17157 2924 17163 2926
rect 17171 2924 17186 2940
rect 17252 2934 17271 2937
rect 16893 2912 16991 2914
rect 17018 2912 17186 2924
rect 17201 2914 17217 2928
rect 17252 2915 17274 2934
rect 17284 2928 17300 2929
rect 17283 2926 17300 2928
rect 17284 2921 17300 2926
rect 17274 2914 17280 2915
rect 17283 2914 17312 2921
rect 17201 2913 17312 2914
rect 17201 2912 17318 2913
rect 16877 2904 16928 2912
rect 16975 2904 17009 2912
rect 16877 2892 16902 2904
rect 16909 2892 16928 2904
rect 16982 2902 17009 2904
rect 17018 2902 17239 2912
rect 17274 2909 17280 2912
rect 16982 2898 17239 2902
rect 16877 2884 16928 2892
rect 16975 2884 17239 2898
rect 17283 2904 17318 2912
rect 16829 2836 16848 2870
rect 16893 2876 16922 2884
rect 16893 2870 16910 2876
rect 16893 2868 16927 2870
rect 16975 2868 16991 2884
rect 16992 2874 17200 2884
rect 17201 2874 17217 2884
rect 17265 2880 17280 2895
rect 17283 2892 17284 2904
rect 17291 2892 17318 2904
rect 17283 2884 17318 2892
rect 17283 2883 17312 2884
rect 17003 2870 17217 2874
rect 17018 2868 17217 2870
rect 17252 2870 17265 2880
rect 17283 2870 17300 2883
rect 17252 2868 17300 2870
rect 16894 2864 16927 2868
rect 16890 2862 16927 2864
rect 16890 2861 16957 2862
rect 16890 2856 16921 2861
rect 16927 2856 16957 2861
rect 16890 2852 16957 2856
rect 16863 2849 16957 2852
rect 16863 2842 16912 2849
rect 16863 2836 16893 2842
rect 16912 2837 16917 2842
rect 16829 2820 16909 2836
rect 16921 2828 16957 2849
rect 17018 2844 17207 2868
rect 17252 2867 17299 2868
rect 17265 2862 17299 2867
rect 17033 2841 17207 2844
rect 17026 2838 17207 2841
rect 17235 2861 17299 2862
rect 16829 2818 16848 2820
rect 16863 2818 16897 2820
rect 16829 2802 16909 2818
rect 16829 2796 16848 2802
rect 16545 2770 16648 2780
rect 16499 2768 16648 2770
rect 16669 2768 16704 2780
rect 16338 2766 16500 2768
rect 16350 2746 16369 2766
rect 16384 2764 16414 2766
rect 16233 2738 16274 2746
rect 16356 2742 16369 2746
rect 16421 2750 16500 2766
rect 16532 2766 16704 2768
rect 16532 2750 16611 2766
rect 16618 2764 16648 2766
rect 16196 2728 16225 2738
rect 16239 2728 16268 2738
rect 16283 2728 16313 2742
rect 16356 2728 16399 2742
rect 16421 2738 16611 2750
rect 16676 2746 16682 2766
rect 16406 2728 16436 2738
rect 16437 2728 16595 2738
rect 16599 2728 16629 2738
rect 16633 2728 16663 2742
rect 16691 2728 16704 2766
rect 16776 2780 16805 2796
rect 16819 2780 16848 2796
rect 16863 2786 16893 2802
rect 16921 2780 16927 2828
rect 16930 2822 16949 2828
rect 16964 2822 16994 2830
rect 16930 2814 16994 2822
rect 16930 2798 17010 2814
rect 17026 2807 17088 2838
rect 17104 2807 17166 2838
rect 17235 2836 17284 2861
rect 17299 2836 17329 2852
rect 17198 2822 17228 2830
rect 17235 2828 17345 2836
rect 17198 2814 17243 2822
rect 16930 2796 16949 2798
rect 16964 2796 17010 2798
rect 16930 2780 17010 2796
rect 17037 2794 17072 2807
rect 17113 2804 17150 2807
rect 17113 2802 17155 2804
rect 17042 2791 17072 2794
rect 17051 2787 17058 2791
rect 17058 2786 17059 2787
rect 17017 2780 17027 2786
rect 16776 2772 16811 2780
rect 16776 2746 16777 2772
rect 16784 2746 16811 2772
rect 16719 2728 16749 2742
rect 16776 2738 16811 2746
rect 16813 2772 16854 2780
rect 16813 2746 16828 2772
rect 16835 2746 16854 2772
rect 16918 2768 16949 2780
rect 16964 2768 17067 2780
rect 17079 2770 17105 2796
rect 17120 2791 17150 2802
rect 17182 2798 17244 2814
rect 17182 2796 17228 2798
rect 17182 2780 17244 2796
rect 17256 2780 17262 2828
rect 17265 2820 17345 2828
rect 17265 2818 17284 2820
rect 17299 2818 17333 2820
rect 17265 2802 17345 2818
rect 17265 2780 17284 2802
rect 17299 2786 17329 2802
rect 17357 2796 17363 2870
rect 17366 2796 17385 2940
rect 17400 2796 17406 2940
rect 17415 2870 17428 2940
rect 17480 2936 17502 2940
rect 17473 2914 17502 2928
rect 17555 2914 17571 2928
rect 17609 2924 17615 2926
rect 17622 2924 17730 2940
rect 17737 2924 17743 2926
rect 17751 2924 17766 2940
rect 17832 2934 17851 2937
rect 17473 2912 17571 2914
rect 17598 2912 17766 2924
rect 17781 2914 17797 2928
rect 17832 2915 17854 2934
rect 17864 2928 17880 2929
rect 17863 2926 17880 2928
rect 17864 2921 17880 2926
rect 17854 2914 17860 2915
rect 17863 2914 17892 2921
rect 17781 2913 17892 2914
rect 17781 2912 17898 2913
rect 17457 2904 17508 2912
rect 17555 2904 17589 2912
rect 17457 2892 17482 2904
rect 17489 2892 17508 2904
rect 17562 2902 17589 2904
rect 17598 2902 17819 2912
rect 17854 2909 17860 2912
rect 17562 2898 17819 2902
rect 17457 2884 17508 2892
rect 17555 2884 17819 2898
rect 17863 2904 17898 2912
rect 17409 2836 17428 2870
rect 17473 2876 17502 2884
rect 17473 2870 17490 2876
rect 17473 2868 17507 2870
rect 17555 2868 17571 2884
rect 17572 2874 17780 2884
rect 17781 2874 17797 2884
rect 17845 2880 17860 2895
rect 17863 2892 17864 2904
rect 17871 2892 17898 2904
rect 17863 2884 17898 2892
rect 17863 2883 17892 2884
rect 17583 2870 17797 2874
rect 17598 2868 17797 2870
rect 17832 2870 17845 2880
rect 17863 2870 17880 2883
rect 17832 2868 17880 2870
rect 17474 2864 17507 2868
rect 17470 2862 17507 2864
rect 17470 2861 17537 2862
rect 17470 2856 17501 2861
rect 17507 2856 17537 2861
rect 17470 2852 17537 2856
rect 17443 2849 17537 2852
rect 17443 2842 17492 2849
rect 17443 2836 17473 2842
rect 17492 2837 17497 2842
rect 17409 2820 17489 2836
rect 17501 2828 17537 2849
rect 17598 2844 17787 2868
rect 17832 2867 17879 2868
rect 17845 2862 17879 2867
rect 17613 2841 17787 2844
rect 17606 2838 17787 2841
rect 17815 2861 17879 2862
rect 17409 2818 17428 2820
rect 17443 2818 17477 2820
rect 17409 2802 17489 2818
rect 17409 2796 17428 2802
rect 17125 2770 17228 2780
rect 17079 2768 17228 2770
rect 17249 2768 17284 2780
rect 16918 2766 17080 2768
rect 16930 2746 16949 2766
rect 16964 2764 16994 2766
rect 16813 2738 16854 2746
rect 16936 2742 16949 2746
rect 17001 2750 17080 2766
rect 17112 2766 17284 2768
rect 17112 2750 17191 2766
rect 17198 2764 17228 2766
rect 16776 2728 16805 2738
rect 16819 2728 16848 2738
rect 16863 2728 16893 2742
rect 16936 2728 16979 2742
rect 17001 2738 17191 2750
rect 17256 2746 17262 2766
rect 16986 2728 17016 2738
rect 17017 2728 17175 2738
rect 17179 2728 17209 2738
rect 17213 2728 17243 2742
rect 17271 2728 17284 2766
rect 17356 2780 17385 2796
rect 17399 2780 17428 2796
rect 17443 2786 17473 2802
rect 17501 2780 17507 2828
rect 17510 2822 17529 2828
rect 17544 2822 17574 2830
rect 17510 2814 17574 2822
rect 17510 2798 17590 2814
rect 17606 2807 17668 2838
rect 17684 2807 17746 2838
rect 17815 2836 17864 2861
rect 17879 2836 17909 2852
rect 17778 2822 17808 2830
rect 17815 2828 17925 2836
rect 17778 2814 17823 2822
rect 17510 2796 17529 2798
rect 17544 2796 17590 2798
rect 17510 2780 17590 2796
rect 17617 2794 17652 2807
rect 17693 2804 17730 2807
rect 17693 2802 17735 2804
rect 17622 2791 17652 2794
rect 17631 2787 17638 2791
rect 17638 2786 17639 2787
rect 17597 2780 17607 2786
rect 17356 2772 17391 2780
rect 17356 2746 17357 2772
rect 17364 2746 17391 2772
rect 17299 2728 17329 2742
rect 17356 2738 17391 2746
rect 17393 2772 17434 2780
rect 17393 2746 17408 2772
rect 17415 2746 17434 2772
rect 17498 2768 17529 2780
rect 17544 2768 17647 2780
rect 17659 2770 17685 2796
rect 17700 2791 17730 2802
rect 17762 2798 17824 2814
rect 17762 2796 17808 2798
rect 17762 2780 17824 2796
rect 17836 2780 17842 2828
rect 17845 2820 17925 2828
rect 17845 2818 17864 2820
rect 17879 2818 17913 2820
rect 17845 2802 17925 2818
rect 17845 2780 17864 2802
rect 17879 2786 17909 2802
rect 17937 2796 17943 2870
rect 17946 2796 17965 2940
rect 17980 2796 17986 2940
rect 17995 2870 18008 2940
rect 18060 2936 18082 2940
rect 18053 2914 18082 2928
rect 18135 2914 18151 2928
rect 18189 2924 18195 2926
rect 18202 2924 18310 2940
rect 18317 2924 18323 2926
rect 18331 2924 18346 2940
rect 18412 2934 18431 2937
rect 18053 2912 18151 2914
rect 18178 2912 18346 2924
rect 18361 2914 18377 2928
rect 18412 2915 18434 2934
rect 18444 2928 18460 2929
rect 18443 2926 18460 2928
rect 18444 2921 18460 2926
rect 18434 2914 18440 2915
rect 18443 2914 18472 2921
rect 18361 2913 18472 2914
rect 18361 2912 18478 2913
rect 18037 2904 18088 2912
rect 18135 2904 18169 2912
rect 18037 2892 18062 2904
rect 18069 2892 18088 2904
rect 18142 2902 18169 2904
rect 18178 2902 18399 2912
rect 18434 2909 18440 2912
rect 18142 2898 18399 2902
rect 18037 2884 18088 2892
rect 18135 2884 18399 2898
rect 18443 2904 18478 2912
rect 17989 2836 18008 2870
rect 18053 2876 18082 2884
rect 18053 2870 18070 2876
rect 18053 2868 18087 2870
rect 18135 2868 18151 2884
rect 18152 2874 18360 2884
rect 18361 2874 18377 2884
rect 18425 2880 18440 2895
rect 18443 2892 18444 2904
rect 18451 2892 18478 2904
rect 18443 2884 18478 2892
rect 18443 2883 18472 2884
rect 18163 2870 18377 2874
rect 18178 2868 18377 2870
rect 18412 2870 18425 2880
rect 18443 2870 18460 2883
rect 18412 2868 18460 2870
rect 18054 2864 18087 2868
rect 18050 2862 18087 2864
rect 18050 2861 18117 2862
rect 18050 2856 18081 2861
rect 18087 2856 18117 2861
rect 18050 2852 18117 2856
rect 18023 2849 18117 2852
rect 18023 2842 18072 2849
rect 18023 2836 18053 2842
rect 18072 2837 18077 2842
rect 17989 2820 18069 2836
rect 18081 2828 18117 2849
rect 18178 2844 18367 2868
rect 18412 2867 18459 2868
rect 18425 2862 18459 2867
rect 18193 2841 18367 2844
rect 18186 2838 18367 2841
rect 18395 2861 18459 2862
rect 17989 2818 18008 2820
rect 18023 2818 18057 2820
rect 17989 2802 18069 2818
rect 17989 2796 18008 2802
rect 17705 2770 17808 2780
rect 17659 2768 17808 2770
rect 17829 2768 17864 2780
rect 17498 2766 17660 2768
rect 17510 2746 17529 2766
rect 17544 2764 17574 2766
rect 17393 2738 17434 2746
rect 17516 2742 17529 2746
rect 17581 2750 17660 2766
rect 17692 2766 17864 2768
rect 17692 2750 17771 2766
rect 17778 2764 17808 2766
rect 17356 2728 17385 2738
rect 17399 2728 17428 2738
rect 17443 2728 17473 2742
rect 17516 2728 17559 2742
rect 17581 2738 17771 2750
rect 17836 2746 17842 2766
rect 17566 2728 17596 2738
rect 17597 2728 17755 2738
rect 17759 2728 17789 2738
rect 17793 2728 17823 2742
rect 17851 2728 17864 2766
rect 17936 2780 17965 2796
rect 17979 2780 18008 2796
rect 18023 2786 18053 2802
rect 18081 2780 18087 2828
rect 18090 2822 18109 2828
rect 18124 2822 18154 2830
rect 18090 2814 18154 2822
rect 18090 2798 18170 2814
rect 18186 2807 18248 2838
rect 18264 2807 18326 2838
rect 18395 2836 18444 2861
rect 18459 2836 18489 2852
rect 18358 2822 18388 2830
rect 18395 2828 18505 2836
rect 18358 2814 18403 2822
rect 18090 2796 18109 2798
rect 18124 2796 18170 2798
rect 18090 2780 18170 2796
rect 18197 2794 18232 2807
rect 18273 2804 18310 2807
rect 18273 2802 18315 2804
rect 18202 2791 18232 2794
rect 18211 2787 18218 2791
rect 18218 2786 18219 2787
rect 18177 2780 18187 2786
rect 17936 2772 17971 2780
rect 17936 2746 17937 2772
rect 17944 2746 17971 2772
rect 17879 2728 17909 2742
rect 17936 2738 17971 2746
rect 17973 2772 18014 2780
rect 17973 2746 17988 2772
rect 17995 2746 18014 2772
rect 18078 2768 18109 2780
rect 18124 2768 18227 2780
rect 18239 2770 18265 2796
rect 18280 2791 18310 2802
rect 18342 2798 18404 2814
rect 18342 2796 18388 2798
rect 18342 2780 18404 2796
rect 18416 2780 18422 2828
rect 18425 2820 18505 2828
rect 18425 2818 18444 2820
rect 18459 2818 18493 2820
rect 18425 2802 18505 2818
rect 18425 2780 18444 2802
rect 18459 2786 18489 2802
rect 18517 2796 18523 2870
rect 18532 2796 18545 2940
rect 18285 2770 18388 2780
rect 18239 2768 18388 2770
rect 18409 2768 18444 2780
rect 18078 2766 18240 2768
rect 18090 2746 18109 2766
rect 18124 2764 18154 2766
rect 17973 2738 18014 2746
rect 18096 2742 18109 2746
rect 18161 2750 18240 2766
rect 18272 2766 18444 2768
rect 18272 2750 18351 2766
rect 18358 2764 18388 2766
rect 17936 2728 17965 2738
rect 17979 2728 18008 2738
rect 18023 2728 18053 2742
rect 18096 2728 18139 2742
rect 18161 2738 18351 2750
rect 18416 2746 18422 2766
rect 18146 2728 18176 2738
rect 18177 2728 18335 2738
rect 18339 2728 18369 2738
rect 18373 2728 18403 2742
rect 18431 2728 18444 2766
rect 18516 2780 18545 2796
rect 18516 2772 18551 2780
rect 18516 2746 18517 2772
rect 18524 2746 18551 2772
rect 18459 2728 18489 2742
rect 18516 2738 18551 2746
rect 18516 2728 18545 2738
rect -1 2722 18545 2728
rect 0 2714 18545 2722
rect 15 2684 28 2714
rect 43 2700 73 2714
rect 116 2700 159 2714
rect 166 2700 386 2714
rect 393 2700 423 2714
rect 83 2686 98 2698
rect 117 2686 130 2700
rect 198 2696 351 2700
rect 80 2684 102 2686
rect 180 2684 372 2696
rect 451 2684 464 2714
rect 479 2700 509 2714
rect 546 2684 565 2714
rect 580 2684 586 2714
rect 595 2684 608 2714
rect 623 2700 653 2714
rect 696 2700 739 2714
rect 746 2700 966 2714
rect 973 2700 1003 2714
rect 663 2686 678 2698
rect 697 2686 710 2700
rect 778 2696 931 2700
rect 660 2684 682 2686
rect 760 2684 952 2696
rect 1031 2684 1044 2714
rect 1059 2700 1089 2714
rect 1126 2684 1145 2714
rect 1160 2684 1166 2714
rect 1175 2684 1188 2714
rect 1203 2700 1233 2714
rect 1276 2700 1319 2714
rect 1326 2700 1546 2714
rect 1553 2700 1583 2714
rect 1243 2686 1258 2698
rect 1277 2686 1290 2700
rect 1358 2696 1511 2700
rect 1240 2684 1262 2686
rect 1340 2684 1532 2696
rect 1611 2684 1624 2714
rect 1639 2700 1669 2714
rect 1706 2684 1725 2714
rect 1740 2684 1746 2714
rect 1755 2684 1768 2714
rect 1783 2700 1813 2714
rect 1856 2700 1899 2714
rect 1906 2700 2126 2714
rect 2133 2700 2163 2714
rect 1823 2686 1838 2698
rect 1857 2686 1870 2700
rect 1938 2696 2091 2700
rect 1820 2684 1842 2686
rect 1920 2684 2112 2696
rect 2191 2684 2204 2714
rect 2219 2700 2249 2714
rect 2286 2684 2305 2714
rect 2320 2684 2326 2714
rect 2335 2684 2348 2714
rect 2363 2700 2393 2714
rect 2436 2700 2479 2714
rect 2486 2700 2706 2714
rect 2713 2700 2743 2714
rect 2403 2686 2418 2698
rect 2437 2686 2450 2700
rect 2518 2696 2671 2700
rect 2400 2684 2422 2686
rect 2500 2684 2692 2696
rect 2771 2684 2784 2714
rect 2799 2700 2829 2714
rect 2866 2684 2885 2714
rect 2900 2684 2906 2714
rect 2915 2684 2928 2714
rect 2943 2700 2973 2714
rect 3016 2700 3059 2714
rect 3066 2700 3286 2714
rect 3293 2700 3323 2714
rect 2983 2686 2998 2698
rect 3017 2686 3030 2700
rect 3098 2696 3251 2700
rect 2980 2684 3002 2686
rect 3080 2684 3272 2696
rect 3351 2684 3364 2714
rect 3379 2700 3409 2714
rect 3446 2684 3465 2714
rect 3480 2684 3486 2714
rect 3495 2684 3508 2714
rect 3523 2700 3553 2714
rect 3596 2700 3639 2714
rect 3646 2700 3866 2714
rect 3873 2700 3903 2714
rect 3563 2686 3578 2698
rect 3597 2686 3610 2700
rect 3678 2696 3831 2700
rect 3560 2684 3582 2686
rect 3660 2684 3852 2696
rect 3931 2684 3944 2714
rect 3959 2700 3989 2714
rect 4026 2684 4045 2714
rect 4060 2684 4066 2714
rect 4075 2684 4088 2714
rect 4103 2700 4133 2714
rect 4176 2700 4219 2714
rect 4226 2700 4446 2714
rect 4453 2700 4483 2714
rect 4143 2686 4158 2698
rect 4177 2686 4190 2700
rect 4258 2696 4411 2700
rect 4140 2684 4162 2686
rect 4240 2684 4432 2696
rect 4511 2684 4524 2714
rect 4539 2700 4569 2714
rect 4606 2684 4625 2714
rect 4640 2684 4646 2714
rect 4655 2684 4668 2714
rect 4683 2700 4713 2714
rect 4756 2700 4799 2714
rect 4806 2700 5026 2714
rect 5033 2700 5063 2714
rect 4723 2686 4738 2698
rect 4757 2686 4770 2700
rect 4838 2696 4991 2700
rect 4720 2684 4742 2686
rect 4820 2684 5012 2696
rect 5091 2684 5104 2714
rect 5119 2700 5149 2714
rect 5186 2684 5205 2714
rect 5220 2684 5226 2714
rect 5235 2684 5248 2714
rect 5263 2700 5293 2714
rect 5336 2700 5379 2714
rect 5386 2700 5606 2714
rect 5613 2700 5643 2714
rect 5303 2686 5318 2698
rect 5337 2686 5350 2700
rect 5418 2696 5571 2700
rect 5300 2684 5322 2686
rect 5400 2684 5592 2696
rect 5671 2684 5684 2714
rect 5699 2700 5729 2714
rect 5766 2684 5785 2714
rect 5800 2684 5806 2714
rect 5815 2684 5828 2714
rect 5843 2700 5873 2714
rect 5916 2700 5959 2714
rect 5966 2700 6186 2714
rect 6193 2700 6223 2714
rect 5883 2686 5898 2698
rect 5917 2686 5930 2700
rect 5998 2696 6151 2700
rect 5880 2684 5902 2686
rect 5980 2684 6172 2696
rect 6251 2684 6264 2714
rect 6279 2700 6309 2714
rect 6346 2684 6365 2714
rect 6380 2684 6386 2714
rect 6395 2684 6408 2714
rect 6423 2700 6453 2714
rect 6496 2700 6539 2714
rect 6546 2700 6766 2714
rect 6773 2700 6803 2714
rect 6463 2686 6478 2698
rect 6497 2686 6510 2700
rect 6578 2696 6731 2700
rect 6460 2684 6482 2686
rect 6560 2684 6752 2696
rect 6831 2684 6844 2714
rect 6859 2700 6889 2714
rect 6926 2684 6945 2714
rect 6960 2684 6966 2714
rect 6975 2684 6988 2714
rect 7003 2700 7033 2714
rect 7076 2700 7119 2714
rect 7126 2700 7346 2714
rect 7353 2700 7383 2714
rect 7043 2686 7058 2698
rect 7077 2686 7090 2700
rect 7158 2696 7311 2700
rect 7040 2684 7062 2686
rect 7140 2684 7332 2696
rect 7411 2684 7424 2714
rect 7439 2700 7469 2714
rect 7506 2684 7525 2714
rect 7540 2684 7546 2714
rect 7555 2684 7568 2714
rect 7583 2700 7613 2714
rect 7656 2700 7699 2714
rect 7706 2700 7926 2714
rect 7933 2700 7963 2714
rect 7623 2686 7638 2698
rect 7657 2686 7670 2700
rect 7738 2696 7891 2700
rect 7620 2684 7642 2686
rect 7720 2684 7912 2696
rect 7991 2684 8004 2714
rect 8019 2700 8049 2714
rect 8086 2684 8105 2714
rect 8120 2684 8126 2714
rect 8135 2684 8148 2714
rect 8163 2700 8193 2714
rect 8236 2700 8279 2714
rect 8286 2700 8506 2714
rect 8513 2700 8543 2714
rect 8203 2686 8218 2698
rect 8237 2686 8250 2700
rect 8318 2696 8471 2700
rect 8200 2684 8222 2686
rect 8300 2684 8492 2696
rect 8571 2684 8584 2714
rect 8599 2700 8629 2714
rect 8666 2684 8685 2714
rect 8700 2684 8706 2714
rect 8715 2684 8728 2714
rect 8743 2700 8773 2714
rect 8816 2700 8859 2714
rect 8866 2700 9086 2714
rect 9093 2700 9123 2714
rect 8783 2686 8798 2698
rect 8817 2686 8830 2700
rect 8898 2696 9051 2700
rect 8780 2684 8802 2686
rect 8880 2684 9072 2696
rect 9151 2684 9164 2714
rect 9179 2700 9209 2714
rect 9246 2684 9265 2714
rect 9280 2684 9286 2714
rect 9295 2684 9308 2714
rect 9323 2700 9353 2714
rect 9396 2700 9439 2714
rect 9446 2700 9666 2714
rect 9673 2700 9703 2714
rect 9363 2686 9378 2698
rect 9397 2686 9410 2700
rect 9478 2696 9631 2700
rect 9360 2684 9382 2686
rect 9460 2684 9652 2696
rect 9731 2684 9744 2714
rect 9759 2700 9789 2714
rect 9826 2684 9845 2714
rect 9860 2684 9866 2714
rect 9875 2684 9888 2714
rect 9903 2700 9933 2714
rect 9976 2700 10019 2714
rect 10026 2700 10246 2714
rect 10253 2700 10283 2714
rect 9943 2686 9958 2698
rect 9977 2686 9990 2700
rect 10058 2696 10211 2700
rect 9940 2684 9962 2686
rect 10040 2684 10232 2696
rect 10311 2684 10324 2714
rect 10339 2700 10369 2714
rect 10406 2684 10425 2714
rect 10440 2684 10446 2714
rect 10455 2684 10468 2714
rect 10483 2700 10513 2714
rect 10556 2700 10599 2714
rect 10606 2700 10826 2714
rect 10833 2700 10863 2714
rect 10523 2686 10538 2698
rect 10557 2686 10570 2700
rect 10638 2696 10791 2700
rect 10520 2684 10542 2686
rect 10620 2684 10812 2696
rect 10891 2684 10904 2714
rect 10919 2700 10949 2714
rect 10986 2684 11005 2714
rect 11020 2684 11026 2714
rect 11035 2684 11048 2714
rect 11063 2700 11093 2714
rect 11136 2700 11179 2714
rect 11186 2700 11406 2714
rect 11413 2700 11443 2714
rect 11103 2686 11118 2698
rect 11137 2686 11150 2700
rect 11218 2696 11371 2700
rect 11100 2684 11122 2686
rect 11200 2684 11392 2696
rect 11471 2684 11484 2714
rect 11499 2700 11529 2714
rect 11566 2684 11585 2714
rect 11600 2684 11606 2714
rect 11615 2684 11628 2714
rect 11643 2700 11673 2714
rect 11716 2700 11759 2714
rect 11766 2700 11986 2714
rect 11993 2700 12023 2714
rect 11683 2686 11698 2698
rect 11717 2686 11730 2700
rect 11798 2696 11951 2700
rect 11680 2684 11702 2686
rect 11780 2684 11972 2696
rect 12051 2684 12064 2714
rect 12079 2700 12109 2714
rect 12146 2684 12165 2714
rect 12180 2684 12186 2714
rect 12195 2684 12208 2714
rect 12223 2700 12253 2714
rect 12296 2700 12339 2714
rect 12346 2700 12566 2714
rect 12573 2700 12603 2714
rect 12263 2686 12278 2698
rect 12297 2686 12310 2700
rect 12378 2696 12531 2700
rect 12260 2684 12282 2686
rect 12360 2684 12552 2696
rect 12631 2684 12644 2714
rect 12659 2700 12689 2714
rect 12726 2684 12745 2714
rect 12760 2684 12766 2714
rect 12775 2684 12788 2714
rect 12803 2700 12833 2714
rect 12876 2700 12919 2714
rect 12926 2700 13146 2714
rect 13153 2700 13183 2714
rect 12843 2686 12858 2698
rect 12877 2686 12890 2700
rect 12958 2696 13111 2700
rect 12840 2684 12862 2686
rect 12940 2684 13132 2696
rect 13211 2684 13224 2714
rect 13239 2700 13269 2714
rect 13306 2684 13325 2714
rect 13340 2684 13346 2714
rect 13355 2684 13368 2714
rect 13383 2700 13413 2714
rect 13456 2700 13499 2714
rect 13506 2700 13726 2714
rect 13733 2700 13763 2714
rect 13423 2686 13438 2698
rect 13457 2686 13470 2700
rect 13538 2696 13691 2700
rect 13420 2684 13442 2686
rect 13520 2684 13712 2696
rect 13791 2684 13804 2714
rect 13819 2700 13849 2714
rect 13886 2684 13905 2714
rect 13920 2684 13926 2714
rect 13935 2684 13948 2714
rect 13963 2700 13993 2714
rect 14036 2700 14079 2714
rect 14086 2700 14306 2714
rect 14313 2700 14343 2714
rect 14003 2686 14018 2698
rect 14037 2686 14050 2700
rect 14118 2696 14271 2700
rect 14000 2684 14022 2686
rect 14100 2684 14292 2696
rect 14371 2684 14384 2714
rect 14399 2700 14429 2714
rect 14466 2684 14485 2714
rect 14500 2684 14506 2714
rect 14515 2684 14528 2714
rect 14543 2700 14573 2714
rect 14616 2700 14659 2714
rect 14666 2700 14886 2714
rect 14893 2700 14923 2714
rect 14583 2686 14598 2698
rect 14617 2686 14630 2700
rect 14698 2696 14851 2700
rect 14580 2684 14602 2686
rect 14680 2684 14872 2696
rect 14951 2684 14964 2714
rect 14979 2700 15009 2714
rect 15046 2684 15065 2714
rect 15080 2684 15086 2714
rect 15095 2684 15108 2714
rect 15123 2700 15153 2714
rect 15196 2700 15239 2714
rect 15246 2700 15466 2714
rect 15473 2700 15503 2714
rect 15163 2686 15178 2698
rect 15197 2686 15210 2700
rect 15278 2696 15431 2700
rect 15160 2684 15182 2686
rect 15260 2684 15452 2696
rect 15531 2684 15544 2714
rect 15559 2700 15589 2714
rect 15626 2684 15645 2714
rect 15660 2684 15666 2714
rect 15675 2684 15688 2714
rect 15703 2700 15733 2714
rect 15776 2700 15819 2714
rect 15826 2700 16046 2714
rect 16053 2700 16083 2714
rect 15743 2686 15758 2698
rect 15777 2686 15790 2700
rect 15858 2696 16011 2700
rect 15740 2684 15762 2686
rect 15840 2684 16032 2696
rect 16111 2684 16124 2714
rect 16139 2700 16169 2714
rect 16206 2684 16225 2714
rect 16240 2684 16246 2714
rect 16255 2684 16268 2714
rect 16283 2700 16313 2714
rect 16356 2700 16399 2714
rect 16406 2700 16626 2714
rect 16633 2700 16663 2714
rect 16323 2686 16338 2698
rect 16357 2686 16370 2700
rect 16438 2696 16591 2700
rect 16320 2684 16342 2686
rect 16420 2684 16612 2696
rect 16691 2684 16704 2714
rect 16719 2700 16749 2714
rect 16786 2684 16805 2714
rect 16820 2684 16826 2714
rect 16835 2684 16848 2714
rect 16863 2700 16893 2714
rect 16936 2700 16979 2714
rect 16986 2700 17206 2714
rect 17213 2700 17243 2714
rect 16903 2686 16918 2698
rect 16937 2686 16950 2700
rect 17018 2696 17171 2700
rect 16900 2684 16922 2686
rect 17000 2684 17192 2696
rect 17271 2684 17284 2714
rect 17299 2700 17329 2714
rect 17366 2684 17385 2714
rect 17400 2684 17406 2714
rect 17415 2684 17428 2714
rect 17443 2700 17473 2714
rect 17516 2700 17559 2714
rect 17566 2700 17786 2714
rect 17793 2700 17823 2714
rect 17483 2686 17498 2698
rect 17517 2686 17530 2700
rect 17598 2696 17751 2700
rect 17480 2684 17502 2686
rect 17580 2684 17772 2696
rect 17851 2684 17864 2714
rect 17879 2700 17909 2714
rect 17946 2684 17965 2714
rect 17980 2684 17986 2714
rect 17995 2684 18008 2714
rect 18023 2700 18053 2714
rect 18096 2700 18139 2714
rect 18146 2700 18366 2714
rect 18373 2700 18403 2714
rect 18063 2686 18078 2698
rect 18097 2686 18110 2700
rect 18178 2696 18331 2700
rect 18060 2684 18082 2686
rect 18160 2684 18352 2696
rect 18431 2684 18444 2714
rect 18459 2700 18489 2714
rect 18532 2684 18545 2714
rect 0 2670 18545 2684
rect 15 2600 28 2670
rect 80 2666 102 2670
rect 73 2644 102 2658
rect 155 2644 171 2658
rect 209 2654 215 2656
rect 222 2654 330 2670
rect 337 2654 343 2656
rect 351 2654 366 2670
rect 432 2664 451 2667
rect 73 2642 171 2644
rect 198 2642 366 2654
rect 381 2644 397 2658
rect 432 2645 454 2664
rect 464 2658 480 2659
rect 463 2656 480 2658
rect 464 2651 480 2656
rect 454 2644 460 2645
rect 463 2644 492 2651
rect 381 2643 492 2644
rect 381 2642 498 2643
rect 57 2634 108 2642
rect 155 2634 189 2642
rect 57 2622 82 2634
rect 89 2622 108 2634
rect 162 2632 189 2634
rect 198 2632 419 2642
rect 454 2639 460 2642
rect 162 2628 419 2632
rect 57 2614 108 2622
rect 155 2614 419 2628
rect 463 2634 498 2642
rect 9 2566 28 2600
rect 73 2606 102 2614
rect 73 2600 90 2606
rect 73 2598 107 2600
rect 155 2598 171 2614
rect 172 2604 380 2614
rect 381 2604 397 2614
rect 445 2610 460 2625
rect 463 2622 464 2634
rect 471 2622 498 2634
rect 463 2614 498 2622
rect 463 2613 492 2614
rect 183 2600 397 2604
rect 198 2598 397 2600
rect 432 2600 445 2610
rect 463 2600 480 2613
rect 432 2598 480 2600
rect 74 2594 107 2598
rect 70 2592 107 2594
rect 70 2591 137 2592
rect 70 2586 101 2591
rect 107 2586 137 2591
rect 70 2582 137 2586
rect 43 2579 137 2582
rect 43 2572 92 2579
rect 43 2566 73 2572
rect 92 2567 97 2572
rect 9 2550 89 2566
rect 101 2558 137 2579
rect 198 2574 387 2598
rect 432 2597 479 2598
rect 445 2592 479 2597
rect 213 2571 387 2574
rect 206 2568 387 2571
rect 415 2591 479 2592
rect 9 2548 28 2550
rect 43 2548 77 2550
rect 9 2532 89 2548
rect 9 2526 28 2532
rect -1 2510 28 2526
rect 43 2516 73 2532
rect 101 2510 107 2558
rect 110 2552 129 2558
rect 144 2552 174 2560
rect 110 2544 174 2552
rect 110 2528 190 2544
rect 206 2537 268 2568
rect 284 2537 346 2568
rect 415 2566 464 2591
rect 479 2566 509 2582
rect 378 2552 408 2560
rect 415 2558 525 2566
rect 378 2544 423 2552
rect 110 2526 129 2528
rect 144 2526 190 2528
rect 110 2510 190 2526
rect 217 2524 252 2537
rect 293 2534 330 2537
rect 293 2532 335 2534
rect 222 2521 252 2524
rect 231 2517 238 2521
rect 238 2516 239 2517
rect 197 2510 207 2516
rect -7 2502 34 2510
rect -7 2476 8 2502
rect 15 2476 34 2502
rect 98 2498 129 2510
rect 144 2498 247 2510
rect 259 2500 285 2526
rect 300 2521 330 2532
rect 362 2528 424 2544
rect 362 2526 408 2528
rect 362 2510 424 2526
rect 436 2510 442 2558
rect 445 2550 525 2558
rect 445 2548 464 2550
rect 479 2548 513 2550
rect 445 2532 525 2548
rect 445 2510 464 2532
rect 479 2516 509 2532
rect 537 2526 543 2600
rect 546 2526 565 2670
rect 580 2526 586 2670
rect 595 2600 608 2670
rect 660 2666 682 2670
rect 653 2644 682 2658
rect 735 2644 751 2658
rect 789 2654 795 2656
rect 802 2654 910 2670
rect 917 2654 923 2656
rect 931 2654 946 2670
rect 1012 2664 1031 2667
rect 653 2642 751 2644
rect 778 2642 946 2654
rect 961 2644 977 2658
rect 1012 2645 1034 2664
rect 1044 2658 1060 2659
rect 1043 2656 1060 2658
rect 1044 2651 1060 2656
rect 1034 2644 1040 2645
rect 1043 2644 1072 2651
rect 961 2643 1072 2644
rect 961 2642 1078 2643
rect 637 2634 688 2642
rect 735 2634 769 2642
rect 637 2622 662 2634
rect 669 2622 688 2634
rect 742 2632 769 2634
rect 778 2632 999 2642
rect 1034 2639 1040 2642
rect 742 2628 999 2632
rect 637 2614 688 2622
rect 735 2614 999 2628
rect 1043 2634 1078 2642
rect 589 2566 608 2600
rect 653 2606 682 2614
rect 653 2600 670 2606
rect 653 2598 687 2600
rect 735 2598 751 2614
rect 752 2604 960 2614
rect 961 2604 977 2614
rect 1025 2610 1040 2625
rect 1043 2622 1044 2634
rect 1051 2622 1078 2634
rect 1043 2614 1078 2622
rect 1043 2613 1072 2614
rect 763 2600 977 2604
rect 778 2598 977 2600
rect 1012 2600 1025 2610
rect 1043 2600 1060 2613
rect 1012 2598 1060 2600
rect 654 2594 687 2598
rect 650 2592 687 2594
rect 650 2591 717 2592
rect 650 2586 681 2591
rect 687 2586 717 2591
rect 650 2582 717 2586
rect 623 2579 717 2582
rect 623 2572 672 2579
rect 623 2566 653 2572
rect 672 2567 677 2572
rect 589 2550 669 2566
rect 681 2558 717 2579
rect 778 2574 967 2598
rect 1012 2597 1059 2598
rect 1025 2592 1059 2597
rect 793 2571 967 2574
rect 786 2568 967 2571
rect 995 2591 1059 2592
rect 589 2548 608 2550
rect 623 2548 657 2550
rect 589 2532 669 2548
rect 589 2526 608 2532
rect 305 2500 408 2510
rect 259 2498 408 2500
rect 429 2498 464 2510
rect 98 2496 260 2498
rect 110 2476 129 2496
rect 144 2494 174 2496
rect -7 2468 34 2476
rect 116 2472 129 2476
rect 181 2480 260 2496
rect 292 2496 464 2498
rect 292 2480 371 2496
rect 378 2494 408 2496
rect -1 2458 28 2468
rect 43 2458 73 2472
rect 116 2458 159 2472
rect 181 2468 371 2480
rect 436 2476 442 2496
rect 166 2458 196 2468
rect 197 2458 355 2468
rect 359 2458 389 2468
rect 393 2458 423 2472
rect 451 2458 464 2496
rect 536 2510 565 2526
rect 579 2510 608 2526
rect 623 2516 653 2532
rect 681 2510 687 2558
rect 690 2552 709 2558
rect 724 2552 754 2560
rect 690 2544 754 2552
rect 690 2528 770 2544
rect 786 2537 848 2568
rect 864 2537 926 2568
rect 995 2566 1044 2591
rect 1059 2566 1089 2582
rect 958 2552 988 2560
rect 995 2558 1105 2566
rect 958 2544 1003 2552
rect 690 2526 709 2528
rect 724 2526 770 2528
rect 690 2510 770 2526
rect 797 2524 832 2537
rect 873 2534 910 2537
rect 873 2532 915 2534
rect 802 2521 832 2524
rect 811 2517 818 2521
rect 818 2516 819 2517
rect 777 2510 787 2516
rect 536 2502 571 2510
rect 536 2476 537 2502
rect 544 2476 571 2502
rect 479 2458 509 2472
rect 536 2468 571 2476
rect 573 2502 614 2510
rect 573 2476 588 2502
rect 595 2476 614 2502
rect 678 2498 709 2510
rect 724 2498 827 2510
rect 839 2500 865 2526
rect 880 2521 910 2532
rect 942 2528 1004 2544
rect 942 2526 988 2528
rect 942 2510 1004 2526
rect 1016 2510 1022 2558
rect 1025 2550 1105 2558
rect 1025 2548 1044 2550
rect 1059 2548 1093 2550
rect 1025 2532 1105 2548
rect 1025 2510 1044 2532
rect 1059 2516 1089 2532
rect 1117 2526 1123 2600
rect 1126 2526 1145 2670
rect 1160 2526 1166 2670
rect 1175 2600 1188 2670
rect 1240 2666 1262 2670
rect 1233 2644 1262 2658
rect 1315 2644 1331 2658
rect 1369 2654 1375 2656
rect 1382 2654 1490 2670
rect 1497 2654 1503 2656
rect 1511 2654 1526 2670
rect 1592 2664 1611 2667
rect 1233 2642 1331 2644
rect 1358 2642 1526 2654
rect 1541 2644 1557 2658
rect 1592 2645 1614 2664
rect 1624 2658 1640 2659
rect 1623 2656 1640 2658
rect 1624 2651 1640 2656
rect 1614 2644 1620 2645
rect 1623 2644 1652 2651
rect 1541 2643 1652 2644
rect 1541 2642 1658 2643
rect 1217 2634 1268 2642
rect 1315 2634 1349 2642
rect 1217 2622 1242 2634
rect 1249 2622 1268 2634
rect 1322 2632 1349 2634
rect 1358 2632 1579 2642
rect 1614 2639 1620 2642
rect 1322 2628 1579 2632
rect 1217 2614 1268 2622
rect 1315 2614 1579 2628
rect 1623 2634 1658 2642
rect 1169 2566 1188 2600
rect 1233 2606 1262 2614
rect 1233 2600 1250 2606
rect 1233 2598 1267 2600
rect 1315 2598 1331 2614
rect 1332 2604 1540 2614
rect 1541 2604 1557 2614
rect 1605 2610 1620 2625
rect 1623 2622 1624 2634
rect 1631 2622 1658 2634
rect 1623 2614 1658 2622
rect 1623 2613 1652 2614
rect 1343 2600 1557 2604
rect 1358 2598 1557 2600
rect 1592 2600 1605 2610
rect 1623 2600 1640 2613
rect 1592 2598 1640 2600
rect 1234 2594 1267 2598
rect 1230 2592 1267 2594
rect 1230 2591 1297 2592
rect 1230 2586 1261 2591
rect 1267 2586 1297 2591
rect 1230 2582 1297 2586
rect 1203 2579 1297 2582
rect 1203 2572 1252 2579
rect 1203 2566 1233 2572
rect 1252 2567 1257 2572
rect 1169 2550 1249 2566
rect 1261 2558 1297 2579
rect 1358 2574 1547 2598
rect 1592 2597 1639 2598
rect 1605 2592 1639 2597
rect 1373 2571 1547 2574
rect 1366 2568 1547 2571
rect 1575 2591 1639 2592
rect 1169 2548 1188 2550
rect 1203 2548 1237 2550
rect 1169 2532 1249 2548
rect 1169 2526 1188 2532
rect 885 2500 988 2510
rect 839 2498 988 2500
rect 1009 2498 1044 2510
rect 678 2496 840 2498
rect 690 2476 709 2496
rect 724 2494 754 2496
rect 573 2468 614 2476
rect 696 2472 709 2476
rect 761 2480 840 2496
rect 872 2496 1044 2498
rect 872 2480 951 2496
rect 958 2494 988 2496
rect 536 2458 565 2468
rect 579 2458 608 2468
rect 623 2458 653 2472
rect 696 2458 739 2472
rect 761 2468 951 2480
rect 1016 2476 1022 2496
rect 746 2458 776 2468
rect 777 2458 935 2468
rect 939 2458 969 2468
rect 973 2458 1003 2472
rect 1031 2458 1044 2496
rect 1116 2510 1145 2526
rect 1159 2510 1188 2526
rect 1203 2516 1233 2532
rect 1261 2510 1267 2558
rect 1270 2552 1289 2558
rect 1304 2552 1334 2560
rect 1270 2544 1334 2552
rect 1270 2528 1350 2544
rect 1366 2537 1428 2568
rect 1444 2537 1506 2568
rect 1575 2566 1624 2591
rect 1639 2566 1669 2582
rect 1538 2552 1568 2560
rect 1575 2558 1685 2566
rect 1538 2544 1583 2552
rect 1270 2526 1289 2528
rect 1304 2526 1350 2528
rect 1270 2510 1350 2526
rect 1377 2524 1412 2537
rect 1453 2534 1490 2537
rect 1453 2532 1495 2534
rect 1382 2521 1412 2524
rect 1391 2517 1398 2521
rect 1398 2516 1399 2517
rect 1357 2510 1367 2516
rect 1116 2502 1151 2510
rect 1116 2476 1117 2502
rect 1124 2476 1151 2502
rect 1059 2458 1089 2472
rect 1116 2468 1151 2476
rect 1153 2502 1194 2510
rect 1153 2476 1168 2502
rect 1175 2476 1194 2502
rect 1258 2498 1289 2510
rect 1304 2498 1407 2510
rect 1419 2500 1445 2526
rect 1460 2521 1490 2532
rect 1522 2528 1584 2544
rect 1522 2526 1568 2528
rect 1522 2510 1584 2526
rect 1596 2510 1602 2558
rect 1605 2550 1685 2558
rect 1605 2548 1624 2550
rect 1639 2548 1673 2550
rect 1605 2532 1685 2548
rect 1605 2510 1624 2532
rect 1639 2516 1669 2532
rect 1697 2526 1703 2600
rect 1706 2526 1725 2670
rect 1740 2526 1746 2670
rect 1755 2600 1768 2670
rect 1820 2666 1842 2670
rect 1813 2644 1842 2658
rect 1895 2644 1911 2658
rect 1949 2654 1955 2656
rect 1962 2654 2070 2670
rect 2077 2654 2083 2656
rect 2091 2654 2106 2670
rect 2172 2664 2191 2667
rect 1813 2642 1911 2644
rect 1938 2642 2106 2654
rect 2121 2644 2137 2658
rect 2172 2645 2194 2664
rect 2204 2658 2220 2659
rect 2203 2656 2220 2658
rect 2204 2651 2220 2656
rect 2194 2644 2200 2645
rect 2203 2644 2232 2651
rect 2121 2643 2232 2644
rect 2121 2642 2238 2643
rect 1797 2634 1848 2642
rect 1895 2634 1929 2642
rect 1797 2622 1822 2634
rect 1829 2622 1848 2634
rect 1902 2632 1929 2634
rect 1938 2632 2159 2642
rect 2194 2639 2200 2642
rect 1902 2628 2159 2632
rect 1797 2614 1848 2622
rect 1895 2614 2159 2628
rect 2203 2634 2238 2642
rect 1749 2566 1768 2600
rect 1813 2606 1842 2614
rect 1813 2600 1830 2606
rect 1813 2598 1847 2600
rect 1895 2598 1911 2614
rect 1912 2604 2120 2614
rect 2121 2604 2137 2614
rect 2185 2610 2200 2625
rect 2203 2622 2204 2634
rect 2211 2622 2238 2634
rect 2203 2614 2238 2622
rect 2203 2613 2232 2614
rect 1923 2600 2137 2604
rect 1938 2598 2137 2600
rect 2172 2600 2185 2610
rect 2203 2600 2220 2613
rect 2172 2598 2220 2600
rect 1814 2594 1847 2598
rect 1810 2592 1847 2594
rect 1810 2591 1877 2592
rect 1810 2586 1841 2591
rect 1847 2586 1877 2591
rect 1810 2582 1877 2586
rect 1783 2579 1877 2582
rect 1783 2572 1832 2579
rect 1783 2566 1813 2572
rect 1832 2567 1837 2572
rect 1749 2550 1829 2566
rect 1841 2558 1877 2579
rect 1938 2574 2127 2598
rect 2172 2597 2219 2598
rect 2185 2592 2219 2597
rect 1953 2571 2127 2574
rect 1946 2568 2127 2571
rect 2155 2591 2219 2592
rect 1749 2548 1768 2550
rect 1783 2548 1817 2550
rect 1749 2532 1829 2548
rect 1749 2526 1768 2532
rect 1465 2500 1568 2510
rect 1419 2498 1568 2500
rect 1589 2498 1624 2510
rect 1258 2496 1420 2498
rect 1270 2476 1289 2496
rect 1304 2494 1334 2496
rect 1153 2468 1194 2476
rect 1276 2472 1289 2476
rect 1341 2480 1420 2496
rect 1452 2496 1624 2498
rect 1452 2480 1531 2496
rect 1538 2494 1568 2496
rect 1116 2458 1145 2468
rect 1159 2458 1188 2468
rect 1203 2458 1233 2472
rect 1276 2458 1319 2472
rect 1341 2468 1531 2480
rect 1596 2476 1602 2496
rect 1326 2458 1356 2468
rect 1357 2458 1515 2468
rect 1519 2458 1549 2468
rect 1553 2458 1583 2472
rect 1611 2458 1624 2496
rect 1696 2510 1725 2526
rect 1739 2510 1768 2526
rect 1783 2516 1813 2532
rect 1841 2510 1847 2558
rect 1850 2552 1869 2558
rect 1884 2552 1914 2560
rect 1850 2544 1914 2552
rect 1850 2528 1930 2544
rect 1946 2537 2008 2568
rect 2024 2537 2086 2568
rect 2155 2566 2204 2591
rect 2219 2566 2249 2582
rect 2118 2552 2148 2560
rect 2155 2558 2265 2566
rect 2118 2544 2163 2552
rect 1850 2526 1869 2528
rect 1884 2526 1930 2528
rect 1850 2510 1930 2526
rect 1957 2524 1992 2537
rect 2033 2534 2070 2537
rect 2033 2532 2075 2534
rect 1962 2521 1992 2524
rect 1971 2517 1978 2521
rect 1978 2516 1979 2517
rect 1937 2510 1947 2516
rect 1696 2502 1731 2510
rect 1696 2476 1697 2502
rect 1704 2476 1731 2502
rect 1639 2458 1669 2472
rect 1696 2468 1731 2476
rect 1733 2502 1774 2510
rect 1733 2476 1748 2502
rect 1755 2476 1774 2502
rect 1838 2498 1869 2510
rect 1884 2498 1987 2510
rect 1999 2500 2025 2526
rect 2040 2521 2070 2532
rect 2102 2528 2164 2544
rect 2102 2526 2148 2528
rect 2102 2510 2164 2526
rect 2176 2510 2182 2558
rect 2185 2550 2265 2558
rect 2185 2548 2204 2550
rect 2219 2548 2253 2550
rect 2185 2532 2265 2548
rect 2185 2510 2204 2532
rect 2219 2516 2249 2532
rect 2277 2526 2283 2600
rect 2286 2526 2305 2670
rect 2320 2526 2326 2670
rect 2335 2600 2348 2670
rect 2400 2666 2422 2670
rect 2393 2644 2422 2658
rect 2475 2644 2491 2658
rect 2529 2654 2535 2656
rect 2542 2654 2650 2670
rect 2657 2654 2663 2656
rect 2671 2654 2686 2670
rect 2752 2664 2771 2667
rect 2393 2642 2491 2644
rect 2518 2642 2686 2654
rect 2701 2644 2717 2658
rect 2752 2645 2774 2664
rect 2784 2658 2800 2659
rect 2783 2656 2800 2658
rect 2784 2651 2800 2656
rect 2774 2644 2780 2645
rect 2783 2644 2812 2651
rect 2701 2643 2812 2644
rect 2701 2642 2818 2643
rect 2377 2634 2428 2642
rect 2475 2634 2509 2642
rect 2377 2622 2402 2634
rect 2409 2622 2428 2634
rect 2482 2632 2509 2634
rect 2518 2632 2739 2642
rect 2774 2639 2780 2642
rect 2482 2628 2739 2632
rect 2377 2614 2428 2622
rect 2475 2614 2739 2628
rect 2783 2634 2818 2642
rect 2329 2566 2348 2600
rect 2393 2606 2422 2614
rect 2393 2600 2410 2606
rect 2393 2598 2427 2600
rect 2475 2598 2491 2614
rect 2492 2604 2700 2614
rect 2701 2604 2717 2614
rect 2765 2610 2780 2625
rect 2783 2622 2784 2634
rect 2791 2622 2818 2634
rect 2783 2614 2818 2622
rect 2783 2613 2812 2614
rect 2503 2600 2717 2604
rect 2518 2598 2717 2600
rect 2752 2600 2765 2610
rect 2783 2600 2800 2613
rect 2752 2598 2800 2600
rect 2394 2594 2427 2598
rect 2390 2592 2427 2594
rect 2390 2591 2457 2592
rect 2390 2586 2421 2591
rect 2427 2586 2457 2591
rect 2390 2582 2457 2586
rect 2363 2579 2457 2582
rect 2363 2572 2412 2579
rect 2363 2566 2393 2572
rect 2412 2567 2417 2572
rect 2329 2550 2409 2566
rect 2421 2558 2457 2579
rect 2518 2574 2707 2598
rect 2752 2597 2799 2598
rect 2765 2592 2799 2597
rect 2533 2571 2707 2574
rect 2526 2568 2707 2571
rect 2735 2591 2799 2592
rect 2329 2548 2348 2550
rect 2363 2548 2397 2550
rect 2329 2532 2409 2548
rect 2329 2526 2348 2532
rect 2045 2500 2148 2510
rect 1999 2498 2148 2500
rect 2169 2498 2204 2510
rect 1838 2496 2000 2498
rect 1850 2476 1869 2496
rect 1884 2494 1914 2496
rect 1733 2468 1774 2476
rect 1856 2472 1869 2476
rect 1921 2480 2000 2496
rect 2032 2496 2204 2498
rect 2032 2480 2111 2496
rect 2118 2494 2148 2496
rect 1696 2458 1725 2468
rect 1739 2458 1768 2468
rect 1783 2458 1813 2472
rect 1856 2458 1899 2472
rect 1921 2468 2111 2480
rect 2176 2476 2182 2496
rect 1906 2458 1936 2468
rect 1937 2458 2095 2468
rect 2099 2458 2129 2468
rect 2133 2458 2163 2472
rect 2191 2458 2204 2496
rect 2276 2510 2305 2526
rect 2319 2510 2348 2526
rect 2363 2516 2393 2532
rect 2421 2510 2427 2558
rect 2430 2552 2449 2558
rect 2464 2552 2494 2560
rect 2430 2544 2494 2552
rect 2430 2528 2510 2544
rect 2526 2537 2588 2568
rect 2604 2537 2666 2568
rect 2735 2566 2784 2591
rect 2799 2566 2829 2582
rect 2698 2552 2728 2560
rect 2735 2558 2845 2566
rect 2698 2544 2743 2552
rect 2430 2526 2449 2528
rect 2464 2526 2510 2528
rect 2430 2510 2510 2526
rect 2537 2524 2572 2537
rect 2613 2534 2650 2537
rect 2613 2532 2655 2534
rect 2542 2521 2572 2524
rect 2551 2517 2558 2521
rect 2558 2516 2559 2517
rect 2517 2510 2527 2516
rect 2276 2502 2311 2510
rect 2276 2476 2277 2502
rect 2284 2476 2311 2502
rect 2219 2458 2249 2472
rect 2276 2468 2311 2476
rect 2313 2502 2354 2510
rect 2313 2476 2328 2502
rect 2335 2476 2354 2502
rect 2418 2498 2449 2510
rect 2464 2498 2567 2510
rect 2579 2500 2605 2526
rect 2620 2521 2650 2532
rect 2682 2528 2744 2544
rect 2682 2526 2728 2528
rect 2682 2510 2744 2526
rect 2756 2510 2762 2558
rect 2765 2550 2845 2558
rect 2765 2548 2784 2550
rect 2799 2548 2833 2550
rect 2765 2532 2845 2548
rect 2765 2510 2784 2532
rect 2799 2516 2829 2532
rect 2857 2526 2863 2600
rect 2866 2526 2885 2670
rect 2900 2526 2906 2670
rect 2915 2600 2928 2670
rect 2980 2666 3002 2670
rect 2973 2644 3002 2658
rect 3055 2644 3071 2658
rect 3109 2654 3115 2656
rect 3122 2654 3230 2670
rect 3237 2654 3243 2656
rect 3251 2654 3266 2670
rect 3332 2664 3351 2667
rect 2973 2642 3071 2644
rect 3098 2642 3266 2654
rect 3281 2644 3297 2658
rect 3332 2645 3354 2664
rect 3364 2658 3380 2659
rect 3363 2656 3380 2658
rect 3364 2651 3380 2656
rect 3354 2644 3360 2645
rect 3363 2644 3392 2651
rect 3281 2643 3392 2644
rect 3281 2642 3398 2643
rect 2957 2634 3008 2642
rect 3055 2634 3089 2642
rect 2957 2622 2982 2634
rect 2989 2622 3008 2634
rect 3062 2632 3089 2634
rect 3098 2632 3319 2642
rect 3354 2639 3360 2642
rect 3062 2628 3319 2632
rect 2957 2614 3008 2622
rect 3055 2614 3319 2628
rect 3363 2634 3398 2642
rect 2909 2566 2928 2600
rect 2973 2606 3002 2614
rect 2973 2600 2990 2606
rect 2973 2598 3007 2600
rect 3055 2598 3071 2614
rect 3072 2604 3280 2614
rect 3281 2604 3297 2614
rect 3345 2610 3360 2625
rect 3363 2622 3364 2634
rect 3371 2622 3398 2634
rect 3363 2614 3398 2622
rect 3363 2613 3392 2614
rect 3083 2600 3297 2604
rect 3098 2598 3297 2600
rect 3332 2600 3345 2610
rect 3363 2600 3380 2613
rect 3332 2598 3380 2600
rect 2974 2594 3007 2598
rect 2970 2592 3007 2594
rect 2970 2591 3037 2592
rect 2970 2586 3001 2591
rect 3007 2586 3037 2591
rect 2970 2582 3037 2586
rect 2943 2579 3037 2582
rect 2943 2572 2992 2579
rect 2943 2566 2973 2572
rect 2992 2567 2997 2572
rect 2909 2550 2989 2566
rect 3001 2558 3037 2579
rect 3098 2574 3287 2598
rect 3332 2597 3379 2598
rect 3345 2592 3379 2597
rect 3113 2571 3287 2574
rect 3106 2568 3287 2571
rect 3315 2591 3379 2592
rect 2909 2548 2928 2550
rect 2943 2548 2977 2550
rect 2909 2532 2989 2548
rect 2909 2526 2928 2532
rect 2625 2500 2728 2510
rect 2579 2498 2728 2500
rect 2749 2498 2784 2510
rect 2418 2496 2580 2498
rect 2430 2476 2449 2496
rect 2464 2494 2494 2496
rect 2313 2468 2354 2476
rect 2436 2472 2449 2476
rect 2501 2480 2580 2496
rect 2612 2496 2784 2498
rect 2612 2480 2691 2496
rect 2698 2494 2728 2496
rect 2276 2458 2305 2468
rect 2319 2458 2348 2468
rect 2363 2458 2393 2472
rect 2436 2458 2479 2472
rect 2501 2468 2691 2480
rect 2756 2476 2762 2496
rect 2486 2458 2516 2468
rect 2517 2458 2675 2468
rect 2679 2458 2709 2468
rect 2713 2458 2743 2472
rect 2771 2458 2784 2496
rect 2856 2510 2885 2526
rect 2899 2510 2928 2526
rect 2943 2516 2973 2532
rect 3001 2510 3007 2558
rect 3010 2552 3029 2558
rect 3044 2552 3074 2560
rect 3010 2544 3074 2552
rect 3010 2528 3090 2544
rect 3106 2537 3168 2568
rect 3184 2537 3246 2568
rect 3315 2566 3364 2591
rect 3379 2566 3409 2582
rect 3278 2552 3308 2560
rect 3315 2558 3425 2566
rect 3278 2544 3323 2552
rect 3010 2526 3029 2528
rect 3044 2526 3090 2528
rect 3010 2510 3090 2526
rect 3117 2524 3152 2537
rect 3193 2534 3230 2537
rect 3193 2532 3235 2534
rect 3122 2521 3152 2524
rect 3131 2517 3138 2521
rect 3138 2516 3139 2517
rect 3097 2510 3107 2516
rect 2856 2502 2891 2510
rect 2856 2476 2857 2502
rect 2864 2476 2891 2502
rect 2799 2458 2829 2472
rect 2856 2468 2891 2476
rect 2893 2502 2934 2510
rect 2893 2476 2908 2502
rect 2915 2476 2934 2502
rect 2998 2498 3029 2510
rect 3044 2498 3147 2510
rect 3159 2500 3185 2526
rect 3200 2521 3230 2532
rect 3262 2528 3324 2544
rect 3262 2526 3308 2528
rect 3262 2510 3324 2526
rect 3336 2510 3342 2558
rect 3345 2550 3425 2558
rect 3345 2548 3364 2550
rect 3379 2548 3413 2550
rect 3345 2532 3425 2548
rect 3345 2510 3364 2532
rect 3379 2516 3409 2532
rect 3437 2526 3443 2600
rect 3446 2526 3465 2670
rect 3480 2526 3486 2670
rect 3495 2600 3508 2670
rect 3560 2666 3582 2670
rect 3553 2644 3582 2658
rect 3635 2644 3651 2658
rect 3689 2654 3695 2656
rect 3702 2654 3810 2670
rect 3817 2654 3823 2656
rect 3831 2654 3846 2670
rect 3912 2664 3931 2667
rect 3553 2642 3651 2644
rect 3678 2642 3846 2654
rect 3861 2644 3877 2658
rect 3912 2645 3934 2664
rect 3944 2658 3960 2659
rect 3943 2656 3960 2658
rect 3944 2651 3960 2656
rect 3934 2644 3940 2645
rect 3943 2644 3972 2651
rect 3861 2643 3972 2644
rect 3861 2642 3978 2643
rect 3537 2634 3588 2642
rect 3635 2634 3669 2642
rect 3537 2622 3562 2634
rect 3569 2622 3588 2634
rect 3642 2632 3669 2634
rect 3678 2632 3899 2642
rect 3934 2639 3940 2642
rect 3642 2628 3899 2632
rect 3537 2614 3588 2622
rect 3635 2614 3899 2628
rect 3943 2634 3978 2642
rect 3489 2566 3508 2600
rect 3553 2606 3582 2614
rect 3553 2600 3570 2606
rect 3553 2598 3587 2600
rect 3635 2598 3651 2614
rect 3652 2604 3860 2614
rect 3861 2604 3877 2614
rect 3925 2610 3940 2625
rect 3943 2622 3944 2634
rect 3951 2622 3978 2634
rect 3943 2614 3978 2622
rect 3943 2613 3972 2614
rect 3663 2600 3877 2604
rect 3678 2598 3877 2600
rect 3912 2600 3925 2610
rect 3943 2600 3960 2613
rect 3912 2598 3960 2600
rect 3554 2594 3587 2598
rect 3550 2592 3587 2594
rect 3550 2591 3617 2592
rect 3550 2586 3581 2591
rect 3587 2586 3617 2591
rect 3550 2582 3617 2586
rect 3523 2579 3617 2582
rect 3523 2572 3572 2579
rect 3523 2566 3553 2572
rect 3572 2567 3577 2572
rect 3489 2550 3569 2566
rect 3581 2558 3617 2579
rect 3678 2574 3867 2598
rect 3912 2597 3959 2598
rect 3925 2592 3959 2597
rect 3693 2571 3867 2574
rect 3686 2568 3867 2571
rect 3895 2591 3959 2592
rect 3489 2548 3508 2550
rect 3523 2548 3557 2550
rect 3489 2532 3569 2548
rect 3489 2526 3508 2532
rect 3205 2500 3308 2510
rect 3159 2498 3308 2500
rect 3329 2498 3364 2510
rect 2998 2496 3160 2498
rect 3010 2476 3029 2496
rect 3044 2494 3074 2496
rect 2893 2468 2934 2476
rect 3016 2472 3029 2476
rect 3081 2480 3160 2496
rect 3192 2496 3364 2498
rect 3192 2480 3271 2496
rect 3278 2494 3308 2496
rect 2856 2458 2885 2468
rect 2899 2458 2928 2468
rect 2943 2458 2973 2472
rect 3016 2458 3059 2472
rect 3081 2468 3271 2480
rect 3336 2476 3342 2496
rect 3066 2458 3096 2468
rect 3097 2458 3255 2468
rect 3259 2458 3289 2468
rect 3293 2458 3323 2472
rect 3351 2458 3364 2496
rect 3436 2510 3465 2526
rect 3479 2510 3508 2526
rect 3523 2516 3553 2532
rect 3581 2510 3587 2558
rect 3590 2552 3609 2558
rect 3624 2552 3654 2560
rect 3590 2544 3654 2552
rect 3590 2528 3670 2544
rect 3686 2537 3748 2568
rect 3764 2537 3826 2568
rect 3895 2566 3944 2591
rect 3959 2566 3989 2582
rect 3858 2552 3888 2560
rect 3895 2558 4005 2566
rect 3858 2544 3903 2552
rect 3590 2526 3609 2528
rect 3624 2526 3670 2528
rect 3590 2510 3670 2526
rect 3697 2524 3732 2537
rect 3773 2534 3810 2537
rect 3773 2532 3815 2534
rect 3702 2521 3732 2524
rect 3711 2517 3718 2521
rect 3718 2516 3719 2517
rect 3677 2510 3687 2516
rect 3436 2502 3471 2510
rect 3436 2476 3437 2502
rect 3444 2476 3471 2502
rect 3379 2458 3409 2472
rect 3436 2468 3471 2476
rect 3473 2502 3514 2510
rect 3473 2476 3488 2502
rect 3495 2476 3514 2502
rect 3578 2498 3609 2510
rect 3624 2498 3727 2510
rect 3739 2500 3765 2526
rect 3780 2521 3810 2532
rect 3842 2528 3904 2544
rect 3842 2526 3888 2528
rect 3842 2510 3904 2526
rect 3916 2510 3922 2558
rect 3925 2550 4005 2558
rect 3925 2548 3944 2550
rect 3959 2548 3993 2550
rect 3925 2532 4005 2548
rect 3925 2510 3944 2532
rect 3959 2516 3989 2532
rect 4017 2526 4023 2600
rect 4026 2526 4045 2670
rect 4060 2526 4066 2670
rect 4075 2600 4088 2670
rect 4140 2666 4162 2670
rect 4133 2644 4162 2658
rect 4215 2644 4231 2658
rect 4269 2654 4275 2656
rect 4282 2654 4390 2670
rect 4397 2654 4403 2656
rect 4411 2654 4426 2670
rect 4492 2664 4511 2667
rect 4133 2642 4231 2644
rect 4258 2642 4426 2654
rect 4441 2644 4457 2658
rect 4492 2645 4514 2664
rect 4524 2658 4540 2659
rect 4523 2656 4540 2658
rect 4524 2651 4540 2656
rect 4514 2644 4520 2645
rect 4523 2644 4552 2651
rect 4441 2643 4552 2644
rect 4441 2642 4558 2643
rect 4117 2634 4168 2642
rect 4215 2634 4249 2642
rect 4117 2622 4142 2634
rect 4149 2622 4168 2634
rect 4222 2632 4249 2634
rect 4258 2632 4479 2642
rect 4514 2639 4520 2642
rect 4222 2628 4479 2632
rect 4117 2614 4168 2622
rect 4215 2614 4479 2628
rect 4523 2634 4558 2642
rect 4069 2566 4088 2600
rect 4133 2606 4162 2614
rect 4133 2600 4150 2606
rect 4133 2598 4167 2600
rect 4215 2598 4231 2614
rect 4232 2604 4440 2614
rect 4441 2604 4457 2614
rect 4505 2610 4520 2625
rect 4523 2622 4524 2634
rect 4531 2622 4558 2634
rect 4523 2614 4558 2622
rect 4523 2613 4552 2614
rect 4243 2600 4457 2604
rect 4258 2598 4457 2600
rect 4492 2600 4505 2610
rect 4523 2600 4540 2613
rect 4492 2598 4540 2600
rect 4134 2594 4167 2598
rect 4130 2592 4167 2594
rect 4130 2591 4197 2592
rect 4130 2586 4161 2591
rect 4167 2586 4197 2591
rect 4130 2582 4197 2586
rect 4103 2579 4197 2582
rect 4103 2572 4152 2579
rect 4103 2566 4133 2572
rect 4152 2567 4157 2572
rect 4069 2550 4149 2566
rect 4161 2558 4197 2579
rect 4258 2574 4447 2598
rect 4492 2597 4539 2598
rect 4505 2592 4539 2597
rect 4273 2571 4447 2574
rect 4266 2568 4447 2571
rect 4475 2591 4539 2592
rect 4069 2548 4088 2550
rect 4103 2548 4137 2550
rect 4069 2532 4149 2548
rect 4069 2526 4088 2532
rect 3785 2500 3888 2510
rect 3739 2498 3888 2500
rect 3909 2498 3944 2510
rect 3578 2496 3740 2498
rect 3590 2476 3609 2496
rect 3624 2494 3654 2496
rect 3473 2468 3514 2476
rect 3596 2472 3609 2476
rect 3661 2480 3740 2496
rect 3772 2496 3944 2498
rect 3772 2480 3851 2496
rect 3858 2494 3888 2496
rect 3436 2458 3465 2468
rect 3479 2458 3508 2468
rect 3523 2458 3553 2472
rect 3596 2458 3639 2472
rect 3661 2468 3851 2480
rect 3916 2476 3922 2496
rect 3646 2458 3676 2468
rect 3677 2458 3835 2468
rect 3839 2458 3869 2468
rect 3873 2458 3903 2472
rect 3931 2458 3944 2496
rect 4016 2510 4045 2526
rect 4059 2510 4088 2526
rect 4103 2516 4133 2532
rect 4161 2510 4167 2558
rect 4170 2552 4189 2558
rect 4204 2552 4234 2560
rect 4170 2544 4234 2552
rect 4170 2528 4250 2544
rect 4266 2537 4328 2568
rect 4344 2537 4406 2568
rect 4475 2566 4524 2591
rect 4539 2566 4569 2582
rect 4438 2552 4468 2560
rect 4475 2558 4585 2566
rect 4438 2544 4483 2552
rect 4170 2526 4189 2528
rect 4204 2526 4250 2528
rect 4170 2510 4250 2526
rect 4277 2524 4312 2537
rect 4353 2534 4390 2537
rect 4353 2532 4395 2534
rect 4282 2521 4312 2524
rect 4291 2517 4298 2521
rect 4298 2516 4299 2517
rect 4257 2510 4267 2516
rect 4016 2502 4051 2510
rect 4016 2476 4017 2502
rect 4024 2476 4051 2502
rect 3959 2458 3989 2472
rect 4016 2468 4051 2476
rect 4053 2502 4094 2510
rect 4053 2476 4068 2502
rect 4075 2476 4094 2502
rect 4158 2498 4189 2510
rect 4204 2498 4307 2510
rect 4319 2500 4345 2526
rect 4360 2521 4390 2532
rect 4422 2528 4484 2544
rect 4422 2526 4468 2528
rect 4422 2510 4484 2526
rect 4496 2510 4502 2558
rect 4505 2550 4585 2558
rect 4505 2548 4524 2550
rect 4539 2548 4573 2550
rect 4505 2532 4585 2548
rect 4505 2510 4524 2532
rect 4539 2516 4569 2532
rect 4597 2526 4603 2600
rect 4606 2526 4625 2670
rect 4640 2526 4646 2670
rect 4655 2600 4668 2670
rect 4720 2666 4742 2670
rect 4713 2644 4742 2658
rect 4795 2644 4811 2658
rect 4849 2654 4855 2656
rect 4862 2654 4970 2670
rect 4977 2654 4983 2656
rect 4991 2654 5006 2670
rect 5072 2664 5091 2667
rect 4713 2642 4811 2644
rect 4838 2642 5006 2654
rect 5021 2644 5037 2658
rect 5072 2645 5094 2664
rect 5104 2658 5120 2659
rect 5103 2656 5120 2658
rect 5104 2651 5120 2656
rect 5094 2644 5100 2645
rect 5103 2644 5132 2651
rect 5021 2643 5132 2644
rect 5021 2642 5138 2643
rect 4697 2634 4748 2642
rect 4795 2634 4829 2642
rect 4697 2622 4722 2634
rect 4729 2622 4748 2634
rect 4802 2632 4829 2634
rect 4838 2632 5059 2642
rect 5094 2639 5100 2642
rect 4802 2628 5059 2632
rect 4697 2614 4748 2622
rect 4795 2614 5059 2628
rect 5103 2634 5138 2642
rect 4649 2566 4668 2600
rect 4713 2606 4742 2614
rect 4713 2600 4730 2606
rect 4713 2598 4747 2600
rect 4795 2598 4811 2614
rect 4812 2604 5020 2614
rect 5021 2604 5037 2614
rect 5085 2610 5100 2625
rect 5103 2622 5104 2634
rect 5111 2622 5138 2634
rect 5103 2614 5138 2622
rect 5103 2613 5132 2614
rect 4823 2600 5037 2604
rect 4838 2598 5037 2600
rect 5072 2600 5085 2610
rect 5103 2600 5120 2613
rect 5072 2598 5120 2600
rect 4714 2594 4747 2598
rect 4710 2592 4747 2594
rect 4710 2591 4777 2592
rect 4710 2586 4741 2591
rect 4747 2586 4777 2591
rect 4710 2582 4777 2586
rect 4683 2579 4777 2582
rect 4683 2572 4732 2579
rect 4683 2566 4713 2572
rect 4732 2567 4737 2572
rect 4649 2550 4729 2566
rect 4741 2558 4777 2579
rect 4838 2574 5027 2598
rect 5072 2597 5119 2598
rect 5085 2592 5119 2597
rect 4853 2571 5027 2574
rect 4846 2568 5027 2571
rect 5055 2591 5119 2592
rect 4649 2548 4668 2550
rect 4683 2548 4717 2550
rect 4649 2532 4729 2548
rect 4649 2526 4668 2532
rect 4365 2500 4468 2510
rect 4319 2498 4468 2500
rect 4489 2498 4524 2510
rect 4158 2496 4320 2498
rect 4170 2476 4189 2496
rect 4204 2494 4234 2496
rect 4053 2468 4094 2476
rect 4176 2472 4189 2476
rect 4241 2480 4320 2496
rect 4352 2496 4524 2498
rect 4352 2480 4431 2496
rect 4438 2494 4468 2496
rect 4016 2458 4045 2468
rect 4059 2458 4088 2468
rect 4103 2458 4133 2472
rect 4176 2458 4219 2472
rect 4241 2468 4431 2480
rect 4496 2476 4502 2496
rect 4226 2458 4256 2468
rect 4257 2458 4415 2468
rect 4419 2458 4449 2468
rect 4453 2458 4483 2472
rect 4511 2458 4524 2496
rect 4596 2510 4625 2526
rect 4639 2510 4668 2526
rect 4683 2516 4713 2532
rect 4741 2510 4747 2558
rect 4750 2552 4769 2558
rect 4784 2552 4814 2560
rect 4750 2544 4814 2552
rect 4750 2528 4830 2544
rect 4846 2537 4908 2568
rect 4924 2537 4986 2568
rect 5055 2566 5104 2591
rect 5119 2566 5149 2582
rect 5018 2552 5048 2560
rect 5055 2558 5165 2566
rect 5018 2544 5063 2552
rect 4750 2526 4769 2528
rect 4784 2526 4830 2528
rect 4750 2510 4830 2526
rect 4857 2524 4892 2537
rect 4933 2534 4970 2537
rect 4933 2532 4975 2534
rect 4862 2521 4892 2524
rect 4871 2517 4878 2521
rect 4878 2516 4879 2517
rect 4837 2510 4847 2516
rect 4596 2502 4631 2510
rect 4596 2476 4597 2502
rect 4604 2476 4631 2502
rect 4539 2458 4569 2472
rect 4596 2468 4631 2476
rect 4633 2502 4674 2510
rect 4633 2476 4648 2502
rect 4655 2476 4674 2502
rect 4738 2498 4769 2510
rect 4784 2498 4887 2510
rect 4899 2500 4925 2526
rect 4940 2521 4970 2532
rect 5002 2528 5064 2544
rect 5002 2526 5048 2528
rect 5002 2510 5064 2526
rect 5076 2510 5082 2558
rect 5085 2550 5165 2558
rect 5085 2548 5104 2550
rect 5119 2548 5153 2550
rect 5085 2532 5165 2548
rect 5085 2510 5104 2532
rect 5119 2516 5149 2532
rect 5177 2526 5183 2600
rect 5186 2526 5205 2670
rect 5220 2526 5226 2670
rect 5235 2600 5248 2670
rect 5300 2666 5322 2670
rect 5293 2644 5322 2658
rect 5375 2644 5391 2658
rect 5429 2654 5435 2656
rect 5442 2654 5550 2670
rect 5557 2654 5563 2656
rect 5571 2654 5586 2670
rect 5652 2664 5671 2667
rect 5293 2642 5391 2644
rect 5418 2642 5586 2654
rect 5601 2644 5617 2658
rect 5652 2645 5674 2664
rect 5684 2658 5700 2659
rect 5683 2656 5700 2658
rect 5684 2651 5700 2656
rect 5674 2644 5680 2645
rect 5683 2644 5712 2651
rect 5601 2643 5712 2644
rect 5601 2642 5718 2643
rect 5277 2634 5328 2642
rect 5375 2634 5409 2642
rect 5277 2622 5302 2634
rect 5309 2622 5328 2634
rect 5382 2632 5409 2634
rect 5418 2632 5639 2642
rect 5674 2639 5680 2642
rect 5382 2628 5639 2632
rect 5277 2614 5328 2622
rect 5375 2614 5639 2628
rect 5683 2634 5718 2642
rect 5229 2566 5248 2600
rect 5293 2606 5322 2614
rect 5293 2600 5310 2606
rect 5293 2598 5327 2600
rect 5375 2598 5391 2614
rect 5392 2604 5600 2614
rect 5601 2604 5617 2614
rect 5665 2610 5680 2625
rect 5683 2622 5684 2634
rect 5691 2622 5718 2634
rect 5683 2614 5718 2622
rect 5683 2613 5712 2614
rect 5403 2600 5617 2604
rect 5418 2598 5617 2600
rect 5652 2600 5665 2610
rect 5683 2600 5700 2613
rect 5652 2598 5700 2600
rect 5294 2594 5327 2598
rect 5290 2592 5327 2594
rect 5290 2591 5357 2592
rect 5290 2586 5321 2591
rect 5327 2586 5357 2591
rect 5290 2582 5357 2586
rect 5263 2579 5357 2582
rect 5263 2572 5312 2579
rect 5263 2566 5293 2572
rect 5312 2567 5317 2572
rect 5229 2550 5309 2566
rect 5321 2558 5357 2579
rect 5418 2574 5607 2598
rect 5652 2597 5699 2598
rect 5665 2592 5699 2597
rect 5433 2571 5607 2574
rect 5426 2568 5607 2571
rect 5635 2591 5699 2592
rect 5229 2548 5248 2550
rect 5263 2548 5297 2550
rect 5229 2532 5309 2548
rect 5229 2526 5248 2532
rect 4945 2500 5048 2510
rect 4899 2498 5048 2500
rect 5069 2498 5104 2510
rect 4738 2496 4900 2498
rect 4750 2476 4769 2496
rect 4784 2494 4814 2496
rect 4633 2468 4674 2476
rect 4756 2472 4769 2476
rect 4821 2480 4900 2496
rect 4932 2496 5104 2498
rect 4932 2480 5011 2496
rect 5018 2494 5048 2496
rect 4596 2458 4625 2468
rect 4639 2458 4668 2468
rect 4683 2458 4713 2472
rect 4756 2458 4799 2472
rect 4821 2468 5011 2480
rect 5076 2476 5082 2496
rect 4806 2458 4836 2468
rect 4837 2458 4995 2468
rect 4999 2458 5029 2468
rect 5033 2458 5063 2472
rect 5091 2458 5104 2496
rect 5176 2510 5205 2526
rect 5219 2510 5248 2526
rect 5263 2516 5293 2532
rect 5321 2510 5327 2558
rect 5330 2552 5349 2558
rect 5364 2552 5394 2560
rect 5330 2544 5394 2552
rect 5330 2528 5410 2544
rect 5426 2537 5488 2568
rect 5504 2537 5566 2568
rect 5635 2566 5684 2591
rect 5699 2566 5729 2582
rect 5598 2552 5628 2560
rect 5635 2558 5745 2566
rect 5598 2544 5643 2552
rect 5330 2526 5349 2528
rect 5364 2526 5410 2528
rect 5330 2510 5410 2526
rect 5437 2524 5472 2537
rect 5513 2534 5550 2537
rect 5513 2532 5555 2534
rect 5442 2521 5472 2524
rect 5451 2517 5458 2521
rect 5458 2516 5459 2517
rect 5417 2510 5427 2516
rect 5176 2502 5211 2510
rect 5176 2476 5177 2502
rect 5184 2476 5211 2502
rect 5119 2458 5149 2472
rect 5176 2468 5211 2476
rect 5213 2502 5254 2510
rect 5213 2476 5228 2502
rect 5235 2476 5254 2502
rect 5318 2498 5349 2510
rect 5364 2498 5467 2510
rect 5479 2500 5505 2526
rect 5520 2521 5550 2532
rect 5582 2528 5644 2544
rect 5582 2526 5628 2528
rect 5582 2510 5644 2526
rect 5656 2510 5662 2558
rect 5665 2550 5745 2558
rect 5665 2548 5684 2550
rect 5699 2548 5733 2550
rect 5665 2532 5745 2548
rect 5665 2510 5684 2532
rect 5699 2516 5729 2532
rect 5757 2526 5763 2600
rect 5766 2526 5785 2670
rect 5800 2526 5806 2670
rect 5815 2600 5828 2670
rect 5880 2666 5902 2670
rect 5873 2644 5902 2658
rect 5955 2644 5971 2658
rect 6009 2654 6015 2656
rect 6022 2654 6130 2670
rect 6137 2654 6143 2656
rect 6151 2654 6166 2670
rect 6232 2664 6251 2667
rect 5873 2642 5971 2644
rect 5998 2642 6166 2654
rect 6181 2644 6197 2658
rect 6232 2645 6254 2664
rect 6264 2658 6280 2659
rect 6263 2656 6280 2658
rect 6264 2651 6280 2656
rect 6254 2644 6260 2645
rect 6263 2644 6292 2651
rect 6181 2643 6292 2644
rect 6181 2642 6298 2643
rect 5857 2634 5908 2642
rect 5955 2634 5989 2642
rect 5857 2622 5882 2634
rect 5889 2622 5908 2634
rect 5962 2632 5989 2634
rect 5998 2632 6219 2642
rect 6254 2639 6260 2642
rect 5962 2628 6219 2632
rect 5857 2614 5908 2622
rect 5955 2614 6219 2628
rect 6263 2634 6298 2642
rect 5809 2566 5828 2600
rect 5873 2606 5902 2614
rect 5873 2600 5890 2606
rect 5873 2598 5907 2600
rect 5955 2598 5971 2614
rect 5972 2604 6180 2614
rect 6181 2604 6197 2614
rect 6245 2610 6260 2625
rect 6263 2622 6264 2634
rect 6271 2622 6298 2634
rect 6263 2614 6298 2622
rect 6263 2613 6292 2614
rect 5983 2600 6197 2604
rect 5998 2598 6197 2600
rect 6232 2600 6245 2610
rect 6263 2600 6280 2613
rect 6232 2598 6280 2600
rect 5874 2594 5907 2598
rect 5870 2592 5907 2594
rect 5870 2591 5937 2592
rect 5870 2586 5901 2591
rect 5907 2586 5937 2591
rect 5870 2582 5937 2586
rect 5843 2579 5937 2582
rect 5843 2572 5892 2579
rect 5843 2566 5873 2572
rect 5892 2567 5897 2572
rect 5809 2550 5889 2566
rect 5901 2558 5937 2579
rect 5998 2574 6187 2598
rect 6232 2597 6279 2598
rect 6245 2592 6279 2597
rect 6013 2571 6187 2574
rect 6006 2568 6187 2571
rect 6215 2591 6279 2592
rect 5809 2548 5828 2550
rect 5843 2548 5877 2550
rect 5809 2532 5889 2548
rect 5809 2526 5828 2532
rect 5525 2500 5628 2510
rect 5479 2498 5628 2500
rect 5649 2498 5684 2510
rect 5318 2496 5480 2498
rect 5330 2476 5349 2496
rect 5364 2494 5394 2496
rect 5213 2468 5254 2476
rect 5336 2472 5349 2476
rect 5401 2480 5480 2496
rect 5512 2496 5684 2498
rect 5512 2480 5591 2496
rect 5598 2494 5628 2496
rect 5176 2458 5205 2468
rect 5219 2458 5248 2468
rect 5263 2458 5293 2472
rect 5336 2458 5379 2472
rect 5401 2468 5591 2480
rect 5656 2476 5662 2496
rect 5386 2458 5416 2468
rect 5417 2458 5575 2468
rect 5579 2458 5609 2468
rect 5613 2458 5643 2472
rect 5671 2458 5684 2496
rect 5756 2510 5785 2526
rect 5799 2510 5828 2526
rect 5843 2516 5873 2532
rect 5901 2510 5907 2558
rect 5910 2552 5929 2558
rect 5944 2552 5974 2560
rect 5910 2544 5974 2552
rect 5910 2528 5990 2544
rect 6006 2537 6068 2568
rect 6084 2537 6146 2568
rect 6215 2566 6264 2591
rect 6279 2566 6309 2582
rect 6178 2552 6208 2560
rect 6215 2558 6325 2566
rect 6178 2544 6223 2552
rect 5910 2526 5929 2528
rect 5944 2526 5990 2528
rect 5910 2510 5990 2526
rect 6017 2524 6052 2537
rect 6093 2534 6130 2537
rect 6093 2532 6135 2534
rect 6022 2521 6052 2524
rect 6031 2517 6038 2521
rect 6038 2516 6039 2517
rect 5997 2510 6007 2516
rect 5756 2502 5791 2510
rect 5756 2476 5757 2502
rect 5764 2476 5791 2502
rect 5699 2458 5729 2472
rect 5756 2468 5791 2476
rect 5793 2502 5834 2510
rect 5793 2476 5808 2502
rect 5815 2476 5834 2502
rect 5898 2498 5929 2510
rect 5944 2498 6047 2510
rect 6059 2500 6085 2526
rect 6100 2521 6130 2532
rect 6162 2528 6224 2544
rect 6162 2526 6208 2528
rect 6162 2510 6224 2526
rect 6236 2510 6242 2558
rect 6245 2550 6325 2558
rect 6245 2548 6264 2550
rect 6279 2548 6313 2550
rect 6245 2532 6325 2548
rect 6245 2510 6264 2532
rect 6279 2516 6309 2532
rect 6337 2526 6343 2600
rect 6346 2526 6365 2670
rect 6380 2526 6386 2670
rect 6395 2600 6408 2670
rect 6460 2666 6482 2670
rect 6453 2644 6482 2658
rect 6535 2644 6551 2658
rect 6589 2654 6595 2656
rect 6602 2654 6710 2670
rect 6717 2654 6723 2656
rect 6731 2654 6746 2670
rect 6812 2664 6831 2667
rect 6453 2642 6551 2644
rect 6578 2642 6746 2654
rect 6761 2644 6777 2658
rect 6812 2645 6834 2664
rect 6844 2658 6860 2659
rect 6843 2656 6860 2658
rect 6844 2651 6860 2656
rect 6834 2644 6840 2645
rect 6843 2644 6872 2651
rect 6761 2643 6872 2644
rect 6761 2642 6878 2643
rect 6437 2634 6488 2642
rect 6535 2634 6569 2642
rect 6437 2622 6462 2634
rect 6469 2622 6488 2634
rect 6542 2632 6569 2634
rect 6578 2632 6799 2642
rect 6834 2639 6840 2642
rect 6542 2628 6799 2632
rect 6437 2614 6488 2622
rect 6535 2614 6799 2628
rect 6843 2634 6878 2642
rect 6389 2566 6408 2600
rect 6453 2606 6482 2614
rect 6453 2600 6470 2606
rect 6453 2598 6487 2600
rect 6535 2598 6551 2614
rect 6552 2604 6760 2614
rect 6761 2604 6777 2614
rect 6825 2610 6840 2625
rect 6843 2622 6844 2634
rect 6851 2622 6878 2634
rect 6843 2614 6878 2622
rect 6843 2613 6872 2614
rect 6563 2600 6777 2604
rect 6578 2598 6777 2600
rect 6812 2600 6825 2610
rect 6843 2600 6860 2613
rect 6812 2598 6860 2600
rect 6454 2594 6487 2598
rect 6450 2592 6487 2594
rect 6450 2591 6517 2592
rect 6450 2586 6481 2591
rect 6487 2586 6517 2591
rect 6450 2582 6517 2586
rect 6423 2579 6517 2582
rect 6423 2572 6472 2579
rect 6423 2566 6453 2572
rect 6472 2567 6477 2572
rect 6389 2550 6469 2566
rect 6481 2558 6517 2579
rect 6578 2574 6767 2598
rect 6812 2597 6859 2598
rect 6825 2592 6859 2597
rect 6593 2571 6767 2574
rect 6586 2568 6767 2571
rect 6795 2591 6859 2592
rect 6389 2548 6408 2550
rect 6423 2548 6457 2550
rect 6389 2532 6469 2548
rect 6389 2526 6408 2532
rect 6105 2500 6208 2510
rect 6059 2498 6208 2500
rect 6229 2498 6264 2510
rect 5898 2496 6060 2498
rect 5910 2476 5929 2496
rect 5944 2494 5974 2496
rect 5793 2468 5834 2476
rect 5916 2472 5929 2476
rect 5981 2480 6060 2496
rect 6092 2496 6264 2498
rect 6092 2480 6171 2496
rect 6178 2494 6208 2496
rect 5756 2458 5785 2468
rect 5799 2458 5828 2468
rect 5843 2458 5873 2472
rect 5916 2458 5959 2472
rect 5981 2468 6171 2480
rect 6236 2476 6242 2496
rect 5966 2458 5996 2468
rect 5997 2458 6155 2468
rect 6159 2458 6189 2468
rect 6193 2458 6223 2472
rect 6251 2458 6264 2496
rect 6336 2510 6365 2526
rect 6379 2510 6408 2526
rect 6423 2516 6453 2532
rect 6481 2510 6487 2558
rect 6490 2552 6509 2558
rect 6524 2552 6554 2560
rect 6490 2544 6554 2552
rect 6490 2528 6570 2544
rect 6586 2537 6648 2568
rect 6664 2537 6726 2568
rect 6795 2566 6844 2591
rect 6859 2566 6889 2582
rect 6758 2552 6788 2560
rect 6795 2558 6905 2566
rect 6758 2544 6803 2552
rect 6490 2526 6509 2528
rect 6524 2526 6570 2528
rect 6490 2510 6570 2526
rect 6597 2524 6632 2537
rect 6673 2534 6710 2537
rect 6673 2532 6715 2534
rect 6602 2521 6632 2524
rect 6611 2517 6618 2521
rect 6618 2516 6619 2517
rect 6577 2510 6587 2516
rect 6336 2502 6371 2510
rect 6336 2476 6337 2502
rect 6344 2476 6371 2502
rect 6279 2458 6309 2472
rect 6336 2468 6371 2476
rect 6373 2502 6414 2510
rect 6373 2476 6388 2502
rect 6395 2476 6414 2502
rect 6478 2498 6509 2510
rect 6524 2498 6627 2510
rect 6639 2500 6665 2526
rect 6680 2521 6710 2532
rect 6742 2528 6804 2544
rect 6742 2526 6788 2528
rect 6742 2510 6804 2526
rect 6816 2510 6822 2558
rect 6825 2550 6905 2558
rect 6825 2548 6844 2550
rect 6859 2548 6893 2550
rect 6825 2532 6905 2548
rect 6825 2510 6844 2532
rect 6859 2516 6889 2532
rect 6917 2526 6923 2600
rect 6926 2526 6945 2670
rect 6960 2526 6966 2670
rect 6975 2600 6988 2670
rect 7040 2666 7062 2670
rect 7033 2644 7062 2658
rect 7115 2644 7131 2658
rect 7169 2654 7175 2656
rect 7182 2654 7290 2670
rect 7297 2654 7303 2656
rect 7311 2654 7326 2670
rect 7392 2664 7411 2667
rect 7033 2642 7131 2644
rect 7158 2642 7326 2654
rect 7341 2644 7357 2658
rect 7392 2645 7414 2664
rect 7424 2658 7440 2659
rect 7423 2656 7440 2658
rect 7424 2651 7440 2656
rect 7414 2644 7420 2645
rect 7423 2644 7452 2651
rect 7341 2643 7452 2644
rect 7341 2642 7458 2643
rect 7017 2634 7068 2642
rect 7115 2634 7149 2642
rect 7017 2622 7042 2634
rect 7049 2622 7068 2634
rect 7122 2632 7149 2634
rect 7158 2632 7379 2642
rect 7414 2639 7420 2642
rect 7122 2628 7379 2632
rect 7017 2614 7068 2622
rect 7115 2614 7379 2628
rect 7423 2634 7458 2642
rect 6969 2566 6988 2600
rect 7033 2606 7062 2614
rect 7033 2600 7050 2606
rect 7033 2598 7067 2600
rect 7115 2598 7131 2614
rect 7132 2604 7340 2614
rect 7341 2604 7357 2614
rect 7405 2610 7420 2625
rect 7423 2622 7424 2634
rect 7431 2622 7458 2634
rect 7423 2614 7458 2622
rect 7423 2613 7452 2614
rect 7151 2600 7357 2604
rect 7158 2598 7357 2600
rect 7392 2600 7405 2610
rect 7423 2600 7440 2613
rect 7392 2598 7440 2600
rect 7034 2594 7067 2598
rect 7030 2592 7067 2594
rect 7030 2591 7097 2592
rect 7030 2586 7061 2591
rect 7067 2586 7097 2591
rect 7030 2582 7097 2586
rect 7003 2579 7097 2582
rect 7003 2572 7052 2579
rect 7003 2566 7033 2572
rect 7052 2567 7057 2572
rect 6969 2550 7049 2566
rect 7061 2558 7097 2579
rect 7158 2574 7347 2598
rect 7392 2597 7439 2598
rect 7405 2592 7439 2597
rect 7173 2571 7347 2574
rect 7166 2568 7347 2571
rect 7375 2591 7439 2592
rect 6969 2548 6988 2550
rect 7003 2548 7037 2550
rect 6969 2532 7049 2548
rect 6969 2526 6988 2532
rect 6685 2500 6788 2510
rect 6639 2498 6788 2500
rect 6809 2498 6844 2510
rect 6478 2496 6640 2498
rect 6490 2476 6509 2496
rect 6524 2494 6554 2496
rect 6373 2468 6414 2476
rect 6496 2472 6509 2476
rect 6561 2480 6640 2496
rect 6672 2496 6844 2498
rect 6672 2480 6751 2496
rect 6758 2494 6788 2496
rect 6336 2458 6365 2468
rect 6379 2458 6408 2468
rect 6423 2458 6453 2472
rect 6496 2458 6539 2472
rect 6561 2468 6751 2480
rect 6816 2476 6822 2496
rect 6546 2458 6576 2468
rect 6577 2458 6735 2468
rect 6739 2458 6769 2468
rect 6773 2458 6803 2472
rect 6831 2458 6844 2496
rect 6916 2510 6945 2526
rect 6959 2510 6988 2526
rect 7003 2516 7033 2532
rect 7061 2510 7067 2558
rect 7070 2552 7089 2558
rect 7104 2552 7134 2560
rect 7070 2544 7134 2552
rect 7070 2528 7150 2544
rect 7166 2537 7228 2568
rect 7244 2537 7306 2568
rect 7375 2566 7424 2591
rect 7439 2566 7469 2582
rect 7338 2552 7368 2560
rect 7375 2558 7485 2566
rect 7338 2544 7383 2552
rect 7070 2526 7089 2528
rect 7104 2526 7150 2528
rect 7070 2510 7150 2526
rect 7177 2524 7212 2537
rect 7253 2534 7290 2537
rect 7253 2532 7295 2534
rect 7182 2521 7212 2524
rect 7191 2517 7198 2521
rect 7198 2516 7199 2517
rect 7157 2510 7167 2516
rect 6916 2502 6951 2510
rect 6916 2476 6917 2502
rect 6924 2476 6951 2502
rect 6859 2458 6889 2472
rect 6916 2468 6951 2476
rect 6953 2502 6994 2510
rect 6953 2476 6968 2502
rect 6975 2476 6994 2502
rect 7058 2498 7089 2510
rect 7104 2498 7207 2510
rect 7219 2500 7245 2526
rect 7260 2521 7290 2532
rect 7322 2528 7384 2544
rect 7322 2526 7368 2528
rect 7322 2510 7384 2526
rect 7396 2510 7402 2558
rect 7405 2550 7485 2558
rect 7405 2548 7424 2550
rect 7439 2548 7473 2550
rect 7405 2532 7485 2548
rect 7405 2510 7424 2532
rect 7439 2516 7469 2532
rect 7497 2526 7503 2600
rect 7506 2526 7525 2670
rect 7540 2526 7546 2670
rect 7555 2600 7568 2670
rect 7620 2666 7642 2670
rect 7613 2644 7642 2658
rect 7695 2644 7711 2658
rect 7749 2654 7755 2656
rect 7762 2654 7870 2670
rect 7877 2654 7883 2656
rect 7891 2654 7906 2670
rect 7972 2664 7991 2667
rect 7613 2642 7711 2644
rect 7738 2642 7906 2654
rect 7921 2644 7937 2658
rect 7972 2645 7994 2664
rect 8004 2658 8020 2659
rect 8003 2656 8020 2658
rect 8004 2651 8020 2656
rect 7994 2644 8000 2645
rect 8003 2644 8032 2651
rect 7921 2643 8032 2644
rect 7921 2642 8038 2643
rect 7597 2634 7648 2642
rect 7695 2634 7729 2642
rect 7597 2622 7622 2634
rect 7629 2622 7648 2634
rect 7702 2632 7729 2634
rect 7738 2632 7959 2642
rect 7994 2639 8000 2642
rect 7702 2628 7959 2632
rect 7597 2614 7648 2622
rect 7695 2614 7959 2628
rect 8003 2634 8038 2642
rect 7549 2566 7568 2600
rect 7613 2606 7642 2614
rect 7613 2600 7630 2606
rect 7613 2598 7647 2600
rect 7695 2598 7711 2614
rect 7712 2604 7920 2614
rect 7921 2604 7937 2614
rect 7985 2610 8000 2625
rect 8003 2622 8004 2634
rect 8011 2622 8038 2634
rect 8003 2614 8038 2622
rect 8003 2613 8032 2614
rect 7723 2600 7937 2604
rect 7738 2598 7937 2600
rect 7972 2600 7985 2610
rect 8003 2600 8020 2613
rect 7972 2598 8020 2600
rect 7614 2594 7647 2598
rect 7610 2592 7647 2594
rect 7610 2591 7677 2592
rect 7610 2586 7641 2591
rect 7647 2586 7677 2591
rect 7610 2582 7677 2586
rect 7583 2579 7677 2582
rect 7583 2572 7632 2579
rect 7583 2566 7613 2572
rect 7632 2567 7637 2572
rect 7549 2550 7629 2566
rect 7641 2558 7677 2579
rect 7738 2574 7927 2598
rect 7972 2597 8019 2598
rect 7985 2592 8019 2597
rect 7753 2571 7927 2574
rect 7746 2568 7927 2571
rect 7955 2591 8019 2592
rect 7549 2548 7568 2550
rect 7583 2548 7617 2550
rect 7549 2532 7629 2548
rect 7549 2526 7568 2532
rect 7265 2500 7368 2510
rect 7219 2498 7368 2500
rect 7389 2498 7424 2510
rect 7058 2496 7220 2498
rect 7070 2476 7089 2496
rect 7104 2494 7134 2496
rect 6953 2468 6994 2476
rect 7076 2472 7089 2476
rect 7141 2480 7220 2496
rect 7252 2496 7424 2498
rect 7252 2480 7331 2496
rect 7338 2494 7368 2496
rect 6916 2458 6945 2468
rect 6959 2458 6988 2468
rect 7003 2458 7033 2472
rect 7076 2458 7119 2472
rect 7141 2468 7331 2480
rect 7396 2476 7402 2496
rect 7126 2458 7156 2468
rect 7157 2458 7315 2468
rect 7319 2458 7349 2468
rect 7353 2458 7383 2472
rect 7411 2458 7424 2496
rect 7496 2510 7525 2526
rect 7539 2510 7568 2526
rect 7583 2516 7613 2532
rect 7641 2510 7647 2558
rect 7650 2552 7669 2558
rect 7684 2552 7714 2560
rect 7650 2544 7714 2552
rect 7650 2528 7730 2544
rect 7746 2537 7808 2568
rect 7824 2537 7886 2568
rect 7955 2566 8004 2591
rect 8019 2566 8049 2582
rect 7918 2552 7948 2560
rect 7955 2558 8065 2566
rect 7918 2544 7963 2552
rect 7650 2526 7669 2528
rect 7684 2526 7730 2528
rect 7650 2510 7730 2526
rect 7757 2524 7792 2537
rect 7833 2534 7870 2537
rect 7833 2532 7875 2534
rect 7762 2521 7792 2524
rect 7771 2517 7778 2521
rect 7778 2516 7779 2517
rect 7737 2510 7747 2516
rect 7496 2502 7531 2510
rect 7496 2476 7497 2502
rect 7504 2476 7531 2502
rect 7439 2458 7469 2472
rect 7496 2468 7531 2476
rect 7533 2502 7574 2510
rect 7533 2476 7548 2502
rect 7555 2476 7574 2502
rect 7638 2498 7669 2510
rect 7684 2498 7787 2510
rect 7799 2500 7825 2526
rect 7840 2521 7870 2532
rect 7902 2528 7964 2544
rect 7902 2526 7948 2528
rect 7902 2510 7964 2526
rect 7976 2510 7982 2558
rect 7985 2550 8065 2558
rect 7985 2548 8004 2550
rect 8019 2548 8053 2550
rect 7985 2532 8065 2548
rect 7985 2510 8004 2532
rect 8019 2516 8049 2532
rect 8077 2526 8083 2600
rect 8086 2526 8105 2670
rect 8120 2526 8126 2670
rect 8135 2600 8148 2670
rect 8200 2666 8222 2670
rect 8193 2644 8222 2658
rect 8275 2644 8291 2658
rect 8329 2654 8335 2656
rect 8342 2654 8450 2670
rect 8457 2654 8463 2656
rect 8471 2654 8486 2670
rect 8552 2664 8571 2667
rect 8193 2642 8291 2644
rect 8318 2642 8486 2654
rect 8501 2644 8517 2658
rect 8552 2645 8574 2664
rect 8584 2658 8600 2659
rect 8583 2656 8600 2658
rect 8584 2651 8600 2656
rect 8574 2644 8580 2645
rect 8583 2644 8612 2651
rect 8501 2643 8612 2644
rect 8501 2642 8618 2643
rect 8177 2634 8228 2642
rect 8275 2634 8309 2642
rect 8177 2622 8202 2634
rect 8209 2622 8228 2634
rect 8282 2632 8309 2634
rect 8318 2632 8539 2642
rect 8574 2639 8580 2642
rect 8282 2628 8539 2632
rect 8177 2614 8228 2622
rect 8275 2614 8539 2628
rect 8583 2634 8618 2642
rect 8129 2566 8148 2600
rect 8193 2606 8222 2614
rect 8193 2600 8210 2606
rect 8193 2598 8227 2600
rect 8275 2598 8291 2614
rect 8292 2604 8500 2614
rect 8501 2604 8517 2614
rect 8565 2610 8580 2625
rect 8583 2622 8584 2634
rect 8591 2622 8618 2634
rect 8583 2614 8618 2622
rect 8583 2613 8612 2614
rect 8303 2600 8517 2604
rect 8318 2598 8517 2600
rect 8552 2600 8565 2610
rect 8583 2600 8600 2613
rect 8552 2598 8600 2600
rect 8194 2594 8227 2598
rect 8190 2592 8227 2594
rect 8190 2591 8257 2592
rect 8190 2586 8221 2591
rect 8227 2586 8257 2591
rect 8190 2582 8257 2586
rect 8163 2579 8257 2582
rect 8163 2572 8212 2579
rect 8163 2566 8193 2572
rect 8212 2567 8217 2572
rect 8129 2550 8209 2566
rect 8221 2558 8257 2579
rect 8318 2574 8507 2598
rect 8552 2597 8599 2598
rect 8565 2592 8599 2597
rect 8333 2571 8507 2574
rect 8326 2568 8507 2571
rect 8535 2591 8599 2592
rect 8129 2548 8148 2550
rect 8163 2548 8197 2550
rect 8129 2532 8209 2548
rect 8129 2526 8148 2532
rect 7845 2500 7948 2510
rect 7799 2498 7948 2500
rect 7969 2498 8004 2510
rect 7638 2496 7800 2498
rect 7650 2476 7669 2496
rect 7684 2494 7714 2496
rect 7533 2468 7574 2476
rect 7656 2472 7669 2476
rect 7721 2480 7800 2496
rect 7832 2496 8004 2498
rect 7832 2480 7911 2496
rect 7918 2494 7948 2496
rect 7496 2458 7525 2468
rect 7539 2458 7568 2468
rect 7583 2458 7613 2472
rect 7656 2458 7699 2472
rect 7721 2468 7911 2480
rect 7976 2476 7982 2496
rect 7706 2458 7736 2468
rect 7737 2458 7895 2468
rect 7899 2458 7929 2468
rect 7933 2458 7963 2472
rect 7991 2458 8004 2496
rect 8076 2510 8105 2526
rect 8119 2510 8148 2526
rect 8163 2516 8193 2532
rect 8221 2510 8227 2558
rect 8230 2552 8249 2558
rect 8264 2552 8294 2560
rect 8230 2544 8294 2552
rect 8230 2528 8310 2544
rect 8326 2537 8388 2568
rect 8404 2537 8466 2568
rect 8535 2566 8584 2591
rect 8599 2566 8629 2582
rect 8498 2552 8528 2560
rect 8535 2558 8645 2566
rect 8498 2544 8543 2552
rect 8230 2526 8249 2528
rect 8264 2526 8310 2528
rect 8230 2510 8310 2526
rect 8337 2524 8372 2537
rect 8413 2534 8450 2537
rect 8413 2532 8455 2534
rect 8342 2521 8372 2524
rect 8351 2517 8358 2521
rect 8358 2516 8359 2517
rect 8317 2510 8327 2516
rect 8076 2502 8111 2510
rect 8076 2476 8077 2502
rect 8084 2476 8111 2502
rect 8019 2458 8049 2472
rect 8076 2468 8111 2476
rect 8113 2502 8154 2510
rect 8113 2476 8128 2502
rect 8135 2476 8154 2502
rect 8218 2498 8249 2510
rect 8264 2498 8367 2510
rect 8379 2500 8405 2526
rect 8420 2521 8450 2532
rect 8482 2528 8544 2544
rect 8482 2526 8528 2528
rect 8482 2510 8544 2526
rect 8556 2510 8562 2558
rect 8565 2550 8645 2558
rect 8565 2548 8584 2550
rect 8599 2548 8633 2550
rect 8565 2532 8645 2548
rect 8565 2510 8584 2532
rect 8599 2516 8629 2532
rect 8657 2526 8663 2600
rect 8666 2526 8685 2670
rect 8700 2526 8706 2670
rect 8715 2600 8728 2670
rect 8780 2666 8802 2670
rect 8773 2644 8802 2658
rect 8855 2644 8871 2658
rect 8909 2654 8915 2656
rect 8922 2654 9030 2670
rect 9037 2654 9043 2656
rect 9051 2654 9066 2670
rect 9132 2664 9151 2667
rect 8773 2642 8871 2644
rect 8898 2642 9066 2654
rect 9081 2644 9097 2658
rect 9132 2645 9154 2664
rect 9164 2658 9180 2659
rect 9163 2656 9180 2658
rect 9164 2651 9180 2656
rect 9154 2644 9160 2645
rect 9163 2644 9192 2651
rect 9081 2643 9192 2644
rect 9081 2642 9198 2643
rect 8757 2634 8808 2642
rect 8855 2634 8889 2642
rect 8757 2622 8782 2634
rect 8789 2622 8808 2634
rect 8862 2632 8889 2634
rect 8898 2632 9119 2642
rect 9154 2639 9160 2642
rect 8862 2628 9119 2632
rect 8757 2614 8808 2622
rect 8855 2614 9119 2628
rect 9163 2634 9198 2642
rect 8709 2566 8728 2600
rect 8773 2606 8802 2614
rect 8773 2600 8790 2606
rect 8773 2598 8807 2600
rect 8855 2598 8871 2614
rect 8872 2604 9080 2614
rect 9081 2604 9097 2614
rect 9145 2610 9160 2625
rect 9163 2622 9164 2634
rect 9171 2622 9198 2634
rect 9163 2614 9198 2622
rect 9163 2613 9192 2614
rect 8883 2600 9097 2604
rect 8898 2598 9097 2600
rect 9132 2600 9145 2610
rect 9163 2600 9180 2613
rect 9132 2598 9180 2600
rect 8774 2594 8807 2598
rect 8770 2592 8807 2594
rect 8770 2591 8837 2592
rect 8770 2586 8801 2591
rect 8807 2586 8837 2591
rect 8770 2582 8837 2586
rect 8743 2579 8837 2582
rect 8743 2572 8792 2579
rect 8743 2566 8773 2572
rect 8792 2567 8797 2572
rect 8709 2550 8789 2566
rect 8801 2558 8837 2579
rect 8898 2574 9087 2598
rect 9132 2597 9179 2598
rect 9145 2592 9179 2597
rect 8913 2571 9087 2574
rect 8906 2568 9087 2571
rect 9115 2591 9179 2592
rect 8709 2548 8728 2550
rect 8743 2548 8777 2550
rect 8709 2532 8789 2548
rect 8709 2526 8728 2532
rect 8425 2500 8528 2510
rect 8379 2498 8528 2500
rect 8549 2498 8584 2510
rect 8218 2496 8380 2498
rect 8230 2476 8249 2496
rect 8264 2494 8294 2496
rect 8113 2468 8154 2476
rect 8236 2472 8249 2476
rect 8301 2480 8380 2496
rect 8412 2496 8584 2498
rect 8412 2480 8491 2496
rect 8498 2494 8528 2496
rect 8076 2458 8105 2468
rect 8119 2458 8148 2468
rect 8163 2458 8193 2472
rect 8236 2458 8279 2472
rect 8301 2468 8491 2480
rect 8556 2476 8562 2496
rect 8286 2458 8316 2468
rect 8317 2458 8475 2468
rect 8479 2458 8509 2468
rect 8513 2458 8543 2472
rect 8571 2458 8584 2496
rect 8656 2510 8685 2526
rect 8699 2510 8728 2526
rect 8743 2516 8773 2532
rect 8801 2510 8807 2558
rect 8810 2552 8829 2558
rect 8844 2552 8874 2560
rect 8810 2544 8874 2552
rect 8810 2528 8890 2544
rect 8906 2537 8968 2568
rect 8984 2537 9046 2568
rect 9115 2566 9164 2591
rect 9179 2566 9209 2582
rect 9078 2552 9108 2560
rect 9115 2558 9225 2566
rect 9078 2544 9123 2552
rect 8810 2526 8829 2528
rect 8844 2526 8890 2528
rect 8810 2510 8890 2526
rect 8917 2524 8952 2537
rect 8993 2534 9030 2537
rect 8993 2532 9035 2534
rect 8922 2521 8952 2524
rect 8931 2517 8938 2521
rect 8938 2516 8939 2517
rect 8897 2510 8907 2516
rect 8656 2502 8691 2510
rect 8656 2476 8657 2502
rect 8664 2476 8691 2502
rect 8599 2458 8629 2472
rect 8656 2468 8691 2476
rect 8693 2502 8734 2510
rect 8693 2476 8708 2502
rect 8715 2476 8734 2502
rect 8798 2498 8829 2510
rect 8844 2498 8947 2510
rect 8959 2500 8985 2526
rect 9000 2521 9030 2532
rect 9062 2528 9124 2544
rect 9062 2526 9108 2528
rect 9062 2510 9124 2526
rect 9136 2510 9142 2558
rect 9145 2550 9225 2558
rect 9145 2548 9164 2550
rect 9179 2548 9213 2550
rect 9145 2532 9225 2548
rect 9145 2510 9164 2532
rect 9179 2516 9209 2532
rect 9237 2526 9243 2600
rect 9246 2526 9265 2670
rect 9280 2526 9286 2670
rect 9295 2600 9308 2670
rect 9360 2666 9382 2670
rect 9353 2644 9382 2658
rect 9435 2644 9451 2658
rect 9489 2654 9495 2656
rect 9502 2654 9610 2670
rect 9617 2654 9623 2656
rect 9631 2654 9646 2670
rect 9712 2664 9731 2667
rect 9353 2642 9451 2644
rect 9478 2642 9646 2654
rect 9661 2644 9677 2658
rect 9712 2645 9734 2664
rect 9744 2658 9760 2659
rect 9743 2656 9760 2658
rect 9744 2651 9760 2656
rect 9734 2644 9740 2645
rect 9743 2644 9772 2651
rect 9661 2643 9772 2644
rect 9661 2642 9778 2643
rect 9337 2634 9388 2642
rect 9435 2634 9469 2642
rect 9337 2622 9362 2634
rect 9369 2622 9388 2634
rect 9442 2632 9469 2634
rect 9478 2632 9699 2642
rect 9734 2639 9740 2642
rect 9442 2628 9699 2632
rect 9337 2614 9388 2622
rect 9435 2614 9699 2628
rect 9743 2634 9778 2642
rect 9289 2566 9308 2600
rect 9353 2606 9382 2614
rect 9353 2600 9370 2606
rect 9353 2598 9387 2600
rect 9435 2598 9451 2614
rect 9452 2604 9660 2614
rect 9661 2604 9677 2614
rect 9725 2610 9740 2625
rect 9743 2622 9744 2634
rect 9751 2622 9778 2634
rect 9743 2614 9778 2622
rect 9743 2613 9772 2614
rect 9463 2600 9677 2604
rect 9478 2598 9677 2600
rect 9712 2600 9725 2610
rect 9743 2600 9760 2613
rect 9712 2598 9760 2600
rect 9354 2594 9387 2598
rect 9350 2592 9387 2594
rect 9350 2591 9417 2592
rect 9350 2586 9381 2591
rect 9387 2586 9417 2591
rect 9350 2582 9417 2586
rect 9323 2579 9417 2582
rect 9323 2572 9372 2579
rect 9323 2566 9353 2572
rect 9372 2567 9377 2572
rect 9289 2550 9369 2566
rect 9381 2558 9417 2579
rect 9478 2574 9667 2598
rect 9712 2597 9759 2598
rect 9725 2592 9759 2597
rect 9493 2571 9667 2574
rect 9486 2568 9667 2571
rect 9695 2591 9759 2592
rect 9289 2548 9308 2550
rect 9323 2548 9357 2550
rect 9289 2532 9369 2548
rect 9289 2526 9308 2532
rect 9005 2500 9108 2510
rect 8959 2498 9108 2500
rect 9129 2498 9164 2510
rect 8798 2496 8960 2498
rect 8810 2476 8829 2496
rect 8844 2494 8874 2496
rect 8693 2468 8734 2476
rect 8816 2472 8829 2476
rect 8881 2480 8960 2496
rect 8992 2496 9164 2498
rect 8992 2480 9071 2496
rect 9078 2494 9108 2496
rect 8656 2458 8685 2468
rect 8699 2458 8728 2468
rect 8743 2458 8773 2472
rect 8816 2458 8859 2472
rect 8881 2468 9071 2480
rect 9136 2476 9142 2496
rect 8866 2458 8896 2468
rect 8897 2458 9055 2468
rect 9059 2458 9089 2468
rect 9093 2458 9123 2472
rect 9151 2458 9164 2496
rect 9236 2510 9265 2526
rect 9279 2510 9308 2526
rect 9323 2516 9353 2532
rect 9381 2510 9387 2558
rect 9390 2552 9409 2558
rect 9424 2552 9454 2560
rect 9390 2544 9454 2552
rect 9390 2528 9470 2544
rect 9486 2537 9548 2568
rect 9564 2537 9626 2568
rect 9695 2566 9744 2591
rect 9759 2566 9789 2582
rect 9658 2552 9688 2560
rect 9695 2558 9805 2566
rect 9658 2544 9703 2552
rect 9390 2526 9409 2528
rect 9424 2526 9470 2528
rect 9390 2510 9470 2526
rect 9497 2524 9532 2537
rect 9573 2534 9610 2537
rect 9573 2532 9615 2534
rect 9502 2521 9532 2524
rect 9511 2517 9518 2521
rect 9518 2516 9519 2517
rect 9477 2510 9487 2516
rect 9236 2502 9271 2510
rect 9236 2476 9237 2502
rect 9244 2476 9271 2502
rect 9179 2458 9209 2472
rect 9236 2468 9271 2476
rect 9273 2502 9314 2510
rect 9273 2476 9288 2502
rect 9295 2476 9314 2502
rect 9378 2498 9409 2510
rect 9424 2498 9527 2510
rect 9539 2500 9565 2526
rect 9580 2521 9610 2532
rect 9642 2528 9704 2544
rect 9642 2526 9688 2528
rect 9642 2510 9704 2526
rect 9716 2510 9722 2558
rect 9725 2550 9805 2558
rect 9725 2548 9744 2550
rect 9759 2548 9793 2550
rect 9725 2532 9805 2548
rect 9725 2510 9744 2532
rect 9759 2516 9789 2532
rect 9817 2526 9823 2600
rect 9826 2526 9845 2670
rect 9860 2526 9866 2670
rect 9875 2600 9888 2670
rect 9940 2666 9962 2670
rect 9933 2644 9962 2658
rect 10015 2644 10031 2658
rect 10069 2654 10075 2656
rect 10082 2654 10190 2670
rect 10197 2654 10203 2656
rect 10211 2654 10226 2670
rect 10292 2664 10311 2667
rect 9933 2642 10031 2644
rect 10058 2642 10226 2654
rect 10241 2644 10257 2658
rect 10292 2645 10314 2664
rect 10324 2658 10340 2659
rect 10323 2656 10340 2658
rect 10324 2651 10340 2656
rect 10314 2644 10320 2645
rect 10323 2644 10352 2651
rect 10241 2643 10352 2644
rect 10241 2642 10358 2643
rect 9917 2634 9968 2642
rect 10015 2634 10049 2642
rect 9917 2622 9942 2634
rect 9949 2622 9968 2634
rect 10022 2632 10049 2634
rect 10058 2632 10279 2642
rect 10314 2639 10320 2642
rect 10022 2628 10279 2632
rect 9917 2614 9968 2622
rect 10015 2614 10279 2628
rect 10323 2634 10358 2642
rect 9869 2566 9888 2600
rect 9933 2606 9962 2614
rect 9933 2600 9950 2606
rect 9933 2598 9967 2600
rect 10015 2598 10031 2614
rect 10032 2604 10240 2614
rect 10241 2604 10257 2614
rect 10305 2610 10320 2625
rect 10323 2622 10324 2634
rect 10331 2622 10358 2634
rect 10323 2614 10358 2622
rect 10323 2613 10352 2614
rect 10043 2600 10257 2604
rect 10058 2598 10257 2600
rect 10292 2600 10305 2610
rect 10323 2600 10340 2613
rect 10292 2598 10340 2600
rect 9934 2594 9967 2598
rect 9930 2592 9967 2594
rect 9930 2591 9997 2592
rect 9930 2586 9961 2591
rect 9967 2586 9997 2591
rect 9930 2582 9997 2586
rect 9903 2579 9997 2582
rect 9903 2572 9952 2579
rect 9903 2566 9933 2572
rect 9952 2567 9957 2572
rect 9869 2550 9949 2566
rect 9961 2558 9997 2579
rect 10058 2574 10247 2598
rect 10292 2597 10339 2598
rect 10305 2592 10339 2597
rect 10073 2571 10247 2574
rect 10066 2568 10247 2571
rect 10275 2591 10339 2592
rect 9869 2548 9888 2550
rect 9903 2548 9937 2550
rect 9869 2532 9949 2548
rect 9869 2526 9888 2532
rect 9585 2500 9688 2510
rect 9539 2498 9688 2500
rect 9709 2498 9744 2510
rect 9378 2496 9540 2498
rect 9390 2476 9409 2496
rect 9424 2494 9454 2496
rect 9273 2468 9314 2476
rect 9396 2472 9409 2476
rect 9461 2480 9540 2496
rect 9572 2496 9744 2498
rect 9572 2480 9651 2496
rect 9658 2494 9688 2496
rect 9236 2458 9265 2468
rect 9279 2458 9308 2468
rect 9323 2458 9353 2472
rect 9396 2458 9439 2472
rect 9461 2468 9651 2480
rect 9716 2476 9722 2496
rect 9446 2458 9476 2468
rect 9477 2458 9635 2468
rect 9639 2458 9669 2468
rect 9673 2458 9703 2472
rect 9731 2458 9744 2496
rect 9816 2510 9845 2526
rect 9859 2510 9888 2526
rect 9903 2516 9933 2532
rect 9961 2510 9967 2558
rect 9970 2552 9989 2558
rect 10004 2552 10034 2560
rect 9970 2544 10034 2552
rect 9970 2528 10050 2544
rect 10066 2537 10128 2568
rect 10144 2537 10206 2568
rect 10275 2566 10324 2591
rect 10339 2566 10369 2582
rect 10238 2552 10268 2560
rect 10275 2558 10385 2566
rect 10238 2544 10283 2552
rect 9970 2526 9989 2528
rect 10004 2526 10050 2528
rect 9970 2510 10050 2526
rect 10077 2524 10112 2537
rect 10153 2534 10190 2537
rect 10153 2532 10195 2534
rect 10082 2521 10112 2524
rect 10091 2517 10098 2521
rect 10098 2516 10099 2517
rect 10057 2510 10067 2516
rect 9816 2502 9851 2510
rect 9816 2476 9817 2502
rect 9824 2476 9851 2502
rect 9759 2458 9789 2472
rect 9816 2468 9851 2476
rect 9853 2502 9894 2510
rect 9853 2476 9868 2502
rect 9875 2476 9894 2502
rect 9958 2498 9989 2510
rect 10004 2498 10107 2510
rect 10119 2500 10145 2526
rect 10160 2521 10190 2532
rect 10222 2528 10284 2544
rect 10222 2526 10268 2528
rect 10222 2510 10284 2526
rect 10296 2510 10302 2558
rect 10305 2550 10385 2558
rect 10305 2548 10324 2550
rect 10339 2548 10373 2550
rect 10305 2532 10385 2548
rect 10305 2510 10324 2532
rect 10339 2516 10369 2532
rect 10397 2526 10403 2600
rect 10406 2526 10425 2670
rect 10440 2526 10446 2670
rect 10455 2600 10468 2670
rect 10520 2666 10542 2670
rect 10513 2644 10542 2658
rect 10595 2644 10611 2658
rect 10649 2654 10655 2656
rect 10662 2654 10770 2670
rect 10777 2654 10783 2656
rect 10791 2654 10806 2670
rect 10872 2664 10891 2667
rect 10513 2642 10611 2644
rect 10638 2642 10806 2654
rect 10821 2644 10837 2658
rect 10872 2645 10894 2664
rect 10904 2658 10920 2659
rect 10903 2656 10920 2658
rect 10904 2651 10920 2656
rect 10894 2644 10900 2645
rect 10903 2644 10932 2651
rect 10821 2643 10932 2644
rect 10821 2642 10938 2643
rect 10497 2634 10548 2642
rect 10595 2634 10629 2642
rect 10497 2622 10522 2634
rect 10529 2622 10548 2634
rect 10602 2632 10629 2634
rect 10638 2632 10859 2642
rect 10894 2639 10900 2642
rect 10602 2628 10859 2632
rect 10497 2614 10548 2622
rect 10595 2614 10859 2628
rect 10903 2634 10938 2642
rect 10449 2566 10468 2600
rect 10513 2606 10542 2614
rect 10513 2600 10530 2606
rect 10513 2598 10547 2600
rect 10595 2598 10611 2614
rect 10612 2604 10820 2614
rect 10821 2604 10837 2614
rect 10885 2610 10900 2625
rect 10903 2622 10904 2634
rect 10911 2622 10938 2634
rect 10903 2614 10938 2622
rect 10903 2613 10932 2614
rect 10623 2600 10837 2604
rect 10638 2598 10837 2600
rect 10872 2600 10885 2610
rect 10903 2600 10920 2613
rect 10872 2598 10920 2600
rect 10514 2594 10547 2598
rect 10510 2592 10547 2594
rect 10510 2591 10577 2592
rect 10510 2586 10541 2591
rect 10547 2586 10577 2591
rect 10510 2582 10577 2586
rect 10483 2579 10577 2582
rect 10483 2572 10532 2579
rect 10483 2566 10513 2572
rect 10532 2567 10537 2572
rect 10449 2550 10529 2566
rect 10541 2558 10577 2579
rect 10638 2574 10827 2598
rect 10872 2597 10919 2598
rect 10885 2592 10919 2597
rect 10653 2571 10827 2574
rect 10646 2568 10827 2571
rect 10855 2591 10919 2592
rect 10449 2548 10468 2550
rect 10483 2548 10517 2550
rect 10449 2532 10529 2548
rect 10449 2526 10468 2532
rect 10165 2500 10268 2510
rect 10119 2498 10268 2500
rect 10289 2498 10324 2510
rect 9958 2496 10120 2498
rect 9970 2476 9989 2496
rect 10004 2494 10034 2496
rect 9853 2468 9894 2476
rect 9976 2472 9989 2476
rect 10041 2480 10120 2496
rect 10152 2496 10324 2498
rect 10152 2480 10231 2496
rect 10238 2494 10268 2496
rect 9816 2458 9845 2468
rect 9859 2458 9888 2468
rect 9903 2458 9933 2472
rect 9976 2458 10019 2472
rect 10041 2468 10231 2480
rect 10296 2476 10302 2496
rect 10026 2458 10056 2468
rect 10057 2458 10215 2468
rect 10219 2458 10249 2468
rect 10253 2458 10283 2472
rect 10311 2458 10324 2496
rect 10396 2510 10425 2526
rect 10439 2510 10468 2526
rect 10483 2516 10513 2532
rect 10541 2510 10547 2558
rect 10550 2552 10569 2558
rect 10584 2552 10614 2560
rect 10550 2544 10614 2552
rect 10550 2528 10630 2544
rect 10646 2537 10708 2568
rect 10724 2537 10786 2568
rect 10855 2566 10904 2591
rect 10919 2566 10949 2582
rect 10818 2552 10848 2560
rect 10855 2558 10965 2566
rect 10818 2544 10863 2552
rect 10550 2526 10569 2528
rect 10584 2526 10630 2528
rect 10550 2510 10630 2526
rect 10657 2524 10692 2537
rect 10733 2534 10770 2537
rect 10733 2532 10775 2534
rect 10662 2521 10692 2524
rect 10671 2517 10678 2521
rect 10678 2516 10679 2517
rect 10637 2510 10647 2516
rect 10396 2502 10431 2510
rect 10396 2476 10397 2502
rect 10404 2476 10431 2502
rect 10339 2458 10369 2472
rect 10396 2468 10431 2476
rect 10433 2502 10474 2510
rect 10433 2476 10448 2502
rect 10455 2476 10474 2502
rect 10538 2498 10569 2510
rect 10584 2498 10687 2510
rect 10699 2500 10725 2526
rect 10740 2521 10770 2532
rect 10802 2528 10864 2544
rect 10802 2526 10848 2528
rect 10802 2510 10864 2526
rect 10876 2510 10882 2558
rect 10885 2550 10965 2558
rect 10885 2548 10904 2550
rect 10919 2548 10953 2550
rect 10885 2532 10965 2548
rect 10885 2510 10904 2532
rect 10919 2516 10949 2532
rect 10977 2526 10983 2600
rect 10986 2526 11005 2670
rect 11020 2526 11026 2670
rect 11035 2600 11048 2670
rect 11100 2666 11122 2670
rect 11093 2644 11122 2658
rect 11175 2644 11191 2658
rect 11229 2654 11235 2656
rect 11242 2654 11350 2670
rect 11357 2654 11363 2656
rect 11371 2654 11386 2670
rect 11452 2664 11471 2667
rect 11093 2642 11191 2644
rect 11218 2642 11386 2654
rect 11401 2644 11417 2658
rect 11452 2645 11474 2664
rect 11484 2658 11500 2659
rect 11483 2656 11500 2658
rect 11484 2651 11500 2656
rect 11474 2644 11480 2645
rect 11483 2644 11512 2651
rect 11401 2643 11512 2644
rect 11401 2642 11518 2643
rect 11077 2634 11128 2642
rect 11175 2634 11209 2642
rect 11077 2622 11102 2634
rect 11109 2622 11128 2634
rect 11182 2632 11209 2634
rect 11218 2632 11439 2642
rect 11474 2639 11480 2642
rect 11182 2628 11439 2632
rect 11077 2614 11128 2622
rect 11175 2614 11439 2628
rect 11483 2634 11518 2642
rect 11029 2566 11048 2600
rect 11093 2606 11122 2614
rect 11093 2600 11110 2606
rect 11093 2598 11127 2600
rect 11175 2598 11191 2614
rect 11192 2604 11400 2614
rect 11401 2604 11417 2614
rect 11465 2610 11480 2625
rect 11483 2622 11484 2634
rect 11491 2622 11518 2634
rect 11483 2614 11518 2622
rect 11483 2613 11512 2614
rect 11203 2600 11417 2604
rect 11218 2598 11417 2600
rect 11452 2600 11465 2610
rect 11483 2600 11500 2613
rect 11452 2598 11500 2600
rect 11094 2594 11127 2598
rect 11090 2592 11127 2594
rect 11090 2591 11157 2592
rect 11090 2586 11121 2591
rect 11127 2586 11157 2591
rect 11090 2582 11157 2586
rect 11063 2579 11157 2582
rect 11063 2572 11112 2579
rect 11063 2566 11093 2572
rect 11112 2567 11117 2572
rect 11029 2550 11109 2566
rect 11121 2558 11157 2579
rect 11218 2574 11407 2598
rect 11452 2597 11499 2598
rect 11465 2592 11499 2597
rect 11233 2571 11407 2574
rect 11226 2568 11407 2571
rect 11435 2591 11499 2592
rect 11029 2548 11048 2550
rect 11063 2548 11097 2550
rect 11029 2532 11109 2548
rect 11029 2526 11048 2532
rect 10745 2500 10848 2510
rect 10699 2498 10848 2500
rect 10869 2498 10904 2510
rect 10538 2496 10700 2498
rect 10550 2476 10569 2496
rect 10584 2494 10614 2496
rect 10433 2468 10474 2476
rect 10556 2472 10569 2476
rect 10621 2480 10700 2496
rect 10732 2496 10904 2498
rect 10732 2480 10811 2496
rect 10818 2494 10848 2496
rect 10396 2458 10425 2468
rect 10439 2458 10468 2468
rect 10483 2458 10513 2472
rect 10556 2458 10599 2472
rect 10621 2468 10811 2480
rect 10876 2476 10882 2496
rect 10606 2458 10636 2468
rect 10637 2458 10795 2468
rect 10799 2458 10829 2468
rect 10833 2458 10863 2472
rect 10891 2458 10904 2496
rect 10976 2510 11005 2526
rect 11019 2510 11048 2526
rect 11063 2516 11093 2532
rect 11121 2510 11127 2558
rect 11130 2552 11149 2558
rect 11164 2552 11194 2560
rect 11130 2544 11194 2552
rect 11130 2528 11210 2544
rect 11226 2537 11288 2568
rect 11304 2537 11366 2568
rect 11435 2566 11484 2591
rect 11499 2566 11529 2582
rect 11398 2552 11428 2560
rect 11435 2558 11545 2566
rect 11398 2544 11443 2552
rect 11130 2526 11149 2528
rect 11164 2526 11210 2528
rect 11130 2510 11210 2526
rect 11237 2524 11272 2537
rect 11313 2534 11350 2537
rect 11313 2532 11355 2534
rect 11242 2521 11272 2524
rect 11251 2517 11258 2521
rect 11258 2516 11259 2517
rect 11217 2510 11227 2516
rect 10976 2502 11011 2510
rect 10976 2476 10977 2502
rect 10984 2476 11011 2502
rect 10919 2458 10949 2472
rect 10976 2468 11011 2476
rect 11013 2502 11054 2510
rect 11013 2476 11028 2502
rect 11035 2476 11054 2502
rect 11118 2498 11149 2510
rect 11164 2498 11267 2510
rect 11279 2500 11305 2526
rect 11320 2521 11350 2532
rect 11382 2528 11444 2544
rect 11382 2526 11428 2528
rect 11382 2510 11444 2526
rect 11456 2510 11462 2558
rect 11465 2550 11545 2558
rect 11465 2548 11484 2550
rect 11499 2548 11533 2550
rect 11465 2532 11545 2548
rect 11465 2510 11484 2532
rect 11499 2516 11529 2532
rect 11557 2526 11563 2600
rect 11566 2526 11585 2670
rect 11600 2526 11606 2670
rect 11615 2600 11628 2670
rect 11680 2666 11702 2670
rect 11673 2644 11702 2658
rect 11755 2644 11771 2658
rect 11809 2654 11815 2656
rect 11822 2654 11930 2670
rect 11937 2654 11943 2656
rect 11951 2654 11966 2670
rect 12032 2664 12051 2667
rect 11673 2642 11771 2644
rect 11798 2642 11966 2654
rect 11981 2644 11997 2658
rect 12032 2645 12054 2664
rect 12064 2658 12080 2659
rect 12063 2656 12080 2658
rect 12064 2651 12080 2656
rect 12054 2644 12060 2645
rect 12063 2644 12092 2651
rect 11981 2643 12092 2644
rect 11981 2642 12098 2643
rect 11657 2634 11708 2642
rect 11755 2634 11789 2642
rect 11657 2622 11682 2634
rect 11689 2622 11708 2634
rect 11762 2632 11789 2634
rect 11798 2632 12019 2642
rect 12054 2639 12060 2642
rect 11762 2628 12019 2632
rect 11657 2614 11708 2622
rect 11755 2614 12019 2628
rect 12063 2634 12098 2642
rect 11609 2566 11628 2600
rect 11673 2606 11702 2614
rect 11673 2600 11690 2606
rect 11673 2598 11707 2600
rect 11755 2598 11771 2614
rect 11772 2604 11980 2614
rect 11981 2604 11997 2614
rect 12045 2610 12060 2625
rect 12063 2622 12064 2634
rect 12071 2622 12098 2634
rect 12063 2614 12098 2622
rect 12063 2613 12092 2614
rect 11783 2600 11997 2604
rect 11798 2598 11997 2600
rect 12032 2600 12045 2610
rect 12063 2600 12080 2613
rect 12032 2598 12080 2600
rect 11674 2594 11707 2598
rect 11670 2592 11707 2594
rect 11670 2591 11737 2592
rect 11670 2586 11701 2591
rect 11707 2586 11737 2591
rect 11670 2582 11737 2586
rect 11643 2579 11737 2582
rect 11643 2572 11692 2579
rect 11643 2566 11673 2572
rect 11692 2567 11697 2572
rect 11609 2550 11689 2566
rect 11701 2558 11737 2579
rect 11798 2574 11987 2598
rect 12032 2597 12079 2598
rect 12045 2592 12079 2597
rect 11813 2571 11987 2574
rect 11806 2568 11987 2571
rect 12015 2591 12079 2592
rect 11609 2548 11628 2550
rect 11643 2548 11677 2550
rect 11609 2532 11689 2548
rect 11609 2526 11628 2532
rect 11325 2500 11428 2510
rect 11279 2498 11428 2500
rect 11449 2498 11484 2510
rect 11118 2496 11280 2498
rect 11130 2476 11149 2496
rect 11164 2494 11194 2496
rect 11013 2468 11054 2476
rect 11136 2472 11149 2476
rect 11201 2480 11280 2496
rect 11312 2496 11484 2498
rect 11312 2480 11391 2496
rect 11398 2494 11428 2496
rect 10976 2458 11005 2468
rect 11019 2458 11048 2468
rect 11063 2458 11093 2472
rect 11136 2458 11179 2472
rect 11201 2468 11391 2480
rect 11456 2476 11462 2496
rect 11186 2458 11216 2468
rect 11217 2458 11375 2468
rect 11379 2458 11409 2468
rect 11413 2458 11443 2472
rect 11471 2458 11484 2496
rect 11556 2510 11585 2526
rect 11599 2510 11628 2526
rect 11643 2516 11673 2532
rect 11701 2510 11707 2558
rect 11710 2552 11729 2558
rect 11744 2552 11774 2560
rect 11710 2544 11774 2552
rect 11710 2528 11790 2544
rect 11806 2537 11868 2568
rect 11884 2537 11946 2568
rect 12015 2566 12064 2591
rect 12079 2566 12109 2582
rect 11978 2552 12008 2560
rect 12015 2558 12125 2566
rect 11978 2544 12023 2552
rect 11710 2526 11729 2528
rect 11744 2526 11790 2528
rect 11710 2510 11790 2526
rect 11817 2524 11852 2537
rect 11893 2534 11930 2537
rect 11893 2532 11935 2534
rect 11822 2521 11852 2524
rect 11831 2517 11838 2521
rect 11838 2516 11839 2517
rect 11797 2510 11807 2516
rect 11556 2502 11591 2510
rect 11556 2476 11557 2502
rect 11564 2476 11591 2502
rect 11499 2458 11529 2472
rect 11556 2468 11591 2476
rect 11593 2502 11634 2510
rect 11593 2476 11608 2502
rect 11615 2476 11634 2502
rect 11698 2498 11729 2510
rect 11744 2498 11847 2510
rect 11859 2500 11885 2526
rect 11900 2521 11930 2532
rect 11962 2528 12024 2544
rect 11962 2526 12008 2528
rect 11962 2510 12024 2526
rect 12036 2510 12042 2558
rect 12045 2550 12125 2558
rect 12045 2548 12064 2550
rect 12079 2548 12113 2550
rect 12045 2532 12125 2548
rect 12045 2510 12064 2532
rect 12079 2516 12109 2532
rect 12137 2526 12143 2600
rect 12146 2526 12165 2670
rect 12180 2526 12186 2670
rect 12195 2600 12208 2670
rect 12260 2666 12282 2670
rect 12253 2644 12282 2658
rect 12335 2644 12351 2658
rect 12389 2654 12395 2656
rect 12402 2654 12510 2670
rect 12517 2654 12523 2656
rect 12531 2654 12546 2670
rect 12612 2664 12631 2667
rect 12253 2642 12351 2644
rect 12378 2642 12546 2654
rect 12561 2644 12577 2658
rect 12612 2645 12634 2664
rect 12644 2658 12660 2659
rect 12643 2656 12660 2658
rect 12644 2651 12660 2656
rect 12634 2644 12640 2645
rect 12643 2644 12672 2651
rect 12561 2643 12672 2644
rect 12561 2642 12678 2643
rect 12237 2634 12288 2642
rect 12335 2634 12369 2642
rect 12237 2622 12262 2634
rect 12269 2622 12288 2634
rect 12342 2632 12369 2634
rect 12378 2632 12599 2642
rect 12634 2639 12640 2642
rect 12342 2628 12599 2632
rect 12237 2614 12288 2622
rect 12335 2614 12599 2628
rect 12643 2634 12678 2642
rect 12189 2566 12208 2600
rect 12253 2606 12282 2614
rect 12253 2600 12270 2606
rect 12253 2598 12287 2600
rect 12335 2598 12351 2614
rect 12352 2604 12560 2614
rect 12561 2604 12577 2614
rect 12625 2610 12640 2625
rect 12643 2622 12644 2634
rect 12651 2622 12678 2634
rect 12643 2614 12678 2622
rect 12643 2613 12672 2614
rect 12363 2600 12577 2604
rect 12378 2598 12577 2600
rect 12612 2600 12625 2610
rect 12643 2600 12660 2613
rect 12612 2598 12660 2600
rect 12254 2594 12287 2598
rect 12250 2592 12287 2594
rect 12250 2591 12317 2592
rect 12250 2586 12281 2591
rect 12287 2586 12317 2591
rect 12250 2582 12317 2586
rect 12223 2579 12317 2582
rect 12223 2572 12272 2579
rect 12223 2566 12253 2572
rect 12272 2567 12277 2572
rect 12189 2550 12269 2566
rect 12281 2558 12317 2579
rect 12378 2574 12567 2598
rect 12612 2597 12659 2598
rect 12625 2592 12659 2597
rect 12393 2571 12567 2574
rect 12386 2568 12567 2571
rect 12595 2591 12659 2592
rect 12189 2548 12208 2550
rect 12223 2548 12257 2550
rect 12189 2532 12269 2548
rect 12189 2526 12208 2532
rect 11905 2500 12008 2510
rect 11859 2498 12008 2500
rect 12029 2498 12064 2510
rect 11698 2496 11860 2498
rect 11710 2476 11729 2496
rect 11744 2494 11774 2496
rect 11593 2468 11634 2476
rect 11716 2472 11729 2476
rect 11781 2480 11860 2496
rect 11892 2496 12064 2498
rect 11892 2480 11971 2496
rect 11978 2494 12008 2496
rect 11556 2458 11585 2468
rect 11599 2458 11628 2468
rect 11643 2458 11673 2472
rect 11716 2458 11759 2472
rect 11781 2468 11971 2480
rect 12036 2476 12042 2496
rect 11766 2458 11796 2468
rect 11797 2458 11955 2468
rect 11959 2458 11989 2468
rect 11993 2458 12023 2472
rect 12051 2458 12064 2496
rect 12136 2510 12165 2526
rect 12179 2510 12208 2526
rect 12223 2516 12253 2532
rect 12281 2510 12287 2558
rect 12290 2552 12309 2558
rect 12324 2552 12354 2560
rect 12290 2544 12354 2552
rect 12290 2528 12370 2544
rect 12386 2537 12448 2568
rect 12464 2537 12526 2568
rect 12595 2566 12644 2591
rect 12659 2566 12689 2582
rect 12558 2552 12588 2560
rect 12595 2558 12705 2566
rect 12558 2544 12603 2552
rect 12290 2526 12309 2528
rect 12324 2526 12370 2528
rect 12290 2510 12370 2526
rect 12397 2524 12432 2537
rect 12473 2534 12510 2537
rect 12473 2532 12515 2534
rect 12402 2521 12432 2524
rect 12411 2517 12418 2521
rect 12418 2516 12419 2517
rect 12377 2510 12387 2516
rect 12136 2502 12171 2510
rect 12136 2476 12137 2502
rect 12144 2476 12171 2502
rect 12079 2458 12109 2472
rect 12136 2468 12171 2476
rect 12173 2502 12214 2510
rect 12173 2476 12188 2502
rect 12195 2476 12214 2502
rect 12278 2498 12309 2510
rect 12324 2498 12427 2510
rect 12439 2500 12465 2526
rect 12480 2521 12510 2532
rect 12542 2528 12604 2544
rect 12542 2526 12588 2528
rect 12542 2510 12604 2526
rect 12616 2510 12622 2558
rect 12625 2550 12705 2558
rect 12625 2548 12644 2550
rect 12659 2548 12693 2550
rect 12625 2532 12705 2548
rect 12625 2510 12644 2532
rect 12659 2516 12689 2532
rect 12717 2526 12723 2600
rect 12726 2526 12745 2670
rect 12760 2526 12766 2670
rect 12775 2600 12788 2670
rect 12840 2666 12862 2670
rect 12833 2644 12862 2658
rect 12915 2644 12931 2658
rect 12969 2654 12975 2656
rect 12982 2654 13090 2670
rect 13097 2654 13103 2656
rect 13111 2654 13126 2670
rect 13192 2664 13211 2667
rect 12833 2642 12931 2644
rect 12958 2642 13126 2654
rect 13141 2644 13157 2658
rect 13192 2645 13214 2664
rect 13224 2658 13240 2659
rect 13223 2656 13240 2658
rect 13224 2651 13240 2656
rect 13214 2644 13220 2645
rect 13223 2644 13252 2651
rect 13141 2643 13252 2644
rect 13141 2642 13258 2643
rect 12817 2634 12868 2642
rect 12915 2634 12949 2642
rect 12817 2622 12842 2634
rect 12849 2622 12868 2634
rect 12922 2632 12949 2634
rect 12958 2632 13179 2642
rect 13214 2639 13220 2642
rect 12922 2628 13179 2632
rect 12817 2614 12868 2622
rect 12915 2614 13179 2628
rect 13223 2634 13258 2642
rect 12769 2566 12788 2600
rect 12833 2606 12862 2614
rect 12833 2600 12850 2606
rect 12833 2598 12867 2600
rect 12915 2598 12931 2614
rect 12932 2604 13140 2614
rect 13141 2604 13157 2614
rect 13205 2610 13220 2625
rect 13223 2622 13224 2634
rect 13231 2622 13258 2634
rect 13223 2614 13258 2622
rect 13223 2613 13252 2614
rect 12943 2600 13157 2604
rect 12958 2598 13157 2600
rect 13192 2600 13205 2610
rect 13223 2600 13240 2613
rect 13192 2598 13240 2600
rect 12834 2594 12867 2598
rect 12830 2592 12867 2594
rect 12830 2591 12897 2592
rect 12830 2586 12861 2591
rect 12867 2586 12897 2591
rect 12830 2582 12897 2586
rect 12803 2579 12897 2582
rect 12803 2572 12852 2579
rect 12803 2566 12833 2572
rect 12852 2567 12857 2572
rect 12769 2550 12849 2566
rect 12861 2558 12897 2579
rect 12958 2574 13147 2598
rect 13192 2597 13239 2598
rect 13205 2592 13239 2597
rect 12973 2571 13147 2574
rect 12966 2568 13147 2571
rect 13175 2591 13239 2592
rect 12769 2548 12788 2550
rect 12803 2548 12837 2550
rect 12769 2532 12849 2548
rect 12769 2526 12788 2532
rect 12485 2500 12588 2510
rect 12439 2498 12588 2500
rect 12609 2498 12644 2510
rect 12278 2496 12440 2498
rect 12290 2476 12309 2496
rect 12324 2494 12354 2496
rect 12173 2468 12214 2476
rect 12296 2472 12309 2476
rect 12361 2480 12440 2496
rect 12472 2496 12644 2498
rect 12472 2480 12551 2496
rect 12558 2494 12588 2496
rect 12136 2458 12165 2468
rect 12179 2458 12208 2468
rect 12223 2458 12253 2472
rect 12296 2458 12339 2472
rect 12361 2468 12551 2480
rect 12616 2476 12622 2496
rect 12346 2458 12376 2468
rect 12377 2458 12535 2468
rect 12539 2458 12569 2468
rect 12573 2458 12603 2472
rect 12631 2458 12644 2496
rect 12716 2510 12745 2526
rect 12759 2510 12788 2526
rect 12803 2516 12833 2532
rect 12861 2510 12867 2558
rect 12870 2552 12889 2558
rect 12904 2552 12934 2560
rect 12870 2544 12934 2552
rect 12870 2528 12950 2544
rect 12966 2537 13028 2568
rect 13044 2537 13106 2568
rect 13175 2566 13224 2591
rect 13239 2566 13269 2582
rect 13138 2552 13168 2560
rect 13175 2558 13285 2566
rect 13138 2544 13183 2552
rect 12870 2526 12889 2528
rect 12904 2526 12950 2528
rect 12870 2510 12950 2526
rect 12977 2524 13012 2537
rect 13053 2534 13090 2537
rect 13053 2532 13095 2534
rect 12982 2521 13012 2524
rect 12991 2517 12998 2521
rect 12998 2516 12999 2517
rect 12957 2510 12967 2516
rect 12716 2502 12751 2510
rect 12716 2476 12717 2502
rect 12724 2476 12751 2502
rect 12659 2458 12689 2472
rect 12716 2468 12751 2476
rect 12753 2502 12794 2510
rect 12753 2476 12768 2502
rect 12775 2476 12794 2502
rect 12858 2498 12889 2510
rect 12904 2498 13007 2510
rect 13019 2500 13045 2526
rect 13060 2521 13090 2532
rect 13122 2528 13184 2544
rect 13122 2526 13168 2528
rect 13122 2510 13184 2526
rect 13196 2510 13202 2558
rect 13205 2550 13285 2558
rect 13205 2548 13224 2550
rect 13239 2548 13273 2550
rect 13205 2532 13285 2548
rect 13205 2510 13224 2532
rect 13239 2516 13269 2532
rect 13297 2526 13303 2600
rect 13306 2526 13325 2670
rect 13340 2526 13346 2670
rect 13355 2600 13368 2670
rect 13420 2666 13442 2670
rect 13413 2644 13442 2658
rect 13495 2644 13511 2658
rect 13549 2654 13555 2656
rect 13562 2654 13670 2670
rect 13677 2654 13683 2656
rect 13691 2654 13706 2670
rect 13772 2664 13791 2667
rect 13413 2642 13511 2644
rect 13538 2642 13706 2654
rect 13721 2644 13737 2658
rect 13772 2645 13794 2664
rect 13804 2658 13820 2659
rect 13803 2656 13820 2658
rect 13804 2651 13820 2656
rect 13794 2644 13800 2645
rect 13803 2644 13832 2651
rect 13721 2643 13832 2644
rect 13721 2642 13838 2643
rect 13397 2634 13448 2642
rect 13495 2634 13529 2642
rect 13397 2622 13422 2634
rect 13429 2622 13448 2634
rect 13502 2632 13529 2634
rect 13538 2632 13759 2642
rect 13794 2639 13800 2642
rect 13502 2628 13759 2632
rect 13397 2614 13448 2622
rect 13495 2614 13759 2628
rect 13803 2634 13838 2642
rect 13349 2566 13368 2600
rect 13413 2606 13442 2614
rect 13413 2600 13430 2606
rect 13413 2598 13447 2600
rect 13495 2598 13511 2614
rect 13512 2604 13720 2614
rect 13721 2604 13737 2614
rect 13785 2610 13800 2625
rect 13803 2622 13804 2634
rect 13811 2622 13838 2634
rect 13803 2614 13838 2622
rect 13803 2613 13832 2614
rect 13523 2600 13737 2604
rect 13538 2598 13737 2600
rect 13772 2600 13785 2610
rect 13803 2600 13820 2613
rect 13772 2598 13820 2600
rect 13414 2594 13447 2598
rect 13410 2592 13447 2594
rect 13410 2591 13477 2592
rect 13410 2586 13441 2591
rect 13447 2586 13477 2591
rect 13410 2582 13477 2586
rect 13383 2579 13477 2582
rect 13383 2572 13432 2579
rect 13383 2566 13413 2572
rect 13432 2567 13437 2572
rect 13349 2550 13429 2566
rect 13441 2558 13477 2579
rect 13538 2574 13727 2598
rect 13772 2597 13819 2598
rect 13785 2592 13819 2597
rect 13553 2571 13727 2574
rect 13546 2568 13727 2571
rect 13755 2591 13819 2592
rect 13349 2548 13368 2550
rect 13383 2548 13417 2550
rect 13349 2532 13429 2548
rect 13349 2526 13368 2532
rect 13065 2500 13168 2510
rect 13019 2498 13168 2500
rect 13189 2498 13224 2510
rect 12858 2496 13020 2498
rect 12870 2476 12889 2496
rect 12904 2494 12934 2496
rect 12753 2468 12794 2476
rect 12876 2472 12889 2476
rect 12941 2480 13020 2496
rect 13052 2496 13224 2498
rect 13052 2480 13131 2496
rect 13138 2494 13168 2496
rect 12716 2458 12745 2468
rect 12759 2458 12788 2468
rect 12803 2458 12833 2472
rect 12876 2458 12919 2472
rect 12941 2468 13131 2480
rect 13196 2476 13202 2496
rect 12926 2458 12956 2468
rect 12957 2458 13115 2468
rect 13119 2458 13149 2468
rect 13153 2458 13183 2472
rect 13211 2458 13224 2496
rect 13296 2510 13325 2526
rect 13339 2510 13368 2526
rect 13383 2516 13413 2532
rect 13441 2510 13447 2558
rect 13450 2552 13469 2558
rect 13484 2552 13514 2560
rect 13450 2544 13514 2552
rect 13450 2528 13530 2544
rect 13546 2537 13608 2568
rect 13624 2537 13686 2568
rect 13755 2566 13804 2591
rect 13819 2566 13849 2582
rect 13718 2552 13748 2560
rect 13755 2558 13865 2566
rect 13718 2544 13763 2552
rect 13450 2526 13469 2528
rect 13484 2526 13530 2528
rect 13450 2510 13530 2526
rect 13557 2524 13592 2537
rect 13633 2534 13670 2537
rect 13633 2532 13675 2534
rect 13562 2521 13592 2524
rect 13571 2517 13578 2521
rect 13578 2516 13579 2517
rect 13537 2510 13547 2516
rect 13296 2502 13331 2510
rect 13296 2476 13297 2502
rect 13304 2476 13331 2502
rect 13239 2458 13269 2472
rect 13296 2468 13331 2476
rect 13333 2502 13374 2510
rect 13333 2476 13348 2502
rect 13355 2476 13374 2502
rect 13438 2498 13469 2510
rect 13484 2498 13587 2510
rect 13599 2500 13625 2526
rect 13640 2521 13670 2532
rect 13702 2528 13764 2544
rect 13702 2526 13748 2528
rect 13702 2510 13764 2526
rect 13776 2510 13782 2558
rect 13785 2550 13865 2558
rect 13785 2548 13804 2550
rect 13819 2548 13853 2550
rect 13785 2532 13865 2548
rect 13785 2510 13804 2532
rect 13819 2516 13849 2532
rect 13877 2526 13883 2600
rect 13886 2526 13905 2670
rect 13920 2526 13926 2670
rect 13935 2600 13948 2670
rect 14000 2666 14022 2670
rect 13993 2644 14022 2658
rect 14075 2644 14091 2658
rect 14129 2654 14135 2656
rect 14142 2654 14250 2670
rect 14257 2654 14263 2656
rect 14271 2654 14286 2670
rect 14352 2664 14371 2667
rect 13993 2642 14091 2644
rect 14118 2642 14286 2654
rect 14301 2644 14317 2658
rect 14352 2645 14374 2664
rect 14384 2658 14400 2659
rect 14383 2656 14400 2658
rect 14384 2651 14400 2656
rect 14374 2644 14380 2645
rect 14383 2644 14412 2651
rect 14301 2643 14412 2644
rect 14301 2642 14418 2643
rect 13977 2634 14028 2642
rect 14075 2634 14109 2642
rect 13977 2622 14002 2634
rect 14009 2622 14028 2634
rect 14082 2632 14109 2634
rect 14118 2632 14339 2642
rect 14374 2639 14380 2642
rect 14082 2628 14339 2632
rect 13977 2614 14028 2622
rect 14075 2614 14339 2628
rect 14383 2634 14418 2642
rect 13929 2566 13948 2600
rect 13993 2606 14022 2614
rect 13993 2600 14010 2606
rect 13993 2598 14027 2600
rect 14075 2598 14091 2614
rect 14092 2604 14300 2614
rect 14301 2604 14317 2614
rect 14365 2610 14380 2625
rect 14383 2622 14384 2634
rect 14391 2622 14418 2634
rect 14383 2614 14418 2622
rect 14383 2613 14412 2614
rect 14103 2600 14317 2604
rect 14118 2598 14317 2600
rect 14352 2600 14365 2610
rect 14383 2600 14400 2613
rect 14352 2598 14400 2600
rect 13994 2594 14027 2598
rect 13990 2592 14027 2594
rect 13990 2591 14057 2592
rect 13990 2586 14021 2591
rect 14027 2586 14057 2591
rect 13990 2582 14057 2586
rect 13963 2579 14057 2582
rect 13963 2572 14012 2579
rect 13963 2566 13993 2572
rect 14012 2567 14017 2572
rect 13929 2550 14009 2566
rect 14021 2558 14057 2579
rect 14118 2574 14307 2598
rect 14352 2597 14399 2598
rect 14365 2592 14399 2597
rect 14133 2571 14307 2574
rect 14126 2568 14307 2571
rect 14335 2591 14399 2592
rect 13929 2548 13948 2550
rect 13963 2548 13997 2550
rect 13929 2532 14009 2548
rect 13929 2526 13948 2532
rect 13645 2500 13748 2510
rect 13599 2498 13748 2500
rect 13769 2498 13804 2510
rect 13438 2496 13600 2498
rect 13450 2476 13469 2496
rect 13484 2494 13514 2496
rect 13333 2468 13374 2476
rect 13456 2472 13469 2476
rect 13521 2480 13600 2496
rect 13632 2496 13804 2498
rect 13632 2480 13711 2496
rect 13718 2494 13748 2496
rect 13296 2458 13325 2468
rect 13339 2458 13368 2468
rect 13383 2458 13413 2472
rect 13456 2458 13499 2472
rect 13521 2468 13711 2480
rect 13776 2476 13782 2496
rect 13506 2458 13536 2468
rect 13537 2458 13695 2468
rect 13699 2458 13729 2468
rect 13733 2458 13763 2472
rect 13791 2458 13804 2496
rect 13876 2510 13905 2526
rect 13919 2510 13948 2526
rect 13963 2516 13993 2532
rect 14021 2510 14027 2558
rect 14030 2552 14049 2558
rect 14064 2552 14094 2560
rect 14030 2544 14094 2552
rect 14030 2528 14110 2544
rect 14126 2537 14188 2568
rect 14204 2537 14266 2568
rect 14335 2566 14384 2591
rect 14399 2566 14429 2582
rect 14298 2552 14328 2560
rect 14335 2558 14445 2566
rect 14298 2544 14343 2552
rect 14030 2526 14049 2528
rect 14064 2526 14110 2528
rect 14030 2510 14110 2526
rect 14137 2524 14172 2537
rect 14213 2534 14250 2537
rect 14213 2532 14255 2534
rect 14142 2521 14172 2524
rect 14151 2517 14158 2521
rect 14158 2516 14159 2517
rect 14117 2510 14127 2516
rect 13876 2502 13911 2510
rect 13876 2476 13877 2502
rect 13884 2476 13911 2502
rect 13819 2458 13849 2472
rect 13876 2468 13911 2476
rect 13913 2502 13954 2510
rect 13913 2476 13928 2502
rect 13935 2476 13954 2502
rect 14018 2498 14049 2510
rect 14064 2498 14167 2510
rect 14179 2500 14205 2526
rect 14220 2521 14250 2532
rect 14282 2528 14344 2544
rect 14282 2526 14328 2528
rect 14282 2510 14344 2526
rect 14356 2510 14362 2558
rect 14365 2550 14445 2558
rect 14365 2548 14384 2550
rect 14399 2548 14433 2550
rect 14365 2532 14445 2548
rect 14365 2510 14384 2532
rect 14399 2516 14429 2532
rect 14457 2526 14463 2600
rect 14466 2526 14485 2670
rect 14500 2526 14506 2670
rect 14515 2600 14528 2670
rect 14580 2666 14602 2670
rect 14573 2644 14602 2658
rect 14655 2644 14671 2658
rect 14709 2654 14715 2656
rect 14722 2654 14830 2670
rect 14837 2654 14843 2656
rect 14851 2654 14866 2670
rect 14932 2664 14951 2667
rect 14573 2642 14671 2644
rect 14698 2642 14866 2654
rect 14881 2644 14897 2658
rect 14932 2645 14954 2664
rect 14964 2658 14980 2659
rect 14963 2656 14980 2658
rect 14964 2651 14980 2656
rect 14954 2644 14960 2645
rect 14963 2644 14992 2651
rect 14881 2643 14992 2644
rect 14881 2642 14998 2643
rect 14557 2634 14608 2642
rect 14655 2634 14689 2642
rect 14557 2622 14582 2634
rect 14589 2622 14608 2634
rect 14662 2632 14689 2634
rect 14698 2632 14919 2642
rect 14954 2639 14960 2642
rect 14662 2628 14919 2632
rect 14557 2614 14608 2622
rect 14655 2614 14919 2628
rect 14963 2634 14998 2642
rect 14509 2566 14528 2600
rect 14573 2606 14602 2614
rect 14573 2600 14590 2606
rect 14573 2598 14607 2600
rect 14655 2598 14671 2614
rect 14672 2604 14880 2614
rect 14881 2604 14897 2614
rect 14945 2610 14960 2625
rect 14963 2622 14964 2634
rect 14971 2622 14998 2634
rect 14963 2614 14998 2622
rect 14963 2613 14992 2614
rect 14683 2600 14897 2604
rect 14698 2598 14897 2600
rect 14932 2600 14945 2610
rect 14963 2600 14980 2613
rect 14932 2598 14980 2600
rect 14574 2594 14607 2598
rect 14570 2592 14607 2594
rect 14570 2591 14637 2592
rect 14570 2586 14601 2591
rect 14607 2586 14637 2591
rect 14570 2582 14637 2586
rect 14543 2579 14637 2582
rect 14543 2572 14592 2579
rect 14543 2566 14573 2572
rect 14592 2567 14597 2572
rect 14509 2550 14589 2566
rect 14601 2558 14637 2579
rect 14698 2574 14887 2598
rect 14932 2597 14979 2598
rect 14945 2592 14979 2597
rect 14713 2571 14887 2574
rect 14706 2568 14887 2571
rect 14915 2591 14979 2592
rect 14509 2548 14528 2550
rect 14543 2548 14577 2550
rect 14509 2532 14589 2548
rect 14509 2526 14528 2532
rect 14225 2500 14328 2510
rect 14179 2498 14328 2500
rect 14349 2498 14384 2510
rect 14018 2496 14180 2498
rect 14030 2476 14049 2496
rect 14064 2494 14094 2496
rect 13913 2468 13954 2476
rect 14036 2472 14049 2476
rect 14101 2480 14180 2496
rect 14212 2496 14384 2498
rect 14212 2480 14291 2496
rect 14298 2494 14328 2496
rect 13876 2458 13905 2468
rect 13919 2458 13948 2468
rect 13963 2458 13993 2472
rect 14036 2458 14079 2472
rect 14101 2468 14291 2480
rect 14356 2476 14362 2496
rect 14086 2458 14116 2468
rect 14117 2458 14275 2468
rect 14279 2458 14309 2468
rect 14313 2458 14343 2472
rect 14371 2458 14384 2496
rect 14456 2510 14485 2526
rect 14499 2510 14528 2526
rect 14543 2516 14573 2532
rect 14601 2510 14607 2558
rect 14610 2552 14629 2558
rect 14644 2552 14674 2560
rect 14610 2544 14674 2552
rect 14610 2528 14690 2544
rect 14706 2537 14768 2568
rect 14784 2537 14846 2568
rect 14915 2566 14964 2591
rect 14979 2566 15009 2582
rect 14878 2552 14908 2560
rect 14915 2558 15025 2566
rect 14878 2544 14923 2552
rect 14610 2526 14629 2528
rect 14644 2526 14690 2528
rect 14610 2510 14690 2526
rect 14717 2524 14752 2537
rect 14793 2534 14830 2537
rect 14793 2532 14835 2534
rect 14722 2521 14752 2524
rect 14731 2517 14738 2521
rect 14738 2516 14739 2517
rect 14697 2510 14707 2516
rect 14456 2502 14491 2510
rect 14456 2476 14457 2502
rect 14464 2476 14491 2502
rect 14399 2458 14429 2472
rect 14456 2468 14491 2476
rect 14493 2502 14534 2510
rect 14493 2476 14508 2502
rect 14515 2476 14534 2502
rect 14598 2498 14629 2510
rect 14644 2498 14747 2510
rect 14759 2500 14785 2526
rect 14800 2521 14830 2532
rect 14862 2528 14924 2544
rect 14862 2526 14908 2528
rect 14862 2510 14924 2526
rect 14936 2510 14942 2558
rect 14945 2550 15025 2558
rect 14945 2548 14964 2550
rect 14979 2548 15013 2550
rect 14945 2532 15025 2548
rect 14945 2510 14964 2532
rect 14979 2516 15009 2532
rect 15037 2526 15043 2600
rect 15046 2526 15065 2670
rect 15080 2526 15086 2670
rect 15095 2600 15108 2670
rect 15160 2666 15182 2670
rect 15153 2644 15182 2658
rect 15235 2644 15251 2658
rect 15289 2654 15295 2656
rect 15302 2654 15410 2670
rect 15417 2654 15423 2656
rect 15431 2654 15446 2670
rect 15512 2664 15531 2667
rect 15153 2642 15251 2644
rect 15278 2642 15446 2654
rect 15461 2644 15477 2658
rect 15512 2645 15534 2664
rect 15544 2658 15560 2659
rect 15543 2656 15560 2658
rect 15544 2651 15560 2656
rect 15534 2644 15540 2645
rect 15543 2644 15572 2651
rect 15461 2643 15572 2644
rect 15461 2642 15578 2643
rect 15137 2634 15188 2642
rect 15235 2634 15269 2642
rect 15137 2622 15162 2634
rect 15169 2622 15188 2634
rect 15242 2632 15269 2634
rect 15278 2632 15499 2642
rect 15534 2639 15540 2642
rect 15242 2628 15499 2632
rect 15137 2614 15188 2622
rect 15235 2614 15499 2628
rect 15543 2634 15578 2642
rect 15089 2566 15108 2600
rect 15153 2606 15182 2614
rect 15153 2600 15170 2606
rect 15153 2598 15187 2600
rect 15235 2598 15251 2614
rect 15252 2604 15460 2614
rect 15461 2604 15477 2614
rect 15525 2610 15540 2625
rect 15543 2622 15544 2634
rect 15551 2622 15578 2634
rect 15543 2614 15578 2622
rect 15543 2613 15572 2614
rect 15263 2600 15477 2604
rect 15278 2598 15477 2600
rect 15512 2600 15525 2610
rect 15543 2600 15560 2613
rect 15512 2598 15560 2600
rect 15154 2594 15187 2598
rect 15150 2592 15187 2594
rect 15150 2591 15217 2592
rect 15150 2586 15181 2591
rect 15187 2586 15217 2591
rect 15150 2582 15217 2586
rect 15123 2579 15217 2582
rect 15123 2572 15172 2579
rect 15123 2566 15153 2572
rect 15172 2567 15177 2572
rect 15089 2550 15169 2566
rect 15181 2558 15217 2579
rect 15278 2574 15467 2598
rect 15512 2597 15559 2598
rect 15525 2592 15559 2597
rect 15293 2571 15467 2574
rect 15286 2568 15467 2571
rect 15495 2591 15559 2592
rect 15089 2548 15108 2550
rect 15123 2548 15157 2550
rect 15089 2532 15169 2548
rect 15089 2526 15108 2532
rect 14805 2500 14908 2510
rect 14759 2498 14908 2500
rect 14929 2498 14964 2510
rect 14598 2496 14760 2498
rect 14610 2476 14629 2496
rect 14644 2494 14674 2496
rect 14493 2468 14534 2476
rect 14616 2472 14629 2476
rect 14681 2480 14760 2496
rect 14792 2496 14964 2498
rect 14792 2480 14871 2496
rect 14878 2494 14908 2496
rect 14456 2458 14485 2468
rect 14499 2458 14528 2468
rect 14543 2458 14573 2472
rect 14616 2458 14659 2472
rect 14681 2468 14871 2480
rect 14936 2476 14942 2496
rect 14666 2458 14696 2468
rect 14697 2458 14855 2468
rect 14859 2458 14889 2468
rect 14893 2458 14923 2472
rect 14951 2458 14964 2496
rect 15036 2510 15065 2526
rect 15079 2510 15108 2526
rect 15123 2516 15153 2532
rect 15181 2510 15187 2558
rect 15190 2552 15209 2558
rect 15224 2552 15254 2560
rect 15190 2544 15254 2552
rect 15190 2528 15270 2544
rect 15286 2537 15348 2568
rect 15364 2537 15426 2568
rect 15495 2566 15544 2591
rect 15559 2566 15589 2582
rect 15458 2552 15488 2560
rect 15495 2558 15605 2566
rect 15458 2544 15503 2552
rect 15190 2526 15209 2528
rect 15224 2526 15270 2528
rect 15190 2510 15270 2526
rect 15297 2524 15332 2537
rect 15373 2534 15410 2537
rect 15373 2532 15415 2534
rect 15302 2521 15332 2524
rect 15311 2517 15318 2521
rect 15318 2516 15319 2517
rect 15277 2510 15287 2516
rect 15036 2502 15071 2510
rect 15036 2476 15037 2502
rect 15044 2476 15071 2502
rect 14979 2458 15009 2472
rect 15036 2468 15071 2476
rect 15073 2502 15114 2510
rect 15073 2476 15088 2502
rect 15095 2476 15114 2502
rect 15178 2498 15209 2510
rect 15224 2498 15327 2510
rect 15339 2500 15365 2526
rect 15380 2521 15410 2532
rect 15442 2528 15504 2544
rect 15442 2526 15488 2528
rect 15442 2510 15504 2526
rect 15516 2510 15522 2558
rect 15525 2550 15605 2558
rect 15525 2548 15544 2550
rect 15559 2548 15593 2550
rect 15525 2532 15605 2548
rect 15525 2510 15544 2532
rect 15559 2516 15589 2532
rect 15617 2526 15623 2600
rect 15626 2526 15645 2670
rect 15660 2526 15666 2670
rect 15675 2600 15688 2670
rect 15740 2666 15762 2670
rect 15733 2644 15762 2658
rect 15815 2644 15831 2658
rect 15869 2654 15875 2656
rect 15882 2654 15990 2670
rect 15997 2654 16003 2656
rect 16011 2654 16026 2670
rect 16092 2664 16111 2667
rect 15733 2642 15831 2644
rect 15858 2642 16026 2654
rect 16041 2644 16057 2658
rect 16092 2645 16114 2664
rect 16124 2658 16140 2659
rect 16123 2656 16140 2658
rect 16124 2651 16140 2656
rect 16114 2644 16120 2645
rect 16123 2644 16152 2651
rect 16041 2643 16152 2644
rect 16041 2642 16158 2643
rect 15717 2634 15768 2642
rect 15815 2634 15849 2642
rect 15717 2622 15742 2634
rect 15749 2622 15768 2634
rect 15822 2632 15849 2634
rect 15858 2632 16079 2642
rect 16114 2639 16120 2642
rect 15822 2628 16079 2632
rect 15717 2614 15768 2622
rect 15815 2614 16079 2628
rect 16123 2634 16158 2642
rect 15669 2566 15688 2600
rect 15733 2606 15762 2614
rect 15733 2600 15750 2606
rect 15733 2598 15767 2600
rect 15815 2598 15831 2614
rect 15832 2604 16040 2614
rect 16041 2604 16057 2614
rect 16105 2610 16120 2625
rect 16123 2622 16124 2634
rect 16131 2622 16158 2634
rect 16123 2614 16158 2622
rect 16123 2613 16152 2614
rect 15843 2600 16057 2604
rect 15858 2598 16057 2600
rect 16092 2600 16105 2610
rect 16123 2600 16140 2613
rect 16092 2598 16140 2600
rect 15734 2594 15767 2598
rect 15730 2592 15767 2594
rect 15730 2591 15797 2592
rect 15730 2586 15761 2591
rect 15767 2586 15797 2591
rect 15730 2582 15797 2586
rect 15703 2579 15797 2582
rect 15703 2572 15752 2579
rect 15703 2566 15733 2572
rect 15752 2567 15757 2572
rect 15669 2550 15749 2566
rect 15761 2558 15797 2579
rect 15858 2574 16047 2598
rect 16092 2597 16139 2598
rect 16105 2592 16139 2597
rect 15873 2571 16047 2574
rect 15866 2568 16047 2571
rect 16075 2591 16139 2592
rect 15669 2548 15688 2550
rect 15703 2548 15737 2550
rect 15669 2532 15749 2548
rect 15669 2526 15688 2532
rect 15385 2500 15488 2510
rect 15339 2498 15488 2500
rect 15509 2498 15544 2510
rect 15178 2496 15340 2498
rect 15190 2476 15209 2496
rect 15224 2494 15254 2496
rect 15073 2468 15114 2476
rect 15196 2472 15209 2476
rect 15261 2480 15340 2496
rect 15372 2496 15544 2498
rect 15372 2480 15451 2496
rect 15458 2494 15488 2496
rect 15036 2458 15065 2468
rect 15079 2458 15108 2468
rect 15123 2458 15153 2472
rect 15196 2458 15239 2472
rect 15261 2468 15451 2480
rect 15516 2476 15522 2496
rect 15246 2458 15276 2468
rect 15277 2458 15435 2468
rect 15439 2458 15469 2468
rect 15473 2458 15503 2472
rect 15531 2458 15544 2496
rect 15616 2510 15645 2526
rect 15659 2510 15688 2526
rect 15703 2516 15733 2532
rect 15761 2510 15767 2558
rect 15770 2552 15789 2558
rect 15804 2552 15834 2560
rect 15770 2544 15834 2552
rect 15770 2528 15850 2544
rect 15866 2537 15928 2568
rect 15944 2537 16006 2568
rect 16075 2566 16124 2591
rect 16139 2566 16169 2582
rect 16038 2552 16068 2560
rect 16075 2558 16185 2566
rect 16038 2544 16083 2552
rect 15770 2526 15789 2528
rect 15804 2526 15850 2528
rect 15770 2510 15850 2526
rect 15877 2524 15912 2537
rect 15953 2534 15990 2537
rect 15953 2532 15995 2534
rect 15882 2521 15912 2524
rect 15891 2517 15898 2521
rect 15898 2516 15899 2517
rect 15857 2510 15867 2516
rect 15616 2502 15651 2510
rect 15616 2476 15617 2502
rect 15624 2476 15651 2502
rect 15559 2458 15589 2472
rect 15616 2468 15651 2476
rect 15653 2502 15694 2510
rect 15653 2476 15668 2502
rect 15675 2476 15694 2502
rect 15758 2498 15789 2510
rect 15804 2498 15907 2510
rect 15919 2500 15945 2526
rect 15960 2521 15990 2532
rect 16022 2528 16084 2544
rect 16022 2526 16068 2528
rect 16022 2510 16084 2526
rect 16096 2510 16102 2558
rect 16105 2550 16185 2558
rect 16105 2548 16124 2550
rect 16139 2548 16173 2550
rect 16105 2532 16185 2548
rect 16105 2510 16124 2532
rect 16139 2516 16169 2532
rect 16197 2526 16203 2600
rect 16206 2526 16225 2670
rect 16240 2526 16246 2670
rect 16255 2600 16268 2670
rect 16320 2666 16342 2670
rect 16313 2644 16342 2658
rect 16395 2644 16411 2658
rect 16449 2654 16455 2656
rect 16462 2654 16570 2670
rect 16577 2654 16583 2656
rect 16591 2654 16606 2670
rect 16672 2664 16691 2667
rect 16313 2642 16411 2644
rect 16438 2642 16606 2654
rect 16621 2644 16637 2658
rect 16672 2645 16694 2664
rect 16704 2658 16720 2659
rect 16703 2656 16720 2658
rect 16704 2651 16720 2656
rect 16694 2644 16700 2645
rect 16703 2644 16732 2651
rect 16621 2643 16732 2644
rect 16621 2642 16738 2643
rect 16297 2634 16348 2642
rect 16395 2634 16429 2642
rect 16297 2622 16322 2634
rect 16329 2622 16348 2634
rect 16402 2632 16429 2634
rect 16438 2632 16659 2642
rect 16694 2639 16700 2642
rect 16402 2628 16659 2632
rect 16297 2614 16348 2622
rect 16395 2614 16659 2628
rect 16703 2634 16738 2642
rect 16249 2566 16268 2600
rect 16313 2606 16342 2614
rect 16313 2600 16330 2606
rect 16313 2598 16347 2600
rect 16395 2598 16411 2614
rect 16412 2604 16620 2614
rect 16621 2604 16637 2614
rect 16685 2610 16700 2625
rect 16703 2622 16704 2634
rect 16711 2622 16738 2634
rect 16703 2614 16738 2622
rect 16703 2613 16732 2614
rect 16423 2600 16637 2604
rect 16438 2598 16637 2600
rect 16672 2600 16685 2610
rect 16703 2600 16720 2613
rect 16672 2598 16720 2600
rect 16314 2594 16347 2598
rect 16310 2592 16347 2594
rect 16310 2591 16377 2592
rect 16310 2586 16341 2591
rect 16347 2586 16377 2591
rect 16310 2582 16377 2586
rect 16283 2579 16377 2582
rect 16283 2572 16332 2579
rect 16283 2566 16313 2572
rect 16332 2567 16337 2572
rect 16249 2550 16329 2566
rect 16341 2558 16377 2579
rect 16438 2574 16627 2598
rect 16672 2597 16719 2598
rect 16685 2592 16719 2597
rect 16453 2571 16627 2574
rect 16446 2568 16627 2571
rect 16655 2591 16719 2592
rect 16249 2548 16268 2550
rect 16283 2548 16317 2550
rect 16249 2532 16329 2548
rect 16249 2526 16268 2532
rect 15965 2500 16068 2510
rect 15919 2498 16068 2500
rect 16089 2498 16124 2510
rect 15758 2496 15920 2498
rect 15770 2476 15789 2496
rect 15804 2494 15834 2496
rect 15653 2468 15694 2476
rect 15776 2472 15789 2476
rect 15841 2480 15920 2496
rect 15952 2496 16124 2498
rect 15952 2480 16031 2496
rect 16038 2494 16068 2496
rect 15616 2458 15645 2468
rect 15659 2458 15688 2468
rect 15703 2458 15733 2472
rect 15776 2458 15819 2472
rect 15841 2468 16031 2480
rect 16096 2476 16102 2496
rect 15826 2458 15856 2468
rect 15857 2458 16015 2468
rect 16019 2458 16049 2468
rect 16053 2458 16083 2472
rect 16111 2458 16124 2496
rect 16196 2510 16225 2526
rect 16239 2510 16268 2526
rect 16283 2516 16313 2532
rect 16341 2510 16347 2558
rect 16350 2552 16369 2558
rect 16384 2552 16414 2560
rect 16350 2544 16414 2552
rect 16350 2528 16430 2544
rect 16446 2537 16508 2568
rect 16524 2537 16586 2568
rect 16655 2566 16704 2591
rect 16719 2566 16749 2582
rect 16618 2552 16648 2560
rect 16655 2558 16765 2566
rect 16618 2544 16663 2552
rect 16350 2526 16369 2528
rect 16384 2526 16430 2528
rect 16350 2510 16430 2526
rect 16457 2524 16492 2537
rect 16533 2534 16570 2537
rect 16533 2532 16575 2534
rect 16462 2521 16492 2524
rect 16471 2517 16478 2521
rect 16478 2516 16479 2517
rect 16437 2510 16447 2516
rect 16196 2502 16231 2510
rect 16196 2476 16197 2502
rect 16204 2476 16231 2502
rect 16139 2458 16169 2472
rect 16196 2468 16231 2476
rect 16233 2502 16274 2510
rect 16233 2476 16248 2502
rect 16255 2476 16274 2502
rect 16338 2498 16369 2510
rect 16384 2498 16487 2510
rect 16499 2500 16525 2526
rect 16540 2521 16570 2532
rect 16602 2528 16664 2544
rect 16602 2526 16648 2528
rect 16602 2510 16664 2526
rect 16676 2510 16682 2558
rect 16685 2550 16765 2558
rect 16685 2548 16704 2550
rect 16719 2548 16753 2550
rect 16685 2532 16765 2548
rect 16685 2510 16704 2532
rect 16719 2516 16749 2532
rect 16777 2526 16783 2600
rect 16786 2526 16805 2670
rect 16820 2526 16826 2670
rect 16835 2600 16848 2670
rect 16900 2666 16922 2670
rect 16893 2644 16922 2658
rect 16975 2644 16991 2658
rect 17029 2654 17035 2656
rect 17042 2654 17150 2670
rect 17157 2654 17163 2656
rect 17171 2654 17186 2670
rect 17252 2664 17271 2667
rect 16893 2642 16991 2644
rect 17018 2642 17186 2654
rect 17201 2644 17217 2658
rect 17252 2645 17274 2664
rect 17284 2658 17300 2659
rect 17283 2656 17300 2658
rect 17284 2651 17300 2656
rect 17274 2644 17280 2645
rect 17283 2644 17312 2651
rect 17201 2643 17312 2644
rect 17201 2642 17318 2643
rect 16877 2634 16928 2642
rect 16975 2634 17009 2642
rect 16877 2622 16902 2634
rect 16909 2622 16928 2634
rect 16982 2632 17009 2634
rect 17018 2632 17239 2642
rect 17274 2639 17280 2642
rect 16982 2628 17239 2632
rect 16877 2614 16928 2622
rect 16975 2614 17239 2628
rect 17283 2634 17318 2642
rect 16829 2566 16848 2600
rect 16893 2606 16922 2614
rect 16893 2600 16910 2606
rect 16893 2598 16927 2600
rect 16975 2598 16991 2614
rect 16992 2604 17200 2614
rect 17201 2604 17217 2614
rect 17265 2610 17280 2625
rect 17283 2622 17284 2634
rect 17291 2622 17318 2634
rect 17283 2614 17318 2622
rect 17283 2613 17312 2614
rect 17003 2600 17217 2604
rect 17018 2598 17217 2600
rect 17252 2600 17265 2610
rect 17283 2600 17300 2613
rect 17252 2598 17300 2600
rect 16894 2594 16927 2598
rect 16890 2592 16927 2594
rect 16890 2591 16957 2592
rect 16890 2586 16921 2591
rect 16927 2586 16957 2591
rect 16890 2582 16957 2586
rect 16863 2579 16957 2582
rect 16863 2572 16912 2579
rect 16863 2566 16893 2572
rect 16912 2567 16917 2572
rect 16829 2550 16909 2566
rect 16921 2558 16957 2579
rect 17018 2574 17207 2598
rect 17252 2597 17299 2598
rect 17265 2592 17299 2597
rect 17033 2571 17207 2574
rect 17026 2568 17207 2571
rect 17235 2591 17299 2592
rect 16829 2548 16848 2550
rect 16863 2548 16897 2550
rect 16829 2532 16909 2548
rect 16829 2526 16848 2532
rect 16545 2500 16648 2510
rect 16499 2498 16648 2500
rect 16669 2498 16704 2510
rect 16338 2496 16500 2498
rect 16350 2476 16369 2496
rect 16384 2494 16414 2496
rect 16233 2468 16274 2476
rect 16356 2472 16369 2476
rect 16421 2480 16500 2496
rect 16532 2496 16704 2498
rect 16532 2480 16611 2496
rect 16618 2494 16648 2496
rect 16196 2458 16225 2468
rect 16239 2458 16268 2468
rect 16283 2458 16313 2472
rect 16356 2458 16399 2472
rect 16421 2468 16611 2480
rect 16676 2476 16682 2496
rect 16406 2458 16436 2468
rect 16437 2458 16595 2468
rect 16599 2458 16629 2468
rect 16633 2458 16663 2472
rect 16691 2458 16704 2496
rect 16776 2510 16805 2526
rect 16819 2510 16848 2526
rect 16863 2516 16893 2532
rect 16921 2510 16927 2558
rect 16930 2552 16949 2558
rect 16964 2552 16994 2560
rect 16930 2544 16994 2552
rect 16930 2528 17010 2544
rect 17026 2537 17088 2568
rect 17104 2537 17166 2568
rect 17235 2566 17284 2591
rect 17299 2566 17329 2582
rect 17198 2552 17228 2560
rect 17235 2558 17345 2566
rect 17198 2544 17243 2552
rect 16930 2526 16949 2528
rect 16964 2526 17010 2528
rect 16930 2510 17010 2526
rect 17037 2524 17072 2537
rect 17113 2534 17150 2537
rect 17113 2532 17155 2534
rect 17042 2521 17072 2524
rect 17051 2517 17058 2521
rect 17058 2516 17059 2517
rect 17017 2510 17027 2516
rect 16776 2502 16811 2510
rect 16776 2476 16777 2502
rect 16784 2476 16811 2502
rect 16719 2458 16749 2472
rect 16776 2468 16811 2476
rect 16813 2502 16854 2510
rect 16813 2476 16828 2502
rect 16835 2476 16854 2502
rect 16918 2498 16949 2510
rect 16964 2498 17067 2510
rect 17079 2500 17105 2526
rect 17120 2521 17150 2532
rect 17182 2528 17244 2544
rect 17182 2526 17228 2528
rect 17182 2510 17244 2526
rect 17256 2510 17262 2558
rect 17265 2550 17345 2558
rect 17265 2548 17284 2550
rect 17299 2548 17333 2550
rect 17265 2532 17345 2548
rect 17265 2510 17284 2532
rect 17299 2516 17329 2532
rect 17357 2526 17363 2600
rect 17366 2526 17385 2670
rect 17400 2526 17406 2670
rect 17415 2600 17428 2670
rect 17480 2666 17502 2670
rect 17473 2644 17502 2658
rect 17555 2644 17571 2658
rect 17609 2654 17615 2656
rect 17622 2654 17730 2670
rect 17737 2654 17743 2656
rect 17751 2654 17766 2670
rect 17832 2664 17851 2667
rect 17473 2642 17571 2644
rect 17598 2642 17766 2654
rect 17781 2644 17797 2658
rect 17832 2645 17854 2664
rect 17864 2658 17880 2659
rect 17863 2656 17880 2658
rect 17864 2651 17880 2656
rect 17854 2644 17860 2645
rect 17863 2644 17892 2651
rect 17781 2643 17892 2644
rect 17781 2642 17898 2643
rect 17457 2634 17508 2642
rect 17555 2634 17589 2642
rect 17457 2622 17482 2634
rect 17489 2622 17508 2634
rect 17562 2632 17589 2634
rect 17598 2632 17819 2642
rect 17854 2639 17860 2642
rect 17562 2628 17819 2632
rect 17457 2614 17508 2622
rect 17555 2614 17819 2628
rect 17863 2634 17898 2642
rect 17409 2566 17428 2600
rect 17473 2606 17502 2614
rect 17473 2600 17490 2606
rect 17473 2598 17507 2600
rect 17555 2598 17571 2614
rect 17572 2604 17780 2614
rect 17781 2604 17797 2614
rect 17845 2610 17860 2625
rect 17863 2622 17864 2634
rect 17871 2622 17898 2634
rect 17863 2614 17898 2622
rect 17863 2613 17892 2614
rect 17583 2600 17797 2604
rect 17598 2598 17797 2600
rect 17832 2600 17845 2610
rect 17863 2600 17880 2613
rect 17832 2598 17880 2600
rect 17474 2594 17507 2598
rect 17470 2592 17507 2594
rect 17470 2591 17537 2592
rect 17470 2586 17501 2591
rect 17507 2586 17537 2591
rect 17470 2582 17537 2586
rect 17443 2579 17537 2582
rect 17443 2572 17492 2579
rect 17443 2566 17473 2572
rect 17492 2567 17497 2572
rect 17409 2550 17489 2566
rect 17501 2558 17537 2579
rect 17598 2574 17787 2598
rect 17832 2597 17879 2598
rect 17845 2592 17879 2597
rect 17613 2571 17787 2574
rect 17606 2568 17787 2571
rect 17815 2591 17879 2592
rect 17409 2548 17428 2550
rect 17443 2548 17477 2550
rect 17409 2532 17489 2548
rect 17409 2526 17428 2532
rect 17125 2500 17228 2510
rect 17079 2498 17228 2500
rect 17249 2498 17284 2510
rect 16918 2496 17080 2498
rect 16930 2476 16949 2496
rect 16964 2494 16994 2496
rect 16813 2468 16854 2476
rect 16936 2472 16949 2476
rect 17001 2480 17080 2496
rect 17112 2496 17284 2498
rect 17112 2480 17191 2496
rect 17198 2494 17228 2496
rect 16776 2458 16805 2468
rect 16819 2458 16848 2468
rect 16863 2458 16893 2472
rect 16936 2458 16979 2472
rect 17001 2468 17191 2480
rect 17256 2476 17262 2496
rect 16986 2458 17016 2468
rect 17017 2458 17175 2468
rect 17179 2458 17209 2468
rect 17213 2458 17243 2472
rect 17271 2458 17284 2496
rect 17356 2510 17385 2526
rect 17399 2510 17428 2526
rect 17443 2516 17473 2532
rect 17501 2510 17507 2558
rect 17510 2552 17529 2558
rect 17544 2552 17574 2560
rect 17510 2544 17574 2552
rect 17510 2528 17590 2544
rect 17606 2537 17668 2568
rect 17684 2537 17746 2568
rect 17815 2566 17864 2591
rect 17879 2566 17909 2582
rect 17778 2552 17808 2560
rect 17815 2558 17925 2566
rect 17778 2544 17823 2552
rect 17510 2526 17529 2528
rect 17544 2526 17590 2528
rect 17510 2510 17590 2526
rect 17617 2524 17652 2537
rect 17693 2534 17730 2537
rect 17693 2532 17735 2534
rect 17622 2521 17652 2524
rect 17631 2517 17638 2521
rect 17638 2516 17639 2517
rect 17597 2510 17607 2516
rect 17356 2502 17391 2510
rect 17356 2476 17357 2502
rect 17364 2476 17391 2502
rect 17299 2458 17329 2472
rect 17356 2468 17391 2476
rect 17393 2502 17434 2510
rect 17393 2476 17408 2502
rect 17415 2476 17434 2502
rect 17498 2498 17529 2510
rect 17544 2498 17647 2510
rect 17659 2500 17685 2526
rect 17700 2521 17730 2532
rect 17762 2528 17824 2544
rect 17762 2526 17808 2528
rect 17762 2510 17824 2526
rect 17836 2510 17842 2558
rect 17845 2550 17925 2558
rect 17845 2548 17864 2550
rect 17879 2548 17913 2550
rect 17845 2532 17925 2548
rect 17845 2510 17864 2532
rect 17879 2516 17909 2532
rect 17937 2526 17943 2600
rect 17946 2526 17965 2670
rect 17980 2526 17986 2670
rect 17995 2600 18008 2670
rect 18060 2666 18082 2670
rect 18053 2644 18082 2658
rect 18135 2644 18151 2658
rect 18189 2654 18195 2656
rect 18202 2654 18310 2670
rect 18317 2654 18323 2656
rect 18331 2654 18346 2670
rect 18412 2664 18431 2667
rect 18053 2642 18151 2644
rect 18178 2642 18346 2654
rect 18361 2644 18377 2658
rect 18412 2645 18434 2664
rect 18444 2658 18460 2659
rect 18443 2656 18460 2658
rect 18444 2651 18460 2656
rect 18434 2644 18440 2645
rect 18443 2644 18472 2651
rect 18361 2643 18472 2644
rect 18361 2642 18478 2643
rect 18037 2634 18088 2642
rect 18135 2634 18169 2642
rect 18037 2622 18062 2634
rect 18069 2622 18088 2634
rect 18142 2632 18169 2634
rect 18178 2632 18399 2642
rect 18434 2639 18440 2642
rect 18142 2628 18399 2632
rect 18037 2614 18088 2622
rect 18135 2614 18399 2628
rect 18443 2634 18478 2642
rect 17989 2566 18008 2600
rect 18053 2606 18082 2614
rect 18053 2600 18070 2606
rect 18053 2598 18087 2600
rect 18135 2598 18151 2614
rect 18152 2604 18360 2614
rect 18361 2604 18377 2614
rect 18425 2610 18440 2625
rect 18443 2622 18444 2634
rect 18451 2622 18478 2634
rect 18443 2614 18478 2622
rect 18443 2613 18472 2614
rect 18163 2600 18377 2604
rect 18178 2598 18377 2600
rect 18412 2600 18425 2610
rect 18443 2600 18460 2613
rect 18412 2598 18460 2600
rect 18054 2594 18087 2598
rect 18050 2592 18087 2594
rect 18050 2591 18117 2592
rect 18050 2586 18081 2591
rect 18087 2586 18117 2591
rect 18050 2582 18117 2586
rect 18023 2579 18117 2582
rect 18023 2572 18072 2579
rect 18023 2566 18053 2572
rect 18072 2567 18077 2572
rect 17989 2550 18069 2566
rect 18081 2558 18117 2579
rect 18178 2574 18367 2598
rect 18412 2597 18459 2598
rect 18425 2592 18459 2597
rect 18193 2571 18367 2574
rect 18186 2568 18367 2571
rect 18395 2591 18459 2592
rect 17989 2548 18008 2550
rect 18023 2548 18057 2550
rect 17989 2532 18069 2548
rect 17989 2526 18008 2532
rect 17705 2500 17808 2510
rect 17659 2498 17808 2500
rect 17829 2498 17864 2510
rect 17498 2496 17660 2498
rect 17510 2476 17529 2496
rect 17544 2494 17574 2496
rect 17393 2468 17434 2476
rect 17516 2472 17529 2476
rect 17581 2480 17660 2496
rect 17692 2496 17864 2498
rect 17692 2480 17771 2496
rect 17778 2494 17808 2496
rect 17356 2458 17385 2468
rect 17399 2458 17428 2468
rect 17443 2458 17473 2472
rect 17516 2458 17559 2472
rect 17581 2468 17771 2480
rect 17836 2476 17842 2496
rect 17566 2458 17596 2468
rect 17597 2458 17755 2468
rect 17759 2458 17789 2468
rect 17793 2458 17823 2472
rect 17851 2458 17864 2496
rect 17936 2510 17965 2526
rect 17979 2510 18008 2526
rect 18023 2516 18053 2532
rect 18081 2510 18087 2558
rect 18090 2552 18109 2558
rect 18124 2552 18154 2560
rect 18090 2544 18154 2552
rect 18090 2528 18170 2544
rect 18186 2537 18248 2568
rect 18264 2537 18326 2568
rect 18395 2566 18444 2591
rect 18459 2566 18489 2582
rect 18358 2552 18388 2560
rect 18395 2558 18505 2566
rect 18358 2544 18403 2552
rect 18090 2526 18109 2528
rect 18124 2526 18170 2528
rect 18090 2510 18170 2526
rect 18197 2524 18232 2537
rect 18273 2534 18310 2537
rect 18273 2532 18315 2534
rect 18202 2521 18232 2524
rect 18211 2517 18218 2521
rect 18218 2516 18219 2517
rect 18177 2510 18187 2516
rect 17936 2502 17971 2510
rect 17936 2476 17937 2502
rect 17944 2476 17971 2502
rect 17879 2458 17909 2472
rect 17936 2468 17971 2476
rect 17973 2502 18014 2510
rect 17973 2476 17988 2502
rect 17995 2476 18014 2502
rect 18078 2498 18109 2510
rect 18124 2498 18227 2510
rect 18239 2500 18265 2526
rect 18280 2521 18310 2532
rect 18342 2528 18404 2544
rect 18342 2526 18388 2528
rect 18342 2510 18404 2526
rect 18416 2510 18422 2558
rect 18425 2550 18505 2558
rect 18425 2548 18444 2550
rect 18459 2548 18493 2550
rect 18425 2532 18505 2548
rect 18425 2510 18444 2532
rect 18459 2516 18489 2532
rect 18517 2526 18523 2600
rect 18532 2526 18545 2670
rect 18285 2500 18388 2510
rect 18239 2498 18388 2500
rect 18409 2498 18444 2510
rect 18078 2496 18240 2498
rect 18090 2476 18109 2496
rect 18124 2494 18154 2496
rect 17973 2468 18014 2476
rect 18096 2472 18109 2476
rect 18161 2480 18240 2496
rect 18272 2496 18444 2498
rect 18272 2480 18351 2496
rect 18358 2494 18388 2496
rect 17936 2458 17965 2468
rect 17979 2458 18008 2468
rect 18023 2458 18053 2472
rect 18096 2458 18139 2472
rect 18161 2468 18351 2480
rect 18416 2476 18422 2496
rect 18146 2458 18176 2468
rect 18177 2458 18335 2468
rect 18339 2458 18369 2468
rect 18373 2458 18403 2472
rect 18431 2458 18444 2496
rect 18516 2510 18545 2526
rect 18516 2502 18551 2510
rect 18516 2476 18517 2502
rect 18524 2476 18551 2502
rect 18459 2458 18489 2472
rect 18516 2468 18551 2476
rect 18516 2458 18545 2468
rect -1 2452 18545 2458
rect 0 2444 18545 2452
rect 15 2414 28 2444
rect 43 2430 73 2444
rect 116 2430 159 2444
rect 166 2430 386 2444
rect 393 2430 423 2444
rect 83 2416 98 2428
rect 117 2416 130 2430
rect 198 2426 351 2430
rect 80 2414 102 2416
rect 180 2414 372 2426
rect 451 2414 464 2444
rect 479 2430 509 2444
rect 546 2414 565 2444
rect 580 2414 586 2444
rect 595 2414 608 2444
rect 623 2430 653 2444
rect 696 2430 739 2444
rect 746 2430 966 2444
rect 973 2430 1003 2444
rect 663 2416 678 2428
rect 697 2416 710 2430
rect 778 2426 931 2430
rect 660 2414 682 2416
rect 760 2414 952 2426
rect 1031 2414 1044 2444
rect 1059 2430 1089 2444
rect 1126 2414 1145 2444
rect 1160 2414 1166 2444
rect 1175 2414 1188 2444
rect 1203 2430 1233 2444
rect 1276 2430 1319 2444
rect 1326 2430 1546 2444
rect 1553 2430 1583 2444
rect 1243 2416 1258 2428
rect 1277 2416 1290 2430
rect 1358 2426 1511 2430
rect 1240 2414 1262 2416
rect 1340 2414 1532 2426
rect 1611 2414 1624 2444
rect 1639 2430 1669 2444
rect 1706 2414 1725 2444
rect 1740 2414 1746 2444
rect 1755 2414 1768 2444
rect 1783 2430 1813 2444
rect 1856 2430 1899 2444
rect 1906 2430 2126 2444
rect 2133 2430 2163 2444
rect 1823 2416 1838 2428
rect 1857 2416 1870 2430
rect 1938 2426 2091 2430
rect 1820 2414 1842 2416
rect 1920 2414 2112 2426
rect 2191 2414 2204 2444
rect 2219 2430 2249 2444
rect 2286 2414 2305 2444
rect 2320 2414 2326 2444
rect 2335 2414 2348 2444
rect 2363 2430 2393 2444
rect 2436 2430 2479 2444
rect 2486 2430 2706 2444
rect 2713 2430 2743 2444
rect 2403 2416 2418 2428
rect 2437 2416 2450 2430
rect 2518 2426 2671 2430
rect 2400 2414 2422 2416
rect 2500 2414 2692 2426
rect 2771 2414 2784 2444
rect 2799 2430 2829 2444
rect 2866 2414 2885 2444
rect 2900 2414 2906 2444
rect 2915 2414 2928 2444
rect 2943 2430 2973 2444
rect 3016 2430 3059 2444
rect 3066 2430 3286 2444
rect 3293 2430 3323 2444
rect 2983 2416 2998 2428
rect 3017 2416 3030 2430
rect 3098 2426 3251 2430
rect 2980 2414 3002 2416
rect 3080 2414 3272 2426
rect 3351 2414 3364 2444
rect 3379 2430 3409 2444
rect 3446 2414 3465 2444
rect 3480 2414 3486 2444
rect 3495 2414 3508 2444
rect 3523 2430 3553 2444
rect 3596 2430 3639 2444
rect 3646 2430 3866 2444
rect 3873 2430 3903 2444
rect 3563 2416 3578 2428
rect 3597 2416 3610 2430
rect 3678 2426 3831 2430
rect 3560 2414 3582 2416
rect 3660 2414 3852 2426
rect 3931 2414 3944 2444
rect 3959 2430 3989 2444
rect 4026 2414 4045 2444
rect 4060 2414 4066 2444
rect 4075 2414 4088 2444
rect 4103 2430 4133 2444
rect 4176 2430 4219 2444
rect 4226 2430 4446 2444
rect 4453 2430 4483 2444
rect 4143 2416 4158 2428
rect 4177 2416 4190 2430
rect 4258 2426 4411 2430
rect 4140 2414 4162 2416
rect 4240 2414 4432 2426
rect 4511 2414 4524 2444
rect 4539 2430 4569 2444
rect 4606 2414 4625 2444
rect 4640 2414 4646 2444
rect 4655 2414 4668 2444
rect 4683 2430 4713 2444
rect 4756 2430 4799 2444
rect 4806 2430 5026 2444
rect 5033 2430 5063 2444
rect 4723 2416 4738 2428
rect 4757 2416 4770 2430
rect 4838 2426 4991 2430
rect 4720 2414 4742 2416
rect 4820 2414 5012 2426
rect 5091 2414 5104 2444
rect 5119 2430 5149 2444
rect 5186 2414 5205 2444
rect 5220 2414 5226 2444
rect 5235 2414 5248 2444
rect 5263 2430 5293 2444
rect 5336 2430 5379 2444
rect 5386 2430 5606 2444
rect 5613 2430 5643 2444
rect 5303 2416 5318 2428
rect 5337 2416 5350 2430
rect 5418 2426 5571 2430
rect 5300 2414 5322 2416
rect 5400 2414 5592 2426
rect 5671 2414 5684 2444
rect 5699 2430 5729 2444
rect 5766 2414 5785 2444
rect 5800 2414 5806 2444
rect 5815 2414 5828 2444
rect 5843 2430 5873 2444
rect 5916 2430 5959 2444
rect 5966 2430 6186 2444
rect 6193 2430 6223 2444
rect 5883 2416 5898 2428
rect 5917 2416 5930 2430
rect 5998 2426 6151 2430
rect 5880 2414 5902 2416
rect 5980 2414 6172 2426
rect 6251 2414 6264 2444
rect 6279 2430 6309 2444
rect 6346 2414 6365 2444
rect 6380 2414 6386 2444
rect 6395 2414 6408 2444
rect 6423 2430 6453 2444
rect 6496 2430 6539 2444
rect 6546 2430 6766 2444
rect 6773 2430 6803 2444
rect 6463 2416 6478 2428
rect 6497 2416 6510 2430
rect 6578 2426 6731 2430
rect 6460 2414 6482 2416
rect 6560 2414 6752 2426
rect 6831 2414 6844 2444
rect 6859 2430 6889 2444
rect 6926 2414 6945 2444
rect 6960 2414 6966 2444
rect 6975 2414 6988 2444
rect 7003 2430 7033 2444
rect 7076 2430 7119 2444
rect 7126 2430 7346 2444
rect 7353 2430 7383 2444
rect 7043 2416 7058 2428
rect 7077 2416 7090 2430
rect 7158 2426 7311 2430
rect 7040 2414 7062 2416
rect 7140 2414 7332 2426
rect 7411 2414 7424 2444
rect 7439 2430 7469 2444
rect 7506 2414 7525 2444
rect 7540 2414 7546 2444
rect 7555 2414 7568 2444
rect 7583 2430 7613 2444
rect 7656 2430 7699 2444
rect 7706 2430 7926 2444
rect 7933 2430 7963 2444
rect 7623 2416 7638 2428
rect 7657 2416 7670 2430
rect 7738 2426 7891 2430
rect 7620 2414 7642 2416
rect 7720 2414 7912 2426
rect 7991 2414 8004 2444
rect 8019 2430 8049 2444
rect 8086 2414 8105 2444
rect 8120 2414 8126 2444
rect 8135 2414 8148 2444
rect 8163 2430 8193 2444
rect 8236 2430 8279 2444
rect 8286 2430 8506 2444
rect 8513 2430 8543 2444
rect 8203 2416 8218 2428
rect 8237 2416 8250 2430
rect 8318 2426 8471 2430
rect 8200 2414 8222 2416
rect 8300 2414 8492 2426
rect 8571 2414 8584 2444
rect 8599 2430 8629 2444
rect 8666 2414 8685 2444
rect 8700 2414 8706 2444
rect 8715 2414 8728 2444
rect 8743 2430 8773 2444
rect 8816 2430 8859 2444
rect 8866 2430 9086 2444
rect 9093 2430 9123 2444
rect 8783 2416 8798 2428
rect 8817 2416 8830 2430
rect 8898 2426 9051 2430
rect 8780 2414 8802 2416
rect 8880 2414 9072 2426
rect 9151 2414 9164 2444
rect 9179 2430 9209 2444
rect 9246 2414 9265 2444
rect 9280 2414 9286 2444
rect 9295 2414 9308 2444
rect 9323 2430 9353 2444
rect 9396 2430 9439 2444
rect 9446 2430 9666 2444
rect 9673 2430 9703 2444
rect 9363 2416 9378 2428
rect 9397 2416 9410 2430
rect 9478 2426 9631 2430
rect 9360 2414 9382 2416
rect 9460 2414 9652 2426
rect 9731 2414 9744 2444
rect 9759 2430 9789 2444
rect 9826 2414 9845 2444
rect 9860 2414 9866 2444
rect 9875 2414 9888 2444
rect 9903 2430 9933 2444
rect 9976 2430 10019 2444
rect 10026 2430 10246 2444
rect 10253 2430 10283 2444
rect 9943 2416 9958 2428
rect 9977 2416 9990 2430
rect 10058 2426 10211 2430
rect 9940 2414 9962 2416
rect 10040 2414 10232 2426
rect 10311 2414 10324 2444
rect 10339 2430 10369 2444
rect 10406 2414 10425 2444
rect 10440 2414 10446 2444
rect 10455 2414 10468 2444
rect 10483 2430 10513 2444
rect 10556 2430 10599 2444
rect 10606 2430 10826 2444
rect 10833 2430 10863 2444
rect 10523 2416 10538 2428
rect 10557 2416 10570 2430
rect 10638 2426 10791 2430
rect 10520 2414 10542 2416
rect 10620 2414 10812 2426
rect 10891 2414 10904 2444
rect 10919 2430 10949 2444
rect 10986 2414 11005 2444
rect 11020 2414 11026 2444
rect 11035 2414 11048 2444
rect 11063 2430 11093 2444
rect 11136 2430 11179 2444
rect 11186 2430 11406 2444
rect 11413 2430 11443 2444
rect 11103 2416 11118 2428
rect 11137 2416 11150 2430
rect 11218 2426 11371 2430
rect 11100 2414 11122 2416
rect 11200 2414 11392 2426
rect 11471 2414 11484 2444
rect 11499 2430 11529 2444
rect 11566 2414 11585 2444
rect 11600 2414 11606 2444
rect 11615 2414 11628 2444
rect 11643 2430 11673 2444
rect 11716 2430 11759 2444
rect 11766 2430 11986 2444
rect 11993 2430 12023 2444
rect 11683 2416 11698 2428
rect 11717 2416 11730 2430
rect 11798 2426 11951 2430
rect 11680 2414 11702 2416
rect 11780 2414 11972 2426
rect 12051 2414 12064 2444
rect 12079 2430 12109 2444
rect 12146 2414 12165 2444
rect 12180 2414 12186 2444
rect 12195 2414 12208 2444
rect 12223 2430 12253 2444
rect 12296 2430 12339 2444
rect 12346 2430 12566 2444
rect 12573 2430 12603 2444
rect 12263 2416 12278 2428
rect 12297 2416 12310 2430
rect 12378 2426 12531 2430
rect 12260 2414 12282 2416
rect 12360 2414 12552 2426
rect 12631 2414 12644 2444
rect 12659 2430 12689 2444
rect 12726 2414 12745 2444
rect 12760 2414 12766 2444
rect 12775 2414 12788 2444
rect 12803 2430 12833 2444
rect 12876 2430 12919 2444
rect 12926 2430 13146 2444
rect 13153 2430 13183 2444
rect 12843 2416 12858 2428
rect 12877 2416 12890 2430
rect 12958 2426 13111 2430
rect 12840 2414 12862 2416
rect 12940 2414 13132 2426
rect 13211 2414 13224 2444
rect 13239 2430 13269 2444
rect 13306 2414 13325 2444
rect 13340 2414 13346 2444
rect 13355 2414 13368 2444
rect 13383 2430 13413 2444
rect 13456 2430 13499 2444
rect 13506 2430 13726 2444
rect 13733 2430 13763 2444
rect 13423 2416 13438 2428
rect 13457 2416 13470 2430
rect 13538 2426 13691 2430
rect 13420 2414 13442 2416
rect 13520 2414 13712 2426
rect 13791 2414 13804 2444
rect 13819 2430 13849 2444
rect 13886 2414 13905 2444
rect 13920 2414 13926 2444
rect 13935 2414 13948 2444
rect 13963 2430 13993 2444
rect 14036 2430 14079 2444
rect 14086 2430 14306 2444
rect 14313 2430 14343 2444
rect 14003 2416 14018 2428
rect 14037 2416 14050 2430
rect 14118 2426 14271 2430
rect 14000 2414 14022 2416
rect 14100 2414 14292 2426
rect 14371 2414 14384 2444
rect 14399 2430 14429 2444
rect 14466 2414 14485 2444
rect 14500 2414 14506 2444
rect 14515 2414 14528 2444
rect 14543 2430 14573 2444
rect 14616 2430 14659 2444
rect 14666 2430 14886 2444
rect 14893 2430 14923 2444
rect 14583 2416 14598 2428
rect 14617 2416 14630 2430
rect 14698 2426 14851 2430
rect 14580 2414 14602 2416
rect 14680 2414 14872 2426
rect 14951 2414 14964 2444
rect 14979 2430 15009 2444
rect 15046 2414 15065 2444
rect 15080 2414 15086 2444
rect 15095 2414 15108 2444
rect 15123 2430 15153 2444
rect 15196 2430 15239 2444
rect 15246 2430 15466 2444
rect 15473 2430 15503 2444
rect 15163 2416 15178 2428
rect 15197 2416 15210 2430
rect 15278 2426 15431 2430
rect 15160 2414 15182 2416
rect 15260 2414 15452 2426
rect 15531 2414 15544 2444
rect 15559 2430 15589 2444
rect 15626 2414 15645 2444
rect 15660 2414 15666 2444
rect 15675 2414 15688 2444
rect 15703 2430 15733 2444
rect 15776 2430 15819 2444
rect 15826 2430 16046 2444
rect 16053 2430 16083 2444
rect 15743 2416 15758 2428
rect 15777 2416 15790 2430
rect 15858 2426 16011 2430
rect 15740 2414 15762 2416
rect 15840 2414 16032 2426
rect 16111 2414 16124 2444
rect 16139 2430 16169 2444
rect 16206 2414 16225 2444
rect 16240 2414 16246 2444
rect 16255 2414 16268 2444
rect 16283 2430 16313 2444
rect 16356 2430 16399 2444
rect 16406 2430 16626 2444
rect 16633 2430 16663 2444
rect 16323 2416 16338 2428
rect 16357 2416 16370 2430
rect 16438 2426 16591 2430
rect 16320 2414 16342 2416
rect 16420 2414 16612 2426
rect 16691 2414 16704 2444
rect 16719 2430 16749 2444
rect 16786 2414 16805 2444
rect 16820 2414 16826 2444
rect 16835 2414 16848 2444
rect 16863 2430 16893 2444
rect 16936 2430 16979 2444
rect 16986 2430 17206 2444
rect 17213 2430 17243 2444
rect 16903 2416 16918 2428
rect 16937 2416 16950 2430
rect 17018 2426 17171 2430
rect 16900 2414 16922 2416
rect 17000 2414 17192 2426
rect 17271 2414 17284 2444
rect 17299 2430 17329 2444
rect 17366 2414 17385 2444
rect 17400 2414 17406 2444
rect 17415 2414 17428 2444
rect 17443 2430 17473 2444
rect 17516 2430 17559 2444
rect 17566 2430 17786 2444
rect 17793 2430 17823 2444
rect 17483 2416 17498 2428
rect 17517 2416 17530 2430
rect 17598 2426 17751 2430
rect 17480 2414 17502 2416
rect 17580 2414 17772 2426
rect 17851 2414 17864 2444
rect 17879 2430 17909 2444
rect 17946 2414 17965 2444
rect 17980 2414 17986 2444
rect 17995 2414 18008 2444
rect 18023 2430 18053 2444
rect 18096 2430 18139 2444
rect 18146 2430 18366 2444
rect 18373 2430 18403 2444
rect 18063 2416 18078 2428
rect 18097 2416 18110 2430
rect 18178 2426 18331 2430
rect 18060 2414 18082 2416
rect 18160 2414 18352 2426
rect 18431 2414 18444 2444
rect 18459 2430 18489 2444
rect 18532 2414 18545 2444
rect 0 2400 18545 2414
rect 15 2330 28 2400
rect 80 2396 102 2400
rect 73 2374 102 2388
rect 155 2374 171 2388
rect 209 2384 215 2386
rect 222 2384 330 2400
rect 337 2384 343 2386
rect 351 2384 366 2400
rect 432 2394 451 2397
rect 73 2372 171 2374
rect 198 2372 366 2384
rect 381 2374 397 2388
rect 432 2375 454 2394
rect 464 2388 480 2389
rect 463 2386 480 2388
rect 464 2381 480 2386
rect 454 2374 460 2375
rect 463 2374 492 2381
rect 381 2373 492 2374
rect 381 2372 498 2373
rect 57 2364 108 2372
rect 155 2364 189 2372
rect 57 2352 82 2364
rect 89 2352 108 2364
rect 162 2362 189 2364
rect 198 2362 419 2372
rect 454 2369 460 2372
rect 162 2358 419 2362
rect 57 2344 108 2352
rect 155 2344 419 2358
rect 463 2364 498 2372
rect 9 2296 28 2330
rect 73 2336 102 2344
rect 73 2330 90 2336
rect 73 2328 107 2330
rect 155 2328 171 2344
rect 172 2334 380 2344
rect 381 2334 397 2344
rect 445 2340 460 2355
rect 463 2352 464 2364
rect 471 2352 498 2364
rect 463 2344 498 2352
rect 463 2343 492 2344
rect 183 2330 397 2334
rect 198 2328 397 2330
rect 432 2330 445 2340
rect 463 2330 480 2343
rect 432 2328 480 2330
rect 74 2324 107 2328
rect 70 2322 107 2324
rect 70 2321 137 2322
rect 70 2316 101 2321
rect 107 2316 137 2321
rect 70 2312 137 2316
rect 43 2309 137 2312
rect 43 2302 92 2309
rect 43 2296 73 2302
rect 92 2297 97 2302
rect 9 2280 89 2296
rect 101 2288 137 2309
rect 198 2304 387 2328
rect 432 2327 479 2328
rect 445 2322 479 2327
rect 213 2301 387 2304
rect 206 2298 387 2301
rect 415 2321 479 2322
rect 9 2278 28 2280
rect 43 2278 77 2280
rect 9 2262 89 2278
rect 9 2256 28 2262
rect -1 2240 28 2256
rect 43 2246 73 2262
rect 101 2240 107 2288
rect 110 2282 129 2288
rect 144 2282 174 2290
rect 110 2274 174 2282
rect 110 2258 190 2274
rect 206 2267 268 2298
rect 284 2267 346 2298
rect 415 2296 464 2321
rect 479 2296 509 2312
rect 378 2282 408 2290
rect 415 2288 525 2296
rect 378 2274 423 2282
rect 110 2256 129 2258
rect 144 2256 190 2258
rect 110 2240 190 2256
rect 217 2254 252 2267
rect 293 2264 330 2267
rect 293 2262 335 2264
rect 222 2251 252 2254
rect 231 2247 238 2251
rect 238 2246 239 2247
rect 197 2240 207 2246
rect -7 2232 34 2240
rect -7 2206 8 2232
rect 15 2206 34 2232
rect 98 2228 129 2240
rect 144 2228 247 2240
rect 259 2230 285 2256
rect 300 2251 330 2262
rect 362 2258 424 2274
rect 362 2256 408 2258
rect 362 2240 424 2256
rect 436 2240 442 2288
rect 445 2280 525 2288
rect 445 2278 464 2280
rect 479 2278 513 2280
rect 445 2262 525 2278
rect 445 2240 464 2262
rect 479 2246 509 2262
rect 537 2256 543 2330
rect 546 2256 565 2400
rect 580 2256 586 2400
rect 595 2330 608 2400
rect 660 2396 682 2400
rect 653 2374 682 2388
rect 735 2374 751 2388
rect 789 2384 795 2386
rect 802 2384 910 2400
rect 917 2384 923 2386
rect 931 2384 946 2400
rect 1012 2394 1031 2397
rect 653 2372 751 2374
rect 778 2372 946 2384
rect 961 2374 977 2388
rect 1012 2375 1034 2394
rect 1044 2388 1060 2389
rect 1043 2386 1060 2388
rect 1044 2381 1060 2386
rect 1034 2374 1040 2375
rect 1043 2374 1072 2381
rect 961 2373 1072 2374
rect 961 2372 1078 2373
rect 637 2364 688 2372
rect 735 2364 769 2372
rect 637 2352 662 2364
rect 669 2352 688 2364
rect 742 2362 769 2364
rect 778 2362 999 2372
rect 1034 2369 1040 2372
rect 742 2358 999 2362
rect 637 2344 688 2352
rect 735 2344 999 2358
rect 1043 2364 1078 2372
rect 589 2296 608 2330
rect 653 2336 682 2344
rect 653 2330 670 2336
rect 653 2328 687 2330
rect 735 2328 751 2344
rect 752 2334 960 2344
rect 961 2334 977 2344
rect 1025 2340 1040 2355
rect 1043 2352 1044 2364
rect 1051 2352 1078 2364
rect 1043 2344 1078 2352
rect 1043 2343 1072 2344
rect 763 2330 977 2334
rect 778 2328 977 2330
rect 1012 2330 1025 2340
rect 1043 2330 1060 2343
rect 1012 2328 1060 2330
rect 654 2324 687 2328
rect 650 2322 687 2324
rect 650 2321 717 2322
rect 650 2316 681 2321
rect 687 2316 717 2321
rect 650 2312 717 2316
rect 623 2309 717 2312
rect 623 2302 672 2309
rect 623 2296 653 2302
rect 672 2297 677 2302
rect 589 2280 669 2296
rect 681 2288 717 2309
rect 778 2304 967 2328
rect 1012 2327 1059 2328
rect 1025 2322 1059 2327
rect 793 2301 967 2304
rect 786 2298 967 2301
rect 995 2321 1059 2322
rect 589 2278 608 2280
rect 623 2278 657 2280
rect 589 2262 669 2278
rect 589 2256 608 2262
rect 305 2230 408 2240
rect 259 2228 408 2230
rect 429 2228 464 2240
rect 98 2226 260 2228
rect 110 2206 129 2226
rect 144 2224 174 2226
rect -7 2198 34 2206
rect 116 2202 129 2206
rect 181 2210 260 2226
rect 292 2226 464 2228
rect 292 2210 371 2226
rect 378 2224 408 2226
rect -1 2188 28 2198
rect 43 2188 73 2202
rect 116 2188 159 2202
rect 181 2198 371 2210
rect 436 2206 442 2226
rect 166 2188 196 2198
rect 197 2188 355 2198
rect 359 2188 389 2198
rect 393 2188 423 2202
rect 451 2188 464 2226
rect 536 2240 565 2256
rect 579 2240 608 2256
rect 623 2246 653 2262
rect 681 2240 687 2288
rect 690 2282 709 2288
rect 724 2282 754 2290
rect 690 2274 754 2282
rect 690 2258 770 2274
rect 786 2267 848 2298
rect 864 2267 926 2298
rect 995 2296 1044 2321
rect 1059 2296 1089 2312
rect 958 2282 988 2290
rect 995 2288 1105 2296
rect 958 2274 1003 2282
rect 690 2256 709 2258
rect 724 2256 770 2258
rect 690 2240 770 2256
rect 797 2254 832 2267
rect 873 2264 910 2267
rect 873 2262 915 2264
rect 802 2251 832 2254
rect 811 2247 818 2251
rect 818 2246 819 2247
rect 777 2240 787 2246
rect 536 2232 571 2240
rect 536 2206 537 2232
rect 544 2206 571 2232
rect 479 2188 509 2202
rect 536 2198 571 2206
rect 573 2232 614 2240
rect 573 2206 588 2232
rect 595 2206 614 2232
rect 678 2228 709 2240
rect 724 2228 827 2240
rect 839 2230 865 2256
rect 880 2251 910 2262
rect 942 2258 1004 2274
rect 942 2256 988 2258
rect 942 2240 1004 2256
rect 1016 2240 1022 2288
rect 1025 2280 1105 2288
rect 1025 2278 1044 2280
rect 1059 2278 1093 2280
rect 1025 2262 1105 2278
rect 1025 2240 1044 2262
rect 1059 2246 1089 2262
rect 1117 2256 1123 2330
rect 1126 2256 1145 2400
rect 1160 2256 1166 2400
rect 1175 2330 1188 2400
rect 1240 2396 1262 2400
rect 1233 2374 1262 2388
rect 1315 2374 1331 2388
rect 1369 2384 1375 2386
rect 1382 2384 1490 2400
rect 1497 2384 1503 2386
rect 1511 2384 1526 2400
rect 1592 2394 1611 2397
rect 1233 2372 1331 2374
rect 1358 2372 1526 2384
rect 1541 2374 1557 2388
rect 1592 2375 1614 2394
rect 1624 2388 1640 2389
rect 1623 2386 1640 2388
rect 1624 2381 1640 2386
rect 1614 2374 1620 2375
rect 1623 2374 1652 2381
rect 1541 2373 1652 2374
rect 1541 2372 1658 2373
rect 1217 2364 1268 2372
rect 1315 2364 1349 2372
rect 1217 2352 1242 2364
rect 1249 2352 1268 2364
rect 1322 2362 1349 2364
rect 1358 2362 1579 2372
rect 1614 2369 1620 2372
rect 1322 2358 1579 2362
rect 1217 2344 1268 2352
rect 1315 2344 1579 2358
rect 1623 2364 1658 2372
rect 1169 2296 1188 2330
rect 1233 2336 1262 2344
rect 1233 2330 1250 2336
rect 1233 2328 1267 2330
rect 1315 2328 1331 2344
rect 1332 2334 1540 2344
rect 1541 2334 1557 2344
rect 1605 2340 1620 2355
rect 1623 2352 1624 2364
rect 1631 2352 1658 2364
rect 1623 2344 1658 2352
rect 1623 2343 1652 2344
rect 1343 2330 1557 2334
rect 1358 2328 1557 2330
rect 1592 2330 1605 2340
rect 1623 2330 1640 2343
rect 1592 2328 1640 2330
rect 1234 2324 1267 2328
rect 1230 2322 1267 2324
rect 1230 2321 1297 2322
rect 1230 2316 1261 2321
rect 1267 2316 1297 2321
rect 1230 2312 1297 2316
rect 1203 2309 1297 2312
rect 1203 2302 1252 2309
rect 1203 2296 1233 2302
rect 1252 2297 1257 2302
rect 1169 2280 1249 2296
rect 1261 2288 1297 2309
rect 1358 2304 1547 2328
rect 1592 2327 1639 2328
rect 1605 2322 1639 2327
rect 1373 2301 1547 2304
rect 1366 2298 1547 2301
rect 1575 2321 1639 2322
rect 1169 2278 1188 2280
rect 1203 2278 1237 2280
rect 1169 2262 1249 2278
rect 1169 2256 1188 2262
rect 885 2230 988 2240
rect 839 2228 988 2230
rect 1009 2228 1044 2240
rect 678 2226 840 2228
rect 690 2206 709 2226
rect 724 2224 754 2226
rect 573 2198 614 2206
rect 696 2202 709 2206
rect 761 2210 840 2226
rect 872 2226 1044 2228
rect 872 2210 951 2226
rect 958 2224 988 2226
rect 536 2188 565 2198
rect 579 2188 608 2198
rect 623 2188 653 2202
rect 696 2188 739 2202
rect 761 2198 951 2210
rect 1016 2206 1022 2226
rect 746 2188 776 2198
rect 777 2188 935 2198
rect 939 2188 969 2198
rect 973 2188 1003 2202
rect 1031 2188 1044 2226
rect 1116 2240 1145 2256
rect 1159 2240 1188 2256
rect 1203 2246 1233 2262
rect 1261 2240 1267 2288
rect 1270 2282 1289 2288
rect 1304 2282 1334 2290
rect 1270 2274 1334 2282
rect 1270 2258 1350 2274
rect 1366 2267 1428 2298
rect 1444 2267 1506 2298
rect 1575 2296 1624 2321
rect 1639 2296 1669 2312
rect 1538 2282 1568 2290
rect 1575 2288 1685 2296
rect 1538 2274 1583 2282
rect 1270 2256 1289 2258
rect 1304 2256 1350 2258
rect 1270 2240 1350 2256
rect 1377 2254 1412 2267
rect 1453 2264 1490 2267
rect 1453 2262 1495 2264
rect 1382 2251 1412 2254
rect 1391 2247 1398 2251
rect 1398 2246 1399 2247
rect 1357 2240 1367 2246
rect 1116 2232 1151 2240
rect 1116 2206 1117 2232
rect 1124 2206 1151 2232
rect 1059 2188 1089 2202
rect 1116 2198 1151 2206
rect 1153 2232 1194 2240
rect 1153 2206 1168 2232
rect 1175 2206 1194 2232
rect 1258 2228 1289 2240
rect 1304 2228 1407 2240
rect 1419 2230 1445 2256
rect 1460 2251 1490 2262
rect 1522 2258 1584 2274
rect 1522 2256 1568 2258
rect 1522 2240 1584 2256
rect 1596 2240 1602 2288
rect 1605 2280 1685 2288
rect 1605 2278 1624 2280
rect 1639 2278 1673 2280
rect 1605 2262 1685 2278
rect 1605 2240 1624 2262
rect 1639 2246 1669 2262
rect 1697 2256 1703 2330
rect 1706 2256 1725 2400
rect 1740 2256 1746 2400
rect 1755 2330 1768 2400
rect 1820 2396 1842 2400
rect 1813 2374 1842 2388
rect 1895 2374 1911 2388
rect 1949 2384 1955 2386
rect 1962 2384 2070 2400
rect 2077 2384 2083 2386
rect 2091 2384 2106 2400
rect 2172 2394 2191 2397
rect 1813 2372 1911 2374
rect 1938 2372 2106 2384
rect 2121 2374 2137 2388
rect 2172 2375 2194 2394
rect 2204 2388 2220 2389
rect 2203 2386 2220 2388
rect 2204 2381 2220 2386
rect 2194 2374 2200 2375
rect 2203 2374 2232 2381
rect 2121 2373 2232 2374
rect 2121 2372 2238 2373
rect 1797 2364 1848 2372
rect 1895 2364 1929 2372
rect 1797 2352 1822 2364
rect 1829 2352 1848 2364
rect 1902 2362 1929 2364
rect 1938 2362 2159 2372
rect 2194 2369 2200 2372
rect 1902 2358 2159 2362
rect 1797 2344 1848 2352
rect 1895 2344 2159 2358
rect 2203 2364 2238 2372
rect 1749 2296 1768 2330
rect 1813 2336 1842 2344
rect 1813 2330 1830 2336
rect 1813 2328 1847 2330
rect 1895 2328 1911 2344
rect 1912 2334 2120 2344
rect 2121 2334 2137 2344
rect 2185 2340 2200 2355
rect 2203 2352 2204 2364
rect 2211 2352 2238 2364
rect 2203 2344 2238 2352
rect 2203 2343 2232 2344
rect 1923 2330 2137 2334
rect 1938 2328 2137 2330
rect 2172 2330 2185 2340
rect 2203 2330 2220 2343
rect 2172 2328 2220 2330
rect 1814 2324 1847 2328
rect 1810 2322 1847 2324
rect 1810 2321 1877 2322
rect 1810 2316 1841 2321
rect 1847 2316 1877 2321
rect 1810 2312 1877 2316
rect 1783 2309 1877 2312
rect 1783 2302 1832 2309
rect 1783 2296 1813 2302
rect 1832 2297 1837 2302
rect 1749 2280 1829 2296
rect 1841 2288 1877 2309
rect 1938 2304 2127 2328
rect 2172 2327 2219 2328
rect 2185 2322 2219 2327
rect 1953 2301 2127 2304
rect 1946 2298 2127 2301
rect 2155 2321 2219 2322
rect 1749 2278 1768 2280
rect 1783 2278 1817 2280
rect 1749 2262 1829 2278
rect 1749 2256 1768 2262
rect 1465 2230 1568 2240
rect 1419 2228 1568 2230
rect 1589 2228 1624 2240
rect 1258 2226 1420 2228
rect 1270 2206 1289 2226
rect 1304 2224 1334 2226
rect 1153 2198 1194 2206
rect 1276 2202 1289 2206
rect 1341 2210 1420 2226
rect 1452 2226 1624 2228
rect 1452 2210 1531 2226
rect 1538 2224 1568 2226
rect 1116 2188 1145 2198
rect 1159 2188 1188 2198
rect 1203 2188 1233 2202
rect 1276 2188 1319 2202
rect 1341 2198 1531 2210
rect 1596 2206 1602 2226
rect 1326 2188 1356 2198
rect 1357 2188 1515 2198
rect 1519 2188 1549 2198
rect 1553 2188 1583 2202
rect 1611 2188 1624 2226
rect 1696 2240 1725 2256
rect 1739 2240 1768 2256
rect 1783 2246 1813 2262
rect 1841 2240 1847 2288
rect 1850 2282 1869 2288
rect 1884 2282 1914 2290
rect 1850 2274 1914 2282
rect 1850 2258 1930 2274
rect 1946 2267 2008 2298
rect 2024 2267 2086 2298
rect 2155 2296 2204 2321
rect 2219 2296 2249 2312
rect 2118 2282 2148 2290
rect 2155 2288 2265 2296
rect 2118 2274 2163 2282
rect 1850 2256 1869 2258
rect 1884 2256 1930 2258
rect 1850 2240 1930 2256
rect 1957 2254 1992 2267
rect 2033 2264 2070 2267
rect 2033 2262 2075 2264
rect 1962 2251 1992 2254
rect 1971 2247 1978 2251
rect 1978 2246 1979 2247
rect 1937 2240 1947 2246
rect 1696 2232 1731 2240
rect 1696 2206 1697 2232
rect 1704 2206 1731 2232
rect 1639 2188 1669 2202
rect 1696 2198 1731 2206
rect 1733 2232 1774 2240
rect 1733 2206 1748 2232
rect 1755 2206 1774 2232
rect 1838 2228 1869 2240
rect 1884 2228 1987 2240
rect 1999 2230 2025 2256
rect 2040 2251 2070 2262
rect 2102 2258 2164 2274
rect 2102 2256 2148 2258
rect 2102 2240 2164 2256
rect 2176 2240 2182 2288
rect 2185 2280 2265 2288
rect 2185 2278 2204 2280
rect 2219 2278 2253 2280
rect 2185 2262 2265 2278
rect 2185 2240 2204 2262
rect 2219 2246 2249 2262
rect 2277 2256 2283 2330
rect 2286 2256 2305 2400
rect 2320 2256 2326 2400
rect 2335 2330 2348 2400
rect 2400 2396 2422 2400
rect 2393 2374 2422 2388
rect 2475 2374 2491 2388
rect 2529 2384 2535 2386
rect 2542 2384 2650 2400
rect 2657 2384 2663 2386
rect 2671 2384 2686 2400
rect 2752 2394 2771 2397
rect 2393 2372 2491 2374
rect 2518 2372 2686 2384
rect 2701 2374 2717 2388
rect 2752 2375 2774 2394
rect 2784 2388 2800 2389
rect 2783 2386 2800 2388
rect 2784 2381 2800 2386
rect 2774 2374 2780 2375
rect 2783 2374 2812 2381
rect 2701 2373 2812 2374
rect 2701 2372 2818 2373
rect 2377 2364 2428 2372
rect 2475 2364 2509 2372
rect 2377 2352 2402 2364
rect 2409 2352 2428 2364
rect 2482 2362 2509 2364
rect 2518 2362 2739 2372
rect 2774 2369 2780 2372
rect 2482 2358 2739 2362
rect 2377 2344 2428 2352
rect 2475 2344 2739 2358
rect 2783 2364 2818 2372
rect 2329 2296 2348 2330
rect 2393 2336 2422 2344
rect 2393 2330 2410 2336
rect 2393 2328 2427 2330
rect 2475 2328 2491 2344
rect 2492 2334 2700 2344
rect 2701 2334 2717 2344
rect 2765 2340 2780 2355
rect 2783 2352 2784 2364
rect 2791 2352 2818 2364
rect 2783 2344 2818 2352
rect 2783 2343 2812 2344
rect 2503 2330 2717 2334
rect 2518 2328 2717 2330
rect 2752 2330 2765 2340
rect 2783 2330 2800 2343
rect 2752 2328 2800 2330
rect 2394 2324 2427 2328
rect 2390 2322 2427 2324
rect 2390 2321 2457 2322
rect 2390 2316 2421 2321
rect 2427 2316 2457 2321
rect 2390 2312 2457 2316
rect 2363 2309 2457 2312
rect 2363 2302 2412 2309
rect 2363 2296 2393 2302
rect 2412 2297 2417 2302
rect 2329 2280 2409 2296
rect 2421 2288 2457 2309
rect 2518 2304 2707 2328
rect 2752 2327 2799 2328
rect 2765 2322 2799 2327
rect 2533 2301 2707 2304
rect 2526 2298 2707 2301
rect 2735 2321 2799 2322
rect 2329 2278 2348 2280
rect 2363 2278 2397 2280
rect 2329 2262 2409 2278
rect 2329 2256 2348 2262
rect 2045 2230 2148 2240
rect 1999 2228 2148 2230
rect 2169 2228 2204 2240
rect 1838 2226 2000 2228
rect 1850 2206 1869 2226
rect 1884 2224 1914 2226
rect 1733 2198 1774 2206
rect 1856 2202 1869 2206
rect 1921 2210 2000 2226
rect 2032 2226 2204 2228
rect 2032 2210 2111 2226
rect 2118 2224 2148 2226
rect 1696 2188 1725 2198
rect 1739 2188 1768 2198
rect 1783 2188 1813 2202
rect 1856 2188 1899 2202
rect 1921 2198 2111 2210
rect 2176 2206 2182 2226
rect 1906 2188 1936 2198
rect 1937 2188 2095 2198
rect 2099 2188 2129 2198
rect 2133 2188 2163 2202
rect 2191 2188 2204 2226
rect 2276 2240 2305 2256
rect 2319 2240 2348 2256
rect 2363 2246 2393 2262
rect 2421 2240 2427 2288
rect 2430 2282 2449 2288
rect 2464 2282 2494 2290
rect 2430 2274 2494 2282
rect 2430 2258 2510 2274
rect 2526 2267 2588 2298
rect 2604 2267 2666 2298
rect 2735 2296 2784 2321
rect 2799 2296 2829 2312
rect 2698 2282 2728 2290
rect 2735 2288 2845 2296
rect 2698 2274 2743 2282
rect 2430 2256 2449 2258
rect 2464 2256 2510 2258
rect 2430 2240 2510 2256
rect 2537 2254 2572 2267
rect 2613 2264 2650 2267
rect 2613 2262 2655 2264
rect 2542 2251 2572 2254
rect 2551 2247 2558 2251
rect 2558 2246 2559 2247
rect 2517 2240 2527 2246
rect 2276 2232 2311 2240
rect 2276 2206 2277 2232
rect 2284 2206 2311 2232
rect 2219 2188 2249 2202
rect 2276 2198 2311 2206
rect 2313 2232 2354 2240
rect 2313 2206 2328 2232
rect 2335 2206 2354 2232
rect 2418 2228 2449 2240
rect 2464 2228 2567 2240
rect 2579 2230 2605 2256
rect 2620 2251 2650 2262
rect 2682 2258 2744 2274
rect 2682 2256 2728 2258
rect 2682 2240 2744 2256
rect 2756 2240 2762 2288
rect 2765 2280 2845 2288
rect 2765 2278 2784 2280
rect 2799 2278 2833 2280
rect 2765 2262 2845 2278
rect 2765 2240 2784 2262
rect 2799 2246 2829 2262
rect 2857 2256 2863 2330
rect 2866 2256 2885 2400
rect 2900 2256 2906 2400
rect 2915 2330 2928 2400
rect 2980 2396 3002 2400
rect 2973 2374 3002 2388
rect 3055 2374 3071 2388
rect 3109 2384 3115 2386
rect 3122 2384 3230 2400
rect 3237 2384 3243 2386
rect 3251 2384 3266 2400
rect 3332 2394 3351 2397
rect 2973 2372 3071 2374
rect 3098 2372 3266 2384
rect 3281 2374 3297 2388
rect 3332 2375 3354 2394
rect 3364 2388 3380 2389
rect 3363 2386 3380 2388
rect 3364 2381 3380 2386
rect 3354 2374 3360 2375
rect 3363 2374 3392 2381
rect 3281 2373 3392 2374
rect 3281 2372 3398 2373
rect 2957 2364 3008 2372
rect 3055 2364 3089 2372
rect 2957 2352 2982 2364
rect 2989 2352 3008 2364
rect 3062 2362 3089 2364
rect 3098 2362 3319 2372
rect 3354 2369 3360 2372
rect 3062 2358 3319 2362
rect 2957 2344 3008 2352
rect 3055 2344 3319 2358
rect 3363 2364 3398 2372
rect 2909 2296 2928 2330
rect 2973 2336 3002 2344
rect 2973 2330 2990 2336
rect 2973 2328 3007 2330
rect 3055 2328 3071 2344
rect 3072 2334 3280 2344
rect 3281 2334 3297 2344
rect 3345 2340 3360 2355
rect 3363 2352 3364 2364
rect 3371 2352 3398 2364
rect 3363 2344 3398 2352
rect 3363 2343 3392 2344
rect 3083 2330 3297 2334
rect 3098 2328 3297 2330
rect 3332 2330 3345 2340
rect 3363 2330 3380 2343
rect 3332 2328 3380 2330
rect 2974 2324 3007 2328
rect 2970 2322 3007 2324
rect 2970 2321 3037 2322
rect 2970 2316 3001 2321
rect 3007 2316 3037 2321
rect 2970 2312 3037 2316
rect 2943 2309 3037 2312
rect 2943 2302 2992 2309
rect 2943 2296 2973 2302
rect 2992 2297 2997 2302
rect 2909 2280 2989 2296
rect 3001 2288 3037 2309
rect 3098 2304 3287 2328
rect 3332 2327 3379 2328
rect 3345 2322 3379 2327
rect 3113 2301 3287 2304
rect 3106 2298 3287 2301
rect 3315 2321 3379 2322
rect 2909 2278 2928 2280
rect 2943 2278 2977 2280
rect 2909 2262 2989 2278
rect 2909 2256 2928 2262
rect 2625 2230 2728 2240
rect 2579 2228 2728 2230
rect 2749 2228 2784 2240
rect 2418 2226 2580 2228
rect 2430 2206 2449 2226
rect 2464 2224 2494 2226
rect 2313 2198 2354 2206
rect 2436 2202 2449 2206
rect 2501 2210 2580 2226
rect 2612 2226 2784 2228
rect 2612 2210 2691 2226
rect 2698 2224 2728 2226
rect 2276 2188 2305 2198
rect 2319 2188 2348 2198
rect 2363 2188 2393 2202
rect 2436 2188 2479 2202
rect 2501 2198 2691 2210
rect 2756 2206 2762 2226
rect 2486 2188 2516 2198
rect 2517 2188 2675 2198
rect 2679 2188 2709 2198
rect 2713 2188 2743 2202
rect 2771 2188 2784 2226
rect 2856 2240 2885 2256
rect 2899 2240 2928 2256
rect 2943 2246 2973 2262
rect 3001 2240 3007 2288
rect 3010 2282 3029 2288
rect 3044 2282 3074 2290
rect 3010 2274 3074 2282
rect 3010 2258 3090 2274
rect 3106 2267 3168 2298
rect 3184 2267 3246 2298
rect 3315 2296 3364 2321
rect 3379 2296 3409 2312
rect 3278 2282 3308 2290
rect 3315 2288 3425 2296
rect 3278 2274 3323 2282
rect 3010 2256 3029 2258
rect 3044 2256 3090 2258
rect 3010 2240 3090 2256
rect 3117 2254 3152 2267
rect 3193 2264 3230 2267
rect 3193 2262 3235 2264
rect 3122 2251 3152 2254
rect 3131 2247 3138 2251
rect 3138 2246 3139 2247
rect 3097 2240 3107 2246
rect 2856 2232 2891 2240
rect 2856 2206 2857 2232
rect 2864 2206 2891 2232
rect 2799 2188 2829 2202
rect 2856 2198 2891 2206
rect 2893 2232 2934 2240
rect 2893 2206 2908 2232
rect 2915 2206 2934 2232
rect 2998 2228 3029 2240
rect 3044 2228 3147 2240
rect 3159 2230 3185 2256
rect 3200 2251 3230 2262
rect 3262 2258 3324 2274
rect 3262 2256 3308 2258
rect 3262 2240 3324 2256
rect 3336 2240 3342 2288
rect 3345 2280 3425 2288
rect 3345 2278 3364 2280
rect 3379 2278 3413 2280
rect 3345 2262 3425 2278
rect 3345 2240 3364 2262
rect 3379 2246 3409 2262
rect 3437 2256 3443 2330
rect 3446 2256 3465 2400
rect 3480 2256 3486 2400
rect 3495 2330 3508 2400
rect 3560 2396 3582 2400
rect 3553 2374 3582 2388
rect 3635 2374 3651 2388
rect 3689 2384 3695 2386
rect 3702 2384 3810 2400
rect 3817 2384 3823 2386
rect 3831 2384 3846 2400
rect 3912 2394 3931 2397
rect 3553 2372 3651 2374
rect 3678 2372 3846 2384
rect 3861 2374 3877 2388
rect 3912 2375 3934 2394
rect 3944 2388 3960 2389
rect 3943 2386 3960 2388
rect 3944 2381 3960 2386
rect 3934 2374 3940 2375
rect 3943 2374 3972 2381
rect 3861 2373 3972 2374
rect 3861 2372 3978 2373
rect 3537 2364 3588 2372
rect 3635 2364 3669 2372
rect 3537 2352 3562 2364
rect 3569 2352 3588 2364
rect 3642 2362 3669 2364
rect 3678 2362 3899 2372
rect 3934 2369 3940 2372
rect 3642 2358 3899 2362
rect 3537 2344 3588 2352
rect 3635 2344 3899 2358
rect 3943 2364 3978 2372
rect 3489 2296 3508 2330
rect 3553 2336 3582 2344
rect 3553 2330 3570 2336
rect 3553 2328 3587 2330
rect 3635 2328 3651 2344
rect 3652 2334 3860 2344
rect 3861 2334 3877 2344
rect 3925 2340 3940 2355
rect 3943 2352 3944 2364
rect 3951 2352 3978 2364
rect 3943 2344 3978 2352
rect 3943 2343 3972 2344
rect 3663 2330 3877 2334
rect 3678 2328 3877 2330
rect 3912 2330 3925 2340
rect 3943 2330 3960 2343
rect 3912 2328 3960 2330
rect 3554 2324 3587 2328
rect 3550 2322 3587 2324
rect 3550 2321 3617 2322
rect 3550 2316 3581 2321
rect 3587 2316 3617 2321
rect 3550 2312 3617 2316
rect 3523 2309 3617 2312
rect 3523 2302 3572 2309
rect 3523 2296 3553 2302
rect 3572 2297 3577 2302
rect 3489 2280 3569 2296
rect 3581 2288 3617 2309
rect 3678 2304 3867 2328
rect 3912 2327 3959 2328
rect 3925 2322 3959 2327
rect 3693 2301 3867 2304
rect 3686 2298 3867 2301
rect 3895 2321 3959 2322
rect 3489 2278 3508 2280
rect 3523 2278 3557 2280
rect 3489 2262 3569 2278
rect 3489 2256 3508 2262
rect 3205 2230 3308 2240
rect 3159 2228 3308 2230
rect 3329 2228 3364 2240
rect 2998 2226 3160 2228
rect 3010 2206 3029 2226
rect 3044 2224 3074 2226
rect 2893 2198 2934 2206
rect 3016 2202 3029 2206
rect 3081 2210 3160 2226
rect 3192 2226 3364 2228
rect 3192 2210 3271 2226
rect 3278 2224 3308 2226
rect 2856 2188 2885 2198
rect 2899 2188 2928 2198
rect 2943 2188 2973 2202
rect 3016 2188 3059 2202
rect 3081 2198 3271 2210
rect 3336 2206 3342 2226
rect 3066 2188 3096 2198
rect 3097 2188 3255 2198
rect 3259 2188 3289 2198
rect 3293 2188 3323 2202
rect 3351 2188 3364 2226
rect 3436 2240 3465 2256
rect 3479 2240 3508 2256
rect 3523 2246 3553 2262
rect 3581 2240 3587 2288
rect 3590 2282 3609 2288
rect 3624 2282 3654 2290
rect 3590 2274 3654 2282
rect 3590 2258 3670 2274
rect 3686 2267 3748 2298
rect 3764 2267 3826 2298
rect 3895 2296 3944 2321
rect 3959 2296 3989 2312
rect 3858 2282 3888 2290
rect 3895 2288 4005 2296
rect 3858 2274 3903 2282
rect 3590 2256 3609 2258
rect 3624 2256 3670 2258
rect 3590 2240 3670 2256
rect 3697 2254 3732 2267
rect 3773 2264 3810 2267
rect 3773 2262 3815 2264
rect 3702 2251 3732 2254
rect 3711 2247 3718 2251
rect 3718 2246 3719 2247
rect 3677 2240 3687 2246
rect 3436 2232 3471 2240
rect 3436 2206 3437 2232
rect 3444 2206 3471 2232
rect 3379 2188 3409 2202
rect 3436 2198 3471 2206
rect 3473 2232 3514 2240
rect 3473 2206 3488 2232
rect 3495 2206 3514 2232
rect 3578 2228 3609 2240
rect 3624 2228 3727 2240
rect 3739 2230 3765 2256
rect 3780 2251 3810 2262
rect 3842 2258 3904 2274
rect 3842 2256 3888 2258
rect 3842 2240 3904 2256
rect 3916 2240 3922 2288
rect 3925 2280 4005 2288
rect 3925 2278 3944 2280
rect 3959 2278 3993 2280
rect 3925 2262 4005 2278
rect 3925 2240 3944 2262
rect 3959 2246 3989 2262
rect 4017 2256 4023 2330
rect 4026 2256 4045 2400
rect 4060 2256 4066 2400
rect 4075 2330 4088 2400
rect 4140 2396 4162 2400
rect 4133 2374 4162 2388
rect 4215 2374 4231 2388
rect 4269 2384 4275 2386
rect 4282 2384 4390 2400
rect 4397 2384 4403 2386
rect 4411 2384 4426 2400
rect 4492 2394 4511 2397
rect 4133 2372 4231 2374
rect 4258 2372 4426 2384
rect 4441 2374 4457 2388
rect 4492 2375 4514 2394
rect 4524 2388 4540 2389
rect 4523 2386 4540 2388
rect 4524 2381 4540 2386
rect 4514 2374 4520 2375
rect 4523 2374 4552 2381
rect 4441 2373 4552 2374
rect 4441 2372 4558 2373
rect 4117 2364 4168 2372
rect 4215 2364 4249 2372
rect 4117 2352 4142 2364
rect 4149 2352 4168 2364
rect 4222 2362 4249 2364
rect 4258 2362 4479 2372
rect 4514 2369 4520 2372
rect 4222 2358 4479 2362
rect 4117 2344 4168 2352
rect 4215 2344 4479 2358
rect 4523 2364 4558 2372
rect 4069 2296 4088 2330
rect 4133 2336 4162 2344
rect 4133 2330 4150 2336
rect 4133 2328 4167 2330
rect 4215 2328 4231 2344
rect 4232 2334 4440 2344
rect 4441 2334 4457 2344
rect 4505 2340 4520 2355
rect 4523 2352 4524 2364
rect 4531 2352 4558 2364
rect 4523 2344 4558 2352
rect 4523 2343 4552 2344
rect 4243 2330 4457 2334
rect 4258 2328 4457 2330
rect 4492 2330 4505 2340
rect 4523 2330 4540 2343
rect 4492 2328 4540 2330
rect 4134 2324 4167 2328
rect 4130 2322 4167 2324
rect 4130 2321 4197 2322
rect 4130 2316 4161 2321
rect 4167 2316 4197 2321
rect 4130 2312 4197 2316
rect 4103 2309 4197 2312
rect 4103 2302 4152 2309
rect 4103 2296 4133 2302
rect 4152 2297 4157 2302
rect 4069 2280 4149 2296
rect 4161 2288 4197 2309
rect 4258 2304 4447 2328
rect 4492 2327 4539 2328
rect 4505 2322 4539 2327
rect 4273 2301 4447 2304
rect 4266 2298 4447 2301
rect 4475 2321 4539 2322
rect 4069 2278 4088 2280
rect 4103 2278 4137 2280
rect 4069 2262 4149 2278
rect 4069 2256 4088 2262
rect 3785 2230 3888 2240
rect 3739 2228 3888 2230
rect 3909 2228 3944 2240
rect 3578 2226 3740 2228
rect 3590 2206 3609 2226
rect 3624 2224 3654 2226
rect 3473 2198 3514 2206
rect 3596 2202 3609 2206
rect 3661 2210 3740 2226
rect 3772 2226 3944 2228
rect 3772 2210 3851 2226
rect 3858 2224 3888 2226
rect 3436 2188 3465 2198
rect 3479 2188 3508 2198
rect 3523 2188 3553 2202
rect 3596 2188 3639 2202
rect 3661 2198 3851 2210
rect 3916 2206 3922 2226
rect 3646 2188 3676 2198
rect 3677 2188 3835 2198
rect 3839 2188 3869 2198
rect 3873 2188 3903 2202
rect 3931 2188 3944 2226
rect 4016 2240 4045 2256
rect 4059 2240 4088 2256
rect 4103 2246 4133 2262
rect 4161 2240 4167 2288
rect 4170 2282 4189 2288
rect 4204 2282 4234 2290
rect 4170 2274 4234 2282
rect 4170 2258 4250 2274
rect 4266 2267 4328 2298
rect 4344 2267 4406 2298
rect 4475 2296 4524 2321
rect 4539 2296 4569 2312
rect 4438 2282 4468 2290
rect 4475 2288 4585 2296
rect 4438 2274 4483 2282
rect 4170 2256 4189 2258
rect 4204 2256 4250 2258
rect 4170 2240 4250 2256
rect 4277 2254 4312 2267
rect 4353 2264 4390 2267
rect 4353 2262 4395 2264
rect 4282 2251 4312 2254
rect 4291 2247 4298 2251
rect 4298 2246 4299 2247
rect 4257 2240 4267 2246
rect 4016 2232 4051 2240
rect 4016 2206 4017 2232
rect 4024 2206 4051 2232
rect 3959 2188 3989 2202
rect 4016 2198 4051 2206
rect 4053 2232 4094 2240
rect 4053 2206 4068 2232
rect 4075 2206 4094 2232
rect 4158 2228 4189 2240
rect 4204 2228 4307 2240
rect 4319 2230 4345 2256
rect 4360 2251 4390 2262
rect 4422 2258 4484 2274
rect 4422 2256 4468 2258
rect 4422 2240 4484 2256
rect 4496 2240 4502 2288
rect 4505 2280 4585 2288
rect 4505 2278 4524 2280
rect 4539 2278 4573 2280
rect 4505 2262 4585 2278
rect 4505 2240 4524 2262
rect 4539 2246 4569 2262
rect 4597 2256 4603 2330
rect 4606 2256 4625 2400
rect 4640 2256 4646 2400
rect 4655 2330 4668 2400
rect 4720 2396 4742 2400
rect 4713 2374 4742 2388
rect 4795 2374 4811 2388
rect 4849 2384 4855 2386
rect 4862 2384 4970 2400
rect 4977 2384 4983 2386
rect 4991 2384 5006 2400
rect 5072 2394 5091 2397
rect 4713 2372 4811 2374
rect 4838 2372 5006 2384
rect 5021 2374 5037 2388
rect 5072 2375 5094 2394
rect 5104 2388 5120 2389
rect 5103 2386 5120 2388
rect 5104 2381 5120 2386
rect 5094 2374 5100 2375
rect 5103 2374 5132 2381
rect 5021 2373 5132 2374
rect 5021 2372 5138 2373
rect 4697 2364 4748 2372
rect 4795 2364 4829 2372
rect 4697 2352 4722 2364
rect 4729 2352 4748 2364
rect 4802 2362 4829 2364
rect 4838 2362 5059 2372
rect 5094 2369 5100 2372
rect 4802 2358 5059 2362
rect 4697 2344 4748 2352
rect 4795 2344 5059 2358
rect 5103 2364 5138 2372
rect 4649 2296 4668 2330
rect 4713 2336 4742 2344
rect 4713 2330 4730 2336
rect 4713 2328 4747 2330
rect 4795 2328 4811 2344
rect 4812 2334 5020 2344
rect 5021 2334 5037 2344
rect 5085 2340 5100 2355
rect 5103 2352 5104 2364
rect 5111 2352 5138 2364
rect 5103 2344 5138 2352
rect 5103 2343 5132 2344
rect 4823 2330 5037 2334
rect 4838 2328 5037 2330
rect 5072 2330 5085 2340
rect 5103 2330 5120 2343
rect 5072 2328 5120 2330
rect 4714 2324 4747 2328
rect 4710 2322 4747 2324
rect 4710 2321 4777 2322
rect 4710 2316 4741 2321
rect 4747 2316 4777 2321
rect 4710 2312 4777 2316
rect 4683 2309 4777 2312
rect 4683 2302 4732 2309
rect 4683 2296 4713 2302
rect 4732 2297 4737 2302
rect 4649 2280 4729 2296
rect 4741 2288 4777 2309
rect 4838 2304 5027 2328
rect 5072 2327 5119 2328
rect 5085 2322 5119 2327
rect 4853 2301 5027 2304
rect 4846 2298 5027 2301
rect 5055 2321 5119 2322
rect 4649 2278 4668 2280
rect 4683 2278 4717 2280
rect 4649 2262 4729 2278
rect 4649 2256 4668 2262
rect 4365 2230 4468 2240
rect 4319 2228 4468 2230
rect 4489 2228 4524 2240
rect 4158 2226 4320 2228
rect 4170 2206 4189 2226
rect 4204 2224 4234 2226
rect 4053 2198 4094 2206
rect 4176 2202 4189 2206
rect 4241 2210 4320 2226
rect 4352 2226 4524 2228
rect 4352 2210 4431 2226
rect 4438 2224 4468 2226
rect 4016 2188 4045 2198
rect 4059 2188 4088 2198
rect 4103 2188 4133 2202
rect 4176 2188 4219 2202
rect 4241 2198 4431 2210
rect 4496 2206 4502 2226
rect 4226 2188 4256 2198
rect 4257 2188 4415 2198
rect 4419 2188 4449 2198
rect 4453 2188 4483 2202
rect 4511 2188 4524 2226
rect 4596 2240 4625 2256
rect 4639 2240 4668 2256
rect 4683 2246 4713 2262
rect 4741 2240 4747 2288
rect 4750 2282 4769 2288
rect 4784 2282 4814 2290
rect 4750 2274 4814 2282
rect 4750 2258 4830 2274
rect 4846 2267 4908 2298
rect 4924 2267 4986 2298
rect 5055 2296 5104 2321
rect 5119 2296 5149 2312
rect 5018 2282 5048 2290
rect 5055 2288 5165 2296
rect 5018 2274 5063 2282
rect 4750 2256 4769 2258
rect 4784 2256 4830 2258
rect 4750 2240 4830 2256
rect 4857 2254 4892 2267
rect 4933 2264 4970 2267
rect 4933 2262 4975 2264
rect 4862 2251 4892 2254
rect 4871 2247 4878 2251
rect 4878 2246 4879 2247
rect 4837 2240 4847 2246
rect 4596 2232 4631 2240
rect 4596 2206 4597 2232
rect 4604 2206 4631 2232
rect 4539 2188 4569 2202
rect 4596 2198 4631 2206
rect 4633 2232 4674 2240
rect 4633 2206 4648 2232
rect 4655 2206 4674 2232
rect 4738 2228 4769 2240
rect 4784 2228 4887 2240
rect 4899 2230 4925 2256
rect 4940 2251 4970 2262
rect 5002 2258 5064 2274
rect 5002 2256 5048 2258
rect 5002 2240 5064 2256
rect 5076 2240 5082 2288
rect 5085 2280 5165 2288
rect 5085 2278 5104 2280
rect 5119 2278 5153 2280
rect 5085 2262 5165 2278
rect 5085 2240 5104 2262
rect 5119 2246 5149 2262
rect 5177 2256 5183 2330
rect 5186 2256 5205 2400
rect 5220 2256 5226 2400
rect 5235 2330 5248 2400
rect 5300 2396 5322 2400
rect 5293 2374 5322 2388
rect 5375 2374 5391 2388
rect 5429 2384 5435 2386
rect 5442 2384 5550 2400
rect 5557 2384 5563 2386
rect 5571 2384 5586 2400
rect 5652 2394 5671 2397
rect 5293 2372 5391 2374
rect 5418 2372 5586 2384
rect 5601 2374 5617 2388
rect 5652 2375 5674 2394
rect 5684 2388 5700 2389
rect 5683 2386 5700 2388
rect 5684 2381 5700 2386
rect 5674 2374 5680 2375
rect 5683 2374 5712 2381
rect 5601 2373 5712 2374
rect 5601 2372 5718 2373
rect 5277 2364 5328 2372
rect 5375 2364 5409 2372
rect 5277 2352 5302 2364
rect 5309 2352 5328 2364
rect 5382 2362 5409 2364
rect 5418 2362 5639 2372
rect 5674 2369 5680 2372
rect 5382 2358 5639 2362
rect 5277 2344 5328 2352
rect 5375 2344 5639 2358
rect 5683 2364 5718 2372
rect 5229 2296 5248 2330
rect 5293 2336 5322 2344
rect 5293 2330 5310 2336
rect 5293 2328 5327 2330
rect 5375 2328 5391 2344
rect 5392 2334 5600 2344
rect 5601 2334 5617 2344
rect 5665 2340 5680 2355
rect 5683 2352 5684 2364
rect 5691 2352 5718 2364
rect 5683 2344 5718 2352
rect 5683 2343 5712 2344
rect 5403 2330 5617 2334
rect 5418 2328 5617 2330
rect 5652 2330 5665 2340
rect 5683 2330 5700 2343
rect 5652 2328 5700 2330
rect 5294 2324 5327 2328
rect 5290 2322 5327 2324
rect 5290 2321 5357 2322
rect 5290 2316 5321 2321
rect 5327 2316 5357 2321
rect 5290 2312 5357 2316
rect 5263 2309 5357 2312
rect 5263 2302 5312 2309
rect 5263 2296 5293 2302
rect 5312 2297 5317 2302
rect 5229 2280 5309 2296
rect 5321 2288 5357 2309
rect 5418 2304 5607 2328
rect 5652 2327 5699 2328
rect 5665 2322 5699 2327
rect 5433 2301 5607 2304
rect 5426 2298 5607 2301
rect 5635 2321 5699 2322
rect 5229 2278 5248 2280
rect 5263 2278 5297 2280
rect 5229 2262 5309 2278
rect 5229 2256 5248 2262
rect 4945 2230 5048 2240
rect 4899 2228 5048 2230
rect 5069 2228 5104 2240
rect 4738 2226 4900 2228
rect 4750 2206 4769 2226
rect 4784 2224 4814 2226
rect 4633 2198 4674 2206
rect 4756 2202 4769 2206
rect 4821 2210 4900 2226
rect 4932 2226 5104 2228
rect 4932 2210 5011 2226
rect 5018 2224 5048 2226
rect 4596 2188 4625 2198
rect 4639 2188 4668 2198
rect 4683 2188 4713 2202
rect 4756 2188 4799 2202
rect 4821 2198 5011 2210
rect 5076 2206 5082 2226
rect 4806 2188 4836 2198
rect 4837 2188 4995 2198
rect 4999 2188 5029 2198
rect 5033 2188 5063 2202
rect 5091 2188 5104 2226
rect 5176 2240 5205 2256
rect 5219 2240 5248 2256
rect 5263 2246 5293 2262
rect 5321 2240 5327 2288
rect 5330 2282 5349 2288
rect 5364 2282 5394 2290
rect 5330 2274 5394 2282
rect 5330 2258 5410 2274
rect 5426 2267 5488 2298
rect 5504 2267 5566 2298
rect 5635 2296 5684 2321
rect 5699 2296 5729 2312
rect 5598 2282 5628 2290
rect 5635 2288 5745 2296
rect 5598 2274 5643 2282
rect 5330 2256 5349 2258
rect 5364 2256 5410 2258
rect 5330 2240 5410 2256
rect 5437 2254 5472 2267
rect 5513 2264 5550 2267
rect 5513 2262 5555 2264
rect 5442 2251 5472 2254
rect 5451 2247 5458 2251
rect 5458 2246 5459 2247
rect 5417 2240 5427 2246
rect 5176 2232 5211 2240
rect 5176 2206 5177 2232
rect 5184 2206 5211 2232
rect 5119 2188 5149 2202
rect 5176 2198 5211 2206
rect 5213 2232 5254 2240
rect 5213 2206 5228 2232
rect 5235 2206 5254 2232
rect 5318 2228 5349 2240
rect 5364 2228 5467 2240
rect 5479 2230 5505 2256
rect 5520 2251 5550 2262
rect 5582 2258 5644 2274
rect 5582 2256 5628 2258
rect 5582 2240 5644 2256
rect 5656 2240 5662 2288
rect 5665 2280 5745 2288
rect 5665 2278 5684 2280
rect 5699 2278 5733 2280
rect 5665 2262 5745 2278
rect 5665 2240 5684 2262
rect 5699 2246 5729 2262
rect 5757 2256 5763 2330
rect 5766 2256 5785 2400
rect 5800 2256 5806 2400
rect 5815 2330 5828 2400
rect 5880 2396 5902 2400
rect 5873 2374 5902 2388
rect 5955 2374 5971 2388
rect 6009 2384 6015 2386
rect 6022 2384 6130 2400
rect 6137 2384 6143 2386
rect 6151 2384 6166 2400
rect 6232 2394 6251 2397
rect 5873 2372 5971 2374
rect 5998 2372 6166 2384
rect 6181 2374 6197 2388
rect 6232 2375 6254 2394
rect 6264 2388 6280 2389
rect 6263 2386 6280 2388
rect 6264 2381 6280 2386
rect 6254 2374 6260 2375
rect 6263 2374 6292 2381
rect 6181 2373 6292 2374
rect 6181 2372 6298 2373
rect 5857 2364 5908 2372
rect 5955 2364 5989 2372
rect 5857 2352 5882 2364
rect 5889 2352 5908 2364
rect 5962 2362 5989 2364
rect 5998 2362 6219 2372
rect 6254 2369 6260 2372
rect 5962 2358 6219 2362
rect 5857 2344 5908 2352
rect 5955 2344 6219 2358
rect 6263 2364 6298 2372
rect 5809 2296 5828 2330
rect 5873 2336 5902 2344
rect 5873 2330 5890 2336
rect 5873 2328 5907 2330
rect 5955 2328 5971 2344
rect 5972 2334 6180 2344
rect 6181 2334 6197 2344
rect 6245 2340 6260 2355
rect 6263 2352 6264 2364
rect 6271 2352 6298 2364
rect 6263 2344 6298 2352
rect 6263 2343 6292 2344
rect 5983 2330 6197 2334
rect 5998 2328 6197 2330
rect 6232 2330 6245 2340
rect 6263 2330 6280 2343
rect 6232 2328 6280 2330
rect 5874 2324 5907 2328
rect 5870 2322 5907 2324
rect 5870 2321 5937 2322
rect 5870 2316 5901 2321
rect 5907 2316 5937 2321
rect 5870 2312 5937 2316
rect 5843 2309 5937 2312
rect 5843 2302 5892 2309
rect 5843 2296 5873 2302
rect 5892 2297 5897 2302
rect 5809 2280 5889 2296
rect 5901 2288 5937 2309
rect 5998 2304 6187 2328
rect 6232 2327 6279 2328
rect 6245 2322 6279 2327
rect 6013 2301 6187 2304
rect 6006 2298 6187 2301
rect 6215 2321 6279 2322
rect 5809 2278 5828 2280
rect 5843 2278 5877 2280
rect 5809 2262 5889 2278
rect 5809 2256 5828 2262
rect 5525 2230 5628 2240
rect 5479 2228 5628 2230
rect 5649 2228 5684 2240
rect 5318 2226 5480 2228
rect 5330 2206 5349 2226
rect 5364 2224 5394 2226
rect 5213 2198 5254 2206
rect 5336 2202 5349 2206
rect 5401 2210 5480 2226
rect 5512 2226 5684 2228
rect 5512 2210 5591 2226
rect 5598 2224 5628 2226
rect 5176 2188 5205 2198
rect 5219 2188 5248 2198
rect 5263 2188 5293 2202
rect 5336 2188 5379 2202
rect 5401 2198 5591 2210
rect 5656 2206 5662 2226
rect 5386 2188 5416 2198
rect 5417 2188 5575 2198
rect 5579 2188 5609 2198
rect 5613 2188 5643 2202
rect 5671 2188 5684 2226
rect 5756 2240 5785 2256
rect 5799 2240 5828 2256
rect 5843 2246 5873 2262
rect 5901 2240 5907 2288
rect 5910 2282 5929 2288
rect 5944 2282 5974 2290
rect 5910 2274 5974 2282
rect 5910 2258 5990 2274
rect 6006 2267 6068 2298
rect 6084 2267 6146 2298
rect 6215 2296 6264 2321
rect 6279 2296 6309 2312
rect 6178 2282 6208 2290
rect 6215 2288 6325 2296
rect 6178 2274 6223 2282
rect 5910 2256 5929 2258
rect 5944 2256 5990 2258
rect 5910 2240 5990 2256
rect 6017 2254 6052 2267
rect 6093 2264 6130 2267
rect 6093 2262 6135 2264
rect 6022 2251 6052 2254
rect 6031 2247 6038 2251
rect 6038 2246 6039 2247
rect 5997 2240 6007 2246
rect 5756 2232 5791 2240
rect 5756 2206 5757 2232
rect 5764 2206 5791 2232
rect 5699 2188 5729 2202
rect 5756 2198 5791 2206
rect 5793 2232 5834 2240
rect 5793 2206 5808 2232
rect 5815 2206 5834 2232
rect 5898 2228 5929 2240
rect 5944 2228 6047 2240
rect 6059 2230 6085 2256
rect 6100 2251 6130 2262
rect 6162 2258 6224 2274
rect 6162 2256 6208 2258
rect 6162 2240 6224 2256
rect 6236 2240 6242 2288
rect 6245 2280 6325 2288
rect 6245 2278 6264 2280
rect 6279 2278 6313 2280
rect 6245 2262 6325 2278
rect 6245 2240 6264 2262
rect 6279 2246 6309 2262
rect 6337 2256 6343 2330
rect 6346 2256 6365 2400
rect 6380 2256 6386 2400
rect 6395 2330 6408 2400
rect 6460 2396 6482 2400
rect 6453 2374 6482 2388
rect 6535 2374 6551 2388
rect 6589 2384 6595 2386
rect 6602 2384 6710 2400
rect 6717 2384 6723 2386
rect 6731 2384 6746 2400
rect 6812 2394 6831 2397
rect 6453 2372 6551 2374
rect 6578 2372 6746 2384
rect 6761 2374 6777 2388
rect 6812 2375 6834 2394
rect 6844 2388 6860 2389
rect 6843 2386 6860 2388
rect 6844 2381 6860 2386
rect 6834 2374 6840 2375
rect 6843 2374 6872 2381
rect 6761 2373 6872 2374
rect 6761 2372 6878 2373
rect 6437 2364 6488 2372
rect 6535 2364 6569 2372
rect 6437 2352 6462 2364
rect 6469 2352 6488 2364
rect 6542 2362 6569 2364
rect 6578 2362 6799 2372
rect 6834 2369 6840 2372
rect 6542 2358 6799 2362
rect 6437 2344 6488 2352
rect 6535 2344 6799 2358
rect 6843 2364 6878 2372
rect 6389 2296 6408 2330
rect 6453 2336 6482 2344
rect 6453 2330 6470 2336
rect 6453 2328 6487 2330
rect 6535 2328 6551 2344
rect 6552 2334 6760 2344
rect 6761 2334 6777 2344
rect 6825 2340 6840 2355
rect 6843 2352 6844 2364
rect 6851 2352 6878 2364
rect 6843 2344 6878 2352
rect 6843 2343 6872 2344
rect 6563 2330 6777 2334
rect 6578 2328 6777 2330
rect 6812 2330 6825 2340
rect 6843 2330 6860 2343
rect 6812 2328 6860 2330
rect 6454 2324 6487 2328
rect 6450 2322 6487 2324
rect 6450 2321 6517 2322
rect 6450 2316 6481 2321
rect 6487 2316 6517 2321
rect 6450 2312 6517 2316
rect 6423 2309 6517 2312
rect 6423 2302 6472 2309
rect 6423 2296 6453 2302
rect 6472 2297 6477 2302
rect 6389 2280 6469 2296
rect 6481 2288 6517 2309
rect 6578 2304 6767 2328
rect 6812 2327 6859 2328
rect 6825 2322 6859 2327
rect 6593 2301 6767 2304
rect 6586 2298 6767 2301
rect 6795 2321 6859 2322
rect 6389 2278 6408 2280
rect 6423 2278 6457 2280
rect 6389 2262 6469 2278
rect 6389 2256 6408 2262
rect 6105 2230 6208 2240
rect 6059 2228 6208 2230
rect 6229 2228 6264 2240
rect 5898 2226 6060 2228
rect 5910 2206 5929 2226
rect 5944 2224 5974 2226
rect 5793 2198 5834 2206
rect 5916 2202 5929 2206
rect 5981 2210 6060 2226
rect 6092 2226 6264 2228
rect 6092 2210 6171 2226
rect 6178 2224 6208 2226
rect 5756 2188 5785 2198
rect 5799 2188 5828 2198
rect 5843 2188 5873 2202
rect 5916 2188 5959 2202
rect 5981 2198 6171 2210
rect 6236 2206 6242 2226
rect 5966 2188 5996 2198
rect 5997 2188 6155 2198
rect 6159 2188 6189 2198
rect 6193 2188 6223 2202
rect 6251 2188 6264 2226
rect 6336 2240 6365 2256
rect 6379 2240 6408 2256
rect 6423 2246 6453 2262
rect 6481 2240 6487 2288
rect 6490 2282 6509 2288
rect 6524 2282 6554 2290
rect 6490 2274 6554 2282
rect 6490 2258 6570 2274
rect 6586 2267 6648 2298
rect 6664 2267 6726 2298
rect 6795 2296 6844 2321
rect 6859 2296 6889 2312
rect 6758 2282 6788 2290
rect 6795 2288 6905 2296
rect 6758 2274 6803 2282
rect 6490 2256 6509 2258
rect 6524 2256 6570 2258
rect 6490 2240 6570 2256
rect 6597 2254 6632 2267
rect 6673 2264 6710 2267
rect 6673 2262 6715 2264
rect 6602 2251 6632 2254
rect 6611 2247 6618 2251
rect 6618 2246 6619 2247
rect 6577 2240 6587 2246
rect 6336 2232 6371 2240
rect 6336 2206 6337 2232
rect 6344 2206 6371 2232
rect 6279 2188 6309 2202
rect 6336 2198 6371 2206
rect 6373 2232 6414 2240
rect 6373 2206 6388 2232
rect 6395 2206 6414 2232
rect 6478 2228 6509 2240
rect 6524 2228 6627 2240
rect 6639 2230 6665 2256
rect 6680 2251 6710 2262
rect 6742 2258 6804 2274
rect 6742 2256 6788 2258
rect 6742 2240 6804 2256
rect 6816 2240 6822 2288
rect 6825 2280 6905 2288
rect 6825 2278 6844 2280
rect 6859 2278 6893 2280
rect 6825 2262 6905 2278
rect 6825 2240 6844 2262
rect 6859 2246 6889 2262
rect 6917 2256 6923 2330
rect 6926 2256 6945 2400
rect 6960 2256 6966 2400
rect 6975 2330 6988 2400
rect 7040 2396 7062 2400
rect 7033 2374 7062 2388
rect 7115 2374 7131 2388
rect 7169 2384 7175 2386
rect 7182 2384 7290 2400
rect 7297 2384 7303 2386
rect 7311 2384 7326 2400
rect 7392 2394 7411 2397
rect 7033 2372 7131 2374
rect 7158 2372 7326 2384
rect 7341 2374 7357 2388
rect 7392 2375 7414 2394
rect 7424 2388 7440 2389
rect 7423 2386 7440 2388
rect 7424 2381 7440 2386
rect 7414 2374 7420 2375
rect 7423 2374 7452 2381
rect 7341 2373 7452 2374
rect 7341 2372 7458 2373
rect 7017 2364 7068 2372
rect 7115 2364 7149 2372
rect 7017 2352 7042 2364
rect 7049 2352 7068 2364
rect 7122 2362 7149 2364
rect 7158 2362 7379 2372
rect 7414 2369 7420 2372
rect 7122 2358 7379 2362
rect 7017 2344 7068 2352
rect 7115 2344 7379 2358
rect 7423 2364 7458 2372
rect 6969 2296 6988 2330
rect 7033 2336 7062 2344
rect 7033 2330 7050 2336
rect 7033 2328 7067 2330
rect 7115 2328 7131 2344
rect 7132 2334 7340 2344
rect 7341 2334 7357 2344
rect 7405 2340 7420 2355
rect 7423 2352 7424 2364
rect 7431 2352 7458 2364
rect 7423 2344 7458 2352
rect 7423 2343 7452 2344
rect 7151 2330 7357 2334
rect 7158 2328 7357 2330
rect 7392 2330 7405 2340
rect 7423 2330 7440 2343
rect 7392 2328 7440 2330
rect 7034 2324 7067 2328
rect 7030 2322 7067 2324
rect 7030 2321 7097 2322
rect 7030 2316 7061 2321
rect 7067 2316 7097 2321
rect 7030 2312 7097 2316
rect 7003 2309 7097 2312
rect 7003 2302 7052 2309
rect 7003 2296 7033 2302
rect 7052 2297 7057 2302
rect 6969 2280 7049 2296
rect 7061 2288 7097 2309
rect 7158 2304 7347 2328
rect 7392 2327 7439 2328
rect 7405 2322 7439 2327
rect 7173 2301 7347 2304
rect 7166 2298 7347 2301
rect 7375 2321 7439 2322
rect 6969 2278 6988 2280
rect 7003 2278 7037 2280
rect 6969 2262 7049 2278
rect 6969 2256 6988 2262
rect 6685 2230 6788 2240
rect 6639 2228 6788 2230
rect 6809 2228 6844 2240
rect 6478 2226 6640 2228
rect 6490 2206 6509 2226
rect 6524 2224 6554 2226
rect 6373 2198 6414 2206
rect 6496 2202 6509 2206
rect 6561 2210 6640 2226
rect 6672 2226 6844 2228
rect 6672 2210 6751 2226
rect 6758 2224 6788 2226
rect 6336 2188 6365 2198
rect 6379 2188 6408 2198
rect 6423 2188 6453 2202
rect 6496 2188 6539 2202
rect 6561 2198 6751 2210
rect 6816 2206 6822 2226
rect 6546 2188 6576 2198
rect 6577 2188 6735 2198
rect 6739 2188 6769 2198
rect 6773 2188 6803 2202
rect 6831 2188 6844 2226
rect 6916 2240 6945 2256
rect 6959 2240 6988 2256
rect 7003 2246 7033 2262
rect 7061 2240 7067 2288
rect 7070 2282 7089 2288
rect 7104 2282 7134 2290
rect 7070 2274 7134 2282
rect 7070 2258 7150 2274
rect 7166 2267 7228 2298
rect 7244 2267 7306 2298
rect 7375 2296 7424 2321
rect 7439 2296 7469 2312
rect 7338 2282 7368 2290
rect 7375 2288 7485 2296
rect 7338 2274 7383 2282
rect 7070 2256 7089 2258
rect 7104 2256 7150 2258
rect 7070 2240 7150 2256
rect 7177 2254 7212 2267
rect 7253 2264 7290 2267
rect 7253 2262 7295 2264
rect 7182 2251 7212 2254
rect 7191 2247 7198 2251
rect 7198 2246 7199 2247
rect 7157 2240 7167 2246
rect 6916 2232 6951 2240
rect 6916 2206 6917 2232
rect 6924 2206 6951 2232
rect 6859 2188 6889 2202
rect 6916 2198 6951 2206
rect 6953 2232 6994 2240
rect 6953 2206 6968 2232
rect 6975 2206 6994 2232
rect 7058 2228 7089 2240
rect 7104 2228 7207 2240
rect 7219 2230 7245 2256
rect 7260 2251 7290 2262
rect 7322 2258 7384 2274
rect 7322 2256 7368 2258
rect 7322 2240 7384 2256
rect 7396 2240 7402 2288
rect 7405 2280 7485 2288
rect 7405 2278 7424 2280
rect 7439 2278 7473 2280
rect 7405 2262 7485 2278
rect 7405 2240 7424 2262
rect 7439 2246 7469 2262
rect 7497 2256 7503 2330
rect 7506 2256 7525 2400
rect 7540 2256 7546 2400
rect 7555 2330 7568 2400
rect 7620 2396 7642 2400
rect 7613 2374 7642 2388
rect 7695 2374 7711 2388
rect 7749 2384 7755 2386
rect 7762 2384 7870 2400
rect 7877 2384 7883 2386
rect 7891 2384 7906 2400
rect 7972 2394 7991 2397
rect 7613 2372 7711 2374
rect 7738 2372 7906 2384
rect 7921 2374 7937 2388
rect 7972 2375 7994 2394
rect 8004 2388 8020 2389
rect 8003 2386 8020 2388
rect 8004 2381 8020 2386
rect 7994 2374 8000 2375
rect 8003 2374 8032 2381
rect 7921 2373 8032 2374
rect 7921 2372 8038 2373
rect 7597 2364 7648 2372
rect 7695 2364 7729 2372
rect 7597 2352 7622 2364
rect 7629 2352 7648 2364
rect 7702 2362 7729 2364
rect 7738 2362 7959 2372
rect 7994 2369 8000 2372
rect 7702 2358 7959 2362
rect 7597 2344 7648 2352
rect 7695 2344 7959 2358
rect 8003 2364 8038 2372
rect 7549 2296 7568 2330
rect 7613 2336 7642 2344
rect 7613 2330 7630 2336
rect 7613 2328 7647 2330
rect 7695 2328 7711 2344
rect 7712 2334 7920 2344
rect 7921 2334 7937 2344
rect 7985 2340 8000 2355
rect 8003 2352 8004 2364
rect 8011 2352 8038 2364
rect 8003 2344 8038 2352
rect 8003 2343 8032 2344
rect 7723 2330 7937 2334
rect 7738 2328 7937 2330
rect 7972 2330 7985 2340
rect 8003 2330 8020 2343
rect 7972 2328 8020 2330
rect 7614 2324 7647 2328
rect 7610 2322 7647 2324
rect 7610 2321 7677 2322
rect 7610 2316 7641 2321
rect 7647 2316 7677 2321
rect 7610 2312 7677 2316
rect 7583 2309 7677 2312
rect 7583 2302 7632 2309
rect 7583 2296 7613 2302
rect 7632 2297 7637 2302
rect 7549 2280 7629 2296
rect 7641 2288 7677 2309
rect 7738 2304 7927 2328
rect 7972 2327 8019 2328
rect 7985 2322 8019 2327
rect 7753 2301 7927 2304
rect 7746 2298 7927 2301
rect 7955 2321 8019 2322
rect 7549 2278 7568 2280
rect 7583 2278 7617 2280
rect 7549 2262 7629 2278
rect 7549 2256 7568 2262
rect 7265 2230 7368 2240
rect 7219 2228 7368 2230
rect 7389 2228 7424 2240
rect 7058 2226 7220 2228
rect 7070 2206 7089 2226
rect 7104 2224 7134 2226
rect 6953 2198 6994 2206
rect 7076 2202 7089 2206
rect 7141 2210 7220 2226
rect 7252 2226 7424 2228
rect 7252 2210 7331 2226
rect 7338 2224 7368 2226
rect 6916 2188 6945 2198
rect 6959 2188 6988 2198
rect 7003 2188 7033 2202
rect 7076 2188 7119 2202
rect 7141 2198 7331 2210
rect 7396 2206 7402 2226
rect 7126 2188 7156 2198
rect 7157 2188 7315 2198
rect 7319 2188 7349 2198
rect 7353 2188 7383 2202
rect 7411 2188 7424 2226
rect 7496 2240 7525 2256
rect 7539 2240 7568 2256
rect 7583 2246 7613 2262
rect 7641 2240 7647 2288
rect 7650 2282 7669 2288
rect 7684 2282 7714 2290
rect 7650 2274 7714 2282
rect 7650 2258 7730 2274
rect 7746 2267 7808 2298
rect 7824 2267 7886 2298
rect 7955 2296 8004 2321
rect 8019 2296 8049 2312
rect 7918 2282 7948 2290
rect 7955 2288 8065 2296
rect 7918 2274 7963 2282
rect 7650 2256 7669 2258
rect 7684 2256 7730 2258
rect 7650 2240 7730 2256
rect 7757 2254 7792 2267
rect 7833 2264 7870 2267
rect 7833 2262 7875 2264
rect 7762 2251 7792 2254
rect 7771 2247 7778 2251
rect 7778 2246 7779 2247
rect 7737 2240 7747 2246
rect 7496 2232 7531 2240
rect 7496 2206 7497 2232
rect 7504 2206 7531 2232
rect 7439 2188 7469 2202
rect 7496 2198 7531 2206
rect 7533 2232 7574 2240
rect 7533 2206 7548 2232
rect 7555 2206 7574 2232
rect 7638 2228 7669 2240
rect 7684 2228 7787 2240
rect 7799 2230 7825 2256
rect 7840 2251 7870 2262
rect 7902 2258 7964 2274
rect 7902 2256 7948 2258
rect 7902 2240 7964 2256
rect 7976 2240 7982 2288
rect 7985 2280 8065 2288
rect 7985 2278 8004 2280
rect 8019 2278 8053 2280
rect 7985 2262 8065 2278
rect 7985 2240 8004 2262
rect 8019 2246 8049 2262
rect 8077 2256 8083 2330
rect 8086 2256 8105 2400
rect 8120 2256 8126 2400
rect 8135 2330 8148 2400
rect 8200 2396 8222 2400
rect 8193 2374 8222 2388
rect 8275 2374 8291 2388
rect 8329 2384 8335 2386
rect 8342 2384 8450 2400
rect 8457 2384 8463 2386
rect 8471 2384 8486 2400
rect 8552 2394 8571 2397
rect 8193 2372 8291 2374
rect 8318 2372 8486 2384
rect 8501 2374 8517 2388
rect 8552 2375 8574 2394
rect 8584 2388 8600 2389
rect 8583 2386 8600 2388
rect 8584 2381 8600 2386
rect 8574 2374 8580 2375
rect 8583 2374 8612 2381
rect 8501 2373 8612 2374
rect 8501 2372 8618 2373
rect 8177 2364 8228 2372
rect 8275 2364 8309 2372
rect 8177 2352 8202 2364
rect 8209 2352 8228 2364
rect 8282 2362 8309 2364
rect 8318 2362 8539 2372
rect 8574 2369 8580 2372
rect 8282 2358 8539 2362
rect 8177 2344 8228 2352
rect 8275 2344 8539 2358
rect 8583 2364 8618 2372
rect 8129 2296 8148 2330
rect 8193 2336 8222 2344
rect 8193 2330 8210 2336
rect 8193 2328 8227 2330
rect 8275 2328 8291 2344
rect 8292 2334 8500 2344
rect 8501 2334 8517 2344
rect 8565 2340 8580 2355
rect 8583 2352 8584 2364
rect 8591 2352 8618 2364
rect 8583 2344 8618 2352
rect 8583 2343 8612 2344
rect 8303 2330 8517 2334
rect 8318 2328 8517 2330
rect 8552 2330 8565 2340
rect 8583 2330 8600 2343
rect 8552 2328 8600 2330
rect 8194 2324 8227 2328
rect 8190 2322 8227 2324
rect 8190 2321 8257 2322
rect 8190 2316 8221 2321
rect 8227 2316 8257 2321
rect 8190 2312 8257 2316
rect 8163 2309 8257 2312
rect 8163 2302 8212 2309
rect 8163 2296 8193 2302
rect 8212 2297 8217 2302
rect 8129 2280 8209 2296
rect 8221 2288 8257 2309
rect 8318 2304 8507 2328
rect 8552 2327 8599 2328
rect 8565 2322 8599 2327
rect 8333 2301 8507 2304
rect 8326 2298 8507 2301
rect 8535 2321 8599 2322
rect 8129 2278 8148 2280
rect 8163 2278 8197 2280
rect 8129 2262 8209 2278
rect 8129 2256 8148 2262
rect 7845 2230 7948 2240
rect 7799 2228 7948 2230
rect 7969 2228 8004 2240
rect 7638 2226 7800 2228
rect 7650 2206 7669 2226
rect 7684 2224 7714 2226
rect 7533 2198 7574 2206
rect 7656 2202 7669 2206
rect 7721 2210 7800 2226
rect 7832 2226 8004 2228
rect 7832 2210 7911 2226
rect 7918 2224 7948 2226
rect 7496 2188 7525 2198
rect 7539 2188 7568 2198
rect 7583 2188 7613 2202
rect 7656 2188 7699 2202
rect 7721 2198 7911 2210
rect 7976 2206 7982 2226
rect 7706 2188 7736 2198
rect 7737 2188 7895 2198
rect 7899 2188 7929 2198
rect 7933 2188 7963 2202
rect 7991 2188 8004 2226
rect 8076 2240 8105 2256
rect 8119 2240 8148 2256
rect 8163 2246 8193 2262
rect 8221 2240 8227 2288
rect 8230 2282 8249 2288
rect 8264 2282 8294 2290
rect 8230 2274 8294 2282
rect 8230 2258 8310 2274
rect 8326 2267 8388 2298
rect 8404 2267 8466 2298
rect 8535 2296 8584 2321
rect 8599 2296 8629 2312
rect 8498 2282 8528 2290
rect 8535 2288 8645 2296
rect 8498 2274 8543 2282
rect 8230 2256 8249 2258
rect 8264 2256 8310 2258
rect 8230 2240 8310 2256
rect 8337 2254 8372 2267
rect 8413 2264 8450 2267
rect 8413 2262 8455 2264
rect 8342 2251 8372 2254
rect 8351 2247 8358 2251
rect 8358 2246 8359 2247
rect 8317 2240 8327 2246
rect 8076 2232 8111 2240
rect 8076 2206 8077 2232
rect 8084 2206 8111 2232
rect 8019 2188 8049 2202
rect 8076 2198 8111 2206
rect 8113 2232 8154 2240
rect 8113 2206 8128 2232
rect 8135 2206 8154 2232
rect 8218 2228 8249 2240
rect 8264 2228 8367 2240
rect 8379 2230 8405 2256
rect 8420 2251 8450 2262
rect 8482 2258 8544 2274
rect 8482 2256 8528 2258
rect 8482 2240 8544 2256
rect 8556 2240 8562 2288
rect 8565 2280 8645 2288
rect 8565 2278 8584 2280
rect 8599 2278 8633 2280
rect 8565 2262 8645 2278
rect 8565 2240 8584 2262
rect 8599 2246 8629 2262
rect 8657 2256 8663 2330
rect 8666 2256 8685 2400
rect 8700 2256 8706 2400
rect 8715 2330 8728 2400
rect 8780 2396 8802 2400
rect 8773 2374 8802 2388
rect 8855 2374 8871 2388
rect 8909 2384 8915 2386
rect 8922 2384 9030 2400
rect 9037 2384 9043 2386
rect 9051 2384 9066 2400
rect 9132 2394 9151 2397
rect 8773 2372 8871 2374
rect 8898 2372 9066 2384
rect 9081 2374 9097 2388
rect 9132 2375 9154 2394
rect 9164 2388 9180 2389
rect 9163 2386 9180 2388
rect 9164 2381 9180 2386
rect 9154 2374 9160 2375
rect 9163 2374 9192 2381
rect 9081 2373 9192 2374
rect 9081 2372 9198 2373
rect 8757 2364 8808 2372
rect 8855 2364 8889 2372
rect 8757 2352 8782 2364
rect 8789 2352 8808 2364
rect 8862 2362 8889 2364
rect 8898 2362 9119 2372
rect 9154 2369 9160 2372
rect 8862 2358 9119 2362
rect 8757 2344 8808 2352
rect 8855 2344 9119 2358
rect 9163 2364 9198 2372
rect 8709 2296 8728 2330
rect 8773 2336 8802 2344
rect 8773 2330 8790 2336
rect 8773 2328 8807 2330
rect 8855 2328 8871 2344
rect 8872 2334 9080 2344
rect 9081 2334 9097 2344
rect 9145 2340 9160 2355
rect 9163 2352 9164 2364
rect 9171 2352 9198 2364
rect 9163 2344 9198 2352
rect 9163 2343 9192 2344
rect 8883 2330 9097 2334
rect 8898 2328 9097 2330
rect 9132 2330 9145 2340
rect 9163 2330 9180 2343
rect 9132 2328 9180 2330
rect 8774 2324 8807 2328
rect 8770 2322 8807 2324
rect 8770 2321 8837 2322
rect 8770 2316 8801 2321
rect 8807 2316 8837 2321
rect 8770 2312 8837 2316
rect 8743 2309 8837 2312
rect 8743 2302 8792 2309
rect 8743 2296 8773 2302
rect 8792 2297 8797 2302
rect 8709 2280 8789 2296
rect 8801 2288 8837 2309
rect 8898 2304 9087 2328
rect 9132 2327 9179 2328
rect 9145 2322 9179 2327
rect 8913 2301 9087 2304
rect 8906 2298 9087 2301
rect 9115 2321 9179 2322
rect 8709 2278 8728 2280
rect 8743 2278 8777 2280
rect 8709 2262 8789 2278
rect 8709 2256 8728 2262
rect 8425 2230 8528 2240
rect 8379 2228 8528 2230
rect 8549 2228 8584 2240
rect 8218 2226 8380 2228
rect 8230 2206 8249 2226
rect 8264 2224 8294 2226
rect 8113 2198 8154 2206
rect 8236 2202 8249 2206
rect 8301 2210 8380 2226
rect 8412 2226 8584 2228
rect 8412 2210 8491 2226
rect 8498 2224 8528 2226
rect 8076 2188 8105 2198
rect 8119 2188 8148 2198
rect 8163 2188 8193 2202
rect 8236 2188 8279 2202
rect 8301 2198 8491 2210
rect 8556 2206 8562 2226
rect 8286 2188 8316 2198
rect 8317 2188 8475 2198
rect 8479 2188 8509 2198
rect 8513 2188 8543 2202
rect 8571 2188 8584 2226
rect 8656 2240 8685 2256
rect 8699 2240 8728 2256
rect 8743 2246 8773 2262
rect 8801 2240 8807 2288
rect 8810 2282 8829 2288
rect 8844 2282 8874 2290
rect 8810 2274 8874 2282
rect 8810 2258 8890 2274
rect 8906 2267 8968 2298
rect 8984 2267 9046 2298
rect 9115 2296 9164 2321
rect 9179 2296 9209 2312
rect 9078 2282 9108 2290
rect 9115 2288 9225 2296
rect 9078 2274 9123 2282
rect 8810 2256 8829 2258
rect 8844 2256 8890 2258
rect 8810 2240 8890 2256
rect 8917 2254 8952 2267
rect 8993 2264 9030 2267
rect 8993 2262 9035 2264
rect 8922 2251 8952 2254
rect 8931 2247 8938 2251
rect 8938 2246 8939 2247
rect 8897 2240 8907 2246
rect 8656 2232 8691 2240
rect 8656 2206 8657 2232
rect 8664 2206 8691 2232
rect 8599 2188 8629 2202
rect 8656 2198 8691 2206
rect 8693 2232 8734 2240
rect 8693 2206 8708 2232
rect 8715 2206 8734 2232
rect 8798 2228 8829 2240
rect 8844 2228 8947 2240
rect 8959 2230 8985 2256
rect 9000 2251 9030 2262
rect 9062 2258 9124 2274
rect 9062 2256 9108 2258
rect 9062 2240 9124 2256
rect 9136 2240 9142 2288
rect 9145 2280 9225 2288
rect 9145 2278 9164 2280
rect 9179 2278 9213 2280
rect 9145 2262 9225 2278
rect 9145 2240 9164 2262
rect 9179 2246 9209 2262
rect 9237 2256 9243 2330
rect 9246 2256 9265 2400
rect 9280 2256 9286 2400
rect 9295 2330 9308 2400
rect 9360 2396 9382 2400
rect 9353 2374 9382 2388
rect 9435 2374 9451 2388
rect 9489 2384 9495 2386
rect 9502 2384 9610 2400
rect 9617 2384 9623 2386
rect 9631 2384 9646 2400
rect 9712 2394 9731 2397
rect 9353 2372 9451 2374
rect 9478 2372 9646 2384
rect 9661 2374 9677 2388
rect 9712 2375 9734 2394
rect 9744 2388 9760 2389
rect 9743 2386 9760 2388
rect 9744 2381 9760 2386
rect 9734 2374 9740 2375
rect 9743 2374 9772 2381
rect 9661 2373 9772 2374
rect 9661 2372 9778 2373
rect 9337 2364 9388 2372
rect 9435 2364 9469 2372
rect 9337 2352 9362 2364
rect 9369 2352 9388 2364
rect 9442 2362 9469 2364
rect 9478 2362 9699 2372
rect 9734 2369 9740 2372
rect 9442 2358 9699 2362
rect 9337 2344 9388 2352
rect 9435 2344 9699 2358
rect 9743 2364 9778 2372
rect 9289 2296 9308 2330
rect 9353 2336 9382 2344
rect 9353 2330 9370 2336
rect 9353 2328 9387 2330
rect 9435 2328 9451 2344
rect 9452 2334 9660 2344
rect 9661 2334 9677 2344
rect 9725 2340 9740 2355
rect 9743 2352 9744 2364
rect 9751 2352 9778 2364
rect 9743 2344 9778 2352
rect 9743 2343 9772 2344
rect 9463 2330 9677 2334
rect 9478 2328 9677 2330
rect 9712 2330 9725 2340
rect 9743 2330 9760 2343
rect 9712 2328 9760 2330
rect 9354 2324 9387 2328
rect 9350 2322 9387 2324
rect 9350 2321 9417 2322
rect 9350 2316 9381 2321
rect 9387 2316 9417 2321
rect 9350 2312 9417 2316
rect 9323 2309 9417 2312
rect 9323 2302 9372 2309
rect 9323 2296 9353 2302
rect 9372 2297 9377 2302
rect 9289 2280 9369 2296
rect 9381 2288 9417 2309
rect 9478 2304 9667 2328
rect 9712 2327 9759 2328
rect 9725 2322 9759 2327
rect 9493 2301 9667 2304
rect 9486 2298 9667 2301
rect 9695 2321 9759 2322
rect 9289 2278 9308 2280
rect 9323 2278 9357 2280
rect 9289 2262 9369 2278
rect 9289 2256 9308 2262
rect 9005 2230 9108 2240
rect 8959 2228 9108 2230
rect 9129 2228 9164 2240
rect 8798 2226 8960 2228
rect 8810 2206 8829 2226
rect 8844 2224 8874 2226
rect 8693 2198 8734 2206
rect 8816 2202 8829 2206
rect 8881 2210 8960 2226
rect 8992 2226 9164 2228
rect 8992 2210 9071 2226
rect 9078 2224 9108 2226
rect 8656 2188 8685 2198
rect 8699 2188 8728 2198
rect 8743 2188 8773 2202
rect 8816 2188 8859 2202
rect 8881 2198 9071 2210
rect 9136 2206 9142 2226
rect 8866 2188 8896 2198
rect 8897 2188 9055 2198
rect 9059 2188 9089 2198
rect 9093 2188 9123 2202
rect 9151 2188 9164 2226
rect 9236 2240 9265 2256
rect 9279 2240 9308 2256
rect 9323 2246 9353 2262
rect 9381 2240 9387 2288
rect 9390 2282 9409 2288
rect 9424 2282 9454 2290
rect 9390 2274 9454 2282
rect 9390 2258 9470 2274
rect 9486 2267 9548 2298
rect 9564 2267 9626 2298
rect 9695 2296 9744 2321
rect 9759 2296 9789 2312
rect 9658 2282 9688 2290
rect 9695 2288 9805 2296
rect 9658 2274 9703 2282
rect 9390 2256 9409 2258
rect 9424 2256 9470 2258
rect 9390 2240 9470 2256
rect 9497 2254 9532 2267
rect 9573 2264 9610 2267
rect 9573 2262 9615 2264
rect 9502 2251 9532 2254
rect 9511 2247 9518 2251
rect 9518 2246 9519 2247
rect 9477 2240 9487 2246
rect 9236 2232 9271 2240
rect 9236 2206 9237 2232
rect 9244 2206 9271 2232
rect 9179 2188 9209 2202
rect 9236 2198 9271 2206
rect 9273 2232 9314 2240
rect 9273 2206 9288 2232
rect 9295 2206 9314 2232
rect 9378 2228 9409 2240
rect 9424 2228 9527 2240
rect 9539 2230 9565 2256
rect 9580 2251 9610 2262
rect 9642 2258 9704 2274
rect 9642 2256 9688 2258
rect 9642 2240 9704 2256
rect 9716 2240 9722 2288
rect 9725 2280 9805 2288
rect 9725 2278 9744 2280
rect 9759 2278 9793 2280
rect 9725 2262 9805 2278
rect 9725 2240 9744 2262
rect 9759 2246 9789 2262
rect 9817 2256 9823 2330
rect 9826 2256 9845 2400
rect 9860 2256 9866 2400
rect 9875 2330 9888 2400
rect 9940 2396 9962 2400
rect 9933 2374 9962 2388
rect 10015 2374 10031 2388
rect 10069 2384 10075 2386
rect 10082 2384 10190 2400
rect 10197 2384 10203 2386
rect 10211 2384 10226 2400
rect 10292 2394 10311 2397
rect 9933 2372 10031 2374
rect 10058 2372 10226 2384
rect 10241 2374 10257 2388
rect 10292 2375 10314 2394
rect 10324 2388 10340 2389
rect 10323 2386 10340 2388
rect 10324 2381 10340 2386
rect 10314 2374 10320 2375
rect 10323 2374 10352 2381
rect 10241 2373 10352 2374
rect 10241 2372 10358 2373
rect 9917 2364 9968 2372
rect 10015 2364 10049 2372
rect 9917 2352 9942 2364
rect 9949 2352 9968 2364
rect 10022 2362 10049 2364
rect 10058 2362 10279 2372
rect 10314 2369 10320 2372
rect 10022 2358 10279 2362
rect 9917 2344 9968 2352
rect 10015 2344 10279 2358
rect 10323 2364 10358 2372
rect 9869 2296 9888 2330
rect 9933 2336 9962 2344
rect 9933 2330 9950 2336
rect 9933 2328 9967 2330
rect 10015 2328 10031 2344
rect 10032 2334 10240 2344
rect 10241 2334 10257 2344
rect 10305 2340 10320 2355
rect 10323 2352 10324 2364
rect 10331 2352 10358 2364
rect 10323 2344 10358 2352
rect 10323 2343 10352 2344
rect 10043 2330 10257 2334
rect 10058 2328 10257 2330
rect 10292 2330 10305 2340
rect 10323 2330 10340 2343
rect 10292 2328 10340 2330
rect 9934 2324 9967 2328
rect 9930 2322 9967 2324
rect 9930 2321 9997 2322
rect 9930 2316 9961 2321
rect 9967 2316 9997 2321
rect 9930 2312 9997 2316
rect 9903 2309 9997 2312
rect 9903 2302 9952 2309
rect 9903 2296 9933 2302
rect 9952 2297 9957 2302
rect 9869 2280 9949 2296
rect 9961 2288 9997 2309
rect 10058 2304 10247 2328
rect 10292 2327 10339 2328
rect 10305 2322 10339 2327
rect 10073 2301 10247 2304
rect 10066 2298 10247 2301
rect 10275 2321 10339 2322
rect 9869 2278 9888 2280
rect 9903 2278 9937 2280
rect 9869 2262 9949 2278
rect 9869 2256 9888 2262
rect 9585 2230 9688 2240
rect 9539 2228 9688 2230
rect 9709 2228 9744 2240
rect 9378 2226 9540 2228
rect 9390 2206 9409 2226
rect 9424 2224 9454 2226
rect 9273 2198 9314 2206
rect 9396 2202 9409 2206
rect 9461 2210 9540 2226
rect 9572 2226 9744 2228
rect 9572 2210 9651 2226
rect 9658 2224 9688 2226
rect 9236 2188 9265 2198
rect 9279 2188 9308 2198
rect 9323 2188 9353 2202
rect 9396 2188 9439 2202
rect 9461 2198 9651 2210
rect 9716 2206 9722 2226
rect 9446 2188 9476 2198
rect 9477 2188 9635 2198
rect 9639 2188 9669 2198
rect 9673 2188 9703 2202
rect 9731 2188 9744 2226
rect 9816 2240 9845 2256
rect 9859 2240 9888 2256
rect 9903 2246 9933 2262
rect 9961 2240 9967 2288
rect 9970 2282 9989 2288
rect 10004 2282 10034 2290
rect 9970 2274 10034 2282
rect 9970 2258 10050 2274
rect 10066 2267 10128 2298
rect 10144 2267 10206 2298
rect 10275 2296 10324 2321
rect 10339 2296 10369 2312
rect 10238 2282 10268 2290
rect 10275 2288 10385 2296
rect 10238 2274 10283 2282
rect 9970 2256 9989 2258
rect 10004 2256 10050 2258
rect 9970 2240 10050 2256
rect 10077 2254 10112 2267
rect 10153 2264 10190 2267
rect 10153 2262 10195 2264
rect 10082 2251 10112 2254
rect 10091 2247 10098 2251
rect 10098 2246 10099 2247
rect 10057 2240 10067 2246
rect 9816 2232 9851 2240
rect 9816 2206 9817 2232
rect 9824 2206 9851 2232
rect 9759 2188 9789 2202
rect 9816 2198 9851 2206
rect 9853 2232 9894 2240
rect 9853 2206 9868 2232
rect 9875 2206 9894 2232
rect 9958 2228 9989 2240
rect 10004 2228 10107 2240
rect 10119 2230 10145 2256
rect 10160 2251 10190 2262
rect 10222 2258 10284 2274
rect 10222 2256 10268 2258
rect 10222 2240 10284 2256
rect 10296 2240 10302 2288
rect 10305 2280 10385 2288
rect 10305 2278 10324 2280
rect 10339 2278 10373 2280
rect 10305 2262 10385 2278
rect 10305 2240 10324 2262
rect 10339 2246 10369 2262
rect 10397 2256 10403 2330
rect 10406 2256 10425 2400
rect 10440 2256 10446 2400
rect 10455 2330 10468 2400
rect 10520 2396 10542 2400
rect 10513 2374 10542 2388
rect 10595 2374 10611 2388
rect 10649 2384 10655 2386
rect 10662 2384 10770 2400
rect 10777 2384 10783 2386
rect 10791 2384 10806 2400
rect 10872 2394 10891 2397
rect 10513 2372 10611 2374
rect 10638 2372 10806 2384
rect 10821 2374 10837 2388
rect 10872 2375 10894 2394
rect 10904 2388 10920 2389
rect 10903 2386 10920 2388
rect 10904 2381 10920 2386
rect 10894 2374 10900 2375
rect 10903 2374 10932 2381
rect 10821 2373 10932 2374
rect 10821 2372 10938 2373
rect 10497 2364 10548 2372
rect 10595 2364 10629 2372
rect 10497 2352 10522 2364
rect 10529 2352 10548 2364
rect 10602 2362 10629 2364
rect 10638 2362 10859 2372
rect 10894 2369 10900 2372
rect 10602 2358 10859 2362
rect 10497 2344 10548 2352
rect 10595 2344 10859 2358
rect 10903 2364 10938 2372
rect 10449 2296 10468 2330
rect 10513 2336 10542 2344
rect 10513 2330 10530 2336
rect 10513 2328 10547 2330
rect 10595 2328 10611 2344
rect 10612 2334 10820 2344
rect 10821 2334 10837 2344
rect 10885 2340 10900 2355
rect 10903 2352 10904 2364
rect 10911 2352 10938 2364
rect 10903 2344 10938 2352
rect 10903 2343 10932 2344
rect 10623 2330 10837 2334
rect 10638 2328 10837 2330
rect 10872 2330 10885 2340
rect 10903 2330 10920 2343
rect 10872 2328 10920 2330
rect 10514 2324 10547 2328
rect 10510 2322 10547 2324
rect 10510 2321 10577 2322
rect 10510 2316 10541 2321
rect 10547 2316 10577 2321
rect 10510 2312 10577 2316
rect 10483 2309 10577 2312
rect 10483 2302 10532 2309
rect 10483 2296 10513 2302
rect 10532 2297 10537 2302
rect 10449 2280 10529 2296
rect 10541 2288 10577 2309
rect 10638 2304 10827 2328
rect 10872 2327 10919 2328
rect 10885 2322 10919 2327
rect 10653 2301 10827 2304
rect 10646 2298 10827 2301
rect 10855 2321 10919 2322
rect 10449 2278 10468 2280
rect 10483 2278 10517 2280
rect 10449 2262 10529 2278
rect 10449 2256 10468 2262
rect 10165 2230 10268 2240
rect 10119 2228 10268 2230
rect 10289 2228 10324 2240
rect 9958 2226 10120 2228
rect 9970 2206 9989 2226
rect 10004 2224 10034 2226
rect 9853 2198 9894 2206
rect 9976 2202 9989 2206
rect 10041 2210 10120 2226
rect 10152 2226 10324 2228
rect 10152 2210 10231 2226
rect 10238 2224 10268 2226
rect 9816 2188 9845 2198
rect 9859 2188 9888 2198
rect 9903 2188 9933 2202
rect 9976 2188 10019 2202
rect 10041 2198 10231 2210
rect 10296 2206 10302 2226
rect 10026 2188 10056 2198
rect 10057 2188 10215 2198
rect 10219 2188 10249 2198
rect 10253 2188 10283 2202
rect 10311 2188 10324 2226
rect 10396 2240 10425 2256
rect 10439 2240 10468 2256
rect 10483 2246 10513 2262
rect 10541 2240 10547 2288
rect 10550 2282 10569 2288
rect 10584 2282 10614 2290
rect 10550 2274 10614 2282
rect 10550 2258 10630 2274
rect 10646 2267 10708 2298
rect 10724 2267 10786 2298
rect 10855 2296 10904 2321
rect 10919 2296 10949 2312
rect 10818 2282 10848 2290
rect 10855 2288 10965 2296
rect 10818 2274 10863 2282
rect 10550 2256 10569 2258
rect 10584 2256 10630 2258
rect 10550 2240 10630 2256
rect 10657 2254 10692 2267
rect 10733 2264 10770 2267
rect 10733 2262 10775 2264
rect 10662 2251 10692 2254
rect 10671 2247 10678 2251
rect 10678 2246 10679 2247
rect 10637 2240 10647 2246
rect 10396 2232 10431 2240
rect 10396 2206 10397 2232
rect 10404 2206 10431 2232
rect 10339 2188 10369 2202
rect 10396 2198 10431 2206
rect 10433 2232 10474 2240
rect 10433 2206 10448 2232
rect 10455 2206 10474 2232
rect 10538 2228 10569 2240
rect 10584 2228 10687 2240
rect 10699 2230 10725 2256
rect 10740 2251 10770 2262
rect 10802 2258 10864 2274
rect 10802 2256 10848 2258
rect 10802 2240 10864 2256
rect 10876 2240 10882 2288
rect 10885 2280 10965 2288
rect 10885 2278 10904 2280
rect 10919 2278 10953 2280
rect 10885 2262 10965 2278
rect 10885 2240 10904 2262
rect 10919 2246 10949 2262
rect 10977 2256 10983 2330
rect 10986 2256 11005 2400
rect 11020 2256 11026 2400
rect 11035 2330 11048 2400
rect 11100 2396 11122 2400
rect 11093 2374 11122 2388
rect 11175 2374 11191 2388
rect 11229 2384 11235 2386
rect 11242 2384 11350 2400
rect 11357 2384 11363 2386
rect 11371 2384 11386 2400
rect 11452 2394 11471 2397
rect 11093 2372 11191 2374
rect 11218 2372 11386 2384
rect 11401 2374 11417 2388
rect 11452 2375 11474 2394
rect 11484 2388 11500 2389
rect 11483 2386 11500 2388
rect 11484 2381 11500 2386
rect 11474 2374 11480 2375
rect 11483 2374 11512 2381
rect 11401 2373 11512 2374
rect 11401 2372 11518 2373
rect 11077 2364 11128 2372
rect 11175 2364 11209 2372
rect 11077 2352 11102 2364
rect 11109 2352 11128 2364
rect 11182 2362 11209 2364
rect 11218 2362 11439 2372
rect 11474 2369 11480 2372
rect 11182 2358 11439 2362
rect 11077 2344 11128 2352
rect 11175 2344 11439 2358
rect 11483 2364 11518 2372
rect 11029 2296 11048 2330
rect 11093 2336 11122 2344
rect 11093 2330 11110 2336
rect 11093 2328 11127 2330
rect 11175 2328 11191 2344
rect 11192 2334 11400 2344
rect 11401 2334 11417 2344
rect 11465 2340 11480 2355
rect 11483 2352 11484 2364
rect 11491 2352 11518 2364
rect 11483 2344 11518 2352
rect 11483 2343 11512 2344
rect 11203 2330 11417 2334
rect 11218 2328 11417 2330
rect 11452 2330 11465 2340
rect 11483 2330 11500 2343
rect 11452 2328 11500 2330
rect 11094 2324 11127 2328
rect 11090 2322 11127 2324
rect 11090 2321 11157 2322
rect 11090 2316 11121 2321
rect 11127 2316 11157 2321
rect 11090 2312 11157 2316
rect 11063 2309 11157 2312
rect 11063 2302 11112 2309
rect 11063 2296 11093 2302
rect 11112 2297 11117 2302
rect 11029 2280 11109 2296
rect 11121 2288 11157 2309
rect 11218 2304 11407 2328
rect 11452 2327 11499 2328
rect 11465 2322 11499 2327
rect 11233 2301 11407 2304
rect 11226 2298 11407 2301
rect 11435 2321 11499 2322
rect 11029 2278 11048 2280
rect 11063 2278 11097 2280
rect 11029 2262 11109 2278
rect 11029 2256 11048 2262
rect 10745 2230 10848 2240
rect 10699 2228 10848 2230
rect 10869 2228 10904 2240
rect 10538 2226 10700 2228
rect 10550 2206 10569 2226
rect 10584 2224 10614 2226
rect 10433 2198 10474 2206
rect 10556 2202 10569 2206
rect 10621 2210 10700 2226
rect 10732 2226 10904 2228
rect 10732 2210 10811 2226
rect 10818 2224 10848 2226
rect 10396 2188 10425 2198
rect 10439 2188 10468 2198
rect 10483 2188 10513 2202
rect 10556 2188 10599 2202
rect 10621 2198 10811 2210
rect 10876 2206 10882 2226
rect 10606 2188 10636 2198
rect 10637 2188 10795 2198
rect 10799 2188 10829 2198
rect 10833 2188 10863 2202
rect 10891 2188 10904 2226
rect 10976 2240 11005 2256
rect 11019 2240 11048 2256
rect 11063 2246 11093 2262
rect 11121 2240 11127 2288
rect 11130 2282 11149 2288
rect 11164 2282 11194 2290
rect 11130 2274 11194 2282
rect 11130 2258 11210 2274
rect 11226 2267 11288 2298
rect 11304 2267 11366 2298
rect 11435 2296 11484 2321
rect 11499 2296 11529 2312
rect 11398 2282 11428 2290
rect 11435 2288 11545 2296
rect 11398 2274 11443 2282
rect 11130 2256 11149 2258
rect 11164 2256 11210 2258
rect 11130 2240 11210 2256
rect 11237 2254 11272 2267
rect 11313 2264 11350 2267
rect 11313 2262 11355 2264
rect 11242 2251 11272 2254
rect 11251 2247 11258 2251
rect 11258 2246 11259 2247
rect 11217 2240 11227 2246
rect 10976 2232 11011 2240
rect 10976 2206 10977 2232
rect 10984 2206 11011 2232
rect 10919 2188 10949 2202
rect 10976 2198 11011 2206
rect 11013 2232 11054 2240
rect 11013 2206 11028 2232
rect 11035 2206 11054 2232
rect 11118 2228 11149 2240
rect 11164 2228 11267 2240
rect 11279 2230 11305 2256
rect 11320 2251 11350 2262
rect 11382 2258 11444 2274
rect 11382 2256 11428 2258
rect 11382 2240 11444 2256
rect 11456 2240 11462 2288
rect 11465 2280 11545 2288
rect 11465 2278 11484 2280
rect 11499 2278 11533 2280
rect 11465 2262 11545 2278
rect 11465 2240 11484 2262
rect 11499 2246 11529 2262
rect 11557 2256 11563 2330
rect 11566 2256 11585 2400
rect 11600 2256 11606 2400
rect 11615 2330 11628 2400
rect 11680 2396 11702 2400
rect 11673 2374 11702 2388
rect 11755 2374 11771 2388
rect 11809 2384 11815 2386
rect 11822 2384 11930 2400
rect 11937 2384 11943 2386
rect 11951 2384 11966 2400
rect 12032 2394 12051 2397
rect 11673 2372 11771 2374
rect 11798 2372 11966 2384
rect 11981 2374 11997 2388
rect 12032 2375 12054 2394
rect 12064 2388 12080 2389
rect 12063 2386 12080 2388
rect 12064 2381 12080 2386
rect 12054 2374 12060 2375
rect 12063 2374 12092 2381
rect 11981 2373 12092 2374
rect 11981 2372 12098 2373
rect 11657 2364 11708 2372
rect 11755 2364 11789 2372
rect 11657 2352 11682 2364
rect 11689 2352 11708 2364
rect 11762 2362 11789 2364
rect 11798 2362 12019 2372
rect 12054 2369 12060 2372
rect 11762 2358 12019 2362
rect 11657 2344 11708 2352
rect 11755 2344 12019 2358
rect 12063 2364 12098 2372
rect 11609 2296 11628 2330
rect 11673 2336 11702 2344
rect 11673 2330 11690 2336
rect 11673 2328 11707 2330
rect 11755 2328 11771 2344
rect 11772 2334 11980 2344
rect 11981 2334 11997 2344
rect 12045 2340 12060 2355
rect 12063 2352 12064 2364
rect 12071 2352 12098 2364
rect 12063 2344 12098 2352
rect 12063 2343 12092 2344
rect 11783 2330 11997 2334
rect 11798 2328 11997 2330
rect 12032 2330 12045 2340
rect 12063 2330 12080 2343
rect 12032 2328 12080 2330
rect 11674 2324 11707 2328
rect 11670 2322 11707 2324
rect 11670 2321 11737 2322
rect 11670 2316 11701 2321
rect 11707 2316 11737 2321
rect 11670 2312 11737 2316
rect 11643 2309 11737 2312
rect 11643 2302 11692 2309
rect 11643 2296 11673 2302
rect 11692 2297 11697 2302
rect 11609 2280 11689 2296
rect 11701 2288 11737 2309
rect 11798 2304 11987 2328
rect 12032 2327 12079 2328
rect 12045 2322 12079 2327
rect 11813 2301 11987 2304
rect 11806 2298 11987 2301
rect 12015 2321 12079 2322
rect 11609 2278 11628 2280
rect 11643 2278 11677 2280
rect 11609 2262 11689 2278
rect 11609 2256 11628 2262
rect 11325 2230 11428 2240
rect 11279 2228 11428 2230
rect 11449 2228 11484 2240
rect 11118 2226 11280 2228
rect 11130 2206 11149 2226
rect 11164 2224 11194 2226
rect 11013 2198 11054 2206
rect 11136 2202 11149 2206
rect 11201 2210 11280 2226
rect 11312 2226 11484 2228
rect 11312 2210 11391 2226
rect 11398 2224 11428 2226
rect 10976 2188 11005 2198
rect 11019 2188 11048 2198
rect 11063 2188 11093 2202
rect 11136 2188 11179 2202
rect 11201 2198 11391 2210
rect 11456 2206 11462 2226
rect 11186 2188 11216 2198
rect 11217 2188 11375 2198
rect 11379 2188 11409 2198
rect 11413 2188 11443 2202
rect 11471 2188 11484 2226
rect 11556 2240 11585 2256
rect 11599 2240 11628 2256
rect 11643 2246 11673 2262
rect 11701 2240 11707 2288
rect 11710 2282 11729 2288
rect 11744 2282 11774 2290
rect 11710 2274 11774 2282
rect 11710 2258 11790 2274
rect 11806 2267 11868 2298
rect 11884 2267 11946 2298
rect 12015 2296 12064 2321
rect 12079 2296 12109 2312
rect 11978 2282 12008 2290
rect 12015 2288 12125 2296
rect 11978 2274 12023 2282
rect 11710 2256 11729 2258
rect 11744 2256 11790 2258
rect 11710 2240 11790 2256
rect 11817 2254 11852 2267
rect 11893 2264 11930 2267
rect 11893 2262 11935 2264
rect 11822 2251 11852 2254
rect 11831 2247 11838 2251
rect 11838 2246 11839 2247
rect 11797 2240 11807 2246
rect 11556 2232 11591 2240
rect 11556 2206 11557 2232
rect 11564 2206 11591 2232
rect 11499 2188 11529 2202
rect 11556 2198 11591 2206
rect 11593 2232 11634 2240
rect 11593 2206 11608 2232
rect 11615 2206 11634 2232
rect 11698 2228 11729 2240
rect 11744 2228 11847 2240
rect 11859 2230 11885 2256
rect 11900 2251 11930 2262
rect 11962 2258 12024 2274
rect 11962 2256 12008 2258
rect 11962 2240 12024 2256
rect 12036 2240 12042 2288
rect 12045 2280 12125 2288
rect 12045 2278 12064 2280
rect 12079 2278 12113 2280
rect 12045 2262 12125 2278
rect 12045 2240 12064 2262
rect 12079 2246 12109 2262
rect 12137 2256 12143 2330
rect 12146 2256 12165 2400
rect 12180 2256 12186 2400
rect 12195 2330 12208 2400
rect 12260 2396 12282 2400
rect 12253 2374 12282 2388
rect 12335 2374 12351 2388
rect 12389 2384 12395 2386
rect 12402 2384 12510 2400
rect 12517 2384 12523 2386
rect 12531 2384 12546 2400
rect 12612 2394 12631 2397
rect 12253 2372 12351 2374
rect 12378 2372 12546 2384
rect 12561 2374 12577 2388
rect 12612 2375 12634 2394
rect 12644 2388 12660 2389
rect 12643 2386 12660 2388
rect 12644 2381 12660 2386
rect 12634 2374 12640 2375
rect 12643 2374 12672 2381
rect 12561 2373 12672 2374
rect 12561 2372 12678 2373
rect 12237 2364 12288 2372
rect 12335 2364 12369 2372
rect 12237 2352 12262 2364
rect 12269 2352 12288 2364
rect 12342 2362 12369 2364
rect 12378 2362 12599 2372
rect 12634 2369 12640 2372
rect 12342 2358 12599 2362
rect 12237 2344 12288 2352
rect 12335 2344 12599 2358
rect 12643 2364 12678 2372
rect 12189 2296 12208 2330
rect 12253 2336 12282 2344
rect 12253 2330 12270 2336
rect 12253 2328 12287 2330
rect 12335 2328 12351 2344
rect 12352 2334 12560 2344
rect 12561 2334 12577 2344
rect 12625 2340 12640 2355
rect 12643 2352 12644 2364
rect 12651 2352 12678 2364
rect 12643 2344 12678 2352
rect 12643 2343 12672 2344
rect 12363 2330 12577 2334
rect 12378 2328 12577 2330
rect 12612 2330 12625 2340
rect 12643 2330 12660 2343
rect 12612 2328 12660 2330
rect 12254 2324 12287 2328
rect 12250 2322 12287 2324
rect 12250 2321 12317 2322
rect 12250 2316 12281 2321
rect 12287 2316 12317 2321
rect 12250 2312 12317 2316
rect 12223 2309 12317 2312
rect 12223 2302 12272 2309
rect 12223 2296 12253 2302
rect 12272 2297 12277 2302
rect 12189 2280 12269 2296
rect 12281 2288 12317 2309
rect 12378 2304 12567 2328
rect 12612 2327 12659 2328
rect 12625 2322 12659 2327
rect 12393 2301 12567 2304
rect 12386 2298 12567 2301
rect 12595 2321 12659 2322
rect 12189 2278 12208 2280
rect 12223 2278 12257 2280
rect 12189 2262 12269 2278
rect 12189 2256 12208 2262
rect 11905 2230 12008 2240
rect 11859 2228 12008 2230
rect 12029 2228 12064 2240
rect 11698 2226 11860 2228
rect 11710 2206 11729 2226
rect 11744 2224 11774 2226
rect 11593 2198 11634 2206
rect 11716 2202 11729 2206
rect 11781 2210 11860 2226
rect 11892 2226 12064 2228
rect 11892 2210 11971 2226
rect 11978 2224 12008 2226
rect 11556 2188 11585 2198
rect 11599 2188 11628 2198
rect 11643 2188 11673 2202
rect 11716 2188 11759 2202
rect 11781 2198 11971 2210
rect 12036 2206 12042 2226
rect 11766 2188 11796 2198
rect 11797 2188 11955 2198
rect 11959 2188 11989 2198
rect 11993 2188 12023 2202
rect 12051 2188 12064 2226
rect 12136 2240 12165 2256
rect 12179 2240 12208 2256
rect 12223 2246 12253 2262
rect 12281 2240 12287 2288
rect 12290 2282 12309 2288
rect 12324 2282 12354 2290
rect 12290 2274 12354 2282
rect 12290 2258 12370 2274
rect 12386 2267 12448 2298
rect 12464 2267 12526 2298
rect 12595 2296 12644 2321
rect 12659 2296 12689 2312
rect 12558 2282 12588 2290
rect 12595 2288 12705 2296
rect 12558 2274 12603 2282
rect 12290 2256 12309 2258
rect 12324 2256 12370 2258
rect 12290 2240 12370 2256
rect 12397 2254 12432 2267
rect 12473 2264 12510 2267
rect 12473 2262 12515 2264
rect 12402 2251 12432 2254
rect 12411 2247 12418 2251
rect 12418 2246 12419 2247
rect 12377 2240 12387 2246
rect 12136 2232 12171 2240
rect 12136 2206 12137 2232
rect 12144 2206 12171 2232
rect 12079 2188 12109 2202
rect 12136 2198 12171 2206
rect 12173 2232 12214 2240
rect 12173 2206 12188 2232
rect 12195 2206 12214 2232
rect 12278 2228 12309 2240
rect 12324 2228 12427 2240
rect 12439 2230 12465 2256
rect 12480 2251 12510 2262
rect 12542 2258 12604 2274
rect 12542 2256 12588 2258
rect 12542 2240 12604 2256
rect 12616 2240 12622 2288
rect 12625 2280 12705 2288
rect 12625 2278 12644 2280
rect 12659 2278 12693 2280
rect 12625 2262 12705 2278
rect 12625 2240 12644 2262
rect 12659 2246 12689 2262
rect 12717 2256 12723 2330
rect 12726 2256 12745 2400
rect 12760 2256 12766 2400
rect 12775 2330 12788 2400
rect 12840 2396 12862 2400
rect 12833 2374 12862 2388
rect 12915 2374 12931 2388
rect 12969 2384 12975 2386
rect 12982 2384 13090 2400
rect 13097 2384 13103 2386
rect 13111 2384 13126 2400
rect 13192 2394 13211 2397
rect 12833 2372 12931 2374
rect 12958 2372 13126 2384
rect 13141 2374 13157 2388
rect 13192 2375 13214 2394
rect 13224 2388 13240 2389
rect 13223 2386 13240 2388
rect 13224 2381 13240 2386
rect 13214 2374 13220 2375
rect 13223 2374 13252 2381
rect 13141 2373 13252 2374
rect 13141 2372 13258 2373
rect 12817 2364 12868 2372
rect 12915 2364 12949 2372
rect 12817 2352 12842 2364
rect 12849 2352 12868 2364
rect 12922 2362 12949 2364
rect 12958 2362 13179 2372
rect 13214 2369 13220 2372
rect 12922 2358 13179 2362
rect 12817 2344 12868 2352
rect 12915 2344 13179 2358
rect 13223 2364 13258 2372
rect 12769 2296 12788 2330
rect 12833 2336 12862 2344
rect 12833 2330 12850 2336
rect 12833 2328 12867 2330
rect 12915 2328 12931 2344
rect 12932 2334 13140 2344
rect 13141 2334 13157 2344
rect 13205 2340 13220 2355
rect 13223 2352 13224 2364
rect 13231 2352 13258 2364
rect 13223 2344 13258 2352
rect 13223 2343 13252 2344
rect 12943 2330 13157 2334
rect 12958 2328 13157 2330
rect 13192 2330 13205 2340
rect 13223 2330 13240 2343
rect 13192 2328 13240 2330
rect 12834 2324 12867 2328
rect 12830 2322 12867 2324
rect 12830 2321 12897 2322
rect 12830 2316 12861 2321
rect 12867 2316 12897 2321
rect 12830 2312 12897 2316
rect 12803 2309 12897 2312
rect 12803 2302 12852 2309
rect 12803 2296 12833 2302
rect 12852 2297 12857 2302
rect 12769 2280 12849 2296
rect 12861 2288 12897 2309
rect 12958 2304 13147 2328
rect 13192 2327 13239 2328
rect 13205 2322 13239 2327
rect 12973 2301 13147 2304
rect 12966 2298 13147 2301
rect 13175 2321 13239 2322
rect 12769 2278 12788 2280
rect 12803 2278 12837 2280
rect 12769 2262 12849 2278
rect 12769 2256 12788 2262
rect 12485 2230 12588 2240
rect 12439 2228 12588 2230
rect 12609 2228 12644 2240
rect 12278 2226 12440 2228
rect 12290 2206 12309 2226
rect 12324 2224 12354 2226
rect 12173 2198 12214 2206
rect 12296 2202 12309 2206
rect 12361 2210 12440 2226
rect 12472 2226 12644 2228
rect 12472 2210 12551 2226
rect 12558 2224 12588 2226
rect 12136 2188 12165 2198
rect 12179 2188 12208 2198
rect 12223 2188 12253 2202
rect 12296 2188 12339 2202
rect 12361 2198 12551 2210
rect 12616 2206 12622 2226
rect 12346 2188 12376 2198
rect 12377 2188 12535 2198
rect 12539 2188 12569 2198
rect 12573 2188 12603 2202
rect 12631 2188 12644 2226
rect 12716 2240 12745 2256
rect 12759 2240 12788 2256
rect 12803 2246 12833 2262
rect 12861 2240 12867 2288
rect 12870 2282 12889 2288
rect 12904 2282 12934 2290
rect 12870 2274 12934 2282
rect 12870 2258 12950 2274
rect 12966 2267 13028 2298
rect 13044 2267 13106 2298
rect 13175 2296 13224 2321
rect 13239 2296 13269 2312
rect 13138 2282 13168 2290
rect 13175 2288 13285 2296
rect 13138 2274 13183 2282
rect 12870 2256 12889 2258
rect 12904 2256 12950 2258
rect 12870 2240 12950 2256
rect 12977 2254 13012 2267
rect 13053 2264 13090 2267
rect 13053 2262 13095 2264
rect 12982 2251 13012 2254
rect 12991 2247 12998 2251
rect 12998 2246 12999 2247
rect 12957 2240 12967 2246
rect 12716 2232 12751 2240
rect 12716 2206 12717 2232
rect 12724 2206 12751 2232
rect 12659 2188 12689 2202
rect 12716 2198 12751 2206
rect 12753 2232 12794 2240
rect 12753 2206 12768 2232
rect 12775 2206 12794 2232
rect 12858 2228 12889 2240
rect 12904 2228 13007 2240
rect 13019 2230 13045 2256
rect 13060 2251 13090 2262
rect 13122 2258 13184 2274
rect 13122 2256 13168 2258
rect 13122 2240 13184 2256
rect 13196 2240 13202 2288
rect 13205 2280 13285 2288
rect 13205 2278 13224 2280
rect 13239 2278 13273 2280
rect 13205 2262 13285 2278
rect 13205 2240 13224 2262
rect 13239 2246 13269 2262
rect 13297 2256 13303 2330
rect 13306 2256 13325 2400
rect 13340 2256 13346 2400
rect 13355 2330 13368 2400
rect 13420 2396 13442 2400
rect 13413 2374 13442 2388
rect 13495 2374 13511 2388
rect 13549 2384 13555 2386
rect 13562 2384 13670 2400
rect 13677 2384 13683 2386
rect 13691 2384 13706 2400
rect 13772 2394 13791 2397
rect 13413 2372 13511 2374
rect 13538 2372 13706 2384
rect 13721 2374 13737 2388
rect 13772 2375 13794 2394
rect 13804 2388 13820 2389
rect 13803 2386 13820 2388
rect 13804 2381 13820 2386
rect 13794 2374 13800 2375
rect 13803 2374 13832 2381
rect 13721 2373 13832 2374
rect 13721 2372 13838 2373
rect 13397 2364 13448 2372
rect 13495 2364 13529 2372
rect 13397 2352 13422 2364
rect 13429 2352 13448 2364
rect 13502 2362 13529 2364
rect 13538 2362 13759 2372
rect 13794 2369 13800 2372
rect 13502 2358 13759 2362
rect 13397 2344 13448 2352
rect 13495 2344 13759 2358
rect 13803 2364 13838 2372
rect 13349 2296 13368 2330
rect 13413 2336 13442 2344
rect 13413 2330 13430 2336
rect 13413 2328 13447 2330
rect 13495 2328 13511 2344
rect 13512 2334 13720 2344
rect 13721 2334 13737 2344
rect 13785 2340 13800 2355
rect 13803 2352 13804 2364
rect 13811 2352 13838 2364
rect 13803 2344 13838 2352
rect 13803 2343 13832 2344
rect 13523 2330 13737 2334
rect 13538 2328 13737 2330
rect 13772 2330 13785 2340
rect 13803 2330 13820 2343
rect 13772 2328 13820 2330
rect 13414 2324 13447 2328
rect 13410 2322 13447 2324
rect 13410 2321 13477 2322
rect 13410 2316 13441 2321
rect 13447 2316 13477 2321
rect 13410 2312 13477 2316
rect 13383 2309 13477 2312
rect 13383 2302 13432 2309
rect 13383 2296 13413 2302
rect 13432 2297 13437 2302
rect 13349 2280 13429 2296
rect 13441 2288 13477 2309
rect 13538 2304 13727 2328
rect 13772 2327 13819 2328
rect 13785 2322 13819 2327
rect 13553 2301 13727 2304
rect 13546 2298 13727 2301
rect 13755 2321 13819 2322
rect 13349 2278 13368 2280
rect 13383 2278 13417 2280
rect 13349 2262 13429 2278
rect 13349 2256 13368 2262
rect 13065 2230 13168 2240
rect 13019 2228 13168 2230
rect 13189 2228 13224 2240
rect 12858 2226 13020 2228
rect 12870 2206 12889 2226
rect 12904 2224 12934 2226
rect 12753 2198 12794 2206
rect 12876 2202 12889 2206
rect 12941 2210 13020 2226
rect 13052 2226 13224 2228
rect 13052 2210 13131 2226
rect 13138 2224 13168 2226
rect 12716 2188 12745 2198
rect 12759 2188 12788 2198
rect 12803 2188 12833 2202
rect 12876 2188 12919 2202
rect 12941 2198 13131 2210
rect 13196 2206 13202 2226
rect 12926 2188 12956 2198
rect 12957 2188 13115 2198
rect 13119 2188 13149 2198
rect 13153 2188 13183 2202
rect 13211 2188 13224 2226
rect 13296 2240 13325 2256
rect 13339 2240 13368 2256
rect 13383 2246 13413 2262
rect 13441 2240 13447 2288
rect 13450 2282 13469 2288
rect 13484 2282 13514 2290
rect 13450 2274 13514 2282
rect 13450 2258 13530 2274
rect 13546 2267 13608 2298
rect 13624 2267 13686 2298
rect 13755 2296 13804 2321
rect 13819 2296 13849 2312
rect 13718 2282 13748 2290
rect 13755 2288 13865 2296
rect 13718 2274 13763 2282
rect 13450 2256 13469 2258
rect 13484 2256 13530 2258
rect 13450 2240 13530 2256
rect 13557 2254 13592 2267
rect 13633 2264 13670 2267
rect 13633 2262 13675 2264
rect 13562 2251 13592 2254
rect 13571 2247 13578 2251
rect 13578 2246 13579 2247
rect 13537 2240 13547 2246
rect 13296 2232 13331 2240
rect 13296 2206 13297 2232
rect 13304 2206 13331 2232
rect 13239 2188 13269 2202
rect 13296 2198 13331 2206
rect 13333 2232 13374 2240
rect 13333 2206 13348 2232
rect 13355 2206 13374 2232
rect 13438 2228 13469 2240
rect 13484 2228 13587 2240
rect 13599 2230 13625 2256
rect 13640 2251 13670 2262
rect 13702 2258 13764 2274
rect 13702 2256 13748 2258
rect 13702 2240 13764 2256
rect 13776 2240 13782 2288
rect 13785 2280 13865 2288
rect 13785 2278 13804 2280
rect 13819 2278 13853 2280
rect 13785 2262 13865 2278
rect 13785 2240 13804 2262
rect 13819 2246 13849 2262
rect 13877 2256 13883 2330
rect 13886 2256 13905 2400
rect 13920 2256 13926 2400
rect 13935 2330 13948 2400
rect 14000 2396 14022 2400
rect 13993 2374 14022 2388
rect 14075 2374 14091 2388
rect 14129 2384 14135 2386
rect 14142 2384 14250 2400
rect 14257 2384 14263 2386
rect 14271 2384 14286 2400
rect 14352 2394 14371 2397
rect 13993 2372 14091 2374
rect 14118 2372 14286 2384
rect 14301 2374 14317 2388
rect 14352 2375 14374 2394
rect 14384 2388 14400 2389
rect 14383 2386 14400 2388
rect 14384 2381 14400 2386
rect 14374 2374 14380 2375
rect 14383 2374 14412 2381
rect 14301 2373 14412 2374
rect 14301 2372 14418 2373
rect 13977 2364 14028 2372
rect 14075 2364 14109 2372
rect 13977 2352 14002 2364
rect 14009 2352 14028 2364
rect 14082 2362 14109 2364
rect 14118 2362 14339 2372
rect 14374 2369 14380 2372
rect 14082 2358 14339 2362
rect 13977 2344 14028 2352
rect 14075 2344 14339 2358
rect 14383 2364 14418 2372
rect 13929 2296 13948 2330
rect 13993 2336 14022 2344
rect 13993 2330 14010 2336
rect 13993 2328 14027 2330
rect 14075 2328 14091 2344
rect 14092 2334 14300 2344
rect 14301 2334 14317 2344
rect 14365 2340 14380 2355
rect 14383 2352 14384 2364
rect 14391 2352 14418 2364
rect 14383 2344 14418 2352
rect 14383 2343 14412 2344
rect 14103 2330 14317 2334
rect 14118 2328 14317 2330
rect 14352 2330 14365 2340
rect 14383 2330 14400 2343
rect 14352 2328 14400 2330
rect 13994 2324 14027 2328
rect 13990 2322 14027 2324
rect 13990 2321 14057 2322
rect 13990 2316 14021 2321
rect 14027 2316 14057 2321
rect 13990 2312 14057 2316
rect 13963 2309 14057 2312
rect 13963 2302 14012 2309
rect 13963 2296 13993 2302
rect 14012 2297 14017 2302
rect 13929 2280 14009 2296
rect 14021 2288 14057 2309
rect 14118 2304 14307 2328
rect 14352 2327 14399 2328
rect 14365 2322 14399 2327
rect 14133 2301 14307 2304
rect 14126 2298 14307 2301
rect 14335 2321 14399 2322
rect 13929 2278 13948 2280
rect 13963 2278 13997 2280
rect 13929 2262 14009 2278
rect 13929 2256 13948 2262
rect 13645 2230 13748 2240
rect 13599 2228 13748 2230
rect 13769 2228 13804 2240
rect 13438 2226 13600 2228
rect 13450 2206 13469 2226
rect 13484 2224 13514 2226
rect 13333 2198 13374 2206
rect 13456 2202 13469 2206
rect 13521 2210 13600 2226
rect 13632 2226 13804 2228
rect 13632 2210 13711 2226
rect 13718 2224 13748 2226
rect 13296 2188 13325 2198
rect 13339 2188 13368 2198
rect 13383 2188 13413 2202
rect 13456 2188 13499 2202
rect 13521 2198 13711 2210
rect 13776 2206 13782 2226
rect 13506 2188 13536 2198
rect 13537 2188 13695 2198
rect 13699 2188 13729 2198
rect 13733 2188 13763 2202
rect 13791 2188 13804 2226
rect 13876 2240 13905 2256
rect 13919 2240 13948 2256
rect 13963 2246 13993 2262
rect 14021 2240 14027 2288
rect 14030 2282 14049 2288
rect 14064 2282 14094 2290
rect 14030 2274 14094 2282
rect 14030 2258 14110 2274
rect 14126 2267 14188 2298
rect 14204 2267 14266 2298
rect 14335 2296 14384 2321
rect 14399 2296 14429 2312
rect 14298 2282 14328 2290
rect 14335 2288 14445 2296
rect 14298 2274 14343 2282
rect 14030 2256 14049 2258
rect 14064 2256 14110 2258
rect 14030 2240 14110 2256
rect 14137 2254 14172 2267
rect 14213 2264 14250 2267
rect 14213 2262 14255 2264
rect 14142 2251 14172 2254
rect 14151 2247 14158 2251
rect 14158 2246 14159 2247
rect 14117 2240 14127 2246
rect 13876 2232 13911 2240
rect 13876 2206 13877 2232
rect 13884 2206 13911 2232
rect 13819 2188 13849 2202
rect 13876 2198 13911 2206
rect 13913 2232 13954 2240
rect 13913 2206 13928 2232
rect 13935 2206 13954 2232
rect 14018 2228 14049 2240
rect 14064 2228 14167 2240
rect 14179 2230 14205 2256
rect 14220 2251 14250 2262
rect 14282 2258 14344 2274
rect 14282 2256 14328 2258
rect 14282 2240 14344 2256
rect 14356 2240 14362 2288
rect 14365 2280 14445 2288
rect 14365 2278 14384 2280
rect 14399 2278 14433 2280
rect 14365 2262 14445 2278
rect 14365 2240 14384 2262
rect 14399 2246 14429 2262
rect 14457 2256 14463 2330
rect 14466 2256 14485 2400
rect 14500 2256 14506 2400
rect 14515 2330 14528 2400
rect 14580 2396 14602 2400
rect 14573 2374 14602 2388
rect 14655 2374 14671 2388
rect 14709 2384 14715 2386
rect 14722 2384 14830 2400
rect 14837 2384 14843 2386
rect 14851 2384 14866 2400
rect 14932 2394 14951 2397
rect 14573 2372 14671 2374
rect 14698 2372 14866 2384
rect 14881 2374 14897 2388
rect 14932 2375 14954 2394
rect 14964 2388 14980 2389
rect 14963 2386 14980 2388
rect 14964 2381 14980 2386
rect 14954 2374 14960 2375
rect 14963 2374 14992 2381
rect 14881 2373 14992 2374
rect 14881 2372 14998 2373
rect 14557 2364 14608 2372
rect 14655 2364 14689 2372
rect 14557 2352 14582 2364
rect 14589 2352 14608 2364
rect 14662 2362 14689 2364
rect 14698 2362 14919 2372
rect 14954 2369 14960 2372
rect 14662 2358 14919 2362
rect 14557 2344 14608 2352
rect 14655 2344 14919 2358
rect 14963 2364 14998 2372
rect 14509 2296 14528 2330
rect 14573 2336 14602 2344
rect 14573 2330 14590 2336
rect 14573 2328 14607 2330
rect 14655 2328 14671 2344
rect 14672 2334 14880 2344
rect 14881 2334 14897 2344
rect 14945 2340 14960 2355
rect 14963 2352 14964 2364
rect 14971 2352 14998 2364
rect 14963 2344 14998 2352
rect 14963 2343 14992 2344
rect 14683 2330 14897 2334
rect 14698 2328 14897 2330
rect 14932 2330 14945 2340
rect 14963 2330 14980 2343
rect 14932 2328 14980 2330
rect 14574 2324 14607 2328
rect 14570 2322 14607 2324
rect 14570 2321 14637 2322
rect 14570 2316 14601 2321
rect 14607 2316 14637 2321
rect 14570 2312 14637 2316
rect 14543 2309 14637 2312
rect 14543 2302 14592 2309
rect 14543 2296 14573 2302
rect 14592 2297 14597 2302
rect 14509 2280 14589 2296
rect 14601 2288 14637 2309
rect 14698 2304 14887 2328
rect 14932 2327 14979 2328
rect 14945 2322 14979 2327
rect 14713 2301 14887 2304
rect 14706 2298 14887 2301
rect 14915 2321 14979 2322
rect 14509 2278 14528 2280
rect 14543 2278 14577 2280
rect 14509 2262 14589 2278
rect 14509 2256 14528 2262
rect 14225 2230 14328 2240
rect 14179 2228 14328 2230
rect 14349 2228 14384 2240
rect 14018 2226 14180 2228
rect 14030 2206 14049 2226
rect 14064 2224 14094 2226
rect 13913 2198 13954 2206
rect 14036 2202 14049 2206
rect 14101 2210 14180 2226
rect 14212 2226 14384 2228
rect 14212 2210 14291 2226
rect 14298 2224 14328 2226
rect 13876 2188 13905 2198
rect 13919 2188 13948 2198
rect 13963 2188 13993 2202
rect 14036 2188 14079 2202
rect 14101 2198 14291 2210
rect 14356 2206 14362 2226
rect 14086 2188 14116 2198
rect 14117 2188 14275 2198
rect 14279 2188 14309 2198
rect 14313 2188 14343 2202
rect 14371 2188 14384 2226
rect 14456 2240 14485 2256
rect 14499 2240 14528 2256
rect 14543 2246 14573 2262
rect 14601 2240 14607 2288
rect 14610 2282 14629 2288
rect 14644 2282 14674 2290
rect 14610 2274 14674 2282
rect 14610 2258 14690 2274
rect 14706 2267 14768 2298
rect 14784 2267 14846 2298
rect 14915 2296 14964 2321
rect 14979 2296 15009 2312
rect 14878 2282 14908 2290
rect 14915 2288 15025 2296
rect 14878 2274 14923 2282
rect 14610 2256 14629 2258
rect 14644 2256 14690 2258
rect 14610 2240 14690 2256
rect 14717 2254 14752 2267
rect 14793 2264 14830 2267
rect 14793 2262 14835 2264
rect 14722 2251 14752 2254
rect 14731 2247 14738 2251
rect 14738 2246 14739 2247
rect 14697 2240 14707 2246
rect 14456 2232 14491 2240
rect 14456 2206 14457 2232
rect 14464 2206 14491 2232
rect 14399 2188 14429 2202
rect 14456 2198 14491 2206
rect 14493 2232 14534 2240
rect 14493 2206 14508 2232
rect 14515 2206 14534 2232
rect 14598 2228 14629 2240
rect 14644 2228 14747 2240
rect 14759 2230 14785 2256
rect 14800 2251 14830 2262
rect 14862 2258 14924 2274
rect 14862 2256 14908 2258
rect 14862 2240 14924 2256
rect 14936 2240 14942 2288
rect 14945 2280 15025 2288
rect 14945 2278 14964 2280
rect 14979 2278 15013 2280
rect 14945 2262 15025 2278
rect 14945 2240 14964 2262
rect 14979 2246 15009 2262
rect 15037 2256 15043 2330
rect 15046 2256 15065 2400
rect 15080 2256 15086 2400
rect 15095 2330 15108 2400
rect 15160 2396 15182 2400
rect 15153 2374 15182 2388
rect 15235 2374 15251 2388
rect 15289 2384 15295 2386
rect 15302 2384 15410 2400
rect 15417 2384 15423 2386
rect 15431 2384 15446 2400
rect 15512 2394 15531 2397
rect 15153 2372 15251 2374
rect 15278 2372 15446 2384
rect 15461 2374 15477 2388
rect 15512 2375 15534 2394
rect 15544 2388 15560 2389
rect 15543 2386 15560 2388
rect 15544 2381 15560 2386
rect 15534 2374 15540 2375
rect 15543 2374 15572 2381
rect 15461 2373 15572 2374
rect 15461 2372 15578 2373
rect 15137 2364 15188 2372
rect 15235 2364 15269 2372
rect 15137 2352 15162 2364
rect 15169 2352 15188 2364
rect 15242 2362 15269 2364
rect 15278 2362 15499 2372
rect 15534 2369 15540 2372
rect 15242 2358 15499 2362
rect 15137 2344 15188 2352
rect 15235 2344 15499 2358
rect 15543 2364 15578 2372
rect 15089 2296 15108 2330
rect 15153 2336 15182 2344
rect 15153 2330 15170 2336
rect 15153 2328 15187 2330
rect 15235 2328 15251 2344
rect 15252 2334 15460 2344
rect 15461 2334 15477 2344
rect 15525 2340 15540 2355
rect 15543 2352 15544 2364
rect 15551 2352 15578 2364
rect 15543 2344 15578 2352
rect 15543 2343 15572 2344
rect 15263 2330 15477 2334
rect 15278 2328 15477 2330
rect 15512 2330 15525 2340
rect 15543 2330 15560 2343
rect 15512 2328 15560 2330
rect 15154 2324 15187 2328
rect 15150 2322 15187 2324
rect 15150 2321 15217 2322
rect 15150 2316 15181 2321
rect 15187 2316 15217 2321
rect 15150 2312 15217 2316
rect 15123 2309 15217 2312
rect 15123 2302 15172 2309
rect 15123 2296 15153 2302
rect 15172 2297 15177 2302
rect 15089 2280 15169 2296
rect 15181 2288 15217 2309
rect 15278 2304 15467 2328
rect 15512 2327 15559 2328
rect 15525 2322 15559 2327
rect 15293 2301 15467 2304
rect 15286 2298 15467 2301
rect 15495 2321 15559 2322
rect 15089 2278 15108 2280
rect 15123 2278 15157 2280
rect 15089 2262 15169 2278
rect 15089 2256 15108 2262
rect 14805 2230 14908 2240
rect 14759 2228 14908 2230
rect 14929 2228 14964 2240
rect 14598 2226 14760 2228
rect 14610 2206 14629 2226
rect 14644 2224 14674 2226
rect 14493 2198 14534 2206
rect 14616 2202 14629 2206
rect 14681 2210 14760 2226
rect 14792 2226 14964 2228
rect 14792 2210 14871 2226
rect 14878 2224 14908 2226
rect 14456 2188 14485 2198
rect 14499 2188 14528 2198
rect 14543 2188 14573 2202
rect 14616 2188 14659 2202
rect 14681 2198 14871 2210
rect 14936 2206 14942 2226
rect 14666 2188 14696 2198
rect 14697 2188 14855 2198
rect 14859 2188 14889 2198
rect 14893 2188 14923 2202
rect 14951 2188 14964 2226
rect 15036 2240 15065 2256
rect 15079 2240 15108 2256
rect 15123 2246 15153 2262
rect 15181 2240 15187 2288
rect 15190 2282 15209 2288
rect 15224 2282 15254 2290
rect 15190 2274 15254 2282
rect 15190 2258 15270 2274
rect 15286 2267 15348 2298
rect 15364 2267 15426 2298
rect 15495 2296 15544 2321
rect 15559 2296 15589 2312
rect 15458 2282 15488 2290
rect 15495 2288 15605 2296
rect 15458 2274 15503 2282
rect 15190 2256 15209 2258
rect 15224 2256 15270 2258
rect 15190 2240 15270 2256
rect 15297 2254 15332 2267
rect 15373 2264 15410 2267
rect 15373 2262 15415 2264
rect 15302 2251 15332 2254
rect 15311 2247 15318 2251
rect 15318 2246 15319 2247
rect 15277 2240 15287 2246
rect 15036 2232 15071 2240
rect 15036 2206 15037 2232
rect 15044 2206 15071 2232
rect 14979 2188 15009 2202
rect 15036 2198 15071 2206
rect 15073 2232 15114 2240
rect 15073 2206 15088 2232
rect 15095 2206 15114 2232
rect 15178 2228 15209 2240
rect 15224 2228 15327 2240
rect 15339 2230 15365 2256
rect 15380 2251 15410 2262
rect 15442 2258 15504 2274
rect 15442 2256 15488 2258
rect 15442 2240 15504 2256
rect 15516 2240 15522 2288
rect 15525 2280 15605 2288
rect 15525 2278 15544 2280
rect 15559 2278 15593 2280
rect 15525 2262 15605 2278
rect 15525 2240 15544 2262
rect 15559 2246 15589 2262
rect 15617 2256 15623 2330
rect 15626 2256 15645 2400
rect 15660 2256 15666 2400
rect 15675 2330 15688 2400
rect 15740 2396 15762 2400
rect 15733 2374 15762 2388
rect 15815 2374 15831 2388
rect 15869 2384 15875 2386
rect 15882 2384 15990 2400
rect 15997 2384 16003 2386
rect 16011 2384 16026 2400
rect 16092 2394 16111 2397
rect 15733 2372 15831 2374
rect 15858 2372 16026 2384
rect 16041 2374 16057 2388
rect 16092 2375 16114 2394
rect 16124 2388 16140 2389
rect 16123 2386 16140 2388
rect 16124 2381 16140 2386
rect 16114 2374 16120 2375
rect 16123 2374 16152 2381
rect 16041 2373 16152 2374
rect 16041 2372 16158 2373
rect 15717 2364 15768 2372
rect 15815 2364 15849 2372
rect 15717 2352 15742 2364
rect 15749 2352 15768 2364
rect 15822 2362 15849 2364
rect 15858 2362 16079 2372
rect 16114 2369 16120 2372
rect 15822 2358 16079 2362
rect 15717 2344 15768 2352
rect 15815 2344 16079 2358
rect 16123 2364 16158 2372
rect 15669 2296 15688 2330
rect 15733 2336 15762 2344
rect 15733 2330 15750 2336
rect 15733 2328 15767 2330
rect 15815 2328 15831 2344
rect 15832 2334 16040 2344
rect 16041 2334 16057 2344
rect 16105 2340 16120 2355
rect 16123 2352 16124 2364
rect 16131 2352 16158 2364
rect 16123 2344 16158 2352
rect 16123 2343 16152 2344
rect 15843 2330 16057 2334
rect 15858 2328 16057 2330
rect 16092 2330 16105 2340
rect 16123 2330 16140 2343
rect 16092 2328 16140 2330
rect 15734 2324 15767 2328
rect 15730 2322 15767 2324
rect 15730 2321 15797 2322
rect 15730 2316 15761 2321
rect 15767 2316 15797 2321
rect 15730 2312 15797 2316
rect 15703 2309 15797 2312
rect 15703 2302 15752 2309
rect 15703 2296 15733 2302
rect 15752 2297 15757 2302
rect 15669 2280 15749 2296
rect 15761 2288 15797 2309
rect 15858 2304 16047 2328
rect 16092 2327 16139 2328
rect 16105 2322 16139 2327
rect 15873 2301 16047 2304
rect 15866 2298 16047 2301
rect 16075 2321 16139 2322
rect 15669 2278 15688 2280
rect 15703 2278 15737 2280
rect 15669 2262 15749 2278
rect 15669 2256 15688 2262
rect 15385 2230 15488 2240
rect 15339 2228 15488 2230
rect 15509 2228 15544 2240
rect 15178 2226 15340 2228
rect 15190 2206 15209 2226
rect 15224 2224 15254 2226
rect 15073 2198 15114 2206
rect 15196 2202 15209 2206
rect 15261 2210 15340 2226
rect 15372 2226 15544 2228
rect 15372 2210 15451 2226
rect 15458 2224 15488 2226
rect 15036 2188 15065 2198
rect 15079 2188 15108 2198
rect 15123 2188 15153 2202
rect 15196 2188 15239 2202
rect 15261 2198 15451 2210
rect 15516 2206 15522 2226
rect 15246 2188 15276 2198
rect 15277 2188 15435 2198
rect 15439 2188 15469 2198
rect 15473 2188 15503 2202
rect 15531 2188 15544 2226
rect 15616 2240 15645 2256
rect 15659 2240 15688 2256
rect 15703 2246 15733 2262
rect 15761 2240 15767 2288
rect 15770 2282 15789 2288
rect 15804 2282 15834 2290
rect 15770 2274 15834 2282
rect 15770 2258 15850 2274
rect 15866 2267 15928 2298
rect 15944 2267 16006 2298
rect 16075 2296 16124 2321
rect 16139 2296 16169 2312
rect 16038 2282 16068 2290
rect 16075 2288 16185 2296
rect 16038 2274 16083 2282
rect 15770 2256 15789 2258
rect 15804 2256 15850 2258
rect 15770 2240 15850 2256
rect 15877 2254 15912 2267
rect 15953 2264 15990 2267
rect 15953 2262 15995 2264
rect 15882 2251 15912 2254
rect 15891 2247 15898 2251
rect 15898 2246 15899 2247
rect 15857 2240 15867 2246
rect 15616 2232 15651 2240
rect 15616 2206 15617 2232
rect 15624 2206 15651 2232
rect 15559 2188 15589 2202
rect 15616 2198 15651 2206
rect 15653 2232 15694 2240
rect 15653 2206 15668 2232
rect 15675 2206 15694 2232
rect 15758 2228 15789 2240
rect 15804 2228 15907 2240
rect 15919 2230 15945 2256
rect 15960 2251 15990 2262
rect 16022 2258 16084 2274
rect 16022 2256 16068 2258
rect 16022 2240 16084 2256
rect 16096 2240 16102 2288
rect 16105 2280 16185 2288
rect 16105 2278 16124 2280
rect 16139 2278 16173 2280
rect 16105 2262 16185 2278
rect 16105 2240 16124 2262
rect 16139 2246 16169 2262
rect 16197 2256 16203 2330
rect 16206 2256 16225 2400
rect 16240 2256 16246 2400
rect 16255 2330 16268 2400
rect 16320 2396 16342 2400
rect 16313 2374 16342 2388
rect 16395 2374 16411 2388
rect 16449 2384 16455 2386
rect 16462 2384 16570 2400
rect 16577 2384 16583 2386
rect 16591 2384 16606 2400
rect 16672 2394 16691 2397
rect 16313 2372 16411 2374
rect 16438 2372 16606 2384
rect 16621 2374 16637 2388
rect 16672 2375 16694 2394
rect 16704 2388 16720 2389
rect 16703 2386 16720 2388
rect 16704 2381 16720 2386
rect 16694 2374 16700 2375
rect 16703 2374 16732 2381
rect 16621 2373 16732 2374
rect 16621 2372 16738 2373
rect 16297 2364 16348 2372
rect 16395 2364 16429 2372
rect 16297 2352 16322 2364
rect 16329 2352 16348 2364
rect 16402 2362 16429 2364
rect 16438 2362 16659 2372
rect 16694 2369 16700 2372
rect 16402 2358 16659 2362
rect 16297 2344 16348 2352
rect 16395 2344 16659 2358
rect 16703 2364 16738 2372
rect 16249 2296 16268 2330
rect 16313 2336 16342 2344
rect 16313 2330 16330 2336
rect 16313 2328 16347 2330
rect 16395 2328 16411 2344
rect 16412 2334 16620 2344
rect 16621 2334 16637 2344
rect 16685 2340 16700 2355
rect 16703 2352 16704 2364
rect 16711 2352 16738 2364
rect 16703 2344 16738 2352
rect 16703 2343 16732 2344
rect 16423 2330 16637 2334
rect 16438 2328 16637 2330
rect 16672 2330 16685 2340
rect 16703 2330 16720 2343
rect 16672 2328 16720 2330
rect 16314 2324 16347 2328
rect 16310 2322 16347 2324
rect 16310 2321 16377 2322
rect 16310 2316 16341 2321
rect 16347 2316 16377 2321
rect 16310 2312 16377 2316
rect 16283 2309 16377 2312
rect 16283 2302 16332 2309
rect 16283 2296 16313 2302
rect 16332 2297 16337 2302
rect 16249 2280 16329 2296
rect 16341 2288 16377 2309
rect 16438 2304 16627 2328
rect 16672 2327 16719 2328
rect 16685 2322 16719 2327
rect 16453 2301 16627 2304
rect 16446 2298 16627 2301
rect 16655 2321 16719 2322
rect 16249 2278 16268 2280
rect 16283 2278 16317 2280
rect 16249 2262 16329 2278
rect 16249 2256 16268 2262
rect 15965 2230 16068 2240
rect 15919 2228 16068 2230
rect 16089 2228 16124 2240
rect 15758 2226 15920 2228
rect 15770 2206 15789 2226
rect 15804 2224 15834 2226
rect 15653 2198 15694 2206
rect 15776 2202 15789 2206
rect 15841 2210 15920 2226
rect 15952 2226 16124 2228
rect 15952 2210 16031 2226
rect 16038 2224 16068 2226
rect 15616 2188 15645 2198
rect 15659 2188 15688 2198
rect 15703 2188 15733 2202
rect 15776 2188 15819 2202
rect 15841 2198 16031 2210
rect 16096 2206 16102 2226
rect 15826 2188 15856 2198
rect 15857 2188 16015 2198
rect 16019 2188 16049 2198
rect 16053 2188 16083 2202
rect 16111 2188 16124 2226
rect 16196 2240 16225 2256
rect 16239 2240 16268 2256
rect 16283 2246 16313 2262
rect 16341 2240 16347 2288
rect 16350 2282 16369 2288
rect 16384 2282 16414 2290
rect 16350 2274 16414 2282
rect 16350 2258 16430 2274
rect 16446 2267 16508 2298
rect 16524 2267 16586 2298
rect 16655 2296 16704 2321
rect 16719 2296 16749 2312
rect 16618 2282 16648 2290
rect 16655 2288 16765 2296
rect 16618 2274 16663 2282
rect 16350 2256 16369 2258
rect 16384 2256 16430 2258
rect 16350 2240 16430 2256
rect 16457 2254 16492 2267
rect 16533 2264 16570 2267
rect 16533 2262 16575 2264
rect 16462 2251 16492 2254
rect 16471 2247 16478 2251
rect 16478 2246 16479 2247
rect 16437 2240 16447 2246
rect 16196 2232 16231 2240
rect 16196 2206 16197 2232
rect 16204 2206 16231 2232
rect 16139 2188 16169 2202
rect 16196 2198 16231 2206
rect 16233 2232 16274 2240
rect 16233 2206 16248 2232
rect 16255 2206 16274 2232
rect 16338 2228 16369 2240
rect 16384 2228 16487 2240
rect 16499 2230 16525 2256
rect 16540 2251 16570 2262
rect 16602 2258 16664 2274
rect 16602 2256 16648 2258
rect 16602 2240 16664 2256
rect 16676 2240 16682 2288
rect 16685 2280 16765 2288
rect 16685 2278 16704 2280
rect 16719 2278 16753 2280
rect 16685 2262 16765 2278
rect 16685 2240 16704 2262
rect 16719 2246 16749 2262
rect 16777 2256 16783 2330
rect 16786 2256 16805 2400
rect 16820 2256 16826 2400
rect 16835 2330 16848 2400
rect 16900 2396 16922 2400
rect 16893 2374 16922 2388
rect 16975 2374 16991 2388
rect 17029 2384 17035 2386
rect 17042 2384 17150 2400
rect 17157 2384 17163 2386
rect 17171 2384 17186 2400
rect 17252 2394 17271 2397
rect 16893 2372 16991 2374
rect 17018 2372 17186 2384
rect 17201 2374 17217 2388
rect 17252 2375 17274 2394
rect 17284 2388 17300 2389
rect 17283 2386 17300 2388
rect 17284 2381 17300 2386
rect 17274 2374 17280 2375
rect 17283 2374 17312 2381
rect 17201 2373 17312 2374
rect 17201 2372 17318 2373
rect 16877 2364 16928 2372
rect 16975 2364 17009 2372
rect 16877 2352 16902 2364
rect 16909 2352 16928 2364
rect 16982 2362 17009 2364
rect 17018 2362 17239 2372
rect 17274 2369 17280 2372
rect 16982 2358 17239 2362
rect 16877 2344 16928 2352
rect 16975 2344 17239 2358
rect 17283 2364 17318 2372
rect 16829 2296 16848 2330
rect 16893 2336 16922 2344
rect 16893 2330 16910 2336
rect 16893 2328 16927 2330
rect 16975 2328 16991 2344
rect 16992 2334 17200 2344
rect 17201 2334 17217 2344
rect 17265 2340 17280 2355
rect 17283 2352 17284 2364
rect 17291 2352 17318 2364
rect 17283 2344 17318 2352
rect 17283 2343 17312 2344
rect 17003 2330 17217 2334
rect 17018 2328 17217 2330
rect 17252 2330 17265 2340
rect 17283 2330 17300 2343
rect 17252 2328 17300 2330
rect 16894 2324 16927 2328
rect 16890 2322 16927 2324
rect 16890 2321 16957 2322
rect 16890 2316 16921 2321
rect 16927 2316 16957 2321
rect 16890 2312 16957 2316
rect 16863 2309 16957 2312
rect 16863 2302 16912 2309
rect 16863 2296 16893 2302
rect 16912 2297 16917 2302
rect 16829 2280 16909 2296
rect 16921 2288 16957 2309
rect 17018 2304 17207 2328
rect 17252 2327 17299 2328
rect 17265 2322 17299 2327
rect 17033 2301 17207 2304
rect 17026 2298 17207 2301
rect 17235 2321 17299 2322
rect 16829 2278 16848 2280
rect 16863 2278 16897 2280
rect 16829 2262 16909 2278
rect 16829 2256 16848 2262
rect 16545 2230 16648 2240
rect 16499 2228 16648 2230
rect 16669 2228 16704 2240
rect 16338 2226 16500 2228
rect 16350 2206 16369 2226
rect 16384 2224 16414 2226
rect 16233 2198 16274 2206
rect 16356 2202 16369 2206
rect 16421 2210 16500 2226
rect 16532 2226 16704 2228
rect 16532 2210 16611 2226
rect 16618 2224 16648 2226
rect 16196 2188 16225 2198
rect 16239 2188 16268 2198
rect 16283 2188 16313 2202
rect 16356 2188 16399 2202
rect 16421 2198 16611 2210
rect 16676 2206 16682 2226
rect 16406 2188 16436 2198
rect 16437 2188 16595 2198
rect 16599 2188 16629 2198
rect 16633 2188 16663 2202
rect 16691 2188 16704 2226
rect 16776 2240 16805 2256
rect 16819 2240 16848 2256
rect 16863 2246 16893 2262
rect 16921 2240 16927 2288
rect 16930 2282 16949 2288
rect 16964 2282 16994 2290
rect 16930 2274 16994 2282
rect 16930 2258 17010 2274
rect 17026 2267 17088 2298
rect 17104 2267 17166 2298
rect 17235 2296 17284 2321
rect 17299 2296 17329 2312
rect 17198 2282 17228 2290
rect 17235 2288 17345 2296
rect 17198 2274 17243 2282
rect 16930 2256 16949 2258
rect 16964 2256 17010 2258
rect 16930 2240 17010 2256
rect 17037 2254 17072 2267
rect 17113 2264 17150 2267
rect 17113 2262 17155 2264
rect 17042 2251 17072 2254
rect 17051 2247 17058 2251
rect 17058 2246 17059 2247
rect 17017 2240 17027 2246
rect 16776 2232 16811 2240
rect 16776 2206 16777 2232
rect 16784 2206 16811 2232
rect 16719 2188 16749 2202
rect 16776 2198 16811 2206
rect 16813 2232 16854 2240
rect 16813 2206 16828 2232
rect 16835 2206 16854 2232
rect 16918 2228 16949 2240
rect 16964 2228 17067 2240
rect 17079 2230 17105 2256
rect 17120 2251 17150 2262
rect 17182 2258 17244 2274
rect 17182 2256 17228 2258
rect 17182 2240 17244 2256
rect 17256 2240 17262 2288
rect 17265 2280 17345 2288
rect 17265 2278 17284 2280
rect 17299 2278 17333 2280
rect 17265 2262 17345 2278
rect 17265 2240 17284 2262
rect 17299 2246 17329 2262
rect 17357 2256 17363 2330
rect 17366 2256 17385 2400
rect 17400 2256 17406 2400
rect 17415 2330 17428 2400
rect 17480 2396 17502 2400
rect 17473 2374 17502 2388
rect 17555 2374 17571 2388
rect 17609 2384 17615 2386
rect 17622 2384 17730 2400
rect 17737 2384 17743 2386
rect 17751 2384 17766 2400
rect 17832 2394 17851 2397
rect 17473 2372 17571 2374
rect 17598 2372 17766 2384
rect 17781 2374 17797 2388
rect 17832 2375 17854 2394
rect 17864 2388 17880 2389
rect 17863 2386 17880 2388
rect 17864 2381 17880 2386
rect 17854 2374 17860 2375
rect 17863 2374 17892 2381
rect 17781 2373 17892 2374
rect 17781 2372 17898 2373
rect 17457 2364 17508 2372
rect 17555 2364 17589 2372
rect 17457 2352 17482 2364
rect 17489 2352 17508 2364
rect 17562 2362 17589 2364
rect 17598 2362 17819 2372
rect 17854 2369 17860 2372
rect 17562 2358 17819 2362
rect 17457 2344 17508 2352
rect 17555 2344 17819 2358
rect 17863 2364 17898 2372
rect 17409 2296 17428 2330
rect 17473 2336 17502 2344
rect 17473 2330 17490 2336
rect 17473 2328 17507 2330
rect 17555 2328 17571 2344
rect 17572 2334 17780 2344
rect 17781 2334 17797 2344
rect 17845 2340 17860 2355
rect 17863 2352 17864 2364
rect 17871 2352 17898 2364
rect 17863 2344 17898 2352
rect 17863 2343 17892 2344
rect 17583 2330 17797 2334
rect 17598 2328 17797 2330
rect 17832 2330 17845 2340
rect 17863 2330 17880 2343
rect 17832 2328 17880 2330
rect 17474 2324 17507 2328
rect 17470 2322 17507 2324
rect 17470 2321 17537 2322
rect 17470 2316 17501 2321
rect 17507 2316 17537 2321
rect 17470 2312 17537 2316
rect 17443 2309 17537 2312
rect 17443 2302 17492 2309
rect 17443 2296 17473 2302
rect 17492 2297 17497 2302
rect 17409 2280 17489 2296
rect 17501 2288 17537 2309
rect 17598 2304 17787 2328
rect 17832 2327 17879 2328
rect 17845 2322 17879 2327
rect 17613 2301 17787 2304
rect 17606 2298 17787 2301
rect 17815 2321 17879 2322
rect 17409 2278 17428 2280
rect 17443 2278 17477 2280
rect 17409 2262 17489 2278
rect 17409 2256 17428 2262
rect 17125 2230 17228 2240
rect 17079 2228 17228 2230
rect 17249 2228 17284 2240
rect 16918 2226 17080 2228
rect 16930 2206 16949 2226
rect 16964 2224 16994 2226
rect 16813 2198 16854 2206
rect 16936 2202 16949 2206
rect 17001 2210 17080 2226
rect 17112 2226 17284 2228
rect 17112 2210 17191 2226
rect 17198 2224 17228 2226
rect 16776 2188 16805 2198
rect 16819 2188 16848 2198
rect 16863 2188 16893 2202
rect 16936 2188 16979 2202
rect 17001 2198 17191 2210
rect 17256 2206 17262 2226
rect 16986 2188 17016 2198
rect 17017 2188 17175 2198
rect 17179 2188 17209 2198
rect 17213 2188 17243 2202
rect 17271 2188 17284 2226
rect 17356 2240 17385 2256
rect 17399 2240 17428 2256
rect 17443 2246 17473 2262
rect 17501 2240 17507 2288
rect 17510 2282 17529 2288
rect 17544 2282 17574 2290
rect 17510 2274 17574 2282
rect 17510 2258 17590 2274
rect 17606 2267 17668 2298
rect 17684 2267 17746 2298
rect 17815 2296 17864 2321
rect 17879 2296 17909 2312
rect 17778 2282 17808 2290
rect 17815 2288 17925 2296
rect 17778 2274 17823 2282
rect 17510 2256 17529 2258
rect 17544 2256 17590 2258
rect 17510 2240 17590 2256
rect 17617 2254 17652 2267
rect 17693 2264 17730 2267
rect 17693 2262 17735 2264
rect 17622 2251 17652 2254
rect 17631 2247 17638 2251
rect 17638 2246 17639 2247
rect 17597 2240 17607 2246
rect 17356 2232 17391 2240
rect 17356 2206 17357 2232
rect 17364 2206 17391 2232
rect 17299 2188 17329 2202
rect 17356 2198 17391 2206
rect 17393 2232 17434 2240
rect 17393 2206 17408 2232
rect 17415 2206 17434 2232
rect 17498 2228 17529 2240
rect 17544 2228 17647 2240
rect 17659 2230 17685 2256
rect 17700 2251 17730 2262
rect 17762 2258 17824 2274
rect 17762 2256 17808 2258
rect 17762 2240 17824 2256
rect 17836 2240 17842 2288
rect 17845 2280 17925 2288
rect 17845 2278 17864 2280
rect 17879 2278 17913 2280
rect 17845 2262 17925 2278
rect 17845 2240 17864 2262
rect 17879 2246 17909 2262
rect 17937 2256 17943 2330
rect 17946 2256 17965 2400
rect 17980 2256 17986 2400
rect 17995 2330 18008 2400
rect 18060 2396 18082 2400
rect 18053 2374 18082 2388
rect 18135 2374 18151 2388
rect 18189 2384 18195 2386
rect 18202 2384 18310 2400
rect 18317 2384 18323 2386
rect 18331 2384 18346 2400
rect 18412 2394 18431 2397
rect 18053 2372 18151 2374
rect 18178 2372 18346 2384
rect 18361 2374 18377 2388
rect 18412 2375 18434 2394
rect 18444 2388 18460 2389
rect 18443 2386 18460 2388
rect 18444 2381 18460 2386
rect 18434 2374 18440 2375
rect 18443 2374 18472 2381
rect 18361 2373 18472 2374
rect 18361 2372 18478 2373
rect 18037 2364 18088 2372
rect 18135 2364 18169 2372
rect 18037 2352 18062 2364
rect 18069 2352 18088 2364
rect 18142 2362 18169 2364
rect 18178 2362 18399 2372
rect 18434 2369 18440 2372
rect 18142 2358 18399 2362
rect 18037 2344 18088 2352
rect 18135 2344 18399 2358
rect 18443 2364 18478 2372
rect 17989 2296 18008 2330
rect 18053 2336 18082 2344
rect 18053 2330 18070 2336
rect 18053 2328 18087 2330
rect 18135 2328 18151 2344
rect 18152 2334 18360 2344
rect 18361 2334 18377 2344
rect 18425 2340 18440 2355
rect 18443 2352 18444 2364
rect 18451 2352 18478 2364
rect 18443 2344 18478 2352
rect 18443 2343 18472 2344
rect 18163 2330 18377 2334
rect 18178 2328 18377 2330
rect 18412 2330 18425 2340
rect 18443 2330 18460 2343
rect 18412 2328 18460 2330
rect 18054 2324 18087 2328
rect 18050 2322 18087 2324
rect 18050 2321 18117 2322
rect 18050 2316 18081 2321
rect 18087 2316 18117 2321
rect 18050 2312 18117 2316
rect 18023 2309 18117 2312
rect 18023 2302 18072 2309
rect 18023 2296 18053 2302
rect 18072 2297 18077 2302
rect 17989 2280 18069 2296
rect 18081 2288 18117 2309
rect 18178 2304 18367 2328
rect 18412 2327 18459 2328
rect 18425 2322 18459 2327
rect 18193 2301 18367 2304
rect 18186 2298 18367 2301
rect 18395 2321 18459 2322
rect 17989 2278 18008 2280
rect 18023 2278 18057 2280
rect 17989 2262 18069 2278
rect 17989 2256 18008 2262
rect 17705 2230 17808 2240
rect 17659 2228 17808 2230
rect 17829 2228 17864 2240
rect 17498 2226 17660 2228
rect 17510 2206 17529 2226
rect 17544 2224 17574 2226
rect 17393 2198 17434 2206
rect 17516 2202 17529 2206
rect 17581 2210 17660 2226
rect 17692 2226 17864 2228
rect 17692 2210 17771 2226
rect 17778 2224 17808 2226
rect 17356 2188 17385 2198
rect 17399 2188 17428 2198
rect 17443 2188 17473 2202
rect 17516 2188 17559 2202
rect 17581 2198 17771 2210
rect 17836 2206 17842 2226
rect 17566 2188 17596 2198
rect 17597 2188 17755 2198
rect 17759 2188 17789 2198
rect 17793 2188 17823 2202
rect 17851 2188 17864 2226
rect 17936 2240 17965 2256
rect 17979 2240 18008 2256
rect 18023 2246 18053 2262
rect 18081 2240 18087 2288
rect 18090 2282 18109 2288
rect 18124 2282 18154 2290
rect 18090 2274 18154 2282
rect 18090 2258 18170 2274
rect 18186 2267 18248 2298
rect 18264 2267 18326 2298
rect 18395 2296 18444 2321
rect 18459 2296 18489 2312
rect 18358 2282 18388 2290
rect 18395 2288 18505 2296
rect 18358 2274 18403 2282
rect 18090 2256 18109 2258
rect 18124 2256 18170 2258
rect 18090 2240 18170 2256
rect 18197 2254 18232 2267
rect 18273 2264 18310 2267
rect 18273 2262 18315 2264
rect 18202 2251 18232 2254
rect 18211 2247 18218 2251
rect 18218 2246 18219 2247
rect 18177 2240 18187 2246
rect 17936 2232 17971 2240
rect 17936 2206 17937 2232
rect 17944 2206 17971 2232
rect 17879 2188 17909 2202
rect 17936 2198 17971 2206
rect 17973 2232 18014 2240
rect 17973 2206 17988 2232
rect 17995 2206 18014 2232
rect 18078 2228 18109 2240
rect 18124 2228 18227 2240
rect 18239 2230 18265 2256
rect 18280 2251 18310 2262
rect 18342 2258 18404 2274
rect 18342 2256 18388 2258
rect 18342 2240 18404 2256
rect 18416 2240 18422 2288
rect 18425 2280 18505 2288
rect 18425 2278 18444 2280
rect 18459 2278 18493 2280
rect 18425 2262 18505 2278
rect 18425 2240 18444 2262
rect 18459 2246 18489 2262
rect 18517 2256 18523 2330
rect 18532 2256 18545 2400
rect 18285 2230 18388 2240
rect 18239 2228 18388 2230
rect 18409 2228 18444 2240
rect 18078 2226 18240 2228
rect 18090 2206 18109 2226
rect 18124 2224 18154 2226
rect 17973 2198 18014 2206
rect 18096 2202 18109 2206
rect 18161 2210 18240 2226
rect 18272 2226 18444 2228
rect 18272 2210 18351 2226
rect 18358 2224 18388 2226
rect 17936 2188 17965 2198
rect 17979 2188 18008 2198
rect 18023 2188 18053 2202
rect 18096 2188 18139 2202
rect 18161 2198 18351 2210
rect 18416 2206 18422 2226
rect 18146 2188 18176 2198
rect 18177 2188 18335 2198
rect 18339 2188 18369 2198
rect 18373 2188 18403 2202
rect 18431 2188 18444 2226
rect 18516 2240 18545 2256
rect 18516 2232 18551 2240
rect 18516 2206 18517 2232
rect 18524 2206 18551 2232
rect 18459 2188 18489 2202
rect 18516 2198 18551 2206
rect 18516 2188 18545 2198
rect -1 2182 18545 2188
rect 0 2174 18545 2182
rect 15 2144 28 2174
rect 43 2160 73 2174
rect 116 2160 159 2174
rect 166 2160 386 2174
rect 393 2160 423 2174
rect 83 2146 98 2158
rect 117 2146 130 2160
rect 198 2156 351 2160
rect 80 2144 102 2146
rect 180 2144 372 2156
rect 451 2144 464 2174
rect 479 2160 509 2174
rect 546 2144 565 2174
rect 580 2144 586 2174
rect 595 2144 608 2174
rect 623 2160 653 2174
rect 696 2160 739 2174
rect 746 2160 966 2174
rect 973 2160 1003 2174
rect 663 2146 678 2158
rect 697 2146 710 2160
rect 778 2156 931 2160
rect 660 2144 682 2146
rect 760 2144 952 2156
rect 1031 2144 1044 2174
rect 1059 2160 1089 2174
rect 1126 2144 1145 2174
rect 1160 2144 1166 2174
rect 1175 2144 1188 2174
rect 1203 2160 1233 2174
rect 1276 2160 1319 2174
rect 1326 2160 1546 2174
rect 1553 2160 1583 2174
rect 1243 2146 1258 2158
rect 1277 2146 1290 2160
rect 1358 2156 1511 2160
rect 1240 2144 1262 2146
rect 1340 2144 1532 2156
rect 1611 2144 1624 2174
rect 1639 2160 1669 2174
rect 1706 2144 1725 2174
rect 1740 2144 1746 2174
rect 1755 2144 1768 2174
rect 1783 2160 1813 2174
rect 1856 2160 1899 2174
rect 1906 2160 2126 2174
rect 2133 2160 2163 2174
rect 1823 2146 1838 2158
rect 1857 2146 1870 2160
rect 1938 2156 2091 2160
rect 1820 2144 1842 2146
rect 1920 2144 2112 2156
rect 2191 2144 2204 2174
rect 2219 2160 2249 2174
rect 2286 2144 2305 2174
rect 2320 2144 2326 2174
rect 2335 2144 2348 2174
rect 2363 2160 2393 2174
rect 2436 2160 2479 2174
rect 2486 2160 2706 2174
rect 2713 2160 2743 2174
rect 2403 2146 2418 2158
rect 2437 2146 2450 2160
rect 2518 2156 2671 2160
rect 2400 2144 2422 2146
rect 2500 2144 2692 2156
rect 2771 2144 2784 2174
rect 2799 2160 2829 2174
rect 2866 2144 2885 2174
rect 2900 2144 2906 2174
rect 2915 2144 2928 2174
rect 2943 2160 2973 2174
rect 3016 2160 3059 2174
rect 3066 2160 3286 2174
rect 3293 2160 3323 2174
rect 2983 2146 2998 2158
rect 3017 2146 3030 2160
rect 3098 2156 3251 2160
rect 2980 2144 3002 2146
rect 3080 2144 3272 2156
rect 3351 2144 3364 2174
rect 3379 2160 3409 2174
rect 3446 2144 3465 2174
rect 3480 2144 3486 2174
rect 3495 2144 3508 2174
rect 3523 2160 3553 2174
rect 3596 2160 3639 2174
rect 3646 2160 3866 2174
rect 3873 2160 3903 2174
rect 3563 2146 3578 2158
rect 3597 2146 3610 2160
rect 3678 2156 3831 2160
rect 3560 2144 3582 2146
rect 3660 2144 3852 2156
rect 3931 2144 3944 2174
rect 3959 2160 3989 2174
rect 4026 2144 4045 2174
rect 4060 2144 4066 2174
rect 4075 2144 4088 2174
rect 4103 2160 4133 2174
rect 4176 2160 4219 2174
rect 4226 2160 4446 2174
rect 4453 2160 4483 2174
rect 4143 2146 4158 2158
rect 4177 2146 4190 2160
rect 4258 2156 4411 2160
rect 4140 2144 4162 2146
rect 4240 2144 4432 2156
rect 4511 2144 4524 2174
rect 4539 2160 4569 2174
rect 4606 2144 4625 2174
rect 4640 2144 4646 2174
rect 4655 2144 4668 2174
rect 4683 2160 4713 2174
rect 4756 2160 4799 2174
rect 4806 2160 5026 2174
rect 5033 2160 5063 2174
rect 4723 2146 4738 2158
rect 4757 2146 4770 2160
rect 4838 2156 4991 2160
rect 4720 2144 4742 2146
rect 4820 2144 5012 2156
rect 5091 2144 5104 2174
rect 5119 2160 5149 2174
rect 5186 2144 5205 2174
rect 5220 2144 5226 2174
rect 5235 2144 5248 2174
rect 5263 2160 5293 2174
rect 5336 2160 5379 2174
rect 5386 2160 5606 2174
rect 5613 2160 5643 2174
rect 5303 2146 5318 2158
rect 5337 2146 5350 2160
rect 5418 2156 5571 2160
rect 5300 2144 5322 2146
rect 5400 2144 5592 2156
rect 5671 2144 5684 2174
rect 5699 2160 5729 2174
rect 5766 2144 5785 2174
rect 5800 2144 5806 2174
rect 5815 2144 5828 2174
rect 5843 2160 5873 2174
rect 5916 2160 5959 2174
rect 5966 2160 6186 2174
rect 6193 2160 6223 2174
rect 5883 2146 5898 2158
rect 5917 2146 5930 2160
rect 5998 2156 6151 2160
rect 5880 2144 5902 2146
rect 5980 2144 6172 2156
rect 6251 2144 6264 2174
rect 6279 2160 6309 2174
rect 6346 2144 6365 2174
rect 6380 2144 6386 2174
rect 6395 2144 6408 2174
rect 6423 2160 6453 2174
rect 6496 2160 6539 2174
rect 6546 2160 6766 2174
rect 6773 2160 6803 2174
rect 6463 2146 6478 2158
rect 6497 2146 6510 2160
rect 6578 2156 6731 2160
rect 6460 2144 6482 2146
rect 6560 2144 6752 2156
rect 6831 2144 6844 2174
rect 6859 2160 6889 2174
rect 6926 2144 6945 2174
rect 6960 2144 6966 2174
rect 6975 2144 6988 2174
rect 7003 2160 7033 2174
rect 7076 2160 7119 2174
rect 7126 2160 7346 2174
rect 7353 2160 7383 2174
rect 7043 2146 7058 2158
rect 7077 2146 7090 2160
rect 7158 2156 7311 2160
rect 7040 2144 7062 2146
rect 7140 2144 7332 2156
rect 7411 2144 7424 2174
rect 7439 2160 7469 2174
rect 7506 2144 7525 2174
rect 7540 2144 7546 2174
rect 7555 2144 7568 2174
rect 7583 2160 7613 2174
rect 7656 2160 7699 2174
rect 7706 2160 7926 2174
rect 7933 2160 7963 2174
rect 7623 2146 7638 2158
rect 7657 2146 7670 2160
rect 7738 2156 7891 2160
rect 7620 2144 7642 2146
rect 7720 2144 7912 2156
rect 7991 2144 8004 2174
rect 8019 2160 8049 2174
rect 8086 2144 8105 2174
rect 8120 2144 8126 2174
rect 8135 2144 8148 2174
rect 8163 2160 8193 2174
rect 8236 2160 8279 2174
rect 8286 2160 8506 2174
rect 8513 2160 8543 2174
rect 8203 2146 8218 2158
rect 8237 2146 8250 2160
rect 8318 2156 8471 2160
rect 8200 2144 8222 2146
rect 8300 2144 8492 2156
rect 8571 2144 8584 2174
rect 8599 2160 8629 2174
rect 8666 2144 8685 2174
rect 8700 2144 8706 2174
rect 8715 2144 8728 2174
rect 8743 2160 8773 2174
rect 8816 2160 8859 2174
rect 8866 2160 9086 2174
rect 9093 2160 9123 2174
rect 8783 2146 8798 2158
rect 8817 2146 8830 2160
rect 8898 2156 9051 2160
rect 8780 2144 8802 2146
rect 8880 2144 9072 2156
rect 9151 2144 9164 2174
rect 9179 2160 9209 2174
rect 9246 2144 9265 2174
rect 9280 2144 9286 2174
rect 9295 2144 9308 2174
rect 9323 2160 9353 2174
rect 9396 2160 9439 2174
rect 9446 2160 9666 2174
rect 9673 2160 9703 2174
rect 9363 2146 9378 2158
rect 9397 2146 9410 2160
rect 9478 2156 9631 2160
rect 9360 2144 9382 2146
rect 9460 2144 9652 2156
rect 9731 2144 9744 2174
rect 9759 2160 9789 2174
rect 9826 2144 9845 2174
rect 9860 2144 9866 2174
rect 9875 2144 9888 2174
rect 9903 2160 9933 2174
rect 9976 2160 10019 2174
rect 10026 2160 10246 2174
rect 10253 2160 10283 2174
rect 9943 2146 9958 2158
rect 9977 2146 9990 2160
rect 10058 2156 10211 2160
rect 9940 2144 9962 2146
rect 10040 2144 10232 2156
rect 10311 2144 10324 2174
rect 10339 2160 10369 2174
rect 10406 2144 10425 2174
rect 10440 2144 10446 2174
rect 10455 2144 10468 2174
rect 10483 2160 10513 2174
rect 10556 2160 10599 2174
rect 10606 2160 10826 2174
rect 10833 2160 10863 2174
rect 10523 2146 10538 2158
rect 10557 2146 10570 2160
rect 10638 2156 10791 2160
rect 10520 2144 10542 2146
rect 10620 2144 10812 2156
rect 10891 2144 10904 2174
rect 10919 2160 10949 2174
rect 10986 2144 11005 2174
rect 11020 2144 11026 2174
rect 11035 2144 11048 2174
rect 11063 2160 11093 2174
rect 11136 2160 11179 2174
rect 11186 2160 11406 2174
rect 11413 2160 11443 2174
rect 11103 2146 11118 2158
rect 11137 2146 11150 2160
rect 11218 2156 11371 2160
rect 11100 2144 11122 2146
rect 11200 2144 11392 2156
rect 11471 2144 11484 2174
rect 11499 2160 11529 2174
rect 11566 2144 11585 2174
rect 11600 2144 11606 2174
rect 11615 2144 11628 2174
rect 11643 2160 11673 2174
rect 11716 2160 11759 2174
rect 11766 2160 11986 2174
rect 11993 2160 12023 2174
rect 11683 2146 11698 2158
rect 11717 2146 11730 2160
rect 11798 2156 11951 2160
rect 11680 2144 11702 2146
rect 11780 2144 11972 2156
rect 12051 2144 12064 2174
rect 12079 2160 12109 2174
rect 12146 2144 12165 2174
rect 12180 2144 12186 2174
rect 12195 2144 12208 2174
rect 12223 2160 12253 2174
rect 12296 2160 12339 2174
rect 12346 2160 12566 2174
rect 12573 2160 12603 2174
rect 12263 2146 12278 2158
rect 12297 2146 12310 2160
rect 12378 2156 12531 2160
rect 12260 2144 12282 2146
rect 12360 2144 12552 2156
rect 12631 2144 12644 2174
rect 12659 2160 12689 2174
rect 12726 2144 12745 2174
rect 12760 2144 12766 2174
rect 12775 2144 12788 2174
rect 12803 2160 12833 2174
rect 12876 2160 12919 2174
rect 12926 2160 13146 2174
rect 13153 2160 13183 2174
rect 12843 2146 12858 2158
rect 12877 2146 12890 2160
rect 12958 2156 13111 2160
rect 12840 2144 12862 2146
rect 12940 2144 13132 2156
rect 13211 2144 13224 2174
rect 13239 2160 13269 2174
rect 13306 2144 13325 2174
rect 13340 2144 13346 2174
rect 13355 2144 13368 2174
rect 13383 2160 13413 2174
rect 13456 2160 13499 2174
rect 13506 2160 13726 2174
rect 13733 2160 13763 2174
rect 13423 2146 13438 2158
rect 13457 2146 13470 2160
rect 13538 2156 13691 2160
rect 13420 2144 13442 2146
rect 13520 2144 13712 2156
rect 13791 2144 13804 2174
rect 13819 2160 13849 2174
rect 13886 2144 13905 2174
rect 13920 2144 13926 2174
rect 13935 2144 13948 2174
rect 13963 2160 13993 2174
rect 14036 2160 14079 2174
rect 14086 2160 14306 2174
rect 14313 2160 14343 2174
rect 14003 2146 14018 2158
rect 14037 2146 14050 2160
rect 14118 2156 14271 2160
rect 14000 2144 14022 2146
rect 14100 2144 14292 2156
rect 14371 2144 14384 2174
rect 14399 2160 14429 2174
rect 14466 2144 14485 2174
rect 14500 2144 14506 2174
rect 14515 2144 14528 2174
rect 14543 2160 14573 2174
rect 14616 2160 14659 2174
rect 14666 2160 14886 2174
rect 14893 2160 14923 2174
rect 14583 2146 14598 2158
rect 14617 2146 14630 2160
rect 14698 2156 14851 2160
rect 14580 2144 14602 2146
rect 14680 2144 14872 2156
rect 14951 2144 14964 2174
rect 14979 2160 15009 2174
rect 15046 2144 15065 2174
rect 15080 2144 15086 2174
rect 15095 2144 15108 2174
rect 15123 2160 15153 2174
rect 15196 2160 15239 2174
rect 15246 2160 15466 2174
rect 15473 2160 15503 2174
rect 15163 2146 15178 2158
rect 15197 2146 15210 2160
rect 15278 2156 15431 2160
rect 15160 2144 15182 2146
rect 15260 2144 15452 2156
rect 15531 2144 15544 2174
rect 15559 2160 15589 2174
rect 15626 2144 15645 2174
rect 15660 2144 15666 2174
rect 15675 2144 15688 2174
rect 15703 2160 15733 2174
rect 15776 2160 15819 2174
rect 15826 2160 16046 2174
rect 16053 2160 16083 2174
rect 15743 2146 15758 2158
rect 15777 2146 15790 2160
rect 15858 2156 16011 2160
rect 15740 2144 15762 2146
rect 15840 2144 16032 2156
rect 16111 2144 16124 2174
rect 16139 2160 16169 2174
rect 16206 2144 16225 2174
rect 16240 2144 16246 2174
rect 16255 2144 16268 2174
rect 16283 2160 16313 2174
rect 16356 2160 16399 2174
rect 16406 2160 16626 2174
rect 16633 2160 16663 2174
rect 16323 2146 16338 2158
rect 16357 2146 16370 2160
rect 16438 2156 16591 2160
rect 16320 2144 16342 2146
rect 16420 2144 16612 2156
rect 16691 2144 16704 2174
rect 16719 2160 16749 2174
rect 16786 2144 16805 2174
rect 16820 2144 16826 2174
rect 16835 2144 16848 2174
rect 16863 2160 16893 2174
rect 16936 2160 16979 2174
rect 16986 2160 17206 2174
rect 17213 2160 17243 2174
rect 16903 2146 16918 2158
rect 16937 2146 16950 2160
rect 17018 2156 17171 2160
rect 16900 2144 16922 2146
rect 17000 2144 17192 2156
rect 17271 2144 17284 2174
rect 17299 2160 17329 2174
rect 17366 2144 17385 2174
rect 17400 2144 17406 2174
rect 17415 2144 17428 2174
rect 17443 2160 17473 2174
rect 17516 2160 17559 2174
rect 17566 2160 17786 2174
rect 17793 2160 17823 2174
rect 17483 2146 17498 2158
rect 17517 2146 17530 2160
rect 17598 2156 17751 2160
rect 17480 2144 17502 2146
rect 17580 2144 17772 2156
rect 17851 2144 17864 2174
rect 17879 2160 17909 2174
rect 17946 2144 17965 2174
rect 17980 2144 17986 2174
rect 17995 2144 18008 2174
rect 18023 2160 18053 2174
rect 18096 2160 18139 2174
rect 18146 2160 18366 2174
rect 18373 2160 18403 2174
rect 18063 2146 18078 2158
rect 18097 2146 18110 2160
rect 18178 2156 18331 2160
rect 18060 2144 18082 2146
rect 18160 2144 18352 2156
rect 18431 2144 18444 2174
rect 18459 2160 18489 2174
rect 18532 2144 18545 2174
rect 0 2130 18545 2144
rect 15 2060 28 2130
rect 80 2126 102 2130
rect 73 2104 102 2118
rect 155 2104 171 2118
rect 209 2114 215 2116
rect 222 2114 330 2130
rect 337 2114 343 2116
rect 351 2114 366 2130
rect 432 2124 451 2127
rect 73 2102 171 2104
rect 198 2102 366 2114
rect 381 2104 397 2118
rect 432 2105 454 2124
rect 464 2118 480 2119
rect 463 2116 480 2118
rect 464 2111 480 2116
rect 454 2104 460 2105
rect 463 2104 492 2111
rect 381 2103 492 2104
rect 381 2102 498 2103
rect 57 2094 108 2102
rect 155 2094 189 2102
rect 57 2082 82 2094
rect 89 2082 108 2094
rect 162 2092 189 2094
rect 198 2092 419 2102
rect 454 2099 460 2102
rect 162 2088 419 2092
rect 57 2074 108 2082
rect 155 2074 419 2088
rect 463 2094 498 2102
rect 9 2026 28 2060
rect 73 2066 102 2074
rect 73 2060 90 2066
rect 73 2058 107 2060
rect 155 2058 171 2074
rect 172 2064 380 2074
rect 381 2064 397 2074
rect 445 2070 460 2085
rect 463 2082 464 2094
rect 471 2082 498 2094
rect 463 2074 498 2082
rect 463 2073 492 2074
rect 183 2060 397 2064
rect 198 2058 397 2060
rect 432 2060 445 2070
rect 463 2060 480 2073
rect 432 2058 480 2060
rect 74 2054 107 2058
rect 70 2052 107 2054
rect 70 2051 137 2052
rect 70 2046 101 2051
rect 107 2046 137 2051
rect 70 2042 137 2046
rect 43 2039 137 2042
rect 43 2032 92 2039
rect 43 2026 73 2032
rect 92 2027 97 2032
rect 9 2010 89 2026
rect 101 2018 137 2039
rect 198 2034 387 2058
rect 432 2057 479 2058
rect 445 2052 479 2057
rect 213 2031 387 2034
rect 206 2028 387 2031
rect 415 2051 479 2052
rect 9 2008 28 2010
rect 43 2008 77 2010
rect 9 1992 89 2008
rect 9 1986 28 1992
rect -1 1970 28 1986
rect 43 1976 73 1992
rect 101 1970 107 2018
rect 110 2012 129 2018
rect 144 2012 174 2020
rect 110 2004 174 2012
rect 110 1988 190 2004
rect 206 1997 268 2028
rect 284 1997 346 2028
rect 415 2026 464 2051
rect 479 2026 509 2042
rect 378 2012 408 2020
rect 415 2018 525 2026
rect 378 2004 423 2012
rect 110 1986 129 1988
rect 144 1986 190 1988
rect 110 1970 190 1986
rect 217 1984 252 1997
rect 293 1994 330 1997
rect 293 1992 335 1994
rect 222 1981 252 1984
rect 231 1977 238 1981
rect 238 1976 239 1977
rect 197 1970 207 1976
rect -7 1962 34 1970
rect -7 1936 8 1962
rect 15 1936 34 1962
rect 98 1958 129 1970
rect 144 1958 247 1970
rect 259 1960 285 1986
rect 300 1981 330 1992
rect 362 1988 424 2004
rect 362 1986 408 1988
rect 362 1970 424 1986
rect 436 1970 442 2018
rect 445 2010 525 2018
rect 445 2008 464 2010
rect 479 2008 513 2010
rect 445 1992 525 2008
rect 445 1970 464 1992
rect 479 1976 509 1992
rect 537 1986 543 2060
rect 546 1986 565 2130
rect 580 1986 586 2130
rect 595 2060 608 2130
rect 660 2126 682 2130
rect 653 2104 682 2118
rect 735 2104 751 2118
rect 789 2114 795 2116
rect 802 2114 910 2130
rect 917 2114 923 2116
rect 931 2114 946 2130
rect 1012 2124 1031 2127
rect 653 2102 751 2104
rect 778 2102 946 2114
rect 961 2104 977 2118
rect 1012 2105 1034 2124
rect 1044 2118 1060 2119
rect 1043 2116 1060 2118
rect 1044 2111 1060 2116
rect 1034 2104 1040 2105
rect 1043 2104 1072 2111
rect 961 2103 1072 2104
rect 961 2102 1078 2103
rect 637 2094 688 2102
rect 735 2094 769 2102
rect 637 2082 662 2094
rect 669 2082 688 2094
rect 742 2092 769 2094
rect 778 2092 999 2102
rect 1034 2099 1040 2102
rect 742 2088 999 2092
rect 637 2074 688 2082
rect 735 2074 999 2088
rect 1043 2094 1078 2102
rect 589 2026 608 2060
rect 653 2066 682 2074
rect 653 2060 670 2066
rect 653 2058 687 2060
rect 735 2058 751 2074
rect 752 2064 960 2074
rect 961 2064 977 2074
rect 1025 2070 1040 2085
rect 1043 2082 1044 2094
rect 1051 2082 1078 2094
rect 1043 2074 1078 2082
rect 1043 2073 1072 2074
rect 763 2060 977 2064
rect 778 2058 977 2060
rect 1012 2060 1025 2070
rect 1043 2060 1060 2073
rect 1012 2058 1060 2060
rect 654 2054 687 2058
rect 650 2052 687 2054
rect 650 2051 717 2052
rect 650 2046 681 2051
rect 687 2046 717 2051
rect 650 2042 717 2046
rect 623 2039 717 2042
rect 623 2032 672 2039
rect 623 2026 653 2032
rect 672 2027 677 2032
rect 589 2010 669 2026
rect 681 2018 717 2039
rect 778 2034 967 2058
rect 1012 2057 1059 2058
rect 1025 2052 1059 2057
rect 793 2031 967 2034
rect 786 2028 967 2031
rect 995 2051 1059 2052
rect 589 2008 608 2010
rect 623 2008 657 2010
rect 589 1992 669 2008
rect 589 1986 608 1992
rect 305 1960 408 1970
rect 259 1958 408 1960
rect 429 1958 464 1970
rect 98 1956 260 1958
rect 110 1936 129 1956
rect 144 1954 174 1956
rect -7 1928 34 1936
rect 116 1932 129 1936
rect 181 1940 260 1956
rect 292 1956 464 1958
rect 292 1940 371 1956
rect 378 1954 408 1956
rect -1 1918 28 1928
rect 43 1918 73 1932
rect 116 1918 159 1932
rect 181 1928 371 1940
rect 436 1936 442 1956
rect 166 1918 196 1928
rect 197 1918 355 1928
rect 359 1918 389 1928
rect 393 1918 423 1932
rect 451 1918 464 1956
rect 536 1970 565 1986
rect 579 1970 608 1986
rect 623 1976 653 1992
rect 681 1970 687 2018
rect 690 2012 709 2018
rect 724 2012 754 2020
rect 690 2004 754 2012
rect 690 1988 770 2004
rect 786 1997 848 2028
rect 864 1997 926 2028
rect 995 2026 1044 2051
rect 1059 2026 1089 2042
rect 958 2012 988 2020
rect 995 2018 1105 2026
rect 958 2004 1003 2012
rect 690 1986 709 1988
rect 724 1986 770 1988
rect 690 1970 770 1986
rect 797 1984 832 1997
rect 873 1994 910 1997
rect 873 1992 915 1994
rect 802 1981 832 1984
rect 811 1977 818 1981
rect 818 1976 819 1977
rect 777 1970 787 1976
rect 536 1962 571 1970
rect 536 1936 537 1962
rect 544 1936 571 1962
rect 479 1918 509 1932
rect 536 1928 571 1936
rect 573 1962 614 1970
rect 573 1936 588 1962
rect 595 1936 614 1962
rect 678 1958 709 1970
rect 724 1958 827 1970
rect 839 1960 865 1986
rect 880 1981 910 1992
rect 942 1988 1004 2004
rect 942 1986 988 1988
rect 942 1970 1004 1986
rect 1016 1970 1022 2018
rect 1025 2010 1105 2018
rect 1025 2008 1044 2010
rect 1059 2008 1093 2010
rect 1025 1992 1105 2008
rect 1025 1970 1044 1992
rect 1059 1976 1089 1992
rect 1117 1986 1123 2060
rect 1126 1986 1145 2130
rect 1160 1986 1166 2130
rect 1175 2060 1188 2130
rect 1240 2126 1262 2130
rect 1233 2104 1262 2118
rect 1315 2104 1331 2118
rect 1369 2114 1375 2116
rect 1382 2114 1490 2130
rect 1497 2114 1503 2116
rect 1511 2114 1526 2130
rect 1592 2124 1611 2127
rect 1233 2102 1331 2104
rect 1358 2102 1526 2114
rect 1541 2104 1557 2118
rect 1592 2105 1614 2124
rect 1624 2118 1640 2119
rect 1623 2116 1640 2118
rect 1624 2111 1640 2116
rect 1614 2104 1620 2105
rect 1623 2104 1652 2111
rect 1541 2103 1652 2104
rect 1541 2102 1658 2103
rect 1217 2094 1268 2102
rect 1315 2094 1349 2102
rect 1217 2082 1242 2094
rect 1249 2082 1268 2094
rect 1322 2092 1349 2094
rect 1358 2092 1579 2102
rect 1614 2099 1620 2102
rect 1322 2088 1579 2092
rect 1217 2074 1268 2082
rect 1315 2074 1579 2088
rect 1623 2094 1658 2102
rect 1169 2026 1188 2060
rect 1233 2066 1262 2074
rect 1233 2060 1250 2066
rect 1233 2058 1267 2060
rect 1315 2058 1331 2074
rect 1332 2064 1540 2074
rect 1541 2064 1557 2074
rect 1605 2070 1620 2085
rect 1623 2082 1624 2094
rect 1631 2082 1658 2094
rect 1623 2074 1658 2082
rect 1623 2073 1652 2074
rect 1343 2060 1557 2064
rect 1358 2058 1557 2060
rect 1592 2060 1605 2070
rect 1623 2060 1640 2073
rect 1592 2058 1640 2060
rect 1234 2054 1267 2058
rect 1230 2052 1267 2054
rect 1230 2051 1297 2052
rect 1230 2046 1261 2051
rect 1267 2046 1297 2051
rect 1230 2042 1297 2046
rect 1203 2039 1297 2042
rect 1203 2032 1252 2039
rect 1203 2026 1233 2032
rect 1252 2027 1257 2032
rect 1169 2010 1249 2026
rect 1261 2018 1297 2039
rect 1358 2034 1547 2058
rect 1592 2057 1639 2058
rect 1605 2052 1639 2057
rect 1373 2031 1547 2034
rect 1366 2028 1547 2031
rect 1575 2051 1639 2052
rect 1169 2008 1188 2010
rect 1203 2008 1237 2010
rect 1169 1992 1249 2008
rect 1169 1986 1188 1992
rect 885 1960 988 1970
rect 839 1958 988 1960
rect 1009 1958 1044 1970
rect 678 1956 840 1958
rect 690 1936 709 1956
rect 724 1954 754 1956
rect 573 1928 614 1936
rect 696 1932 709 1936
rect 761 1940 840 1956
rect 872 1956 1044 1958
rect 872 1940 951 1956
rect 958 1954 988 1956
rect 536 1918 565 1928
rect 579 1918 608 1928
rect 623 1918 653 1932
rect 696 1918 739 1932
rect 761 1928 951 1940
rect 1016 1936 1022 1956
rect 746 1918 776 1928
rect 777 1918 935 1928
rect 939 1918 969 1928
rect 973 1918 1003 1932
rect 1031 1918 1044 1956
rect 1116 1970 1145 1986
rect 1159 1970 1188 1986
rect 1203 1976 1233 1992
rect 1261 1970 1267 2018
rect 1270 2012 1289 2018
rect 1304 2012 1334 2020
rect 1270 2004 1334 2012
rect 1270 1988 1350 2004
rect 1366 1997 1428 2028
rect 1444 1997 1506 2028
rect 1575 2026 1624 2051
rect 1639 2026 1669 2042
rect 1538 2012 1568 2020
rect 1575 2018 1685 2026
rect 1538 2004 1583 2012
rect 1270 1986 1289 1988
rect 1304 1986 1350 1988
rect 1270 1970 1350 1986
rect 1377 1984 1412 1997
rect 1453 1994 1490 1997
rect 1453 1992 1495 1994
rect 1382 1981 1412 1984
rect 1391 1977 1398 1981
rect 1398 1976 1399 1977
rect 1357 1970 1367 1976
rect 1116 1962 1151 1970
rect 1116 1936 1117 1962
rect 1124 1936 1151 1962
rect 1059 1918 1089 1932
rect 1116 1928 1151 1936
rect 1153 1962 1194 1970
rect 1153 1936 1168 1962
rect 1175 1936 1194 1962
rect 1258 1958 1289 1970
rect 1304 1958 1407 1970
rect 1419 1960 1445 1986
rect 1460 1981 1490 1992
rect 1522 1988 1584 2004
rect 1522 1986 1568 1988
rect 1522 1970 1584 1986
rect 1596 1970 1602 2018
rect 1605 2010 1685 2018
rect 1605 2008 1624 2010
rect 1639 2008 1673 2010
rect 1605 1992 1685 2008
rect 1605 1970 1624 1992
rect 1639 1976 1669 1992
rect 1697 1986 1703 2060
rect 1706 1986 1725 2130
rect 1740 1986 1746 2130
rect 1755 2060 1768 2130
rect 1820 2126 1842 2130
rect 1813 2104 1842 2118
rect 1895 2104 1911 2118
rect 1949 2114 1955 2116
rect 1962 2114 2070 2130
rect 2077 2114 2083 2116
rect 2091 2114 2106 2130
rect 2172 2124 2191 2127
rect 1813 2102 1911 2104
rect 1938 2102 2106 2114
rect 2121 2104 2137 2118
rect 2172 2105 2194 2124
rect 2204 2118 2220 2119
rect 2203 2116 2220 2118
rect 2204 2111 2220 2116
rect 2194 2104 2200 2105
rect 2203 2104 2232 2111
rect 2121 2103 2232 2104
rect 2121 2102 2238 2103
rect 1797 2094 1848 2102
rect 1895 2094 1929 2102
rect 1797 2082 1822 2094
rect 1829 2082 1848 2094
rect 1902 2092 1929 2094
rect 1938 2092 2159 2102
rect 2194 2099 2200 2102
rect 1902 2088 2159 2092
rect 1797 2074 1848 2082
rect 1895 2074 2159 2088
rect 2203 2094 2238 2102
rect 1749 2026 1768 2060
rect 1813 2066 1842 2074
rect 1813 2060 1830 2066
rect 1813 2058 1847 2060
rect 1895 2058 1911 2074
rect 1912 2064 2120 2074
rect 2121 2064 2137 2074
rect 2185 2070 2200 2085
rect 2203 2082 2204 2094
rect 2211 2082 2238 2094
rect 2203 2074 2238 2082
rect 2203 2073 2232 2074
rect 1923 2060 2137 2064
rect 1938 2058 2137 2060
rect 2172 2060 2185 2070
rect 2203 2060 2220 2073
rect 2172 2058 2220 2060
rect 1814 2054 1847 2058
rect 1810 2052 1847 2054
rect 1810 2051 1877 2052
rect 1810 2046 1841 2051
rect 1847 2046 1877 2051
rect 1810 2042 1877 2046
rect 1783 2039 1877 2042
rect 1783 2032 1832 2039
rect 1783 2026 1813 2032
rect 1832 2027 1837 2032
rect 1749 2010 1829 2026
rect 1841 2018 1877 2039
rect 1938 2034 2127 2058
rect 2172 2057 2219 2058
rect 2185 2052 2219 2057
rect 1953 2031 2127 2034
rect 1946 2028 2127 2031
rect 2155 2051 2219 2052
rect 1749 2008 1768 2010
rect 1783 2008 1817 2010
rect 1749 1992 1829 2008
rect 1749 1986 1768 1992
rect 1465 1960 1568 1970
rect 1419 1958 1568 1960
rect 1589 1958 1624 1970
rect 1258 1956 1420 1958
rect 1270 1936 1289 1956
rect 1304 1954 1334 1956
rect 1153 1928 1194 1936
rect 1276 1932 1289 1936
rect 1341 1940 1420 1956
rect 1452 1956 1624 1958
rect 1452 1940 1531 1956
rect 1538 1954 1568 1956
rect 1116 1918 1145 1928
rect 1159 1918 1188 1928
rect 1203 1918 1233 1932
rect 1276 1918 1319 1932
rect 1341 1928 1531 1940
rect 1596 1936 1602 1956
rect 1326 1918 1356 1928
rect 1357 1918 1515 1928
rect 1519 1918 1549 1928
rect 1553 1918 1583 1932
rect 1611 1918 1624 1956
rect 1696 1970 1725 1986
rect 1739 1970 1768 1986
rect 1783 1976 1813 1992
rect 1841 1970 1847 2018
rect 1850 2012 1869 2018
rect 1884 2012 1914 2020
rect 1850 2004 1914 2012
rect 1850 1988 1930 2004
rect 1946 1997 2008 2028
rect 2024 1997 2086 2028
rect 2155 2026 2204 2051
rect 2219 2026 2249 2042
rect 2118 2012 2148 2020
rect 2155 2018 2265 2026
rect 2118 2004 2163 2012
rect 1850 1986 1869 1988
rect 1884 1986 1930 1988
rect 1850 1970 1930 1986
rect 1957 1984 1992 1997
rect 2033 1994 2070 1997
rect 2033 1992 2075 1994
rect 1962 1981 1992 1984
rect 1971 1977 1978 1981
rect 1978 1976 1979 1977
rect 1937 1970 1947 1976
rect 1696 1962 1731 1970
rect 1696 1936 1697 1962
rect 1704 1936 1731 1962
rect 1639 1918 1669 1932
rect 1696 1928 1731 1936
rect 1733 1962 1774 1970
rect 1733 1936 1748 1962
rect 1755 1936 1774 1962
rect 1838 1958 1869 1970
rect 1884 1958 1987 1970
rect 1999 1960 2025 1986
rect 2040 1981 2070 1992
rect 2102 1988 2164 2004
rect 2102 1986 2148 1988
rect 2102 1970 2164 1986
rect 2176 1970 2182 2018
rect 2185 2010 2265 2018
rect 2185 2008 2204 2010
rect 2219 2008 2253 2010
rect 2185 1992 2265 2008
rect 2185 1970 2204 1992
rect 2219 1976 2249 1992
rect 2277 1986 2283 2060
rect 2286 1986 2305 2130
rect 2320 1986 2326 2130
rect 2335 2060 2348 2130
rect 2400 2126 2422 2130
rect 2393 2104 2422 2118
rect 2475 2104 2491 2118
rect 2529 2114 2535 2116
rect 2542 2114 2650 2130
rect 2657 2114 2663 2116
rect 2671 2114 2686 2130
rect 2752 2124 2771 2127
rect 2393 2102 2491 2104
rect 2518 2102 2686 2114
rect 2701 2104 2717 2118
rect 2752 2105 2774 2124
rect 2784 2118 2800 2119
rect 2783 2116 2800 2118
rect 2784 2111 2800 2116
rect 2774 2104 2780 2105
rect 2783 2104 2812 2111
rect 2701 2103 2812 2104
rect 2701 2102 2818 2103
rect 2377 2094 2428 2102
rect 2475 2094 2509 2102
rect 2377 2082 2402 2094
rect 2409 2082 2428 2094
rect 2482 2092 2509 2094
rect 2518 2092 2739 2102
rect 2774 2099 2780 2102
rect 2482 2088 2739 2092
rect 2377 2074 2428 2082
rect 2475 2074 2739 2088
rect 2783 2094 2818 2102
rect 2329 2026 2348 2060
rect 2393 2066 2422 2074
rect 2393 2060 2410 2066
rect 2393 2058 2427 2060
rect 2475 2058 2491 2074
rect 2492 2064 2700 2074
rect 2701 2064 2717 2074
rect 2765 2070 2780 2085
rect 2783 2082 2784 2094
rect 2791 2082 2818 2094
rect 2783 2074 2818 2082
rect 2783 2073 2812 2074
rect 2503 2060 2717 2064
rect 2518 2058 2717 2060
rect 2752 2060 2765 2070
rect 2783 2060 2800 2073
rect 2752 2058 2800 2060
rect 2394 2054 2427 2058
rect 2390 2052 2427 2054
rect 2390 2051 2457 2052
rect 2390 2046 2421 2051
rect 2427 2046 2457 2051
rect 2390 2042 2457 2046
rect 2363 2039 2457 2042
rect 2363 2032 2412 2039
rect 2363 2026 2393 2032
rect 2412 2027 2417 2032
rect 2329 2010 2409 2026
rect 2421 2018 2457 2039
rect 2518 2034 2707 2058
rect 2752 2057 2799 2058
rect 2765 2052 2799 2057
rect 2533 2031 2707 2034
rect 2526 2028 2707 2031
rect 2735 2051 2799 2052
rect 2329 2008 2348 2010
rect 2363 2008 2397 2010
rect 2329 1992 2409 2008
rect 2329 1986 2348 1992
rect 2045 1960 2148 1970
rect 1999 1958 2148 1960
rect 2169 1958 2204 1970
rect 1838 1956 2000 1958
rect 1850 1936 1869 1956
rect 1884 1954 1914 1956
rect 1733 1928 1774 1936
rect 1856 1932 1869 1936
rect 1921 1940 2000 1956
rect 2032 1956 2204 1958
rect 2032 1940 2111 1956
rect 2118 1954 2148 1956
rect 1696 1918 1725 1928
rect 1739 1918 1768 1928
rect 1783 1918 1813 1932
rect 1856 1918 1899 1932
rect 1921 1928 2111 1940
rect 2176 1936 2182 1956
rect 1906 1918 1936 1928
rect 1937 1918 2095 1928
rect 2099 1918 2129 1928
rect 2133 1918 2163 1932
rect 2191 1918 2204 1956
rect 2276 1970 2305 1986
rect 2319 1970 2348 1986
rect 2363 1976 2393 1992
rect 2421 1970 2427 2018
rect 2430 2012 2449 2018
rect 2464 2012 2494 2020
rect 2430 2004 2494 2012
rect 2430 1988 2510 2004
rect 2526 1997 2588 2028
rect 2604 1997 2666 2028
rect 2735 2026 2784 2051
rect 2799 2026 2829 2042
rect 2698 2012 2728 2020
rect 2735 2018 2845 2026
rect 2698 2004 2743 2012
rect 2430 1986 2449 1988
rect 2464 1986 2510 1988
rect 2430 1970 2510 1986
rect 2537 1984 2572 1997
rect 2613 1994 2650 1997
rect 2613 1992 2655 1994
rect 2542 1981 2572 1984
rect 2551 1977 2558 1981
rect 2558 1976 2559 1977
rect 2517 1970 2527 1976
rect 2276 1962 2311 1970
rect 2276 1936 2277 1962
rect 2284 1936 2311 1962
rect 2219 1918 2249 1932
rect 2276 1928 2311 1936
rect 2313 1962 2354 1970
rect 2313 1936 2328 1962
rect 2335 1936 2354 1962
rect 2418 1958 2449 1970
rect 2464 1958 2567 1970
rect 2579 1960 2605 1986
rect 2620 1981 2650 1992
rect 2682 1988 2744 2004
rect 2682 1986 2728 1988
rect 2682 1970 2744 1986
rect 2756 1970 2762 2018
rect 2765 2010 2845 2018
rect 2765 2008 2784 2010
rect 2799 2008 2833 2010
rect 2765 1992 2845 2008
rect 2765 1970 2784 1992
rect 2799 1976 2829 1992
rect 2857 1986 2863 2060
rect 2866 1986 2885 2130
rect 2900 1986 2906 2130
rect 2915 2060 2928 2130
rect 2980 2126 3002 2130
rect 2973 2104 3002 2118
rect 3055 2104 3071 2118
rect 3109 2114 3115 2116
rect 3122 2114 3230 2130
rect 3237 2114 3243 2116
rect 3251 2114 3266 2130
rect 3332 2124 3351 2127
rect 2973 2102 3071 2104
rect 3098 2102 3266 2114
rect 3281 2104 3297 2118
rect 3332 2105 3354 2124
rect 3364 2118 3380 2119
rect 3363 2116 3380 2118
rect 3364 2111 3380 2116
rect 3354 2104 3360 2105
rect 3363 2104 3392 2111
rect 3281 2103 3392 2104
rect 3281 2102 3398 2103
rect 2957 2094 3008 2102
rect 3055 2094 3089 2102
rect 2957 2082 2982 2094
rect 2989 2082 3008 2094
rect 3062 2092 3089 2094
rect 3098 2092 3319 2102
rect 3354 2099 3360 2102
rect 3062 2088 3319 2092
rect 2957 2074 3008 2082
rect 3055 2074 3319 2088
rect 3363 2094 3398 2102
rect 2909 2026 2928 2060
rect 2973 2066 3002 2074
rect 2973 2060 2990 2066
rect 2973 2058 3007 2060
rect 3055 2058 3071 2074
rect 3072 2064 3280 2074
rect 3281 2064 3297 2074
rect 3345 2070 3360 2085
rect 3363 2082 3364 2094
rect 3371 2082 3398 2094
rect 3363 2074 3398 2082
rect 3363 2073 3392 2074
rect 3083 2060 3297 2064
rect 3098 2058 3297 2060
rect 3332 2060 3345 2070
rect 3363 2060 3380 2073
rect 3332 2058 3380 2060
rect 2974 2054 3007 2058
rect 2970 2052 3007 2054
rect 2970 2051 3037 2052
rect 2970 2046 3001 2051
rect 3007 2046 3037 2051
rect 2970 2042 3037 2046
rect 2943 2039 3037 2042
rect 2943 2032 2992 2039
rect 2943 2026 2973 2032
rect 2992 2027 2997 2032
rect 2909 2010 2989 2026
rect 3001 2018 3037 2039
rect 3098 2034 3287 2058
rect 3332 2057 3379 2058
rect 3345 2052 3379 2057
rect 3113 2031 3287 2034
rect 3106 2028 3287 2031
rect 3315 2051 3379 2052
rect 2909 2008 2928 2010
rect 2943 2008 2977 2010
rect 2909 1992 2989 2008
rect 2909 1986 2928 1992
rect 2625 1960 2728 1970
rect 2579 1958 2728 1960
rect 2749 1958 2784 1970
rect 2418 1956 2580 1958
rect 2430 1936 2449 1956
rect 2464 1954 2494 1956
rect 2313 1928 2354 1936
rect 2436 1932 2449 1936
rect 2501 1940 2580 1956
rect 2612 1956 2784 1958
rect 2612 1940 2691 1956
rect 2698 1954 2728 1956
rect 2276 1918 2305 1928
rect 2319 1918 2348 1928
rect 2363 1918 2393 1932
rect 2436 1918 2479 1932
rect 2501 1928 2691 1940
rect 2756 1936 2762 1956
rect 2486 1918 2516 1928
rect 2517 1918 2675 1928
rect 2679 1918 2709 1928
rect 2713 1918 2743 1932
rect 2771 1918 2784 1956
rect 2856 1970 2885 1986
rect 2899 1970 2928 1986
rect 2943 1976 2973 1992
rect 3001 1970 3007 2018
rect 3010 2012 3029 2018
rect 3044 2012 3074 2020
rect 3010 2004 3074 2012
rect 3010 1988 3090 2004
rect 3106 1997 3168 2028
rect 3184 1997 3246 2028
rect 3315 2026 3364 2051
rect 3379 2026 3409 2042
rect 3278 2012 3308 2020
rect 3315 2018 3425 2026
rect 3278 2004 3323 2012
rect 3010 1986 3029 1988
rect 3044 1986 3090 1988
rect 3010 1970 3090 1986
rect 3117 1984 3152 1997
rect 3193 1994 3230 1997
rect 3193 1992 3235 1994
rect 3122 1981 3152 1984
rect 3131 1977 3138 1981
rect 3138 1976 3139 1977
rect 3097 1970 3107 1976
rect 2856 1962 2891 1970
rect 2856 1936 2857 1962
rect 2864 1936 2891 1962
rect 2799 1918 2829 1932
rect 2856 1928 2891 1936
rect 2893 1962 2934 1970
rect 2893 1936 2908 1962
rect 2915 1936 2934 1962
rect 2998 1958 3029 1970
rect 3044 1958 3147 1970
rect 3159 1960 3185 1986
rect 3200 1981 3230 1992
rect 3262 1988 3324 2004
rect 3262 1986 3308 1988
rect 3262 1970 3324 1986
rect 3336 1970 3342 2018
rect 3345 2010 3425 2018
rect 3345 2008 3364 2010
rect 3379 2008 3413 2010
rect 3345 1992 3425 2008
rect 3345 1970 3364 1992
rect 3379 1976 3409 1992
rect 3437 1986 3443 2060
rect 3446 1986 3465 2130
rect 3480 1986 3486 2130
rect 3495 2060 3508 2130
rect 3560 2126 3582 2130
rect 3553 2104 3582 2118
rect 3635 2104 3651 2118
rect 3689 2114 3695 2116
rect 3702 2114 3810 2130
rect 3817 2114 3823 2116
rect 3831 2114 3846 2130
rect 3912 2124 3931 2127
rect 3553 2102 3651 2104
rect 3678 2102 3846 2114
rect 3861 2104 3877 2118
rect 3912 2105 3934 2124
rect 3944 2118 3960 2119
rect 3943 2116 3960 2118
rect 3944 2111 3960 2116
rect 3934 2104 3940 2105
rect 3943 2104 3972 2111
rect 3861 2103 3972 2104
rect 3861 2102 3978 2103
rect 3537 2094 3588 2102
rect 3635 2094 3669 2102
rect 3537 2082 3562 2094
rect 3569 2082 3588 2094
rect 3642 2092 3669 2094
rect 3678 2092 3899 2102
rect 3934 2099 3940 2102
rect 3642 2088 3899 2092
rect 3537 2074 3588 2082
rect 3635 2074 3899 2088
rect 3943 2094 3978 2102
rect 3489 2026 3508 2060
rect 3553 2066 3582 2074
rect 3553 2060 3570 2066
rect 3553 2058 3587 2060
rect 3635 2058 3651 2074
rect 3652 2064 3860 2074
rect 3861 2064 3877 2074
rect 3925 2070 3940 2085
rect 3943 2082 3944 2094
rect 3951 2082 3978 2094
rect 3943 2074 3978 2082
rect 3943 2073 3972 2074
rect 3663 2060 3877 2064
rect 3678 2058 3877 2060
rect 3912 2060 3925 2070
rect 3943 2060 3960 2073
rect 3912 2058 3960 2060
rect 3554 2054 3587 2058
rect 3550 2052 3587 2054
rect 3550 2051 3617 2052
rect 3550 2046 3581 2051
rect 3587 2046 3617 2051
rect 3550 2042 3617 2046
rect 3523 2039 3617 2042
rect 3523 2032 3572 2039
rect 3523 2026 3553 2032
rect 3572 2027 3577 2032
rect 3489 2010 3569 2026
rect 3581 2018 3617 2039
rect 3678 2034 3867 2058
rect 3912 2057 3959 2058
rect 3925 2052 3959 2057
rect 3693 2031 3867 2034
rect 3686 2028 3867 2031
rect 3895 2051 3959 2052
rect 3489 2008 3508 2010
rect 3523 2008 3557 2010
rect 3489 1992 3569 2008
rect 3489 1986 3508 1992
rect 3205 1960 3308 1970
rect 3159 1958 3308 1960
rect 3329 1958 3364 1970
rect 2998 1956 3160 1958
rect 3010 1936 3029 1956
rect 3044 1954 3074 1956
rect 2893 1928 2934 1936
rect 3016 1932 3029 1936
rect 3081 1940 3160 1956
rect 3192 1956 3364 1958
rect 3192 1940 3271 1956
rect 3278 1954 3308 1956
rect 2856 1918 2885 1928
rect 2899 1918 2928 1928
rect 2943 1918 2973 1932
rect 3016 1918 3059 1932
rect 3081 1928 3271 1940
rect 3336 1936 3342 1956
rect 3066 1918 3096 1928
rect 3097 1918 3255 1928
rect 3259 1918 3289 1928
rect 3293 1918 3323 1932
rect 3351 1918 3364 1956
rect 3436 1970 3465 1986
rect 3479 1970 3508 1986
rect 3523 1976 3553 1992
rect 3581 1970 3587 2018
rect 3590 2012 3609 2018
rect 3624 2012 3654 2020
rect 3590 2004 3654 2012
rect 3590 1988 3670 2004
rect 3686 1997 3748 2028
rect 3764 1997 3826 2028
rect 3895 2026 3944 2051
rect 3959 2026 3989 2042
rect 3858 2012 3888 2020
rect 3895 2018 4005 2026
rect 3858 2004 3903 2012
rect 3590 1986 3609 1988
rect 3624 1986 3670 1988
rect 3590 1970 3670 1986
rect 3697 1984 3732 1997
rect 3773 1994 3810 1997
rect 3773 1992 3815 1994
rect 3702 1981 3732 1984
rect 3711 1977 3718 1981
rect 3718 1976 3719 1977
rect 3677 1970 3687 1976
rect 3436 1962 3471 1970
rect 3436 1936 3437 1962
rect 3444 1936 3471 1962
rect 3379 1918 3409 1932
rect 3436 1928 3471 1936
rect 3473 1962 3514 1970
rect 3473 1936 3488 1962
rect 3495 1936 3514 1962
rect 3578 1958 3609 1970
rect 3624 1958 3727 1970
rect 3739 1960 3765 1986
rect 3780 1981 3810 1992
rect 3842 1988 3904 2004
rect 3842 1986 3888 1988
rect 3842 1970 3904 1986
rect 3916 1970 3922 2018
rect 3925 2010 4005 2018
rect 3925 2008 3944 2010
rect 3959 2008 3993 2010
rect 3925 1992 4005 2008
rect 3925 1970 3944 1992
rect 3959 1976 3989 1992
rect 4017 1986 4023 2060
rect 4026 1986 4045 2130
rect 4060 1986 4066 2130
rect 4075 2060 4088 2130
rect 4140 2126 4162 2130
rect 4133 2104 4162 2118
rect 4215 2104 4231 2118
rect 4269 2114 4275 2116
rect 4282 2114 4390 2130
rect 4397 2114 4403 2116
rect 4411 2114 4426 2130
rect 4492 2124 4511 2127
rect 4133 2102 4231 2104
rect 4258 2102 4426 2114
rect 4441 2104 4457 2118
rect 4492 2105 4514 2124
rect 4524 2118 4540 2119
rect 4523 2116 4540 2118
rect 4524 2111 4540 2116
rect 4514 2104 4520 2105
rect 4523 2104 4552 2111
rect 4441 2103 4552 2104
rect 4441 2102 4558 2103
rect 4117 2094 4168 2102
rect 4215 2094 4249 2102
rect 4117 2082 4142 2094
rect 4149 2082 4168 2094
rect 4222 2092 4249 2094
rect 4258 2092 4479 2102
rect 4514 2099 4520 2102
rect 4222 2088 4479 2092
rect 4117 2074 4168 2082
rect 4215 2074 4479 2088
rect 4523 2094 4558 2102
rect 4069 2026 4088 2060
rect 4133 2066 4162 2074
rect 4133 2060 4150 2066
rect 4133 2058 4167 2060
rect 4215 2058 4231 2074
rect 4232 2064 4440 2074
rect 4441 2064 4457 2074
rect 4505 2070 4520 2085
rect 4523 2082 4524 2094
rect 4531 2082 4558 2094
rect 4523 2074 4558 2082
rect 4523 2073 4552 2074
rect 4243 2060 4457 2064
rect 4258 2058 4457 2060
rect 4492 2060 4505 2070
rect 4523 2060 4540 2073
rect 4492 2058 4540 2060
rect 4134 2054 4167 2058
rect 4130 2052 4167 2054
rect 4130 2051 4197 2052
rect 4130 2046 4161 2051
rect 4167 2046 4197 2051
rect 4130 2042 4197 2046
rect 4103 2039 4197 2042
rect 4103 2032 4152 2039
rect 4103 2026 4133 2032
rect 4152 2027 4157 2032
rect 4069 2010 4149 2026
rect 4161 2018 4197 2039
rect 4258 2034 4447 2058
rect 4492 2057 4539 2058
rect 4505 2052 4539 2057
rect 4273 2031 4447 2034
rect 4266 2028 4447 2031
rect 4475 2051 4539 2052
rect 4069 2008 4088 2010
rect 4103 2008 4137 2010
rect 4069 1992 4149 2008
rect 4069 1986 4088 1992
rect 3785 1960 3888 1970
rect 3739 1958 3888 1960
rect 3909 1958 3944 1970
rect 3578 1956 3740 1958
rect 3590 1936 3609 1956
rect 3624 1954 3654 1956
rect 3473 1928 3514 1936
rect 3596 1932 3609 1936
rect 3661 1940 3740 1956
rect 3772 1956 3944 1958
rect 3772 1940 3851 1956
rect 3858 1954 3888 1956
rect 3436 1918 3465 1928
rect 3479 1918 3508 1928
rect 3523 1918 3553 1932
rect 3596 1918 3639 1932
rect 3661 1928 3851 1940
rect 3916 1936 3922 1956
rect 3646 1918 3676 1928
rect 3677 1918 3835 1928
rect 3839 1918 3869 1928
rect 3873 1918 3903 1932
rect 3931 1918 3944 1956
rect 4016 1970 4045 1986
rect 4059 1970 4088 1986
rect 4103 1976 4133 1992
rect 4161 1970 4167 2018
rect 4170 2012 4189 2018
rect 4204 2012 4234 2020
rect 4170 2004 4234 2012
rect 4170 1988 4250 2004
rect 4266 1997 4328 2028
rect 4344 1997 4406 2028
rect 4475 2026 4524 2051
rect 4539 2026 4569 2042
rect 4438 2012 4468 2020
rect 4475 2018 4585 2026
rect 4438 2004 4483 2012
rect 4170 1986 4189 1988
rect 4204 1986 4250 1988
rect 4170 1970 4250 1986
rect 4277 1984 4312 1997
rect 4353 1994 4390 1997
rect 4353 1992 4395 1994
rect 4282 1981 4312 1984
rect 4291 1977 4298 1981
rect 4298 1976 4299 1977
rect 4257 1970 4267 1976
rect 4016 1962 4051 1970
rect 4016 1936 4017 1962
rect 4024 1936 4051 1962
rect 3959 1918 3989 1932
rect 4016 1928 4051 1936
rect 4053 1962 4094 1970
rect 4053 1936 4068 1962
rect 4075 1936 4094 1962
rect 4158 1958 4189 1970
rect 4204 1958 4307 1970
rect 4319 1960 4345 1986
rect 4360 1981 4390 1992
rect 4422 1988 4484 2004
rect 4422 1986 4468 1988
rect 4422 1970 4484 1986
rect 4496 1970 4502 2018
rect 4505 2010 4585 2018
rect 4505 2008 4524 2010
rect 4539 2008 4573 2010
rect 4505 1992 4585 2008
rect 4505 1970 4524 1992
rect 4539 1976 4569 1992
rect 4597 1986 4603 2060
rect 4606 1986 4625 2130
rect 4640 1986 4646 2130
rect 4655 2060 4668 2130
rect 4720 2126 4742 2130
rect 4713 2104 4742 2118
rect 4795 2104 4811 2118
rect 4849 2114 4855 2116
rect 4862 2114 4970 2130
rect 4977 2114 4983 2116
rect 4991 2114 5006 2130
rect 5072 2124 5091 2127
rect 4713 2102 4811 2104
rect 4838 2102 5006 2114
rect 5021 2104 5037 2118
rect 5072 2105 5094 2124
rect 5104 2118 5120 2119
rect 5103 2116 5120 2118
rect 5104 2111 5120 2116
rect 5094 2104 5100 2105
rect 5103 2104 5132 2111
rect 5021 2103 5132 2104
rect 5021 2102 5138 2103
rect 4697 2094 4748 2102
rect 4795 2094 4829 2102
rect 4697 2082 4722 2094
rect 4729 2082 4748 2094
rect 4802 2092 4829 2094
rect 4838 2092 5059 2102
rect 5094 2099 5100 2102
rect 4802 2088 5059 2092
rect 4697 2074 4748 2082
rect 4795 2074 5059 2088
rect 5103 2094 5138 2102
rect 4649 2026 4668 2060
rect 4713 2066 4742 2074
rect 4713 2060 4730 2066
rect 4713 2058 4747 2060
rect 4795 2058 4811 2074
rect 4812 2064 5020 2074
rect 5021 2064 5037 2074
rect 5085 2070 5100 2085
rect 5103 2082 5104 2094
rect 5111 2082 5138 2094
rect 5103 2074 5138 2082
rect 5103 2073 5132 2074
rect 4823 2060 5037 2064
rect 4838 2058 5037 2060
rect 5072 2060 5085 2070
rect 5103 2060 5120 2073
rect 5072 2058 5120 2060
rect 4714 2054 4747 2058
rect 4710 2052 4747 2054
rect 4710 2051 4777 2052
rect 4710 2046 4741 2051
rect 4747 2046 4777 2051
rect 4710 2042 4777 2046
rect 4683 2039 4777 2042
rect 4683 2032 4732 2039
rect 4683 2026 4713 2032
rect 4732 2027 4737 2032
rect 4649 2010 4729 2026
rect 4741 2018 4777 2039
rect 4838 2034 5027 2058
rect 5072 2057 5119 2058
rect 5085 2052 5119 2057
rect 4853 2031 5027 2034
rect 4846 2028 5027 2031
rect 5055 2051 5119 2052
rect 4649 2008 4668 2010
rect 4683 2008 4717 2010
rect 4649 1992 4729 2008
rect 4649 1986 4668 1992
rect 4365 1960 4468 1970
rect 4319 1958 4468 1960
rect 4489 1958 4524 1970
rect 4158 1956 4320 1958
rect 4170 1936 4189 1956
rect 4204 1954 4234 1956
rect 4053 1928 4094 1936
rect 4176 1932 4189 1936
rect 4241 1940 4320 1956
rect 4352 1956 4524 1958
rect 4352 1940 4431 1956
rect 4438 1954 4468 1956
rect 4016 1918 4045 1928
rect 4059 1918 4088 1928
rect 4103 1918 4133 1932
rect 4176 1918 4219 1932
rect 4241 1928 4431 1940
rect 4496 1936 4502 1956
rect 4226 1918 4256 1928
rect 4257 1918 4415 1928
rect 4419 1918 4449 1928
rect 4453 1918 4483 1932
rect 4511 1918 4524 1956
rect 4596 1970 4625 1986
rect 4639 1970 4668 1986
rect 4683 1976 4713 1992
rect 4741 1970 4747 2018
rect 4750 2012 4769 2018
rect 4784 2012 4814 2020
rect 4750 2004 4814 2012
rect 4750 1988 4830 2004
rect 4846 1997 4908 2028
rect 4924 1997 4986 2028
rect 5055 2026 5104 2051
rect 5119 2026 5149 2042
rect 5018 2012 5048 2020
rect 5055 2018 5165 2026
rect 5018 2004 5063 2012
rect 4750 1986 4769 1988
rect 4784 1986 4830 1988
rect 4750 1970 4830 1986
rect 4857 1984 4892 1997
rect 4933 1994 4970 1997
rect 4933 1992 4975 1994
rect 4862 1981 4892 1984
rect 4871 1977 4878 1981
rect 4878 1976 4879 1977
rect 4837 1970 4847 1976
rect 4596 1962 4631 1970
rect 4596 1936 4597 1962
rect 4604 1936 4631 1962
rect 4539 1918 4569 1932
rect 4596 1928 4631 1936
rect 4633 1962 4674 1970
rect 4633 1936 4648 1962
rect 4655 1936 4674 1962
rect 4738 1958 4769 1970
rect 4784 1958 4887 1970
rect 4899 1960 4925 1986
rect 4940 1981 4970 1992
rect 5002 1988 5064 2004
rect 5002 1986 5048 1988
rect 5002 1970 5064 1986
rect 5076 1970 5082 2018
rect 5085 2010 5165 2018
rect 5085 2008 5104 2010
rect 5119 2008 5153 2010
rect 5085 1992 5165 2008
rect 5085 1970 5104 1992
rect 5119 1976 5149 1992
rect 5177 1986 5183 2060
rect 5186 1986 5205 2130
rect 5220 1986 5226 2130
rect 5235 2060 5248 2130
rect 5300 2126 5322 2130
rect 5293 2104 5322 2118
rect 5375 2104 5391 2118
rect 5429 2114 5435 2116
rect 5442 2114 5550 2130
rect 5557 2114 5563 2116
rect 5571 2114 5586 2130
rect 5652 2124 5671 2127
rect 5293 2102 5391 2104
rect 5418 2102 5586 2114
rect 5601 2104 5617 2118
rect 5652 2105 5674 2124
rect 5684 2118 5700 2119
rect 5683 2116 5700 2118
rect 5684 2111 5700 2116
rect 5674 2104 5680 2105
rect 5683 2104 5712 2111
rect 5601 2103 5712 2104
rect 5601 2102 5718 2103
rect 5277 2094 5328 2102
rect 5375 2094 5409 2102
rect 5277 2082 5302 2094
rect 5309 2082 5328 2094
rect 5382 2092 5409 2094
rect 5418 2092 5639 2102
rect 5674 2099 5680 2102
rect 5382 2088 5639 2092
rect 5277 2074 5328 2082
rect 5375 2074 5639 2088
rect 5683 2094 5718 2102
rect 5229 2026 5248 2060
rect 5293 2066 5322 2074
rect 5293 2060 5310 2066
rect 5293 2058 5327 2060
rect 5375 2058 5391 2074
rect 5392 2064 5600 2074
rect 5601 2064 5617 2074
rect 5665 2070 5680 2085
rect 5683 2082 5684 2094
rect 5691 2082 5718 2094
rect 5683 2074 5718 2082
rect 5683 2073 5712 2074
rect 5403 2060 5617 2064
rect 5418 2058 5617 2060
rect 5652 2060 5665 2070
rect 5683 2060 5700 2073
rect 5652 2058 5700 2060
rect 5294 2054 5327 2058
rect 5290 2052 5327 2054
rect 5290 2051 5357 2052
rect 5290 2046 5321 2051
rect 5327 2046 5357 2051
rect 5290 2042 5357 2046
rect 5263 2039 5357 2042
rect 5263 2032 5312 2039
rect 5263 2026 5293 2032
rect 5312 2027 5317 2032
rect 5229 2010 5309 2026
rect 5321 2018 5357 2039
rect 5418 2034 5607 2058
rect 5652 2057 5699 2058
rect 5665 2052 5699 2057
rect 5433 2031 5607 2034
rect 5426 2028 5607 2031
rect 5635 2051 5699 2052
rect 5229 2008 5248 2010
rect 5263 2008 5297 2010
rect 5229 1992 5309 2008
rect 5229 1986 5248 1992
rect 4945 1960 5048 1970
rect 4899 1958 5048 1960
rect 5069 1958 5104 1970
rect 4738 1956 4900 1958
rect 4750 1936 4769 1956
rect 4784 1954 4814 1956
rect 4633 1928 4674 1936
rect 4756 1932 4769 1936
rect 4821 1940 4900 1956
rect 4932 1956 5104 1958
rect 4932 1940 5011 1956
rect 5018 1954 5048 1956
rect 4596 1918 4625 1928
rect 4639 1918 4668 1928
rect 4683 1918 4713 1932
rect 4756 1918 4799 1932
rect 4821 1928 5011 1940
rect 5076 1936 5082 1956
rect 4806 1918 4836 1928
rect 4837 1918 4995 1928
rect 4999 1918 5029 1928
rect 5033 1918 5063 1932
rect 5091 1918 5104 1956
rect 5176 1970 5205 1986
rect 5219 1970 5248 1986
rect 5263 1976 5293 1992
rect 5321 1970 5327 2018
rect 5330 2012 5349 2018
rect 5364 2012 5394 2020
rect 5330 2004 5394 2012
rect 5330 1988 5410 2004
rect 5426 1997 5488 2028
rect 5504 1997 5566 2028
rect 5635 2026 5684 2051
rect 5699 2026 5729 2042
rect 5598 2012 5628 2020
rect 5635 2018 5745 2026
rect 5598 2004 5643 2012
rect 5330 1986 5349 1988
rect 5364 1986 5410 1988
rect 5330 1970 5410 1986
rect 5437 1984 5472 1997
rect 5513 1994 5550 1997
rect 5513 1992 5555 1994
rect 5442 1981 5472 1984
rect 5451 1977 5458 1981
rect 5458 1976 5459 1977
rect 5417 1970 5427 1976
rect 5176 1962 5211 1970
rect 5176 1936 5177 1962
rect 5184 1936 5211 1962
rect 5119 1918 5149 1932
rect 5176 1928 5211 1936
rect 5213 1962 5254 1970
rect 5213 1936 5228 1962
rect 5235 1936 5254 1962
rect 5318 1958 5349 1970
rect 5364 1958 5467 1970
rect 5479 1960 5505 1986
rect 5520 1981 5550 1992
rect 5582 1988 5644 2004
rect 5582 1986 5628 1988
rect 5582 1970 5644 1986
rect 5656 1970 5662 2018
rect 5665 2010 5745 2018
rect 5665 2008 5684 2010
rect 5699 2008 5733 2010
rect 5665 1992 5745 2008
rect 5665 1970 5684 1992
rect 5699 1976 5729 1992
rect 5757 1986 5763 2060
rect 5766 1986 5785 2130
rect 5800 1986 5806 2130
rect 5815 2060 5828 2130
rect 5880 2126 5902 2130
rect 5873 2104 5902 2118
rect 5955 2104 5971 2118
rect 6009 2114 6015 2116
rect 6022 2114 6130 2130
rect 6137 2114 6143 2116
rect 6151 2114 6166 2130
rect 6232 2124 6251 2127
rect 5873 2102 5971 2104
rect 5998 2102 6166 2114
rect 6181 2104 6197 2118
rect 6232 2105 6254 2124
rect 6264 2118 6280 2119
rect 6263 2116 6280 2118
rect 6264 2111 6280 2116
rect 6254 2104 6260 2105
rect 6263 2104 6292 2111
rect 6181 2103 6292 2104
rect 6181 2102 6298 2103
rect 5857 2094 5908 2102
rect 5955 2094 5989 2102
rect 5857 2082 5882 2094
rect 5889 2082 5908 2094
rect 5962 2092 5989 2094
rect 5998 2092 6219 2102
rect 6254 2099 6260 2102
rect 5962 2088 6219 2092
rect 5857 2074 5908 2082
rect 5955 2074 6219 2088
rect 6263 2094 6298 2102
rect 5809 2026 5828 2060
rect 5873 2066 5902 2074
rect 5873 2060 5890 2066
rect 5873 2058 5907 2060
rect 5955 2058 5971 2074
rect 5972 2064 6180 2074
rect 6181 2064 6197 2074
rect 6245 2070 6260 2085
rect 6263 2082 6264 2094
rect 6271 2082 6298 2094
rect 6263 2074 6298 2082
rect 6263 2073 6292 2074
rect 5983 2060 6197 2064
rect 5998 2058 6197 2060
rect 6232 2060 6245 2070
rect 6263 2060 6280 2073
rect 6232 2058 6280 2060
rect 5874 2054 5907 2058
rect 5870 2052 5907 2054
rect 5870 2051 5937 2052
rect 5870 2046 5901 2051
rect 5907 2046 5937 2051
rect 5870 2042 5937 2046
rect 5843 2039 5937 2042
rect 5843 2032 5892 2039
rect 5843 2026 5873 2032
rect 5892 2027 5897 2032
rect 5809 2010 5889 2026
rect 5901 2018 5937 2039
rect 5998 2034 6187 2058
rect 6232 2057 6279 2058
rect 6245 2052 6279 2057
rect 6013 2031 6187 2034
rect 6006 2028 6187 2031
rect 6215 2051 6279 2052
rect 5809 2008 5828 2010
rect 5843 2008 5877 2010
rect 5809 1992 5889 2008
rect 5809 1986 5828 1992
rect 5525 1960 5628 1970
rect 5479 1958 5628 1960
rect 5649 1958 5684 1970
rect 5318 1956 5480 1958
rect 5330 1936 5349 1956
rect 5364 1954 5394 1956
rect 5213 1928 5254 1936
rect 5336 1932 5349 1936
rect 5401 1940 5480 1956
rect 5512 1956 5684 1958
rect 5512 1940 5591 1956
rect 5598 1954 5628 1956
rect 5176 1918 5205 1928
rect 5219 1918 5248 1928
rect 5263 1918 5293 1932
rect 5336 1918 5379 1932
rect 5401 1928 5591 1940
rect 5656 1936 5662 1956
rect 5386 1918 5416 1928
rect 5417 1918 5575 1928
rect 5579 1918 5609 1928
rect 5613 1918 5643 1932
rect 5671 1918 5684 1956
rect 5756 1970 5785 1986
rect 5799 1970 5828 1986
rect 5843 1976 5873 1992
rect 5901 1970 5907 2018
rect 5910 2012 5929 2018
rect 5944 2012 5974 2020
rect 5910 2004 5974 2012
rect 5910 1988 5990 2004
rect 6006 1997 6068 2028
rect 6084 1997 6146 2028
rect 6215 2026 6264 2051
rect 6279 2026 6309 2042
rect 6178 2012 6208 2020
rect 6215 2018 6325 2026
rect 6178 2004 6223 2012
rect 5910 1986 5929 1988
rect 5944 1986 5990 1988
rect 5910 1970 5990 1986
rect 6017 1984 6052 1997
rect 6093 1994 6130 1997
rect 6093 1992 6135 1994
rect 6022 1981 6052 1984
rect 6031 1977 6038 1981
rect 6038 1976 6039 1977
rect 5997 1970 6007 1976
rect 5756 1962 5791 1970
rect 5756 1936 5757 1962
rect 5764 1936 5791 1962
rect 5699 1918 5729 1932
rect 5756 1928 5791 1936
rect 5793 1962 5834 1970
rect 5793 1936 5808 1962
rect 5815 1936 5834 1962
rect 5898 1958 5929 1970
rect 5944 1958 6047 1970
rect 6059 1960 6085 1986
rect 6100 1981 6130 1992
rect 6162 1988 6224 2004
rect 6162 1986 6208 1988
rect 6162 1970 6224 1986
rect 6236 1970 6242 2018
rect 6245 2010 6325 2018
rect 6245 2008 6264 2010
rect 6279 2008 6313 2010
rect 6245 1992 6325 2008
rect 6245 1970 6264 1992
rect 6279 1976 6309 1992
rect 6337 1986 6343 2060
rect 6346 1986 6365 2130
rect 6380 1986 6386 2130
rect 6395 2060 6408 2130
rect 6460 2126 6482 2130
rect 6453 2104 6482 2118
rect 6535 2104 6551 2118
rect 6589 2114 6595 2116
rect 6602 2114 6710 2130
rect 6717 2114 6723 2116
rect 6731 2114 6746 2130
rect 6812 2124 6831 2127
rect 6453 2102 6551 2104
rect 6578 2102 6746 2114
rect 6761 2104 6777 2118
rect 6812 2105 6834 2124
rect 6844 2118 6860 2119
rect 6843 2116 6860 2118
rect 6844 2111 6860 2116
rect 6834 2104 6840 2105
rect 6843 2104 6872 2111
rect 6761 2103 6872 2104
rect 6761 2102 6878 2103
rect 6437 2094 6488 2102
rect 6535 2094 6569 2102
rect 6437 2082 6462 2094
rect 6469 2082 6488 2094
rect 6542 2092 6569 2094
rect 6578 2092 6799 2102
rect 6834 2099 6840 2102
rect 6542 2088 6799 2092
rect 6437 2074 6488 2082
rect 6535 2074 6799 2088
rect 6843 2094 6878 2102
rect 6389 2026 6408 2060
rect 6453 2066 6482 2074
rect 6453 2060 6470 2066
rect 6453 2058 6487 2060
rect 6535 2058 6551 2074
rect 6552 2064 6760 2074
rect 6761 2064 6777 2074
rect 6825 2070 6840 2085
rect 6843 2082 6844 2094
rect 6851 2082 6878 2094
rect 6843 2074 6878 2082
rect 6843 2073 6872 2074
rect 6563 2060 6777 2064
rect 6578 2058 6777 2060
rect 6812 2060 6825 2070
rect 6843 2060 6860 2073
rect 6812 2058 6860 2060
rect 6454 2054 6487 2058
rect 6450 2052 6487 2054
rect 6450 2051 6517 2052
rect 6450 2046 6481 2051
rect 6487 2046 6517 2051
rect 6450 2042 6517 2046
rect 6423 2039 6517 2042
rect 6423 2032 6472 2039
rect 6423 2026 6453 2032
rect 6472 2027 6477 2032
rect 6389 2010 6469 2026
rect 6481 2018 6517 2039
rect 6578 2034 6767 2058
rect 6812 2057 6859 2058
rect 6825 2052 6859 2057
rect 6593 2031 6767 2034
rect 6586 2028 6767 2031
rect 6795 2051 6859 2052
rect 6389 2008 6408 2010
rect 6423 2008 6457 2010
rect 6389 1992 6469 2008
rect 6389 1986 6408 1992
rect 6105 1960 6208 1970
rect 6059 1958 6208 1960
rect 6229 1958 6264 1970
rect 5898 1956 6060 1958
rect 5910 1936 5929 1956
rect 5944 1954 5974 1956
rect 5793 1928 5834 1936
rect 5916 1932 5929 1936
rect 5981 1940 6060 1956
rect 6092 1956 6264 1958
rect 6092 1940 6171 1956
rect 6178 1954 6208 1956
rect 5756 1918 5785 1928
rect 5799 1918 5828 1928
rect 5843 1918 5873 1932
rect 5916 1918 5959 1932
rect 5981 1928 6171 1940
rect 6236 1936 6242 1956
rect 5966 1918 5996 1928
rect 5997 1918 6155 1928
rect 6159 1918 6189 1928
rect 6193 1918 6223 1932
rect 6251 1918 6264 1956
rect 6336 1970 6365 1986
rect 6379 1970 6408 1986
rect 6423 1976 6453 1992
rect 6481 1970 6487 2018
rect 6490 2012 6509 2018
rect 6524 2012 6554 2020
rect 6490 2004 6554 2012
rect 6490 1988 6570 2004
rect 6586 1997 6648 2028
rect 6664 1997 6726 2028
rect 6795 2026 6844 2051
rect 6859 2026 6889 2042
rect 6758 2012 6788 2020
rect 6795 2018 6905 2026
rect 6758 2004 6803 2012
rect 6490 1986 6509 1988
rect 6524 1986 6570 1988
rect 6490 1970 6570 1986
rect 6597 1984 6632 1997
rect 6673 1994 6710 1997
rect 6673 1992 6715 1994
rect 6602 1981 6632 1984
rect 6611 1977 6618 1981
rect 6618 1976 6619 1977
rect 6577 1970 6587 1976
rect 6336 1962 6371 1970
rect 6336 1936 6337 1962
rect 6344 1936 6371 1962
rect 6279 1918 6309 1932
rect 6336 1928 6371 1936
rect 6373 1962 6414 1970
rect 6373 1936 6388 1962
rect 6395 1936 6414 1962
rect 6478 1958 6509 1970
rect 6524 1958 6627 1970
rect 6639 1960 6665 1986
rect 6680 1981 6710 1992
rect 6742 1988 6804 2004
rect 6742 1986 6788 1988
rect 6742 1970 6804 1986
rect 6816 1970 6822 2018
rect 6825 2010 6905 2018
rect 6825 2008 6844 2010
rect 6859 2008 6893 2010
rect 6825 1992 6905 2008
rect 6825 1970 6844 1992
rect 6859 1976 6889 1992
rect 6917 1986 6923 2060
rect 6926 1986 6945 2130
rect 6960 1986 6966 2130
rect 6975 2060 6988 2130
rect 7040 2126 7062 2130
rect 7033 2104 7062 2118
rect 7115 2104 7131 2118
rect 7169 2114 7175 2116
rect 7182 2114 7290 2130
rect 7297 2114 7303 2116
rect 7311 2114 7326 2130
rect 7392 2124 7411 2127
rect 7033 2102 7131 2104
rect 7158 2102 7326 2114
rect 7341 2104 7357 2118
rect 7392 2105 7414 2124
rect 7424 2118 7440 2119
rect 7423 2116 7440 2118
rect 7424 2111 7440 2116
rect 7414 2104 7420 2105
rect 7423 2104 7452 2111
rect 7341 2103 7452 2104
rect 7341 2102 7458 2103
rect 7017 2094 7068 2102
rect 7115 2094 7149 2102
rect 7017 2082 7042 2094
rect 7049 2082 7068 2094
rect 7122 2092 7149 2094
rect 7158 2092 7379 2102
rect 7414 2099 7420 2102
rect 7122 2088 7379 2092
rect 7017 2074 7068 2082
rect 7115 2074 7379 2088
rect 7423 2094 7458 2102
rect 6969 2026 6988 2060
rect 7033 2066 7062 2074
rect 7033 2060 7050 2066
rect 7033 2058 7067 2060
rect 7115 2058 7131 2074
rect 7132 2064 7340 2074
rect 7341 2064 7357 2074
rect 7405 2070 7420 2085
rect 7423 2082 7424 2094
rect 7431 2082 7458 2094
rect 7423 2074 7458 2082
rect 7423 2073 7452 2074
rect 7151 2060 7357 2064
rect 7158 2058 7357 2060
rect 7392 2060 7405 2070
rect 7423 2060 7440 2073
rect 7392 2058 7440 2060
rect 7034 2054 7067 2058
rect 7030 2052 7067 2054
rect 7030 2051 7097 2052
rect 7030 2046 7061 2051
rect 7067 2046 7097 2051
rect 7030 2042 7097 2046
rect 7003 2039 7097 2042
rect 7003 2032 7052 2039
rect 7003 2026 7033 2032
rect 7052 2027 7057 2032
rect 6969 2010 7049 2026
rect 7061 2018 7097 2039
rect 7158 2034 7347 2058
rect 7392 2057 7439 2058
rect 7405 2052 7439 2057
rect 7173 2031 7347 2034
rect 7166 2028 7347 2031
rect 7375 2051 7439 2052
rect 6969 2008 6988 2010
rect 7003 2008 7037 2010
rect 6969 1992 7049 2008
rect 6969 1986 6988 1992
rect 6685 1960 6788 1970
rect 6639 1958 6788 1960
rect 6809 1958 6844 1970
rect 6478 1956 6640 1958
rect 6490 1936 6509 1956
rect 6524 1954 6554 1956
rect 6373 1928 6414 1936
rect 6496 1932 6509 1936
rect 6561 1940 6640 1956
rect 6672 1956 6844 1958
rect 6672 1940 6751 1956
rect 6758 1954 6788 1956
rect 6336 1918 6365 1928
rect 6379 1918 6408 1928
rect 6423 1918 6453 1932
rect 6496 1918 6539 1932
rect 6561 1928 6751 1940
rect 6816 1936 6822 1956
rect 6546 1918 6576 1928
rect 6577 1918 6735 1928
rect 6739 1918 6769 1928
rect 6773 1918 6803 1932
rect 6831 1918 6844 1956
rect 6916 1970 6945 1986
rect 6959 1970 6988 1986
rect 7003 1976 7033 1992
rect 7061 1970 7067 2018
rect 7070 2012 7089 2018
rect 7104 2012 7134 2020
rect 7070 2004 7134 2012
rect 7070 1988 7150 2004
rect 7166 1997 7228 2028
rect 7244 1997 7306 2028
rect 7375 2026 7424 2051
rect 7439 2026 7469 2042
rect 7338 2012 7368 2020
rect 7375 2018 7485 2026
rect 7338 2004 7383 2012
rect 7070 1986 7089 1988
rect 7104 1986 7150 1988
rect 7070 1970 7150 1986
rect 7177 1984 7212 1997
rect 7253 1994 7290 1997
rect 7253 1992 7295 1994
rect 7182 1981 7212 1984
rect 7191 1977 7198 1981
rect 7198 1976 7199 1977
rect 7157 1970 7167 1976
rect 6916 1962 6951 1970
rect 6916 1936 6917 1962
rect 6924 1936 6951 1962
rect 6859 1918 6889 1932
rect 6916 1928 6951 1936
rect 6953 1962 6994 1970
rect 6953 1936 6968 1962
rect 6975 1936 6994 1962
rect 7058 1958 7089 1970
rect 7104 1958 7207 1970
rect 7219 1960 7245 1986
rect 7260 1981 7290 1992
rect 7322 1988 7384 2004
rect 7322 1986 7368 1988
rect 7322 1970 7384 1986
rect 7396 1970 7402 2018
rect 7405 2010 7485 2018
rect 7405 2008 7424 2010
rect 7439 2008 7473 2010
rect 7405 1992 7485 2008
rect 7405 1970 7424 1992
rect 7439 1976 7469 1992
rect 7497 1986 7503 2060
rect 7506 1986 7525 2130
rect 7540 1986 7546 2130
rect 7555 2060 7568 2130
rect 7620 2126 7642 2130
rect 7613 2104 7642 2118
rect 7695 2104 7711 2118
rect 7749 2114 7755 2116
rect 7762 2114 7870 2130
rect 7877 2114 7883 2116
rect 7891 2114 7906 2130
rect 7972 2124 7991 2127
rect 7613 2102 7711 2104
rect 7738 2102 7906 2114
rect 7921 2104 7937 2118
rect 7972 2105 7994 2124
rect 8004 2118 8020 2119
rect 8003 2116 8020 2118
rect 8004 2111 8020 2116
rect 7994 2104 8000 2105
rect 8003 2104 8032 2111
rect 7921 2103 8032 2104
rect 7921 2102 8038 2103
rect 7597 2094 7648 2102
rect 7695 2094 7729 2102
rect 7597 2082 7622 2094
rect 7629 2082 7648 2094
rect 7702 2092 7729 2094
rect 7738 2092 7959 2102
rect 7994 2099 8000 2102
rect 7702 2088 7959 2092
rect 7597 2074 7648 2082
rect 7695 2074 7959 2088
rect 8003 2094 8038 2102
rect 7549 2026 7568 2060
rect 7613 2066 7642 2074
rect 7613 2060 7630 2066
rect 7613 2058 7647 2060
rect 7695 2058 7711 2074
rect 7712 2064 7920 2074
rect 7921 2064 7937 2074
rect 7985 2070 8000 2085
rect 8003 2082 8004 2094
rect 8011 2082 8038 2094
rect 8003 2074 8038 2082
rect 8003 2073 8032 2074
rect 7723 2060 7937 2064
rect 7738 2058 7937 2060
rect 7972 2060 7985 2070
rect 8003 2060 8020 2073
rect 7972 2058 8020 2060
rect 7614 2054 7647 2058
rect 7610 2052 7647 2054
rect 7610 2051 7677 2052
rect 7610 2046 7641 2051
rect 7647 2046 7677 2051
rect 7610 2042 7677 2046
rect 7583 2039 7677 2042
rect 7583 2032 7632 2039
rect 7583 2026 7613 2032
rect 7632 2027 7637 2032
rect 7549 2010 7629 2026
rect 7641 2018 7677 2039
rect 7738 2034 7927 2058
rect 7972 2057 8019 2058
rect 7985 2052 8019 2057
rect 7753 2031 7927 2034
rect 7746 2028 7927 2031
rect 7955 2051 8019 2052
rect 7549 2008 7568 2010
rect 7583 2008 7617 2010
rect 7549 1992 7629 2008
rect 7549 1986 7568 1992
rect 7265 1960 7368 1970
rect 7219 1958 7368 1960
rect 7389 1958 7424 1970
rect 7058 1956 7220 1958
rect 7070 1936 7089 1956
rect 7104 1954 7134 1956
rect 6953 1928 6994 1936
rect 7076 1932 7089 1936
rect 7141 1940 7220 1956
rect 7252 1956 7424 1958
rect 7252 1940 7331 1956
rect 7338 1954 7368 1956
rect 6916 1918 6945 1928
rect 6959 1918 6988 1928
rect 7003 1918 7033 1932
rect 7076 1918 7119 1932
rect 7141 1928 7331 1940
rect 7396 1936 7402 1956
rect 7126 1918 7156 1928
rect 7157 1918 7315 1928
rect 7319 1918 7349 1928
rect 7353 1918 7383 1932
rect 7411 1918 7424 1956
rect 7496 1970 7525 1986
rect 7539 1970 7568 1986
rect 7583 1976 7613 1992
rect 7641 1970 7647 2018
rect 7650 2012 7669 2018
rect 7684 2012 7714 2020
rect 7650 2004 7714 2012
rect 7650 1988 7730 2004
rect 7746 1997 7808 2028
rect 7824 1997 7886 2028
rect 7955 2026 8004 2051
rect 8019 2026 8049 2042
rect 7918 2012 7948 2020
rect 7955 2018 8065 2026
rect 7918 2004 7963 2012
rect 7650 1986 7669 1988
rect 7684 1986 7730 1988
rect 7650 1970 7730 1986
rect 7757 1984 7792 1997
rect 7833 1994 7870 1997
rect 7833 1992 7875 1994
rect 7762 1981 7792 1984
rect 7771 1977 7778 1981
rect 7778 1976 7779 1977
rect 7737 1970 7747 1976
rect 7496 1962 7531 1970
rect 7496 1936 7497 1962
rect 7504 1936 7531 1962
rect 7439 1918 7469 1932
rect 7496 1928 7531 1936
rect 7533 1962 7574 1970
rect 7533 1936 7548 1962
rect 7555 1936 7574 1962
rect 7638 1958 7669 1970
rect 7684 1958 7787 1970
rect 7799 1960 7825 1986
rect 7840 1981 7870 1992
rect 7902 1988 7964 2004
rect 7902 1986 7948 1988
rect 7902 1970 7964 1986
rect 7976 1970 7982 2018
rect 7985 2010 8065 2018
rect 7985 2008 8004 2010
rect 8019 2008 8053 2010
rect 7985 1992 8065 2008
rect 7985 1970 8004 1992
rect 8019 1976 8049 1992
rect 8077 1986 8083 2060
rect 8086 1986 8105 2130
rect 8120 1986 8126 2130
rect 8135 2060 8148 2130
rect 8200 2126 8222 2130
rect 8193 2104 8222 2118
rect 8275 2104 8291 2118
rect 8329 2114 8335 2116
rect 8342 2114 8450 2130
rect 8457 2114 8463 2116
rect 8471 2114 8486 2130
rect 8552 2124 8571 2127
rect 8193 2102 8291 2104
rect 8318 2102 8486 2114
rect 8501 2104 8517 2118
rect 8552 2105 8574 2124
rect 8584 2118 8600 2119
rect 8583 2116 8600 2118
rect 8584 2111 8600 2116
rect 8574 2104 8580 2105
rect 8583 2104 8612 2111
rect 8501 2103 8612 2104
rect 8501 2102 8618 2103
rect 8177 2094 8228 2102
rect 8275 2094 8309 2102
rect 8177 2082 8202 2094
rect 8209 2082 8228 2094
rect 8282 2092 8309 2094
rect 8318 2092 8539 2102
rect 8574 2099 8580 2102
rect 8282 2088 8539 2092
rect 8177 2074 8228 2082
rect 8275 2074 8539 2088
rect 8583 2094 8618 2102
rect 8129 2026 8148 2060
rect 8193 2066 8222 2074
rect 8193 2060 8210 2066
rect 8193 2058 8227 2060
rect 8275 2058 8291 2074
rect 8292 2064 8500 2074
rect 8501 2064 8517 2074
rect 8565 2070 8580 2085
rect 8583 2082 8584 2094
rect 8591 2082 8618 2094
rect 8583 2074 8618 2082
rect 8583 2073 8612 2074
rect 8303 2060 8517 2064
rect 8318 2058 8517 2060
rect 8552 2060 8565 2070
rect 8583 2060 8600 2073
rect 8552 2058 8600 2060
rect 8194 2054 8227 2058
rect 8190 2052 8227 2054
rect 8190 2051 8257 2052
rect 8190 2046 8221 2051
rect 8227 2046 8257 2051
rect 8190 2042 8257 2046
rect 8163 2039 8257 2042
rect 8163 2032 8212 2039
rect 8163 2026 8193 2032
rect 8212 2027 8217 2032
rect 8129 2010 8209 2026
rect 8221 2018 8257 2039
rect 8318 2034 8507 2058
rect 8552 2057 8599 2058
rect 8565 2052 8599 2057
rect 8333 2031 8507 2034
rect 8326 2028 8507 2031
rect 8535 2051 8599 2052
rect 8129 2008 8148 2010
rect 8163 2008 8197 2010
rect 8129 1992 8209 2008
rect 8129 1986 8148 1992
rect 7845 1960 7948 1970
rect 7799 1958 7948 1960
rect 7969 1958 8004 1970
rect 7638 1956 7800 1958
rect 7650 1936 7669 1956
rect 7684 1954 7714 1956
rect 7533 1928 7574 1936
rect 7656 1932 7669 1936
rect 7721 1940 7800 1956
rect 7832 1956 8004 1958
rect 7832 1940 7911 1956
rect 7918 1954 7948 1956
rect 7496 1918 7525 1928
rect 7539 1918 7568 1928
rect 7583 1918 7613 1932
rect 7656 1918 7699 1932
rect 7721 1928 7911 1940
rect 7976 1936 7982 1956
rect 7706 1918 7736 1928
rect 7737 1918 7895 1928
rect 7899 1918 7929 1928
rect 7933 1918 7963 1932
rect 7991 1918 8004 1956
rect 8076 1970 8105 1986
rect 8119 1970 8148 1986
rect 8163 1976 8193 1992
rect 8221 1970 8227 2018
rect 8230 2012 8249 2018
rect 8264 2012 8294 2020
rect 8230 2004 8294 2012
rect 8230 1988 8310 2004
rect 8326 1997 8388 2028
rect 8404 1997 8466 2028
rect 8535 2026 8584 2051
rect 8599 2026 8629 2042
rect 8498 2012 8528 2020
rect 8535 2018 8645 2026
rect 8498 2004 8543 2012
rect 8230 1986 8249 1988
rect 8264 1986 8310 1988
rect 8230 1970 8310 1986
rect 8337 1984 8372 1997
rect 8413 1994 8450 1997
rect 8413 1992 8455 1994
rect 8342 1981 8372 1984
rect 8351 1977 8358 1981
rect 8358 1976 8359 1977
rect 8317 1970 8327 1976
rect 8076 1962 8111 1970
rect 8076 1936 8077 1962
rect 8084 1936 8111 1962
rect 8019 1918 8049 1932
rect 8076 1928 8111 1936
rect 8113 1962 8154 1970
rect 8113 1936 8128 1962
rect 8135 1936 8154 1962
rect 8218 1958 8249 1970
rect 8264 1958 8367 1970
rect 8379 1960 8405 1986
rect 8420 1981 8450 1992
rect 8482 1988 8544 2004
rect 8482 1986 8528 1988
rect 8482 1970 8544 1986
rect 8556 1970 8562 2018
rect 8565 2010 8645 2018
rect 8565 2008 8584 2010
rect 8599 2008 8633 2010
rect 8565 1992 8645 2008
rect 8565 1970 8584 1992
rect 8599 1976 8629 1992
rect 8657 1986 8663 2060
rect 8666 1986 8685 2130
rect 8700 1986 8706 2130
rect 8715 2060 8728 2130
rect 8780 2126 8802 2130
rect 8773 2104 8802 2118
rect 8855 2104 8871 2118
rect 8909 2114 8915 2116
rect 8922 2114 9030 2130
rect 9037 2114 9043 2116
rect 9051 2114 9066 2130
rect 9132 2124 9151 2127
rect 8773 2102 8871 2104
rect 8898 2102 9066 2114
rect 9081 2104 9097 2118
rect 9132 2105 9154 2124
rect 9164 2118 9180 2119
rect 9163 2116 9180 2118
rect 9164 2111 9180 2116
rect 9154 2104 9160 2105
rect 9163 2104 9192 2111
rect 9081 2103 9192 2104
rect 9081 2102 9198 2103
rect 8757 2094 8808 2102
rect 8855 2094 8889 2102
rect 8757 2082 8782 2094
rect 8789 2082 8808 2094
rect 8862 2092 8889 2094
rect 8898 2092 9119 2102
rect 9154 2099 9160 2102
rect 8862 2088 9119 2092
rect 8757 2074 8808 2082
rect 8855 2074 9119 2088
rect 9163 2094 9198 2102
rect 8709 2026 8728 2060
rect 8773 2066 8802 2074
rect 8773 2060 8790 2066
rect 8773 2058 8807 2060
rect 8855 2058 8871 2074
rect 8872 2064 9080 2074
rect 9081 2064 9097 2074
rect 9145 2070 9160 2085
rect 9163 2082 9164 2094
rect 9171 2082 9198 2094
rect 9163 2074 9198 2082
rect 9163 2073 9192 2074
rect 8883 2060 9097 2064
rect 8898 2058 9097 2060
rect 9132 2060 9145 2070
rect 9163 2060 9180 2073
rect 9132 2058 9180 2060
rect 8774 2054 8807 2058
rect 8770 2052 8807 2054
rect 8770 2051 8837 2052
rect 8770 2046 8801 2051
rect 8807 2046 8837 2051
rect 8770 2042 8837 2046
rect 8743 2039 8837 2042
rect 8743 2032 8792 2039
rect 8743 2026 8773 2032
rect 8792 2027 8797 2032
rect 8709 2010 8789 2026
rect 8801 2018 8837 2039
rect 8898 2034 9087 2058
rect 9132 2057 9179 2058
rect 9145 2052 9179 2057
rect 8913 2031 9087 2034
rect 8906 2028 9087 2031
rect 9115 2051 9179 2052
rect 8709 2008 8728 2010
rect 8743 2008 8777 2010
rect 8709 1992 8789 2008
rect 8709 1986 8728 1992
rect 8425 1960 8528 1970
rect 8379 1958 8528 1960
rect 8549 1958 8584 1970
rect 8218 1956 8380 1958
rect 8230 1936 8249 1956
rect 8264 1954 8294 1956
rect 8113 1928 8154 1936
rect 8236 1932 8249 1936
rect 8301 1940 8380 1956
rect 8412 1956 8584 1958
rect 8412 1940 8491 1956
rect 8498 1954 8528 1956
rect 8076 1918 8105 1928
rect 8119 1918 8148 1928
rect 8163 1918 8193 1932
rect 8236 1918 8279 1932
rect 8301 1928 8491 1940
rect 8556 1936 8562 1956
rect 8286 1918 8316 1928
rect 8317 1918 8475 1928
rect 8479 1918 8509 1928
rect 8513 1918 8543 1932
rect 8571 1918 8584 1956
rect 8656 1970 8685 1986
rect 8699 1970 8728 1986
rect 8743 1976 8773 1992
rect 8801 1970 8807 2018
rect 8810 2012 8829 2018
rect 8844 2012 8874 2020
rect 8810 2004 8874 2012
rect 8810 1988 8890 2004
rect 8906 1997 8968 2028
rect 8984 1997 9046 2028
rect 9115 2026 9164 2051
rect 9179 2026 9209 2042
rect 9078 2012 9108 2020
rect 9115 2018 9225 2026
rect 9078 2004 9123 2012
rect 8810 1986 8829 1988
rect 8844 1986 8890 1988
rect 8810 1970 8890 1986
rect 8917 1984 8952 1997
rect 8993 1994 9030 1997
rect 8993 1992 9035 1994
rect 8922 1981 8952 1984
rect 8931 1977 8938 1981
rect 8938 1976 8939 1977
rect 8897 1970 8907 1976
rect 8656 1962 8691 1970
rect 8656 1936 8657 1962
rect 8664 1936 8691 1962
rect 8599 1918 8629 1932
rect 8656 1928 8691 1936
rect 8693 1962 8734 1970
rect 8693 1936 8708 1962
rect 8715 1936 8734 1962
rect 8798 1958 8829 1970
rect 8844 1958 8947 1970
rect 8959 1960 8985 1986
rect 9000 1981 9030 1992
rect 9062 1988 9124 2004
rect 9062 1986 9108 1988
rect 9062 1970 9124 1986
rect 9136 1970 9142 2018
rect 9145 2010 9225 2018
rect 9145 2008 9164 2010
rect 9179 2008 9213 2010
rect 9145 1992 9225 2008
rect 9145 1970 9164 1992
rect 9179 1976 9209 1992
rect 9237 1986 9243 2060
rect 9246 1986 9265 2130
rect 9280 1986 9286 2130
rect 9295 2060 9308 2130
rect 9360 2126 9382 2130
rect 9353 2104 9382 2118
rect 9435 2104 9451 2118
rect 9489 2114 9495 2116
rect 9502 2114 9610 2130
rect 9617 2114 9623 2116
rect 9631 2114 9646 2130
rect 9712 2124 9731 2127
rect 9353 2102 9451 2104
rect 9478 2102 9646 2114
rect 9661 2104 9677 2118
rect 9712 2105 9734 2124
rect 9744 2118 9760 2119
rect 9743 2116 9760 2118
rect 9744 2111 9760 2116
rect 9734 2104 9740 2105
rect 9743 2104 9772 2111
rect 9661 2103 9772 2104
rect 9661 2102 9778 2103
rect 9337 2094 9388 2102
rect 9435 2094 9469 2102
rect 9337 2082 9362 2094
rect 9369 2082 9388 2094
rect 9442 2092 9469 2094
rect 9478 2092 9699 2102
rect 9734 2099 9740 2102
rect 9442 2088 9699 2092
rect 9337 2074 9388 2082
rect 9435 2074 9699 2088
rect 9743 2094 9778 2102
rect 9289 2026 9308 2060
rect 9353 2066 9382 2074
rect 9353 2060 9370 2066
rect 9353 2058 9387 2060
rect 9435 2058 9451 2074
rect 9452 2064 9660 2074
rect 9661 2064 9677 2074
rect 9725 2070 9740 2085
rect 9743 2082 9744 2094
rect 9751 2082 9778 2094
rect 9743 2074 9778 2082
rect 9743 2073 9772 2074
rect 9463 2060 9677 2064
rect 9478 2058 9677 2060
rect 9712 2060 9725 2070
rect 9743 2060 9760 2073
rect 9712 2058 9760 2060
rect 9354 2054 9387 2058
rect 9350 2052 9387 2054
rect 9350 2051 9417 2052
rect 9350 2046 9381 2051
rect 9387 2046 9417 2051
rect 9350 2042 9417 2046
rect 9323 2039 9417 2042
rect 9323 2032 9372 2039
rect 9323 2026 9353 2032
rect 9372 2027 9377 2032
rect 9289 2010 9369 2026
rect 9381 2018 9417 2039
rect 9478 2034 9667 2058
rect 9712 2057 9759 2058
rect 9725 2052 9759 2057
rect 9493 2031 9667 2034
rect 9486 2028 9667 2031
rect 9695 2051 9759 2052
rect 9289 2008 9308 2010
rect 9323 2008 9357 2010
rect 9289 1992 9369 2008
rect 9289 1986 9308 1992
rect 9005 1960 9108 1970
rect 8959 1958 9108 1960
rect 9129 1958 9164 1970
rect 8798 1956 8960 1958
rect 8810 1936 8829 1956
rect 8844 1954 8874 1956
rect 8693 1928 8734 1936
rect 8816 1932 8829 1936
rect 8881 1940 8960 1956
rect 8992 1956 9164 1958
rect 8992 1940 9071 1956
rect 9078 1954 9108 1956
rect 8656 1918 8685 1928
rect 8699 1918 8728 1928
rect 8743 1918 8773 1932
rect 8816 1918 8859 1932
rect 8881 1928 9071 1940
rect 9136 1936 9142 1956
rect 8866 1918 8896 1928
rect 8897 1918 9055 1928
rect 9059 1918 9089 1928
rect 9093 1918 9123 1932
rect 9151 1918 9164 1956
rect 9236 1970 9265 1986
rect 9279 1970 9308 1986
rect 9323 1976 9353 1992
rect 9381 1970 9387 2018
rect 9390 2012 9409 2018
rect 9424 2012 9454 2020
rect 9390 2004 9454 2012
rect 9390 1988 9470 2004
rect 9486 1997 9548 2028
rect 9564 1997 9626 2028
rect 9695 2026 9744 2051
rect 9759 2026 9789 2042
rect 9658 2012 9688 2020
rect 9695 2018 9805 2026
rect 9658 2004 9703 2012
rect 9390 1986 9409 1988
rect 9424 1986 9470 1988
rect 9390 1970 9470 1986
rect 9497 1984 9532 1997
rect 9573 1994 9610 1997
rect 9573 1992 9615 1994
rect 9502 1981 9532 1984
rect 9511 1977 9518 1981
rect 9518 1976 9519 1977
rect 9477 1970 9487 1976
rect 9236 1962 9271 1970
rect 9236 1936 9237 1962
rect 9244 1936 9271 1962
rect 9179 1918 9209 1932
rect 9236 1928 9271 1936
rect 9273 1962 9314 1970
rect 9273 1936 9288 1962
rect 9295 1936 9314 1962
rect 9378 1958 9409 1970
rect 9424 1958 9527 1970
rect 9539 1960 9565 1986
rect 9580 1981 9610 1992
rect 9642 1988 9704 2004
rect 9642 1986 9688 1988
rect 9642 1970 9704 1986
rect 9716 1970 9722 2018
rect 9725 2010 9805 2018
rect 9725 2008 9744 2010
rect 9759 2008 9793 2010
rect 9725 1992 9805 2008
rect 9725 1970 9744 1992
rect 9759 1976 9789 1992
rect 9817 1986 9823 2060
rect 9826 1986 9845 2130
rect 9860 1986 9866 2130
rect 9875 2060 9888 2130
rect 9940 2126 9962 2130
rect 9933 2104 9962 2118
rect 10015 2104 10031 2118
rect 10069 2114 10075 2116
rect 10082 2114 10190 2130
rect 10197 2114 10203 2116
rect 10211 2114 10226 2130
rect 10292 2124 10311 2127
rect 9933 2102 10031 2104
rect 10058 2102 10226 2114
rect 10241 2104 10257 2118
rect 10292 2105 10314 2124
rect 10324 2118 10340 2119
rect 10323 2116 10340 2118
rect 10324 2111 10340 2116
rect 10314 2104 10320 2105
rect 10323 2104 10352 2111
rect 10241 2103 10352 2104
rect 10241 2102 10358 2103
rect 9917 2094 9968 2102
rect 10015 2094 10049 2102
rect 9917 2082 9942 2094
rect 9949 2082 9968 2094
rect 10022 2092 10049 2094
rect 10058 2092 10279 2102
rect 10314 2099 10320 2102
rect 10022 2088 10279 2092
rect 9917 2074 9968 2082
rect 10015 2074 10279 2088
rect 10323 2094 10358 2102
rect 9869 2026 9888 2060
rect 9933 2066 9962 2074
rect 9933 2060 9950 2066
rect 9933 2058 9967 2060
rect 10015 2058 10031 2074
rect 10032 2064 10240 2074
rect 10241 2064 10257 2074
rect 10305 2070 10320 2085
rect 10323 2082 10324 2094
rect 10331 2082 10358 2094
rect 10323 2074 10358 2082
rect 10323 2073 10352 2074
rect 10043 2060 10257 2064
rect 10058 2058 10257 2060
rect 10292 2060 10305 2070
rect 10323 2060 10340 2073
rect 10292 2058 10340 2060
rect 9934 2054 9967 2058
rect 9930 2052 9967 2054
rect 9930 2051 9997 2052
rect 9930 2046 9961 2051
rect 9967 2046 9997 2051
rect 9930 2042 9997 2046
rect 9903 2039 9997 2042
rect 9903 2032 9952 2039
rect 9903 2026 9933 2032
rect 9952 2027 9957 2032
rect 9869 2010 9949 2026
rect 9961 2018 9997 2039
rect 10058 2034 10247 2058
rect 10292 2057 10339 2058
rect 10305 2052 10339 2057
rect 10073 2031 10247 2034
rect 10066 2028 10247 2031
rect 10275 2051 10339 2052
rect 9869 2008 9888 2010
rect 9903 2008 9937 2010
rect 9869 1992 9949 2008
rect 9869 1986 9888 1992
rect 9585 1960 9688 1970
rect 9539 1958 9688 1960
rect 9709 1958 9744 1970
rect 9378 1956 9540 1958
rect 9390 1936 9409 1956
rect 9424 1954 9454 1956
rect 9273 1928 9314 1936
rect 9396 1932 9409 1936
rect 9461 1940 9540 1956
rect 9572 1956 9744 1958
rect 9572 1940 9651 1956
rect 9658 1954 9688 1956
rect 9236 1918 9265 1928
rect 9279 1918 9308 1928
rect 9323 1918 9353 1932
rect 9396 1918 9439 1932
rect 9461 1928 9651 1940
rect 9716 1936 9722 1956
rect 9446 1918 9476 1928
rect 9477 1918 9635 1928
rect 9639 1918 9669 1928
rect 9673 1918 9703 1932
rect 9731 1918 9744 1956
rect 9816 1970 9845 1986
rect 9859 1970 9888 1986
rect 9903 1976 9933 1992
rect 9961 1970 9967 2018
rect 9970 2012 9989 2018
rect 10004 2012 10034 2020
rect 9970 2004 10034 2012
rect 9970 1988 10050 2004
rect 10066 1997 10128 2028
rect 10144 1997 10206 2028
rect 10275 2026 10324 2051
rect 10339 2026 10369 2042
rect 10238 2012 10268 2020
rect 10275 2018 10385 2026
rect 10238 2004 10283 2012
rect 9970 1986 9989 1988
rect 10004 1986 10050 1988
rect 9970 1970 10050 1986
rect 10077 1984 10112 1997
rect 10153 1994 10190 1997
rect 10153 1992 10195 1994
rect 10082 1981 10112 1984
rect 10091 1977 10098 1981
rect 10098 1976 10099 1977
rect 10057 1970 10067 1976
rect 9816 1962 9851 1970
rect 9816 1936 9817 1962
rect 9824 1936 9851 1962
rect 9759 1918 9789 1932
rect 9816 1928 9851 1936
rect 9853 1962 9894 1970
rect 9853 1936 9868 1962
rect 9875 1936 9894 1962
rect 9958 1958 9989 1970
rect 10004 1958 10107 1970
rect 10119 1960 10145 1986
rect 10160 1981 10190 1992
rect 10222 1988 10284 2004
rect 10222 1986 10268 1988
rect 10222 1970 10284 1986
rect 10296 1970 10302 2018
rect 10305 2010 10385 2018
rect 10305 2008 10324 2010
rect 10339 2008 10373 2010
rect 10305 1992 10385 2008
rect 10305 1970 10324 1992
rect 10339 1976 10369 1992
rect 10397 1986 10403 2060
rect 10406 1986 10425 2130
rect 10440 1986 10446 2130
rect 10455 2060 10468 2130
rect 10520 2126 10542 2130
rect 10513 2104 10542 2118
rect 10595 2104 10611 2118
rect 10649 2114 10655 2116
rect 10662 2114 10770 2130
rect 10777 2114 10783 2116
rect 10791 2114 10806 2130
rect 10872 2124 10891 2127
rect 10513 2102 10611 2104
rect 10638 2102 10806 2114
rect 10821 2104 10837 2118
rect 10872 2105 10894 2124
rect 10904 2118 10920 2119
rect 10903 2116 10920 2118
rect 10904 2111 10920 2116
rect 10894 2104 10900 2105
rect 10903 2104 10932 2111
rect 10821 2103 10932 2104
rect 10821 2102 10938 2103
rect 10497 2094 10548 2102
rect 10595 2094 10629 2102
rect 10497 2082 10522 2094
rect 10529 2082 10548 2094
rect 10602 2092 10629 2094
rect 10638 2092 10859 2102
rect 10894 2099 10900 2102
rect 10602 2088 10859 2092
rect 10497 2074 10548 2082
rect 10595 2074 10859 2088
rect 10903 2094 10938 2102
rect 10449 2026 10468 2060
rect 10513 2066 10542 2074
rect 10513 2060 10530 2066
rect 10513 2058 10547 2060
rect 10595 2058 10611 2074
rect 10612 2064 10820 2074
rect 10821 2064 10837 2074
rect 10885 2070 10900 2085
rect 10903 2082 10904 2094
rect 10911 2082 10938 2094
rect 10903 2074 10938 2082
rect 10903 2073 10932 2074
rect 10623 2060 10837 2064
rect 10638 2058 10837 2060
rect 10872 2060 10885 2070
rect 10903 2060 10920 2073
rect 10872 2058 10920 2060
rect 10514 2054 10547 2058
rect 10510 2052 10547 2054
rect 10510 2051 10577 2052
rect 10510 2046 10541 2051
rect 10547 2046 10577 2051
rect 10510 2042 10577 2046
rect 10483 2039 10577 2042
rect 10483 2032 10532 2039
rect 10483 2026 10513 2032
rect 10532 2027 10537 2032
rect 10449 2010 10529 2026
rect 10541 2018 10577 2039
rect 10638 2034 10827 2058
rect 10872 2057 10919 2058
rect 10885 2052 10919 2057
rect 10653 2031 10827 2034
rect 10646 2028 10827 2031
rect 10855 2051 10919 2052
rect 10449 2008 10468 2010
rect 10483 2008 10517 2010
rect 10449 1992 10529 2008
rect 10449 1986 10468 1992
rect 10165 1960 10268 1970
rect 10119 1958 10268 1960
rect 10289 1958 10324 1970
rect 9958 1956 10120 1958
rect 9970 1936 9989 1956
rect 10004 1954 10034 1956
rect 9853 1928 9894 1936
rect 9976 1932 9989 1936
rect 10041 1940 10120 1956
rect 10152 1956 10324 1958
rect 10152 1940 10231 1956
rect 10238 1954 10268 1956
rect 9816 1918 9845 1928
rect 9859 1918 9888 1928
rect 9903 1918 9933 1932
rect 9976 1918 10019 1932
rect 10041 1928 10231 1940
rect 10296 1936 10302 1956
rect 10026 1918 10056 1928
rect 10057 1918 10215 1928
rect 10219 1918 10249 1928
rect 10253 1918 10283 1932
rect 10311 1918 10324 1956
rect 10396 1970 10425 1986
rect 10439 1970 10468 1986
rect 10483 1976 10513 1992
rect 10541 1970 10547 2018
rect 10550 2012 10569 2018
rect 10584 2012 10614 2020
rect 10550 2004 10614 2012
rect 10550 1988 10630 2004
rect 10646 1997 10708 2028
rect 10724 1997 10786 2028
rect 10855 2026 10904 2051
rect 10919 2026 10949 2042
rect 10818 2012 10848 2020
rect 10855 2018 10965 2026
rect 10818 2004 10863 2012
rect 10550 1986 10569 1988
rect 10584 1986 10630 1988
rect 10550 1970 10630 1986
rect 10657 1984 10692 1997
rect 10733 1994 10770 1997
rect 10733 1992 10775 1994
rect 10662 1981 10692 1984
rect 10671 1977 10678 1981
rect 10678 1976 10679 1977
rect 10637 1970 10647 1976
rect 10396 1962 10431 1970
rect 10396 1936 10397 1962
rect 10404 1936 10431 1962
rect 10339 1918 10369 1932
rect 10396 1928 10431 1936
rect 10433 1962 10474 1970
rect 10433 1936 10448 1962
rect 10455 1936 10474 1962
rect 10538 1958 10569 1970
rect 10584 1958 10687 1970
rect 10699 1960 10725 1986
rect 10740 1981 10770 1992
rect 10802 1988 10864 2004
rect 10802 1986 10848 1988
rect 10802 1970 10864 1986
rect 10876 1970 10882 2018
rect 10885 2010 10965 2018
rect 10885 2008 10904 2010
rect 10919 2008 10953 2010
rect 10885 1992 10965 2008
rect 10885 1970 10904 1992
rect 10919 1976 10949 1992
rect 10977 1986 10983 2060
rect 10986 1986 11005 2130
rect 11020 1986 11026 2130
rect 11035 2060 11048 2130
rect 11100 2126 11122 2130
rect 11093 2104 11122 2118
rect 11175 2104 11191 2118
rect 11229 2114 11235 2116
rect 11242 2114 11350 2130
rect 11357 2114 11363 2116
rect 11371 2114 11386 2130
rect 11452 2124 11471 2127
rect 11093 2102 11191 2104
rect 11218 2102 11386 2114
rect 11401 2104 11417 2118
rect 11452 2105 11474 2124
rect 11484 2118 11500 2119
rect 11483 2116 11500 2118
rect 11484 2111 11500 2116
rect 11474 2104 11480 2105
rect 11483 2104 11512 2111
rect 11401 2103 11512 2104
rect 11401 2102 11518 2103
rect 11077 2094 11128 2102
rect 11175 2094 11209 2102
rect 11077 2082 11102 2094
rect 11109 2082 11128 2094
rect 11182 2092 11209 2094
rect 11218 2092 11439 2102
rect 11474 2099 11480 2102
rect 11182 2088 11439 2092
rect 11077 2074 11128 2082
rect 11175 2074 11439 2088
rect 11483 2094 11518 2102
rect 11029 2026 11048 2060
rect 11093 2066 11122 2074
rect 11093 2060 11110 2066
rect 11093 2058 11127 2060
rect 11175 2058 11191 2074
rect 11192 2064 11400 2074
rect 11401 2064 11417 2074
rect 11465 2070 11480 2085
rect 11483 2082 11484 2094
rect 11491 2082 11518 2094
rect 11483 2074 11518 2082
rect 11483 2073 11512 2074
rect 11203 2060 11417 2064
rect 11218 2058 11417 2060
rect 11452 2060 11465 2070
rect 11483 2060 11500 2073
rect 11452 2058 11500 2060
rect 11094 2054 11127 2058
rect 11090 2052 11127 2054
rect 11090 2051 11157 2052
rect 11090 2046 11121 2051
rect 11127 2046 11157 2051
rect 11090 2042 11157 2046
rect 11063 2039 11157 2042
rect 11063 2032 11112 2039
rect 11063 2026 11093 2032
rect 11112 2027 11117 2032
rect 11029 2010 11109 2026
rect 11121 2018 11157 2039
rect 11218 2034 11407 2058
rect 11452 2057 11499 2058
rect 11465 2052 11499 2057
rect 11233 2031 11407 2034
rect 11226 2028 11407 2031
rect 11435 2051 11499 2052
rect 11029 2008 11048 2010
rect 11063 2008 11097 2010
rect 11029 1992 11109 2008
rect 11029 1986 11048 1992
rect 10745 1960 10848 1970
rect 10699 1958 10848 1960
rect 10869 1958 10904 1970
rect 10538 1956 10700 1958
rect 10550 1936 10569 1956
rect 10584 1954 10614 1956
rect 10433 1928 10474 1936
rect 10556 1932 10569 1936
rect 10621 1940 10700 1956
rect 10732 1956 10904 1958
rect 10732 1940 10811 1956
rect 10818 1954 10848 1956
rect 10396 1918 10425 1928
rect 10439 1918 10468 1928
rect 10483 1918 10513 1932
rect 10556 1918 10599 1932
rect 10621 1928 10811 1940
rect 10876 1936 10882 1956
rect 10606 1918 10636 1928
rect 10637 1918 10795 1928
rect 10799 1918 10829 1928
rect 10833 1918 10863 1932
rect 10891 1918 10904 1956
rect 10976 1970 11005 1986
rect 11019 1970 11048 1986
rect 11063 1976 11093 1992
rect 11121 1970 11127 2018
rect 11130 2012 11149 2018
rect 11164 2012 11194 2020
rect 11130 2004 11194 2012
rect 11130 1988 11210 2004
rect 11226 1997 11288 2028
rect 11304 1997 11366 2028
rect 11435 2026 11484 2051
rect 11499 2026 11529 2042
rect 11398 2012 11428 2020
rect 11435 2018 11545 2026
rect 11398 2004 11443 2012
rect 11130 1986 11149 1988
rect 11164 1986 11210 1988
rect 11130 1970 11210 1986
rect 11237 1984 11272 1997
rect 11313 1994 11350 1997
rect 11313 1992 11355 1994
rect 11242 1981 11272 1984
rect 11251 1977 11258 1981
rect 11258 1976 11259 1977
rect 11217 1970 11227 1976
rect 10976 1962 11011 1970
rect 10976 1936 10977 1962
rect 10984 1936 11011 1962
rect 10919 1918 10949 1932
rect 10976 1928 11011 1936
rect 11013 1962 11054 1970
rect 11013 1936 11028 1962
rect 11035 1936 11054 1962
rect 11118 1958 11149 1970
rect 11164 1958 11267 1970
rect 11279 1960 11305 1986
rect 11320 1981 11350 1992
rect 11382 1988 11444 2004
rect 11382 1986 11428 1988
rect 11382 1970 11444 1986
rect 11456 1970 11462 2018
rect 11465 2010 11545 2018
rect 11465 2008 11484 2010
rect 11499 2008 11533 2010
rect 11465 1992 11545 2008
rect 11465 1970 11484 1992
rect 11499 1976 11529 1992
rect 11557 1986 11563 2060
rect 11566 1986 11585 2130
rect 11600 1986 11606 2130
rect 11615 2060 11628 2130
rect 11680 2126 11702 2130
rect 11673 2104 11702 2118
rect 11755 2104 11771 2118
rect 11809 2114 11815 2116
rect 11822 2114 11930 2130
rect 11937 2114 11943 2116
rect 11951 2114 11966 2130
rect 12032 2124 12051 2127
rect 11673 2102 11771 2104
rect 11798 2102 11966 2114
rect 11981 2104 11997 2118
rect 12032 2105 12054 2124
rect 12064 2118 12080 2119
rect 12063 2116 12080 2118
rect 12064 2111 12080 2116
rect 12054 2104 12060 2105
rect 12063 2104 12092 2111
rect 11981 2103 12092 2104
rect 11981 2102 12098 2103
rect 11657 2094 11708 2102
rect 11755 2094 11789 2102
rect 11657 2082 11682 2094
rect 11689 2082 11708 2094
rect 11762 2092 11789 2094
rect 11798 2092 12019 2102
rect 12054 2099 12060 2102
rect 11762 2088 12019 2092
rect 11657 2074 11708 2082
rect 11755 2074 12019 2088
rect 12063 2094 12098 2102
rect 11609 2026 11628 2060
rect 11673 2066 11702 2074
rect 11673 2060 11690 2066
rect 11673 2058 11707 2060
rect 11755 2058 11771 2074
rect 11772 2064 11980 2074
rect 11981 2064 11997 2074
rect 12045 2070 12060 2085
rect 12063 2082 12064 2094
rect 12071 2082 12098 2094
rect 12063 2074 12098 2082
rect 12063 2073 12092 2074
rect 11783 2060 11997 2064
rect 11798 2058 11997 2060
rect 12032 2060 12045 2070
rect 12063 2060 12080 2073
rect 12032 2058 12080 2060
rect 11674 2054 11707 2058
rect 11670 2052 11707 2054
rect 11670 2051 11737 2052
rect 11670 2046 11701 2051
rect 11707 2046 11737 2051
rect 11670 2042 11737 2046
rect 11643 2039 11737 2042
rect 11643 2032 11692 2039
rect 11643 2026 11673 2032
rect 11692 2027 11697 2032
rect 11609 2010 11689 2026
rect 11701 2018 11737 2039
rect 11798 2034 11987 2058
rect 12032 2057 12079 2058
rect 12045 2052 12079 2057
rect 11813 2031 11987 2034
rect 11806 2028 11987 2031
rect 12015 2051 12079 2052
rect 11609 2008 11628 2010
rect 11643 2008 11677 2010
rect 11609 1992 11689 2008
rect 11609 1986 11628 1992
rect 11325 1960 11428 1970
rect 11279 1958 11428 1960
rect 11449 1958 11484 1970
rect 11118 1956 11280 1958
rect 11130 1936 11149 1956
rect 11164 1954 11194 1956
rect 11013 1928 11054 1936
rect 11136 1932 11149 1936
rect 11201 1940 11280 1956
rect 11312 1956 11484 1958
rect 11312 1940 11391 1956
rect 11398 1954 11428 1956
rect 10976 1918 11005 1928
rect 11019 1918 11048 1928
rect 11063 1918 11093 1932
rect 11136 1918 11179 1932
rect 11201 1928 11391 1940
rect 11456 1936 11462 1956
rect 11186 1918 11216 1928
rect 11217 1918 11375 1928
rect 11379 1918 11409 1928
rect 11413 1918 11443 1932
rect 11471 1918 11484 1956
rect 11556 1970 11585 1986
rect 11599 1970 11628 1986
rect 11643 1976 11673 1992
rect 11701 1970 11707 2018
rect 11710 2012 11729 2018
rect 11744 2012 11774 2020
rect 11710 2004 11774 2012
rect 11710 1988 11790 2004
rect 11806 1997 11868 2028
rect 11884 1997 11946 2028
rect 12015 2026 12064 2051
rect 12079 2026 12109 2042
rect 11978 2012 12008 2020
rect 12015 2018 12125 2026
rect 11978 2004 12023 2012
rect 11710 1986 11729 1988
rect 11744 1986 11790 1988
rect 11710 1970 11790 1986
rect 11817 1984 11852 1997
rect 11893 1994 11930 1997
rect 11893 1992 11935 1994
rect 11822 1981 11852 1984
rect 11831 1977 11838 1981
rect 11838 1976 11839 1977
rect 11797 1970 11807 1976
rect 11556 1962 11591 1970
rect 11556 1936 11557 1962
rect 11564 1936 11591 1962
rect 11499 1918 11529 1932
rect 11556 1928 11591 1936
rect 11593 1962 11634 1970
rect 11593 1936 11608 1962
rect 11615 1936 11634 1962
rect 11698 1958 11729 1970
rect 11744 1958 11847 1970
rect 11859 1960 11885 1986
rect 11900 1981 11930 1992
rect 11962 1988 12024 2004
rect 11962 1986 12008 1988
rect 11962 1970 12024 1986
rect 12036 1970 12042 2018
rect 12045 2010 12125 2018
rect 12045 2008 12064 2010
rect 12079 2008 12113 2010
rect 12045 1992 12125 2008
rect 12045 1970 12064 1992
rect 12079 1976 12109 1992
rect 12137 1986 12143 2060
rect 12146 1986 12165 2130
rect 12180 1986 12186 2130
rect 12195 2060 12208 2130
rect 12260 2126 12282 2130
rect 12253 2104 12282 2118
rect 12335 2104 12351 2118
rect 12389 2114 12395 2116
rect 12402 2114 12510 2130
rect 12517 2114 12523 2116
rect 12531 2114 12546 2130
rect 12612 2124 12631 2127
rect 12253 2102 12351 2104
rect 12378 2102 12546 2114
rect 12561 2104 12577 2118
rect 12612 2105 12634 2124
rect 12644 2118 12660 2119
rect 12643 2116 12660 2118
rect 12644 2111 12660 2116
rect 12634 2104 12640 2105
rect 12643 2104 12672 2111
rect 12561 2103 12672 2104
rect 12561 2102 12678 2103
rect 12237 2094 12288 2102
rect 12335 2094 12369 2102
rect 12237 2082 12262 2094
rect 12269 2082 12288 2094
rect 12342 2092 12369 2094
rect 12378 2092 12599 2102
rect 12634 2099 12640 2102
rect 12342 2088 12599 2092
rect 12237 2074 12288 2082
rect 12335 2074 12599 2088
rect 12643 2094 12678 2102
rect 12189 2026 12208 2060
rect 12253 2066 12282 2074
rect 12253 2060 12270 2066
rect 12253 2058 12287 2060
rect 12335 2058 12351 2074
rect 12352 2064 12560 2074
rect 12561 2064 12577 2074
rect 12625 2070 12640 2085
rect 12643 2082 12644 2094
rect 12651 2082 12678 2094
rect 12643 2074 12678 2082
rect 12643 2073 12672 2074
rect 12363 2060 12577 2064
rect 12378 2058 12577 2060
rect 12612 2060 12625 2070
rect 12643 2060 12660 2073
rect 12612 2058 12660 2060
rect 12254 2054 12287 2058
rect 12250 2052 12287 2054
rect 12250 2051 12317 2052
rect 12250 2046 12281 2051
rect 12287 2046 12317 2051
rect 12250 2042 12317 2046
rect 12223 2039 12317 2042
rect 12223 2032 12272 2039
rect 12223 2026 12253 2032
rect 12272 2027 12277 2032
rect 12189 2010 12269 2026
rect 12281 2018 12317 2039
rect 12378 2034 12567 2058
rect 12612 2057 12659 2058
rect 12625 2052 12659 2057
rect 12393 2031 12567 2034
rect 12386 2028 12567 2031
rect 12595 2051 12659 2052
rect 12189 2008 12208 2010
rect 12223 2008 12257 2010
rect 12189 1992 12269 2008
rect 12189 1986 12208 1992
rect 11905 1960 12008 1970
rect 11859 1958 12008 1960
rect 12029 1958 12064 1970
rect 11698 1956 11860 1958
rect 11710 1936 11729 1956
rect 11744 1954 11774 1956
rect 11593 1928 11634 1936
rect 11716 1932 11729 1936
rect 11781 1940 11860 1956
rect 11892 1956 12064 1958
rect 11892 1940 11971 1956
rect 11978 1954 12008 1956
rect 11556 1918 11585 1928
rect 11599 1918 11628 1928
rect 11643 1918 11673 1932
rect 11716 1918 11759 1932
rect 11781 1928 11971 1940
rect 12036 1936 12042 1956
rect 11766 1918 11796 1928
rect 11797 1918 11955 1928
rect 11959 1918 11989 1928
rect 11993 1918 12023 1932
rect 12051 1918 12064 1956
rect 12136 1970 12165 1986
rect 12179 1970 12208 1986
rect 12223 1976 12253 1992
rect 12281 1970 12287 2018
rect 12290 2012 12309 2018
rect 12324 2012 12354 2020
rect 12290 2004 12354 2012
rect 12290 1988 12370 2004
rect 12386 1997 12448 2028
rect 12464 1997 12526 2028
rect 12595 2026 12644 2051
rect 12659 2026 12689 2042
rect 12558 2012 12588 2020
rect 12595 2018 12705 2026
rect 12558 2004 12603 2012
rect 12290 1986 12309 1988
rect 12324 1986 12370 1988
rect 12290 1970 12370 1986
rect 12397 1984 12432 1997
rect 12473 1994 12510 1997
rect 12473 1992 12515 1994
rect 12402 1981 12432 1984
rect 12411 1977 12418 1981
rect 12418 1976 12419 1977
rect 12377 1970 12387 1976
rect 12136 1962 12171 1970
rect 12136 1936 12137 1962
rect 12144 1936 12171 1962
rect 12079 1918 12109 1932
rect 12136 1928 12171 1936
rect 12173 1962 12214 1970
rect 12173 1936 12188 1962
rect 12195 1936 12214 1962
rect 12278 1958 12309 1970
rect 12324 1958 12427 1970
rect 12439 1960 12465 1986
rect 12480 1981 12510 1992
rect 12542 1988 12604 2004
rect 12542 1986 12588 1988
rect 12542 1970 12604 1986
rect 12616 1970 12622 2018
rect 12625 2010 12705 2018
rect 12625 2008 12644 2010
rect 12659 2008 12693 2010
rect 12625 1992 12705 2008
rect 12625 1970 12644 1992
rect 12659 1976 12689 1992
rect 12717 1986 12723 2060
rect 12726 1986 12745 2130
rect 12760 1986 12766 2130
rect 12775 2060 12788 2130
rect 12840 2126 12862 2130
rect 12833 2104 12862 2118
rect 12915 2104 12931 2118
rect 12969 2114 12975 2116
rect 12982 2114 13090 2130
rect 13097 2114 13103 2116
rect 13111 2114 13126 2130
rect 13192 2124 13211 2127
rect 12833 2102 12931 2104
rect 12958 2102 13126 2114
rect 13141 2104 13157 2118
rect 13192 2105 13214 2124
rect 13224 2118 13240 2119
rect 13223 2116 13240 2118
rect 13224 2111 13240 2116
rect 13214 2104 13220 2105
rect 13223 2104 13252 2111
rect 13141 2103 13252 2104
rect 13141 2102 13258 2103
rect 12817 2094 12868 2102
rect 12915 2094 12949 2102
rect 12817 2082 12842 2094
rect 12849 2082 12868 2094
rect 12922 2092 12949 2094
rect 12958 2092 13179 2102
rect 13214 2099 13220 2102
rect 12922 2088 13179 2092
rect 12817 2074 12868 2082
rect 12915 2074 13179 2088
rect 13223 2094 13258 2102
rect 12769 2026 12788 2060
rect 12833 2066 12862 2074
rect 12833 2060 12850 2066
rect 12833 2058 12867 2060
rect 12915 2058 12931 2074
rect 12932 2064 13140 2074
rect 13141 2064 13157 2074
rect 13205 2070 13220 2085
rect 13223 2082 13224 2094
rect 13231 2082 13258 2094
rect 13223 2074 13258 2082
rect 13223 2073 13252 2074
rect 12943 2060 13157 2064
rect 12958 2058 13157 2060
rect 13192 2060 13205 2070
rect 13223 2060 13240 2073
rect 13192 2058 13240 2060
rect 12834 2054 12867 2058
rect 12830 2052 12867 2054
rect 12830 2051 12897 2052
rect 12830 2046 12861 2051
rect 12867 2046 12897 2051
rect 12830 2042 12897 2046
rect 12803 2039 12897 2042
rect 12803 2032 12852 2039
rect 12803 2026 12833 2032
rect 12852 2027 12857 2032
rect 12769 2010 12849 2026
rect 12861 2018 12897 2039
rect 12958 2034 13147 2058
rect 13192 2057 13239 2058
rect 13205 2052 13239 2057
rect 12973 2031 13147 2034
rect 12966 2028 13147 2031
rect 13175 2051 13239 2052
rect 12769 2008 12788 2010
rect 12803 2008 12837 2010
rect 12769 1992 12849 2008
rect 12769 1986 12788 1992
rect 12485 1960 12588 1970
rect 12439 1958 12588 1960
rect 12609 1958 12644 1970
rect 12278 1956 12440 1958
rect 12290 1936 12309 1956
rect 12324 1954 12354 1956
rect 12173 1928 12214 1936
rect 12296 1932 12309 1936
rect 12361 1940 12440 1956
rect 12472 1956 12644 1958
rect 12472 1940 12551 1956
rect 12558 1954 12588 1956
rect 12136 1918 12165 1928
rect 12179 1918 12208 1928
rect 12223 1918 12253 1932
rect 12296 1918 12339 1932
rect 12361 1928 12551 1940
rect 12616 1936 12622 1956
rect 12346 1918 12376 1928
rect 12377 1918 12535 1928
rect 12539 1918 12569 1928
rect 12573 1918 12603 1932
rect 12631 1918 12644 1956
rect 12716 1970 12745 1986
rect 12759 1970 12788 1986
rect 12803 1976 12833 1992
rect 12861 1970 12867 2018
rect 12870 2012 12889 2018
rect 12904 2012 12934 2020
rect 12870 2004 12934 2012
rect 12870 1988 12950 2004
rect 12966 1997 13028 2028
rect 13044 1997 13106 2028
rect 13175 2026 13224 2051
rect 13239 2026 13269 2042
rect 13138 2012 13168 2020
rect 13175 2018 13285 2026
rect 13138 2004 13183 2012
rect 12870 1986 12889 1988
rect 12904 1986 12950 1988
rect 12870 1970 12950 1986
rect 12977 1984 13012 1997
rect 13053 1994 13090 1997
rect 13053 1992 13095 1994
rect 12982 1981 13012 1984
rect 12991 1977 12998 1981
rect 12998 1976 12999 1977
rect 12957 1970 12967 1976
rect 12716 1962 12751 1970
rect 12716 1936 12717 1962
rect 12724 1936 12751 1962
rect 12659 1918 12689 1932
rect 12716 1928 12751 1936
rect 12753 1962 12794 1970
rect 12753 1936 12768 1962
rect 12775 1936 12794 1962
rect 12858 1958 12889 1970
rect 12904 1958 13007 1970
rect 13019 1960 13045 1986
rect 13060 1981 13090 1992
rect 13122 1988 13184 2004
rect 13122 1986 13168 1988
rect 13122 1970 13184 1986
rect 13196 1970 13202 2018
rect 13205 2010 13285 2018
rect 13205 2008 13224 2010
rect 13239 2008 13273 2010
rect 13205 1992 13285 2008
rect 13205 1970 13224 1992
rect 13239 1976 13269 1992
rect 13297 1986 13303 2060
rect 13306 1986 13325 2130
rect 13340 1986 13346 2130
rect 13355 2060 13368 2130
rect 13420 2126 13442 2130
rect 13413 2104 13442 2118
rect 13495 2104 13511 2118
rect 13549 2114 13555 2116
rect 13562 2114 13670 2130
rect 13677 2114 13683 2116
rect 13691 2114 13706 2130
rect 13772 2124 13791 2127
rect 13413 2102 13511 2104
rect 13538 2102 13706 2114
rect 13721 2104 13737 2118
rect 13772 2105 13794 2124
rect 13804 2118 13820 2119
rect 13803 2116 13820 2118
rect 13804 2111 13820 2116
rect 13794 2104 13800 2105
rect 13803 2104 13832 2111
rect 13721 2103 13832 2104
rect 13721 2102 13838 2103
rect 13397 2094 13448 2102
rect 13495 2094 13529 2102
rect 13397 2082 13422 2094
rect 13429 2082 13448 2094
rect 13502 2092 13529 2094
rect 13538 2092 13759 2102
rect 13794 2099 13800 2102
rect 13502 2088 13759 2092
rect 13397 2074 13448 2082
rect 13495 2074 13759 2088
rect 13803 2094 13838 2102
rect 13349 2026 13368 2060
rect 13413 2066 13442 2074
rect 13413 2060 13430 2066
rect 13413 2058 13447 2060
rect 13495 2058 13511 2074
rect 13512 2064 13720 2074
rect 13721 2064 13737 2074
rect 13785 2070 13800 2085
rect 13803 2082 13804 2094
rect 13811 2082 13838 2094
rect 13803 2074 13838 2082
rect 13803 2073 13832 2074
rect 13523 2060 13737 2064
rect 13538 2058 13737 2060
rect 13772 2060 13785 2070
rect 13803 2060 13820 2073
rect 13772 2058 13820 2060
rect 13414 2054 13447 2058
rect 13410 2052 13447 2054
rect 13410 2051 13477 2052
rect 13410 2046 13441 2051
rect 13447 2046 13477 2051
rect 13410 2042 13477 2046
rect 13383 2039 13477 2042
rect 13383 2032 13432 2039
rect 13383 2026 13413 2032
rect 13432 2027 13437 2032
rect 13349 2010 13429 2026
rect 13441 2018 13477 2039
rect 13538 2034 13727 2058
rect 13772 2057 13819 2058
rect 13785 2052 13819 2057
rect 13553 2031 13727 2034
rect 13546 2028 13727 2031
rect 13755 2051 13819 2052
rect 13349 2008 13368 2010
rect 13383 2008 13417 2010
rect 13349 1992 13429 2008
rect 13349 1986 13368 1992
rect 13065 1960 13168 1970
rect 13019 1958 13168 1960
rect 13189 1958 13224 1970
rect 12858 1956 13020 1958
rect 12870 1936 12889 1956
rect 12904 1954 12934 1956
rect 12753 1928 12794 1936
rect 12876 1932 12889 1936
rect 12941 1940 13020 1956
rect 13052 1956 13224 1958
rect 13052 1940 13131 1956
rect 13138 1954 13168 1956
rect 12716 1918 12745 1928
rect 12759 1918 12788 1928
rect 12803 1918 12833 1932
rect 12876 1918 12919 1932
rect 12941 1928 13131 1940
rect 13196 1936 13202 1956
rect 12926 1918 12956 1928
rect 12957 1918 13115 1928
rect 13119 1918 13149 1928
rect 13153 1918 13183 1932
rect 13211 1918 13224 1956
rect 13296 1970 13325 1986
rect 13339 1970 13368 1986
rect 13383 1976 13413 1992
rect 13441 1970 13447 2018
rect 13450 2012 13469 2018
rect 13484 2012 13514 2020
rect 13450 2004 13514 2012
rect 13450 1988 13530 2004
rect 13546 1997 13608 2028
rect 13624 1997 13686 2028
rect 13755 2026 13804 2051
rect 13819 2026 13849 2042
rect 13718 2012 13748 2020
rect 13755 2018 13865 2026
rect 13718 2004 13763 2012
rect 13450 1986 13469 1988
rect 13484 1986 13530 1988
rect 13450 1970 13530 1986
rect 13557 1984 13592 1997
rect 13633 1994 13670 1997
rect 13633 1992 13675 1994
rect 13562 1981 13592 1984
rect 13571 1977 13578 1981
rect 13578 1976 13579 1977
rect 13537 1970 13547 1976
rect 13296 1962 13331 1970
rect 13296 1936 13297 1962
rect 13304 1936 13331 1962
rect 13239 1918 13269 1932
rect 13296 1928 13331 1936
rect 13333 1962 13374 1970
rect 13333 1936 13348 1962
rect 13355 1936 13374 1962
rect 13438 1958 13469 1970
rect 13484 1958 13587 1970
rect 13599 1960 13625 1986
rect 13640 1981 13670 1992
rect 13702 1988 13764 2004
rect 13702 1986 13748 1988
rect 13702 1970 13764 1986
rect 13776 1970 13782 2018
rect 13785 2010 13865 2018
rect 13785 2008 13804 2010
rect 13819 2008 13853 2010
rect 13785 1992 13865 2008
rect 13785 1970 13804 1992
rect 13819 1976 13849 1992
rect 13877 1986 13883 2060
rect 13886 1986 13905 2130
rect 13920 1986 13926 2130
rect 13935 2060 13948 2130
rect 14000 2126 14022 2130
rect 13993 2104 14022 2118
rect 14075 2104 14091 2118
rect 14129 2114 14135 2116
rect 14142 2114 14250 2130
rect 14257 2114 14263 2116
rect 14271 2114 14286 2130
rect 14352 2124 14371 2127
rect 13993 2102 14091 2104
rect 14118 2102 14286 2114
rect 14301 2104 14317 2118
rect 14352 2105 14374 2124
rect 14384 2118 14400 2119
rect 14383 2116 14400 2118
rect 14384 2111 14400 2116
rect 14374 2104 14380 2105
rect 14383 2104 14412 2111
rect 14301 2103 14412 2104
rect 14301 2102 14418 2103
rect 13977 2094 14028 2102
rect 14075 2094 14109 2102
rect 13977 2082 14002 2094
rect 14009 2082 14028 2094
rect 14082 2092 14109 2094
rect 14118 2092 14339 2102
rect 14374 2099 14380 2102
rect 14082 2088 14339 2092
rect 13977 2074 14028 2082
rect 14075 2074 14339 2088
rect 14383 2094 14418 2102
rect 13929 2026 13948 2060
rect 13993 2066 14022 2074
rect 13993 2060 14010 2066
rect 13993 2058 14027 2060
rect 14075 2058 14091 2074
rect 14092 2064 14300 2074
rect 14301 2064 14317 2074
rect 14365 2070 14380 2085
rect 14383 2082 14384 2094
rect 14391 2082 14418 2094
rect 14383 2074 14418 2082
rect 14383 2073 14412 2074
rect 14103 2060 14317 2064
rect 14118 2058 14317 2060
rect 14352 2060 14365 2070
rect 14383 2060 14400 2073
rect 14352 2058 14400 2060
rect 13994 2054 14027 2058
rect 13990 2052 14027 2054
rect 13990 2051 14057 2052
rect 13990 2046 14021 2051
rect 14027 2046 14057 2051
rect 13990 2042 14057 2046
rect 13963 2039 14057 2042
rect 13963 2032 14012 2039
rect 13963 2026 13993 2032
rect 14012 2027 14017 2032
rect 13929 2010 14009 2026
rect 14021 2018 14057 2039
rect 14118 2034 14307 2058
rect 14352 2057 14399 2058
rect 14365 2052 14399 2057
rect 14133 2031 14307 2034
rect 14126 2028 14307 2031
rect 14335 2051 14399 2052
rect 13929 2008 13948 2010
rect 13963 2008 13997 2010
rect 13929 1992 14009 2008
rect 13929 1986 13948 1992
rect 13645 1960 13748 1970
rect 13599 1958 13748 1960
rect 13769 1958 13804 1970
rect 13438 1956 13600 1958
rect 13450 1936 13469 1956
rect 13484 1954 13514 1956
rect 13333 1928 13374 1936
rect 13456 1932 13469 1936
rect 13521 1940 13600 1956
rect 13632 1956 13804 1958
rect 13632 1940 13711 1956
rect 13718 1954 13748 1956
rect 13296 1918 13325 1928
rect 13339 1918 13368 1928
rect 13383 1918 13413 1932
rect 13456 1918 13499 1932
rect 13521 1928 13711 1940
rect 13776 1936 13782 1956
rect 13506 1918 13536 1928
rect 13537 1918 13695 1928
rect 13699 1918 13729 1928
rect 13733 1918 13763 1932
rect 13791 1918 13804 1956
rect 13876 1970 13905 1986
rect 13919 1970 13948 1986
rect 13963 1976 13993 1992
rect 14021 1970 14027 2018
rect 14030 2012 14049 2018
rect 14064 2012 14094 2020
rect 14030 2004 14094 2012
rect 14030 1988 14110 2004
rect 14126 1997 14188 2028
rect 14204 1997 14266 2028
rect 14335 2026 14384 2051
rect 14399 2026 14429 2042
rect 14298 2012 14328 2020
rect 14335 2018 14445 2026
rect 14298 2004 14343 2012
rect 14030 1986 14049 1988
rect 14064 1986 14110 1988
rect 14030 1970 14110 1986
rect 14137 1984 14172 1997
rect 14213 1994 14250 1997
rect 14213 1992 14255 1994
rect 14142 1981 14172 1984
rect 14151 1977 14158 1981
rect 14158 1976 14159 1977
rect 14117 1970 14127 1976
rect 13876 1962 13911 1970
rect 13876 1936 13877 1962
rect 13884 1936 13911 1962
rect 13819 1918 13849 1932
rect 13876 1928 13911 1936
rect 13913 1962 13954 1970
rect 13913 1936 13928 1962
rect 13935 1936 13954 1962
rect 14018 1958 14049 1970
rect 14064 1958 14167 1970
rect 14179 1960 14205 1986
rect 14220 1981 14250 1992
rect 14282 1988 14344 2004
rect 14282 1986 14328 1988
rect 14282 1970 14344 1986
rect 14356 1970 14362 2018
rect 14365 2010 14445 2018
rect 14365 2008 14384 2010
rect 14399 2008 14433 2010
rect 14365 1992 14445 2008
rect 14365 1970 14384 1992
rect 14399 1976 14429 1992
rect 14457 1986 14463 2060
rect 14466 1986 14485 2130
rect 14500 1986 14506 2130
rect 14515 2060 14528 2130
rect 14580 2126 14602 2130
rect 14573 2104 14602 2118
rect 14655 2104 14671 2118
rect 14709 2114 14715 2116
rect 14722 2114 14830 2130
rect 14837 2114 14843 2116
rect 14851 2114 14866 2130
rect 14932 2124 14951 2127
rect 14573 2102 14671 2104
rect 14698 2102 14866 2114
rect 14881 2104 14897 2118
rect 14932 2105 14954 2124
rect 14964 2118 14980 2119
rect 14963 2116 14980 2118
rect 14964 2111 14980 2116
rect 14954 2104 14960 2105
rect 14963 2104 14992 2111
rect 14881 2103 14992 2104
rect 14881 2102 14998 2103
rect 14557 2094 14608 2102
rect 14655 2094 14689 2102
rect 14557 2082 14582 2094
rect 14589 2082 14608 2094
rect 14662 2092 14689 2094
rect 14698 2092 14919 2102
rect 14954 2099 14960 2102
rect 14662 2088 14919 2092
rect 14557 2074 14608 2082
rect 14655 2074 14919 2088
rect 14963 2094 14998 2102
rect 14509 2026 14528 2060
rect 14573 2066 14602 2074
rect 14573 2060 14590 2066
rect 14573 2058 14607 2060
rect 14655 2058 14671 2074
rect 14672 2064 14880 2074
rect 14881 2064 14897 2074
rect 14945 2070 14960 2085
rect 14963 2082 14964 2094
rect 14971 2082 14998 2094
rect 14963 2074 14998 2082
rect 14963 2073 14992 2074
rect 14683 2060 14897 2064
rect 14698 2058 14897 2060
rect 14932 2060 14945 2070
rect 14963 2060 14980 2073
rect 14932 2058 14980 2060
rect 14574 2054 14607 2058
rect 14570 2052 14607 2054
rect 14570 2051 14637 2052
rect 14570 2046 14601 2051
rect 14607 2046 14637 2051
rect 14570 2042 14637 2046
rect 14543 2039 14637 2042
rect 14543 2032 14592 2039
rect 14543 2026 14573 2032
rect 14592 2027 14597 2032
rect 14509 2010 14589 2026
rect 14601 2018 14637 2039
rect 14698 2034 14887 2058
rect 14932 2057 14979 2058
rect 14945 2052 14979 2057
rect 14713 2031 14887 2034
rect 14706 2028 14887 2031
rect 14915 2051 14979 2052
rect 14509 2008 14528 2010
rect 14543 2008 14577 2010
rect 14509 1992 14589 2008
rect 14509 1986 14528 1992
rect 14225 1960 14328 1970
rect 14179 1958 14328 1960
rect 14349 1958 14384 1970
rect 14018 1956 14180 1958
rect 14030 1936 14049 1956
rect 14064 1954 14094 1956
rect 13913 1928 13954 1936
rect 14036 1932 14049 1936
rect 14101 1940 14180 1956
rect 14212 1956 14384 1958
rect 14212 1940 14291 1956
rect 14298 1954 14328 1956
rect 13876 1918 13905 1928
rect 13919 1918 13948 1928
rect 13963 1918 13993 1932
rect 14036 1918 14079 1932
rect 14101 1928 14291 1940
rect 14356 1936 14362 1956
rect 14086 1918 14116 1928
rect 14117 1918 14275 1928
rect 14279 1918 14309 1928
rect 14313 1918 14343 1932
rect 14371 1918 14384 1956
rect 14456 1970 14485 1986
rect 14499 1970 14528 1986
rect 14543 1976 14573 1992
rect 14601 1970 14607 2018
rect 14610 2012 14629 2018
rect 14644 2012 14674 2020
rect 14610 2004 14674 2012
rect 14610 1988 14690 2004
rect 14706 1997 14768 2028
rect 14784 1997 14846 2028
rect 14915 2026 14964 2051
rect 14979 2026 15009 2042
rect 14878 2012 14908 2020
rect 14915 2018 15025 2026
rect 14878 2004 14923 2012
rect 14610 1986 14629 1988
rect 14644 1986 14690 1988
rect 14610 1970 14690 1986
rect 14717 1984 14752 1997
rect 14793 1994 14830 1997
rect 14793 1992 14835 1994
rect 14722 1981 14752 1984
rect 14731 1977 14738 1981
rect 14738 1976 14739 1977
rect 14697 1970 14707 1976
rect 14456 1962 14491 1970
rect 14456 1936 14457 1962
rect 14464 1936 14491 1962
rect 14399 1918 14429 1932
rect 14456 1928 14491 1936
rect 14493 1962 14534 1970
rect 14493 1936 14508 1962
rect 14515 1936 14534 1962
rect 14598 1958 14629 1970
rect 14644 1958 14747 1970
rect 14759 1960 14785 1986
rect 14800 1981 14830 1992
rect 14862 1988 14924 2004
rect 14862 1986 14908 1988
rect 14862 1970 14924 1986
rect 14936 1970 14942 2018
rect 14945 2010 15025 2018
rect 14945 2008 14964 2010
rect 14979 2008 15013 2010
rect 14945 1992 15025 2008
rect 14945 1970 14964 1992
rect 14979 1976 15009 1992
rect 15037 1986 15043 2060
rect 15046 1986 15065 2130
rect 15080 1986 15086 2130
rect 15095 2060 15108 2130
rect 15160 2126 15182 2130
rect 15153 2104 15182 2118
rect 15235 2104 15251 2118
rect 15289 2114 15295 2116
rect 15302 2114 15410 2130
rect 15417 2114 15423 2116
rect 15431 2114 15446 2130
rect 15512 2124 15531 2127
rect 15153 2102 15251 2104
rect 15278 2102 15446 2114
rect 15461 2104 15477 2118
rect 15512 2105 15534 2124
rect 15544 2118 15560 2119
rect 15543 2116 15560 2118
rect 15544 2111 15560 2116
rect 15534 2104 15540 2105
rect 15543 2104 15572 2111
rect 15461 2103 15572 2104
rect 15461 2102 15578 2103
rect 15137 2094 15188 2102
rect 15235 2094 15269 2102
rect 15137 2082 15162 2094
rect 15169 2082 15188 2094
rect 15242 2092 15269 2094
rect 15278 2092 15499 2102
rect 15534 2099 15540 2102
rect 15242 2088 15499 2092
rect 15137 2074 15188 2082
rect 15235 2074 15499 2088
rect 15543 2094 15578 2102
rect 15089 2026 15108 2060
rect 15153 2066 15182 2074
rect 15153 2060 15170 2066
rect 15153 2058 15187 2060
rect 15235 2058 15251 2074
rect 15252 2064 15460 2074
rect 15461 2064 15477 2074
rect 15525 2070 15540 2085
rect 15543 2082 15544 2094
rect 15551 2082 15578 2094
rect 15543 2074 15578 2082
rect 15543 2073 15572 2074
rect 15263 2060 15477 2064
rect 15278 2058 15477 2060
rect 15512 2060 15525 2070
rect 15543 2060 15560 2073
rect 15512 2058 15560 2060
rect 15154 2054 15187 2058
rect 15150 2052 15187 2054
rect 15150 2051 15217 2052
rect 15150 2046 15181 2051
rect 15187 2046 15217 2051
rect 15150 2042 15217 2046
rect 15123 2039 15217 2042
rect 15123 2032 15172 2039
rect 15123 2026 15153 2032
rect 15172 2027 15177 2032
rect 15089 2010 15169 2026
rect 15181 2018 15217 2039
rect 15278 2034 15467 2058
rect 15512 2057 15559 2058
rect 15525 2052 15559 2057
rect 15293 2031 15467 2034
rect 15286 2028 15467 2031
rect 15495 2051 15559 2052
rect 15089 2008 15108 2010
rect 15123 2008 15157 2010
rect 15089 1992 15169 2008
rect 15089 1986 15108 1992
rect 14805 1960 14908 1970
rect 14759 1958 14908 1960
rect 14929 1958 14964 1970
rect 14598 1956 14760 1958
rect 14610 1936 14629 1956
rect 14644 1954 14674 1956
rect 14493 1928 14534 1936
rect 14616 1932 14629 1936
rect 14681 1940 14760 1956
rect 14792 1956 14964 1958
rect 14792 1940 14871 1956
rect 14878 1954 14908 1956
rect 14456 1918 14485 1928
rect 14499 1918 14528 1928
rect 14543 1918 14573 1932
rect 14616 1918 14659 1932
rect 14681 1928 14871 1940
rect 14936 1936 14942 1956
rect 14666 1918 14696 1928
rect 14697 1918 14855 1928
rect 14859 1918 14889 1928
rect 14893 1918 14923 1932
rect 14951 1918 14964 1956
rect 15036 1970 15065 1986
rect 15079 1970 15108 1986
rect 15123 1976 15153 1992
rect 15181 1970 15187 2018
rect 15190 2012 15209 2018
rect 15224 2012 15254 2020
rect 15190 2004 15254 2012
rect 15190 1988 15270 2004
rect 15286 1997 15348 2028
rect 15364 1997 15426 2028
rect 15495 2026 15544 2051
rect 15559 2026 15589 2042
rect 15458 2012 15488 2020
rect 15495 2018 15605 2026
rect 15458 2004 15503 2012
rect 15190 1986 15209 1988
rect 15224 1986 15270 1988
rect 15190 1970 15270 1986
rect 15297 1984 15332 1997
rect 15373 1994 15410 1997
rect 15373 1992 15415 1994
rect 15302 1981 15332 1984
rect 15311 1977 15318 1981
rect 15318 1976 15319 1977
rect 15277 1970 15287 1976
rect 15036 1962 15071 1970
rect 15036 1936 15037 1962
rect 15044 1936 15071 1962
rect 14979 1918 15009 1932
rect 15036 1928 15071 1936
rect 15073 1962 15114 1970
rect 15073 1936 15088 1962
rect 15095 1936 15114 1962
rect 15178 1958 15209 1970
rect 15224 1958 15327 1970
rect 15339 1960 15365 1986
rect 15380 1981 15410 1992
rect 15442 1988 15504 2004
rect 15442 1986 15488 1988
rect 15442 1970 15504 1986
rect 15516 1970 15522 2018
rect 15525 2010 15605 2018
rect 15525 2008 15544 2010
rect 15559 2008 15593 2010
rect 15525 1992 15605 2008
rect 15525 1970 15544 1992
rect 15559 1976 15589 1992
rect 15617 1986 15623 2060
rect 15626 1986 15645 2130
rect 15660 1986 15666 2130
rect 15675 2060 15688 2130
rect 15740 2126 15762 2130
rect 15733 2104 15762 2118
rect 15815 2104 15831 2118
rect 15869 2114 15875 2116
rect 15882 2114 15990 2130
rect 15997 2114 16003 2116
rect 16011 2114 16026 2130
rect 16092 2124 16111 2127
rect 15733 2102 15831 2104
rect 15858 2102 16026 2114
rect 16041 2104 16057 2118
rect 16092 2105 16114 2124
rect 16124 2118 16140 2119
rect 16123 2116 16140 2118
rect 16124 2111 16140 2116
rect 16114 2104 16120 2105
rect 16123 2104 16152 2111
rect 16041 2103 16152 2104
rect 16041 2102 16158 2103
rect 15717 2094 15768 2102
rect 15815 2094 15849 2102
rect 15717 2082 15742 2094
rect 15749 2082 15768 2094
rect 15822 2092 15849 2094
rect 15858 2092 16079 2102
rect 16114 2099 16120 2102
rect 15822 2088 16079 2092
rect 15717 2074 15768 2082
rect 15815 2074 16079 2088
rect 16123 2094 16158 2102
rect 15669 2026 15688 2060
rect 15733 2066 15762 2074
rect 15733 2060 15750 2066
rect 15733 2058 15767 2060
rect 15815 2058 15831 2074
rect 15832 2064 16040 2074
rect 16041 2064 16057 2074
rect 16105 2070 16120 2085
rect 16123 2082 16124 2094
rect 16131 2082 16158 2094
rect 16123 2074 16158 2082
rect 16123 2073 16152 2074
rect 15843 2060 16057 2064
rect 15858 2058 16057 2060
rect 16092 2060 16105 2070
rect 16123 2060 16140 2073
rect 16092 2058 16140 2060
rect 15734 2054 15767 2058
rect 15730 2052 15767 2054
rect 15730 2051 15797 2052
rect 15730 2046 15761 2051
rect 15767 2046 15797 2051
rect 15730 2042 15797 2046
rect 15703 2039 15797 2042
rect 15703 2032 15752 2039
rect 15703 2026 15733 2032
rect 15752 2027 15757 2032
rect 15669 2010 15749 2026
rect 15761 2018 15797 2039
rect 15858 2034 16047 2058
rect 16092 2057 16139 2058
rect 16105 2052 16139 2057
rect 15873 2031 16047 2034
rect 15866 2028 16047 2031
rect 16075 2051 16139 2052
rect 15669 2008 15688 2010
rect 15703 2008 15737 2010
rect 15669 1992 15749 2008
rect 15669 1986 15688 1992
rect 15385 1960 15488 1970
rect 15339 1958 15488 1960
rect 15509 1958 15544 1970
rect 15178 1956 15340 1958
rect 15190 1936 15209 1956
rect 15224 1954 15254 1956
rect 15073 1928 15114 1936
rect 15196 1932 15209 1936
rect 15261 1940 15340 1956
rect 15372 1956 15544 1958
rect 15372 1940 15451 1956
rect 15458 1954 15488 1956
rect 15036 1918 15065 1928
rect 15079 1918 15108 1928
rect 15123 1918 15153 1932
rect 15196 1918 15239 1932
rect 15261 1928 15451 1940
rect 15516 1936 15522 1956
rect 15246 1918 15276 1928
rect 15277 1918 15435 1928
rect 15439 1918 15469 1928
rect 15473 1918 15503 1932
rect 15531 1918 15544 1956
rect 15616 1970 15645 1986
rect 15659 1970 15688 1986
rect 15703 1976 15733 1992
rect 15761 1970 15767 2018
rect 15770 2012 15789 2018
rect 15804 2012 15834 2020
rect 15770 2004 15834 2012
rect 15770 1988 15850 2004
rect 15866 1997 15928 2028
rect 15944 1997 16006 2028
rect 16075 2026 16124 2051
rect 16139 2026 16169 2042
rect 16038 2012 16068 2020
rect 16075 2018 16185 2026
rect 16038 2004 16083 2012
rect 15770 1986 15789 1988
rect 15804 1986 15850 1988
rect 15770 1970 15850 1986
rect 15877 1984 15912 1997
rect 15953 1994 15990 1997
rect 15953 1992 15995 1994
rect 15882 1981 15912 1984
rect 15891 1977 15898 1981
rect 15898 1976 15899 1977
rect 15857 1970 15867 1976
rect 15616 1962 15651 1970
rect 15616 1936 15617 1962
rect 15624 1936 15651 1962
rect 15559 1918 15589 1932
rect 15616 1928 15651 1936
rect 15653 1962 15694 1970
rect 15653 1936 15668 1962
rect 15675 1936 15694 1962
rect 15758 1958 15789 1970
rect 15804 1958 15907 1970
rect 15919 1960 15945 1986
rect 15960 1981 15990 1992
rect 16022 1988 16084 2004
rect 16022 1986 16068 1988
rect 16022 1970 16084 1986
rect 16096 1970 16102 2018
rect 16105 2010 16185 2018
rect 16105 2008 16124 2010
rect 16139 2008 16173 2010
rect 16105 1992 16185 2008
rect 16105 1970 16124 1992
rect 16139 1976 16169 1992
rect 16197 1986 16203 2060
rect 16206 1986 16225 2130
rect 16240 1986 16246 2130
rect 16255 2060 16268 2130
rect 16320 2126 16342 2130
rect 16313 2104 16342 2118
rect 16395 2104 16411 2118
rect 16449 2114 16455 2116
rect 16462 2114 16570 2130
rect 16577 2114 16583 2116
rect 16591 2114 16606 2130
rect 16672 2124 16691 2127
rect 16313 2102 16411 2104
rect 16438 2102 16606 2114
rect 16621 2104 16637 2118
rect 16672 2105 16694 2124
rect 16704 2118 16720 2119
rect 16703 2116 16720 2118
rect 16704 2111 16720 2116
rect 16694 2104 16700 2105
rect 16703 2104 16732 2111
rect 16621 2103 16732 2104
rect 16621 2102 16738 2103
rect 16297 2094 16348 2102
rect 16395 2094 16429 2102
rect 16297 2082 16322 2094
rect 16329 2082 16348 2094
rect 16402 2092 16429 2094
rect 16438 2092 16659 2102
rect 16694 2099 16700 2102
rect 16402 2088 16659 2092
rect 16297 2074 16348 2082
rect 16395 2074 16659 2088
rect 16703 2094 16738 2102
rect 16249 2026 16268 2060
rect 16313 2066 16342 2074
rect 16313 2060 16330 2066
rect 16313 2058 16347 2060
rect 16395 2058 16411 2074
rect 16412 2064 16620 2074
rect 16621 2064 16637 2074
rect 16685 2070 16700 2085
rect 16703 2082 16704 2094
rect 16711 2082 16738 2094
rect 16703 2074 16738 2082
rect 16703 2073 16732 2074
rect 16423 2060 16637 2064
rect 16438 2058 16637 2060
rect 16672 2060 16685 2070
rect 16703 2060 16720 2073
rect 16672 2058 16720 2060
rect 16314 2054 16347 2058
rect 16310 2052 16347 2054
rect 16310 2051 16377 2052
rect 16310 2046 16341 2051
rect 16347 2046 16377 2051
rect 16310 2042 16377 2046
rect 16283 2039 16377 2042
rect 16283 2032 16332 2039
rect 16283 2026 16313 2032
rect 16332 2027 16337 2032
rect 16249 2010 16329 2026
rect 16341 2018 16377 2039
rect 16438 2034 16627 2058
rect 16672 2057 16719 2058
rect 16685 2052 16719 2057
rect 16453 2031 16627 2034
rect 16446 2028 16627 2031
rect 16655 2051 16719 2052
rect 16249 2008 16268 2010
rect 16283 2008 16317 2010
rect 16249 1992 16329 2008
rect 16249 1986 16268 1992
rect 15965 1960 16068 1970
rect 15919 1958 16068 1960
rect 16089 1958 16124 1970
rect 15758 1956 15920 1958
rect 15770 1936 15789 1956
rect 15804 1954 15834 1956
rect 15653 1928 15694 1936
rect 15776 1932 15789 1936
rect 15841 1940 15920 1956
rect 15952 1956 16124 1958
rect 15952 1940 16031 1956
rect 16038 1954 16068 1956
rect 15616 1918 15645 1928
rect 15659 1918 15688 1928
rect 15703 1918 15733 1932
rect 15776 1918 15819 1932
rect 15841 1928 16031 1940
rect 16096 1936 16102 1956
rect 15826 1918 15856 1928
rect 15857 1918 16015 1928
rect 16019 1918 16049 1928
rect 16053 1918 16083 1932
rect 16111 1918 16124 1956
rect 16196 1970 16225 1986
rect 16239 1970 16268 1986
rect 16283 1976 16313 1992
rect 16341 1970 16347 2018
rect 16350 2012 16369 2018
rect 16384 2012 16414 2020
rect 16350 2004 16414 2012
rect 16350 1988 16430 2004
rect 16446 1997 16508 2028
rect 16524 1997 16586 2028
rect 16655 2026 16704 2051
rect 16719 2026 16749 2042
rect 16618 2012 16648 2020
rect 16655 2018 16765 2026
rect 16618 2004 16663 2012
rect 16350 1986 16369 1988
rect 16384 1986 16430 1988
rect 16350 1970 16430 1986
rect 16457 1984 16492 1997
rect 16533 1994 16570 1997
rect 16533 1992 16575 1994
rect 16462 1981 16492 1984
rect 16471 1977 16478 1981
rect 16478 1976 16479 1977
rect 16437 1970 16447 1976
rect 16196 1962 16231 1970
rect 16196 1936 16197 1962
rect 16204 1936 16231 1962
rect 16139 1918 16169 1932
rect 16196 1928 16231 1936
rect 16233 1962 16274 1970
rect 16233 1936 16248 1962
rect 16255 1936 16274 1962
rect 16338 1958 16369 1970
rect 16384 1958 16487 1970
rect 16499 1960 16525 1986
rect 16540 1981 16570 1992
rect 16602 1988 16664 2004
rect 16602 1986 16648 1988
rect 16602 1970 16664 1986
rect 16676 1970 16682 2018
rect 16685 2010 16765 2018
rect 16685 2008 16704 2010
rect 16719 2008 16753 2010
rect 16685 1992 16765 2008
rect 16685 1970 16704 1992
rect 16719 1976 16749 1992
rect 16777 1986 16783 2060
rect 16786 1986 16805 2130
rect 16820 1986 16826 2130
rect 16835 2060 16848 2130
rect 16900 2126 16922 2130
rect 16893 2104 16922 2118
rect 16975 2104 16991 2118
rect 17029 2114 17035 2116
rect 17042 2114 17150 2130
rect 17157 2114 17163 2116
rect 17171 2114 17186 2130
rect 17252 2124 17271 2127
rect 16893 2102 16991 2104
rect 17018 2102 17186 2114
rect 17201 2104 17217 2118
rect 17252 2105 17274 2124
rect 17284 2118 17300 2119
rect 17283 2116 17300 2118
rect 17284 2111 17300 2116
rect 17274 2104 17280 2105
rect 17283 2104 17312 2111
rect 17201 2103 17312 2104
rect 17201 2102 17318 2103
rect 16877 2094 16928 2102
rect 16975 2094 17009 2102
rect 16877 2082 16902 2094
rect 16909 2082 16928 2094
rect 16982 2092 17009 2094
rect 17018 2092 17239 2102
rect 17274 2099 17280 2102
rect 16982 2088 17239 2092
rect 16877 2074 16928 2082
rect 16975 2074 17239 2088
rect 17283 2094 17318 2102
rect 16829 2026 16848 2060
rect 16893 2066 16922 2074
rect 16893 2060 16910 2066
rect 16893 2058 16927 2060
rect 16975 2058 16991 2074
rect 16992 2064 17200 2074
rect 17201 2064 17217 2074
rect 17265 2070 17280 2085
rect 17283 2082 17284 2094
rect 17291 2082 17318 2094
rect 17283 2074 17318 2082
rect 17283 2073 17312 2074
rect 17003 2060 17217 2064
rect 17018 2058 17217 2060
rect 17252 2060 17265 2070
rect 17283 2060 17300 2073
rect 17252 2058 17300 2060
rect 16894 2054 16927 2058
rect 16890 2052 16927 2054
rect 16890 2051 16957 2052
rect 16890 2046 16921 2051
rect 16927 2046 16957 2051
rect 16890 2042 16957 2046
rect 16863 2039 16957 2042
rect 16863 2032 16912 2039
rect 16863 2026 16893 2032
rect 16912 2027 16917 2032
rect 16829 2010 16909 2026
rect 16921 2018 16957 2039
rect 17018 2034 17207 2058
rect 17252 2057 17299 2058
rect 17265 2052 17299 2057
rect 17033 2031 17207 2034
rect 17026 2028 17207 2031
rect 17235 2051 17299 2052
rect 16829 2008 16848 2010
rect 16863 2008 16897 2010
rect 16829 1992 16909 2008
rect 16829 1986 16848 1992
rect 16545 1960 16648 1970
rect 16499 1958 16648 1960
rect 16669 1958 16704 1970
rect 16338 1956 16500 1958
rect 16350 1936 16369 1956
rect 16384 1954 16414 1956
rect 16233 1928 16274 1936
rect 16356 1932 16369 1936
rect 16421 1940 16500 1956
rect 16532 1956 16704 1958
rect 16532 1940 16611 1956
rect 16618 1954 16648 1956
rect 16196 1918 16225 1928
rect 16239 1918 16268 1928
rect 16283 1918 16313 1932
rect 16356 1918 16399 1932
rect 16421 1928 16611 1940
rect 16676 1936 16682 1956
rect 16406 1918 16436 1928
rect 16437 1918 16595 1928
rect 16599 1918 16629 1928
rect 16633 1918 16663 1932
rect 16691 1918 16704 1956
rect 16776 1970 16805 1986
rect 16819 1970 16848 1986
rect 16863 1976 16893 1992
rect 16921 1970 16927 2018
rect 16930 2012 16949 2018
rect 16964 2012 16994 2020
rect 16930 2004 16994 2012
rect 16930 1988 17010 2004
rect 17026 1997 17088 2028
rect 17104 1997 17166 2028
rect 17235 2026 17284 2051
rect 17299 2026 17329 2042
rect 17198 2012 17228 2020
rect 17235 2018 17345 2026
rect 17198 2004 17243 2012
rect 16930 1986 16949 1988
rect 16964 1986 17010 1988
rect 16930 1970 17010 1986
rect 17037 1984 17072 1997
rect 17113 1994 17150 1997
rect 17113 1992 17155 1994
rect 17042 1981 17072 1984
rect 17051 1977 17058 1981
rect 17058 1976 17059 1977
rect 17017 1970 17027 1976
rect 16776 1962 16811 1970
rect 16776 1936 16777 1962
rect 16784 1936 16811 1962
rect 16719 1918 16749 1932
rect 16776 1928 16811 1936
rect 16813 1962 16854 1970
rect 16813 1936 16828 1962
rect 16835 1936 16854 1962
rect 16918 1958 16949 1970
rect 16964 1958 17067 1970
rect 17079 1960 17105 1986
rect 17120 1981 17150 1992
rect 17182 1988 17244 2004
rect 17182 1986 17228 1988
rect 17182 1970 17244 1986
rect 17256 1970 17262 2018
rect 17265 2010 17345 2018
rect 17265 2008 17284 2010
rect 17299 2008 17333 2010
rect 17265 1992 17345 2008
rect 17265 1970 17284 1992
rect 17299 1976 17329 1992
rect 17357 1986 17363 2060
rect 17366 1986 17385 2130
rect 17400 1986 17406 2130
rect 17415 2060 17428 2130
rect 17480 2126 17502 2130
rect 17473 2104 17502 2118
rect 17555 2104 17571 2118
rect 17609 2114 17615 2116
rect 17622 2114 17730 2130
rect 17737 2114 17743 2116
rect 17751 2114 17766 2130
rect 17832 2124 17851 2127
rect 17473 2102 17571 2104
rect 17598 2102 17766 2114
rect 17781 2104 17797 2118
rect 17832 2105 17854 2124
rect 17864 2118 17880 2119
rect 17863 2116 17880 2118
rect 17864 2111 17880 2116
rect 17854 2104 17860 2105
rect 17863 2104 17892 2111
rect 17781 2103 17892 2104
rect 17781 2102 17898 2103
rect 17457 2094 17508 2102
rect 17555 2094 17589 2102
rect 17457 2082 17482 2094
rect 17489 2082 17508 2094
rect 17562 2092 17589 2094
rect 17598 2092 17819 2102
rect 17854 2099 17860 2102
rect 17562 2088 17819 2092
rect 17457 2074 17508 2082
rect 17555 2074 17819 2088
rect 17863 2094 17898 2102
rect 17409 2026 17428 2060
rect 17473 2066 17502 2074
rect 17473 2060 17490 2066
rect 17473 2058 17507 2060
rect 17555 2058 17571 2074
rect 17572 2064 17780 2074
rect 17781 2064 17797 2074
rect 17845 2070 17860 2085
rect 17863 2082 17864 2094
rect 17871 2082 17898 2094
rect 17863 2074 17898 2082
rect 17863 2073 17892 2074
rect 17583 2060 17797 2064
rect 17598 2058 17797 2060
rect 17832 2060 17845 2070
rect 17863 2060 17880 2073
rect 17832 2058 17880 2060
rect 17474 2054 17507 2058
rect 17470 2052 17507 2054
rect 17470 2051 17537 2052
rect 17470 2046 17501 2051
rect 17507 2046 17537 2051
rect 17470 2042 17537 2046
rect 17443 2039 17537 2042
rect 17443 2032 17492 2039
rect 17443 2026 17473 2032
rect 17492 2027 17497 2032
rect 17409 2010 17489 2026
rect 17501 2018 17537 2039
rect 17598 2034 17787 2058
rect 17832 2057 17879 2058
rect 17845 2052 17879 2057
rect 17613 2031 17787 2034
rect 17606 2028 17787 2031
rect 17815 2051 17879 2052
rect 17409 2008 17428 2010
rect 17443 2008 17477 2010
rect 17409 1992 17489 2008
rect 17409 1986 17428 1992
rect 17125 1960 17228 1970
rect 17079 1958 17228 1960
rect 17249 1958 17284 1970
rect 16918 1956 17080 1958
rect 16930 1936 16949 1956
rect 16964 1954 16994 1956
rect 16813 1928 16854 1936
rect 16936 1932 16949 1936
rect 17001 1940 17080 1956
rect 17112 1956 17284 1958
rect 17112 1940 17191 1956
rect 17198 1954 17228 1956
rect 16776 1918 16805 1928
rect 16819 1918 16848 1928
rect 16863 1918 16893 1932
rect 16936 1918 16979 1932
rect 17001 1928 17191 1940
rect 17256 1936 17262 1956
rect 16986 1918 17016 1928
rect 17017 1918 17175 1928
rect 17179 1918 17209 1928
rect 17213 1918 17243 1932
rect 17271 1918 17284 1956
rect 17356 1970 17385 1986
rect 17399 1970 17428 1986
rect 17443 1976 17473 1992
rect 17501 1970 17507 2018
rect 17510 2012 17529 2018
rect 17544 2012 17574 2020
rect 17510 2004 17574 2012
rect 17510 1988 17590 2004
rect 17606 1997 17668 2028
rect 17684 1997 17746 2028
rect 17815 2026 17864 2051
rect 17879 2026 17909 2042
rect 17778 2012 17808 2020
rect 17815 2018 17925 2026
rect 17778 2004 17823 2012
rect 17510 1986 17529 1988
rect 17544 1986 17590 1988
rect 17510 1970 17590 1986
rect 17617 1984 17652 1997
rect 17693 1994 17730 1997
rect 17693 1992 17735 1994
rect 17622 1981 17652 1984
rect 17631 1977 17638 1981
rect 17638 1976 17639 1977
rect 17597 1970 17607 1976
rect 17356 1962 17391 1970
rect 17356 1936 17357 1962
rect 17364 1936 17391 1962
rect 17299 1918 17329 1932
rect 17356 1928 17391 1936
rect 17393 1962 17434 1970
rect 17393 1936 17408 1962
rect 17415 1936 17434 1962
rect 17498 1958 17529 1970
rect 17544 1958 17647 1970
rect 17659 1960 17685 1986
rect 17700 1981 17730 1992
rect 17762 1988 17824 2004
rect 17762 1986 17808 1988
rect 17762 1970 17824 1986
rect 17836 1970 17842 2018
rect 17845 2010 17925 2018
rect 17845 2008 17864 2010
rect 17879 2008 17913 2010
rect 17845 1992 17925 2008
rect 17845 1970 17864 1992
rect 17879 1976 17909 1992
rect 17937 1986 17943 2060
rect 17946 1986 17965 2130
rect 17980 1986 17986 2130
rect 17995 2060 18008 2130
rect 18060 2126 18082 2130
rect 18053 2104 18082 2118
rect 18135 2104 18151 2118
rect 18189 2114 18195 2116
rect 18202 2114 18310 2130
rect 18317 2114 18323 2116
rect 18331 2114 18346 2130
rect 18412 2124 18431 2127
rect 18053 2102 18151 2104
rect 18178 2102 18346 2114
rect 18361 2104 18377 2118
rect 18412 2105 18434 2124
rect 18444 2118 18460 2119
rect 18443 2116 18460 2118
rect 18444 2111 18460 2116
rect 18434 2104 18440 2105
rect 18443 2104 18472 2111
rect 18361 2103 18472 2104
rect 18361 2102 18478 2103
rect 18037 2094 18088 2102
rect 18135 2094 18169 2102
rect 18037 2082 18062 2094
rect 18069 2082 18088 2094
rect 18142 2092 18169 2094
rect 18178 2092 18399 2102
rect 18434 2099 18440 2102
rect 18142 2088 18399 2092
rect 18037 2074 18088 2082
rect 18135 2074 18399 2088
rect 18443 2094 18478 2102
rect 17989 2026 18008 2060
rect 18053 2066 18082 2074
rect 18053 2060 18070 2066
rect 18053 2058 18087 2060
rect 18135 2058 18151 2074
rect 18152 2064 18360 2074
rect 18361 2064 18377 2074
rect 18425 2070 18440 2085
rect 18443 2082 18444 2094
rect 18451 2082 18478 2094
rect 18443 2074 18478 2082
rect 18443 2073 18472 2074
rect 18163 2060 18377 2064
rect 18178 2058 18377 2060
rect 18412 2060 18425 2070
rect 18443 2060 18460 2073
rect 18412 2058 18460 2060
rect 18054 2054 18087 2058
rect 18050 2052 18087 2054
rect 18050 2051 18117 2052
rect 18050 2046 18081 2051
rect 18087 2046 18117 2051
rect 18050 2042 18117 2046
rect 18023 2039 18117 2042
rect 18023 2032 18072 2039
rect 18023 2026 18053 2032
rect 18072 2027 18077 2032
rect 17989 2010 18069 2026
rect 18081 2018 18117 2039
rect 18178 2034 18367 2058
rect 18412 2057 18459 2058
rect 18425 2052 18459 2057
rect 18193 2031 18367 2034
rect 18186 2028 18367 2031
rect 18395 2051 18459 2052
rect 17989 2008 18008 2010
rect 18023 2008 18057 2010
rect 17989 1992 18069 2008
rect 17989 1986 18008 1992
rect 17705 1960 17808 1970
rect 17659 1958 17808 1960
rect 17829 1958 17864 1970
rect 17498 1956 17660 1958
rect 17510 1936 17529 1956
rect 17544 1954 17574 1956
rect 17393 1928 17434 1936
rect 17516 1932 17529 1936
rect 17581 1940 17660 1956
rect 17692 1956 17864 1958
rect 17692 1940 17771 1956
rect 17778 1954 17808 1956
rect 17356 1918 17385 1928
rect 17399 1918 17428 1928
rect 17443 1918 17473 1932
rect 17516 1918 17559 1932
rect 17581 1928 17771 1940
rect 17836 1936 17842 1956
rect 17566 1918 17596 1928
rect 17597 1918 17755 1928
rect 17759 1918 17789 1928
rect 17793 1918 17823 1932
rect 17851 1918 17864 1956
rect 17936 1970 17965 1986
rect 17979 1970 18008 1986
rect 18023 1976 18053 1992
rect 18081 1970 18087 2018
rect 18090 2012 18109 2018
rect 18124 2012 18154 2020
rect 18090 2004 18154 2012
rect 18090 1988 18170 2004
rect 18186 1997 18248 2028
rect 18264 1997 18326 2028
rect 18395 2026 18444 2051
rect 18459 2026 18489 2042
rect 18358 2012 18388 2020
rect 18395 2018 18505 2026
rect 18358 2004 18403 2012
rect 18090 1986 18109 1988
rect 18124 1986 18170 1988
rect 18090 1970 18170 1986
rect 18197 1984 18232 1997
rect 18273 1994 18310 1997
rect 18273 1992 18315 1994
rect 18202 1981 18232 1984
rect 18211 1977 18218 1981
rect 18218 1976 18219 1977
rect 18177 1970 18187 1976
rect 17936 1962 17971 1970
rect 17936 1936 17937 1962
rect 17944 1936 17971 1962
rect 17879 1918 17909 1932
rect 17936 1928 17971 1936
rect 17973 1962 18014 1970
rect 17973 1936 17988 1962
rect 17995 1936 18014 1962
rect 18078 1958 18109 1970
rect 18124 1958 18227 1970
rect 18239 1960 18265 1986
rect 18280 1981 18310 1992
rect 18342 1988 18404 2004
rect 18342 1986 18388 1988
rect 18342 1970 18404 1986
rect 18416 1970 18422 2018
rect 18425 2010 18505 2018
rect 18425 2008 18444 2010
rect 18459 2008 18493 2010
rect 18425 1992 18505 2008
rect 18425 1970 18444 1992
rect 18459 1976 18489 1992
rect 18517 1986 18523 2060
rect 18532 1986 18545 2130
rect 18285 1960 18388 1970
rect 18239 1958 18388 1960
rect 18409 1958 18444 1970
rect 18078 1956 18240 1958
rect 18090 1936 18109 1956
rect 18124 1954 18154 1956
rect 17973 1928 18014 1936
rect 18096 1932 18109 1936
rect 18161 1940 18240 1956
rect 18272 1956 18444 1958
rect 18272 1940 18351 1956
rect 18358 1954 18388 1956
rect 17936 1918 17965 1928
rect 17979 1918 18008 1928
rect 18023 1918 18053 1932
rect 18096 1918 18139 1932
rect 18161 1928 18351 1940
rect 18416 1936 18422 1956
rect 18146 1918 18176 1928
rect 18177 1918 18335 1928
rect 18339 1918 18369 1928
rect 18373 1918 18403 1932
rect 18431 1918 18444 1956
rect 18516 1970 18545 1986
rect 18516 1962 18551 1970
rect 18516 1936 18517 1962
rect 18524 1936 18551 1962
rect 18459 1918 18489 1932
rect 18516 1928 18551 1936
rect 18516 1918 18545 1928
rect -1 1912 18545 1918
rect 0 1904 18545 1912
rect 15 1874 28 1904
rect 43 1890 73 1904
rect 116 1890 159 1904
rect 166 1890 386 1904
rect 393 1890 423 1904
rect 83 1876 98 1888
rect 117 1876 130 1890
rect 198 1886 351 1890
rect 80 1874 102 1876
rect 180 1874 372 1886
rect 451 1874 464 1904
rect 479 1890 509 1904
rect 546 1874 565 1904
rect 580 1874 586 1904
rect 595 1874 608 1904
rect 623 1890 653 1904
rect 696 1890 739 1904
rect 746 1890 966 1904
rect 973 1890 1003 1904
rect 663 1876 678 1888
rect 697 1876 710 1890
rect 778 1886 931 1890
rect 660 1874 682 1876
rect 760 1874 952 1886
rect 1031 1874 1044 1904
rect 1059 1890 1089 1904
rect 1126 1874 1145 1904
rect 1160 1874 1166 1904
rect 1175 1874 1188 1904
rect 1203 1890 1233 1904
rect 1276 1890 1319 1904
rect 1326 1890 1546 1904
rect 1553 1890 1583 1904
rect 1243 1876 1258 1888
rect 1277 1876 1290 1890
rect 1358 1886 1511 1890
rect 1240 1874 1262 1876
rect 1340 1874 1532 1886
rect 1611 1874 1624 1904
rect 1639 1890 1669 1904
rect 1706 1874 1725 1904
rect 1740 1874 1746 1904
rect 1755 1874 1768 1904
rect 1783 1890 1813 1904
rect 1856 1890 1899 1904
rect 1906 1890 2126 1904
rect 2133 1890 2163 1904
rect 1823 1876 1838 1888
rect 1857 1876 1870 1890
rect 1938 1886 2091 1890
rect 1820 1874 1842 1876
rect 1920 1874 2112 1886
rect 2191 1874 2204 1904
rect 2219 1890 2249 1904
rect 2286 1874 2305 1904
rect 2320 1874 2326 1904
rect 2335 1874 2348 1904
rect 2363 1890 2393 1904
rect 2436 1890 2479 1904
rect 2486 1890 2706 1904
rect 2713 1890 2743 1904
rect 2403 1876 2418 1888
rect 2437 1876 2450 1890
rect 2518 1886 2671 1890
rect 2400 1874 2422 1876
rect 2500 1874 2692 1886
rect 2771 1874 2784 1904
rect 2799 1890 2829 1904
rect 2866 1874 2885 1904
rect 2900 1874 2906 1904
rect 2915 1874 2928 1904
rect 2943 1890 2973 1904
rect 3016 1890 3059 1904
rect 3066 1890 3286 1904
rect 3293 1890 3323 1904
rect 2983 1876 2998 1888
rect 3017 1876 3030 1890
rect 3098 1886 3251 1890
rect 2980 1874 3002 1876
rect 3080 1874 3272 1886
rect 3351 1874 3364 1904
rect 3379 1890 3409 1904
rect 3446 1874 3465 1904
rect 3480 1874 3486 1904
rect 3495 1874 3508 1904
rect 3523 1890 3553 1904
rect 3596 1890 3639 1904
rect 3646 1890 3866 1904
rect 3873 1890 3903 1904
rect 3563 1876 3578 1888
rect 3597 1876 3610 1890
rect 3678 1886 3831 1890
rect 3560 1874 3582 1876
rect 3660 1874 3852 1886
rect 3931 1874 3944 1904
rect 3959 1890 3989 1904
rect 4026 1874 4045 1904
rect 4060 1874 4066 1904
rect 4075 1874 4088 1904
rect 4103 1890 4133 1904
rect 4176 1890 4219 1904
rect 4226 1890 4446 1904
rect 4453 1890 4483 1904
rect 4143 1876 4158 1888
rect 4177 1876 4190 1890
rect 4258 1886 4411 1890
rect 4140 1874 4162 1876
rect 4240 1874 4432 1886
rect 4511 1874 4524 1904
rect 4539 1890 4569 1904
rect 4606 1874 4625 1904
rect 4640 1874 4646 1904
rect 4655 1874 4668 1904
rect 4683 1890 4713 1904
rect 4756 1890 4799 1904
rect 4806 1890 5026 1904
rect 5033 1890 5063 1904
rect 4723 1876 4738 1888
rect 4757 1876 4770 1890
rect 4838 1886 4991 1890
rect 4720 1874 4742 1876
rect 4820 1874 5012 1886
rect 5091 1874 5104 1904
rect 5119 1890 5149 1904
rect 5186 1874 5205 1904
rect 5220 1874 5226 1904
rect 5235 1874 5248 1904
rect 5263 1890 5293 1904
rect 5336 1890 5379 1904
rect 5386 1890 5606 1904
rect 5613 1890 5643 1904
rect 5303 1876 5318 1888
rect 5337 1876 5350 1890
rect 5418 1886 5571 1890
rect 5300 1874 5322 1876
rect 5400 1874 5592 1886
rect 5671 1874 5684 1904
rect 5699 1890 5729 1904
rect 5766 1874 5785 1904
rect 5800 1874 5806 1904
rect 5815 1874 5828 1904
rect 5843 1890 5873 1904
rect 5916 1890 5959 1904
rect 5966 1890 6186 1904
rect 6193 1890 6223 1904
rect 5883 1876 5898 1888
rect 5917 1876 5930 1890
rect 5998 1886 6151 1890
rect 5880 1874 5902 1876
rect 5980 1874 6172 1886
rect 6251 1874 6264 1904
rect 6279 1890 6309 1904
rect 6346 1874 6365 1904
rect 6380 1874 6386 1904
rect 6395 1874 6408 1904
rect 6423 1890 6453 1904
rect 6496 1890 6539 1904
rect 6546 1890 6766 1904
rect 6773 1890 6803 1904
rect 6463 1876 6478 1888
rect 6497 1876 6510 1890
rect 6578 1886 6731 1890
rect 6460 1874 6482 1876
rect 6560 1874 6752 1886
rect 6831 1874 6844 1904
rect 6859 1890 6889 1904
rect 6926 1874 6945 1904
rect 6960 1874 6966 1904
rect 6975 1874 6988 1904
rect 7003 1890 7033 1904
rect 7076 1890 7119 1904
rect 7126 1890 7346 1904
rect 7353 1890 7383 1904
rect 7043 1876 7058 1888
rect 7077 1876 7090 1890
rect 7158 1886 7311 1890
rect 7040 1874 7062 1876
rect 7140 1874 7332 1886
rect 7411 1874 7424 1904
rect 7439 1890 7469 1904
rect 7506 1874 7525 1904
rect 7540 1874 7546 1904
rect 7555 1874 7568 1904
rect 7583 1890 7613 1904
rect 7656 1890 7699 1904
rect 7706 1890 7926 1904
rect 7933 1890 7963 1904
rect 7623 1876 7638 1888
rect 7657 1876 7670 1890
rect 7738 1886 7891 1890
rect 7620 1874 7642 1876
rect 7720 1874 7912 1886
rect 7991 1874 8004 1904
rect 8019 1890 8049 1904
rect 8086 1874 8105 1904
rect 8120 1874 8126 1904
rect 8135 1874 8148 1904
rect 8163 1890 8193 1904
rect 8236 1890 8279 1904
rect 8286 1890 8506 1904
rect 8513 1890 8543 1904
rect 8203 1876 8218 1888
rect 8237 1876 8250 1890
rect 8318 1886 8471 1890
rect 8200 1874 8222 1876
rect 8300 1874 8492 1886
rect 8571 1874 8584 1904
rect 8599 1890 8629 1904
rect 8666 1874 8685 1904
rect 8700 1874 8706 1904
rect 8715 1874 8728 1904
rect 8743 1890 8773 1904
rect 8816 1890 8859 1904
rect 8866 1890 9086 1904
rect 9093 1890 9123 1904
rect 8783 1876 8798 1888
rect 8817 1876 8830 1890
rect 8898 1886 9051 1890
rect 8780 1874 8802 1876
rect 8880 1874 9072 1886
rect 9151 1874 9164 1904
rect 9179 1890 9209 1904
rect 9246 1874 9265 1904
rect 9280 1874 9286 1904
rect 9295 1874 9308 1904
rect 9323 1890 9353 1904
rect 9396 1890 9439 1904
rect 9446 1890 9666 1904
rect 9673 1890 9703 1904
rect 9363 1876 9378 1888
rect 9397 1876 9410 1890
rect 9478 1886 9631 1890
rect 9360 1874 9382 1876
rect 9460 1874 9652 1886
rect 9731 1874 9744 1904
rect 9759 1890 9789 1904
rect 9826 1874 9845 1904
rect 9860 1874 9866 1904
rect 9875 1874 9888 1904
rect 9903 1890 9933 1904
rect 9976 1890 10019 1904
rect 10026 1890 10246 1904
rect 10253 1890 10283 1904
rect 9943 1876 9958 1888
rect 9977 1876 9990 1890
rect 10058 1886 10211 1890
rect 9940 1874 9962 1876
rect 10040 1874 10232 1886
rect 10311 1874 10324 1904
rect 10339 1890 10369 1904
rect 10406 1874 10425 1904
rect 10440 1874 10446 1904
rect 10455 1874 10468 1904
rect 10483 1890 10513 1904
rect 10556 1890 10599 1904
rect 10606 1890 10826 1904
rect 10833 1890 10863 1904
rect 10523 1876 10538 1888
rect 10557 1876 10570 1890
rect 10638 1886 10791 1890
rect 10520 1874 10542 1876
rect 10620 1874 10812 1886
rect 10891 1874 10904 1904
rect 10919 1890 10949 1904
rect 10986 1874 11005 1904
rect 11020 1874 11026 1904
rect 11035 1874 11048 1904
rect 11063 1890 11093 1904
rect 11136 1890 11179 1904
rect 11186 1890 11406 1904
rect 11413 1890 11443 1904
rect 11103 1876 11118 1888
rect 11137 1876 11150 1890
rect 11218 1886 11371 1890
rect 11100 1874 11122 1876
rect 11200 1874 11392 1886
rect 11471 1874 11484 1904
rect 11499 1890 11529 1904
rect 11566 1874 11585 1904
rect 11600 1874 11606 1904
rect 11615 1874 11628 1904
rect 11643 1890 11673 1904
rect 11716 1890 11759 1904
rect 11766 1890 11986 1904
rect 11993 1890 12023 1904
rect 11683 1876 11698 1888
rect 11717 1876 11730 1890
rect 11798 1886 11951 1890
rect 11680 1874 11702 1876
rect 11780 1874 11972 1886
rect 12051 1874 12064 1904
rect 12079 1890 12109 1904
rect 12146 1874 12165 1904
rect 12180 1874 12186 1904
rect 12195 1874 12208 1904
rect 12223 1890 12253 1904
rect 12296 1890 12339 1904
rect 12346 1890 12566 1904
rect 12573 1890 12603 1904
rect 12263 1876 12278 1888
rect 12297 1876 12310 1890
rect 12378 1886 12531 1890
rect 12260 1874 12282 1876
rect 12360 1874 12552 1886
rect 12631 1874 12644 1904
rect 12659 1890 12689 1904
rect 12726 1874 12745 1904
rect 12760 1874 12766 1904
rect 12775 1874 12788 1904
rect 12803 1890 12833 1904
rect 12876 1890 12919 1904
rect 12926 1890 13146 1904
rect 13153 1890 13183 1904
rect 12843 1876 12858 1888
rect 12877 1876 12890 1890
rect 12958 1886 13111 1890
rect 12840 1874 12862 1876
rect 12940 1874 13132 1886
rect 13211 1874 13224 1904
rect 13239 1890 13269 1904
rect 13306 1874 13325 1904
rect 13340 1874 13346 1904
rect 13355 1874 13368 1904
rect 13383 1890 13413 1904
rect 13456 1890 13499 1904
rect 13506 1890 13726 1904
rect 13733 1890 13763 1904
rect 13423 1876 13438 1888
rect 13457 1876 13470 1890
rect 13538 1886 13691 1890
rect 13420 1874 13442 1876
rect 13520 1874 13712 1886
rect 13791 1874 13804 1904
rect 13819 1890 13849 1904
rect 13886 1874 13905 1904
rect 13920 1874 13926 1904
rect 13935 1874 13948 1904
rect 13963 1890 13993 1904
rect 14036 1890 14079 1904
rect 14086 1890 14306 1904
rect 14313 1890 14343 1904
rect 14003 1876 14018 1888
rect 14037 1876 14050 1890
rect 14118 1886 14271 1890
rect 14000 1874 14022 1876
rect 14100 1874 14292 1886
rect 14371 1874 14384 1904
rect 14399 1890 14429 1904
rect 14466 1874 14485 1904
rect 14500 1874 14506 1904
rect 14515 1874 14528 1904
rect 14543 1890 14573 1904
rect 14616 1890 14659 1904
rect 14666 1890 14886 1904
rect 14893 1890 14923 1904
rect 14583 1876 14598 1888
rect 14617 1876 14630 1890
rect 14698 1886 14851 1890
rect 14580 1874 14602 1876
rect 14680 1874 14872 1886
rect 14951 1874 14964 1904
rect 14979 1890 15009 1904
rect 15046 1874 15065 1904
rect 15080 1874 15086 1904
rect 15095 1874 15108 1904
rect 15123 1890 15153 1904
rect 15196 1890 15239 1904
rect 15246 1890 15466 1904
rect 15473 1890 15503 1904
rect 15163 1876 15178 1888
rect 15197 1876 15210 1890
rect 15278 1886 15431 1890
rect 15160 1874 15182 1876
rect 15260 1874 15452 1886
rect 15531 1874 15544 1904
rect 15559 1890 15589 1904
rect 15626 1874 15645 1904
rect 15660 1874 15666 1904
rect 15675 1874 15688 1904
rect 15703 1890 15733 1904
rect 15776 1890 15819 1904
rect 15826 1890 16046 1904
rect 16053 1890 16083 1904
rect 15743 1876 15758 1888
rect 15777 1876 15790 1890
rect 15858 1886 16011 1890
rect 15740 1874 15762 1876
rect 15840 1874 16032 1886
rect 16111 1874 16124 1904
rect 16139 1890 16169 1904
rect 16206 1874 16225 1904
rect 16240 1874 16246 1904
rect 16255 1874 16268 1904
rect 16283 1890 16313 1904
rect 16356 1890 16399 1904
rect 16406 1890 16626 1904
rect 16633 1890 16663 1904
rect 16323 1876 16338 1888
rect 16357 1876 16370 1890
rect 16438 1886 16591 1890
rect 16320 1874 16342 1876
rect 16420 1874 16612 1886
rect 16691 1874 16704 1904
rect 16719 1890 16749 1904
rect 16786 1874 16805 1904
rect 16820 1874 16826 1904
rect 16835 1874 16848 1904
rect 16863 1890 16893 1904
rect 16936 1890 16979 1904
rect 16986 1890 17206 1904
rect 17213 1890 17243 1904
rect 16903 1876 16918 1888
rect 16937 1876 16950 1890
rect 17018 1886 17171 1890
rect 16900 1874 16922 1876
rect 17000 1874 17192 1886
rect 17271 1874 17284 1904
rect 17299 1890 17329 1904
rect 17366 1874 17385 1904
rect 17400 1874 17406 1904
rect 17415 1874 17428 1904
rect 17443 1890 17473 1904
rect 17516 1890 17559 1904
rect 17566 1890 17786 1904
rect 17793 1890 17823 1904
rect 17483 1876 17498 1888
rect 17517 1876 17530 1890
rect 17598 1886 17751 1890
rect 17480 1874 17502 1876
rect 17580 1874 17772 1886
rect 17851 1874 17864 1904
rect 17879 1890 17909 1904
rect 17946 1874 17965 1904
rect 17980 1874 17986 1904
rect 17995 1874 18008 1904
rect 18023 1890 18053 1904
rect 18096 1890 18139 1904
rect 18146 1890 18366 1904
rect 18373 1890 18403 1904
rect 18063 1876 18078 1888
rect 18097 1876 18110 1890
rect 18178 1886 18331 1890
rect 18060 1874 18082 1876
rect 18160 1874 18352 1886
rect 18431 1874 18444 1904
rect 18459 1890 18489 1904
rect 18532 1874 18545 1904
rect 0 1860 18545 1874
rect 15 1790 28 1860
rect 80 1856 102 1860
rect 73 1834 102 1848
rect 155 1834 171 1848
rect 209 1844 215 1846
rect 222 1844 330 1860
rect 337 1844 343 1846
rect 351 1844 366 1860
rect 432 1854 451 1857
rect 73 1832 171 1834
rect 198 1832 366 1844
rect 381 1834 397 1848
rect 432 1835 454 1854
rect 464 1848 480 1849
rect 463 1846 480 1848
rect 464 1841 480 1846
rect 454 1834 460 1835
rect 463 1834 492 1841
rect 381 1833 492 1834
rect 381 1832 498 1833
rect 57 1824 108 1832
rect 155 1824 189 1832
rect 57 1812 82 1824
rect 89 1812 108 1824
rect 162 1822 189 1824
rect 198 1822 419 1832
rect 454 1829 460 1832
rect 162 1818 419 1822
rect 57 1804 108 1812
rect 155 1804 419 1818
rect 463 1824 498 1832
rect 9 1756 28 1790
rect 73 1796 102 1804
rect 73 1790 90 1796
rect 73 1788 107 1790
rect 155 1788 171 1804
rect 172 1794 380 1804
rect 381 1794 397 1804
rect 445 1800 460 1815
rect 463 1812 464 1824
rect 471 1812 498 1824
rect 463 1804 498 1812
rect 463 1803 492 1804
rect 183 1790 397 1794
rect 198 1788 397 1790
rect 432 1790 445 1800
rect 463 1790 480 1803
rect 432 1788 480 1790
rect 74 1784 107 1788
rect 70 1782 107 1784
rect 70 1781 137 1782
rect 70 1776 101 1781
rect 107 1776 137 1781
rect 70 1772 137 1776
rect 43 1769 137 1772
rect 43 1762 92 1769
rect 43 1756 73 1762
rect 92 1757 97 1762
rect 9 1740 89 1756
rect 101 1748 137 1769
rect 198 1764 387 1788
rect 432 1787 479 1788
rect 445 1782 479 1787
rect 213 1761 387 1764
rect 206 1758 387 1761
rect 415 1781 479 1782
rect 9 1738 28 1740
rect 43 1738 77 1740
rect 9 1722 89 1738
rect 9 1716 28 1722
rect -1 1700 28 1716
rect 43 1706 73 1722
rect 101 1700 107 1748
rect 110 1742 129 1748
rect 144 1742 174 1750
rect 110 1734 174 1742
rect 110 1718 190 1734
rect 206 1727 268 1758
rect 284 1727 346 1758
rect 415 1756 464 1781
rect 479 1756 509 1772
rect 378 1742 408 1750
rect 415 1748 525 1756
rect 378 1734 423 1742
rect 110 1716 129 1718
rect 144 1716 190 1718
rect 110 1700 190 1716
rect 217 1714 252 1727
rect 293 1724 330 1727
rect 293 1722 335 1724
rect 222 1711 252 1714
rect 231 1707 238 1711
rect 238 1706 239 1707
rect 197 1700 207 1706
rect -7 1692 34 1700
rect -7 1666 8 1692
rect 15 1666 34 1692
rect 98 1688 129 1700
rect 144 1688 247 1700
rect 259 1690 285 1716
rect 300 1711 330 1722
rect 362 1718 424 1734
rect 362 1716 408 1718
rect 362 1700 424 1716
rect 436 1700 442 1748
rect 445 1740 525 1748
rect 445 1738 464 1740
rect 479 1738 513 1740
rect 445 1722 525 1738
rect 445 1700 464 1722
rect 479 1706 509 1722
rect 537 1716 543 1790
rect 546 1716 565 1860
rect 580 1716 586 1860
rect 595 1790 608 1860
rect 660 1856 682 1860
rect 653 1834 682 1848
rect 735 1834 751 1848
rect 789 1844 795 1846
rect 802 1844 910 1860
rect 917 1844 923 1846
rect 931 1844 946 1860
rect 1012 1854 1031 1857
rect 653 1832 751 1834
rect 778 1832 946 1844
rect 961 1834 977 1848
rect 1012 1835 1034 1854
rect 1044 1848 1060 1849
rect 1043 1846 1060 1848
rect 1044 1841 1060 1846
rect 1034 1834 1040 1835
rect 1043 1834 1072 1841
rect 961 1833 1072 1834
rect 961 1832 1078 1833
rect 637 1824 688 1832
rect 735 1824 769 1832
rect 637 1812 662 1824
rect 669 1812 688 1824
rect 742 1822 769 1824
rect 778 1822 999 1832
rect 1034 1829 1040 1832
rect 742 1818 999 1822
rect 637 1804 688 1812
rect 735 1804 999 1818
rect 1043 1824 1078 1832
rect 589 1756 608 1790
rect 653 1796 682 1804
rect 653 1790 670 1796
rect 653 1788 687 1790
rect 735 1788 751 1804
rect 752 1794 960 1804
rect 961 1794 977 1804
rect 1025 1800 1040 1815
rect 1043 1812 1044 1824
rect 1051 1812 1078 1824
rect 1043 1804 1078 1812
rect 1043 1803 1072 1804
rect 763 1790 977 1794
rect 778 1788 977 1790
rect 1012 1790 1025 1800
rect 1043 1790 1060 1803
rect 1012 1788 1060 1790
rect 654 1784 687 1788
rect 650 1782 687 1784
rect 650 1781 717 1782
rect 650 1776 681 1781
rect 687 1776 717 1781
rect 650 1772 717 1776
rect 623 1769 717 1772
rect 623 1762 672 1769
rect 623 1756 653 1762
rect 672 1757 677 1762
rect 589 1740 669 1756
rect 681 1748 717 1769
rect 778 1764 967 1788
rect 1012 1787 1059 1788
rect 1025 1782 1059 1787
rect 793 1761 967 1764
rect 786 1758 967 1761
rect 995 1781 1059 1782
rect 589 1738 608 1740
rect 623 1738 657 1740
rect 589 1722 669 1738
rect 589 1716 608 1722
rect 305 1690 408 1700
rect 259 1688 408 1690
rect 429 1688 464 1700
rect 98 1686 260 1688
rect 110 1666 129 1686
rect 144 1684 174 1686
rect -7 1658 34 1666
rect 116 1662 129 1666
rect 181 1670 260 1686
rect 292 1686 464 1688
rect 292 1670 371 1686
rect 378 1684 408 1686
rect -1 1648 28 1658
rect 43 1648 73 1662
rect 116 1648 159 1662
rect 181 1658 371 1670
rect 436 1666 442 1686
rect 166 1648 196 1658
rect 197 1648 355 1658
rect 359 1648 389 1658
rect 393 1648 423 1662
rect 451 1648 464 1686
rect 536 1700 565 1716
rect 579 1700 608 1716
rect 623 1706 653 1722
rect 681 1700 687 1748
rect 690 1742 709 1748
rect 724 1742 754 1750
rect 690 1734 754 1742
rect 690 1718 770 1734
rect 786 1727 848 1758
rect 864 1727 926 1758
rect 995 1756 1044 1781
rect 1059 1756 1089 1772
rect 958 1742 988 1750
rect 995 1748 1105 1756
rect 958 1734 1003 1742
rect 690 1716 709 1718
rect 724 1716 770 1718
rect 690 1700 770 1716
rect 797 1714 832 1727
rect 873 1724 910 1727
rect 873 1722 915 1724
rect 802 1711 832 1714
rect 811 1707 818 1711
rect 818 1706 819 1707
rect 777 1700 787 1706
rect 536 1692 571 1700
rect 536 1666 537 1692
rect 544 1666 571 1692
rect 479 1648 509 1662
rect 536 1658 571 1666
rect 573 1692 614 1700
rect 573 1666 588 1692
rect 595 1666 614 1692
rect 678 1688 709 1700
rect 724 1688 827 1700
rect 839 1690 865 1716
rect 880 1711 910 1722
rect 942 1718 1004 1734
rect 942 1716 988 1718
rect 942 1700 1004 1716
rect 1016 1700 1022 1748
rect 1025 1740 1105 1748
rect 1025 1738 1044 1740
rect 1059 1738 1093 1740
rect 1025 1722 1105 1738
rect 1025 1700 1044 1722
rect 1059 1706 1089 1722
rect 1117 1716 1123 1790
rect 1126 1716 1145 1860
rect 1160 1716 1166 1860
rect 1175 1790 1188 1860
rect 1240 1856 1262 1860
rect 1233 1834 1262 1848
rect 1315 1834 1331 1848
rect 1369 1844 1375 1846
rect 1382 1844 1490 1860
rect 1497 1844 1503 1846
rect 1511 1844 1526 1860
rect 1592 1854 1611 1857
rect 1233 1832 1331 1834
rect 1358 1832 1526 1844
rect 1541 1834 1557 1848
rect 1592 1835 1614 1854
rect 1624 1848 1640 1849
rect 1623 1846 1640 1848
rect 1624 1841 1640 1846
rect 1614 1834 1620 1835
rect 1623 1834 1652 1841
rect 1541 1833 1652 1834
rect 1541 1832 1658 1833
rect 1217 1824 1268 1832
rect 1315 1824 1349 1832
rect 1217 1812 1242 1824
rect 1249 1812 1268 1824
rect 1322 1822 1349 1824
rect 1358 1822 1579 1832
rect 1614 1829 1620 1832
rect 1322 1818 1579 1822
rect 1217 1804 1268 1812
rect 1315 1804 1579 1818
rect 1623 1824 1658 1832
rect 1169 1756 1188 1790
rect 1233 1796 1262 1804
rect 1233 1790 1250 1796
rect 1233 1788 1267 1790
rect 1315 1788 1331 1804
rect 1332 1794 1540 1804
rect 1541 1794 1557 1804
rect 1605 1800 1620 1815
rect 1623 1812 1624 1824
rect 1631 1812 1658 1824
rect 1623 1804 1658 1812
rect 1623 1803 1652 1804
rect 1343 1790 1557 1794
rect 1358 1788 1557 1790
rect 1592 1790 1605 1800
rect 1623 1790 1640 1803
rect 1592 1788 1640 1790
rect 1234 1784 1267 1788
rect 1230 1782 1267 1784
rect 1230 1781 1297 1782
rect 1230 1776 1261 1781
rect 1267 1776 1297 1781
rect 1230 1772 1297 1776
rect 1203 1769 1297 1772
rect 1203 1762 1252 1769
rect 1203 1756 1233 1762
rect 1252 1757 1257 1762
rect 1169 1740 1249 1756
rect 1261 1748 1297 1769
rect 1358 1764 1547 1788
rect 1592 1787 1639 1788
rect 1605 1782 1639 1787
rect 1373 1761 1547 1764
rect 1366 1758 1547 1761
rect 1575 1781 1639 1782
rect 1169 1738 1188 1740
rect 1203 1738 1237 1740
rect 1169 1722 1249 1738
rect 1169 1716 1188 1722
rect 885 1690 988 1700
rect 839 1688 988 1690
rect 1009 1688 1044 1700
rect 678 1686 840 1688
rect 690 1666 709 1686
rect 724 1684 754 1686
rect 573 1658 614 1666
rect 696 1662 709 1666
rect 761 1670 840 1686
rect 872 1686 1044 1688
rect 872 1670 951 1686
rect 958 1684 988 1686
rect 536 1648 565 1658
rect 579 1648 608 1658
rect 623 1648 653 1662
rect 696 1648 739 1662
rect 761 1658 951 1670
rect 1016 1666 1022 1686
rect 746 1648 776 1658
rect 777 1648 935 1658
rect 939 1648 969 1658
rect 973 1648 1003 1662
rect 1031 1648 1044 1686
rect 1116 1700 1145 1716
rect 1159 1700 1188 1716
rect 1203 1706 1233 1722
rect 1261 1700 1267 1748
rect 1270 1742 1289 1748
rect 1304 1742 1334 1750
rect 1270 1734 1334 1742
rect 1270 1718 1350 1734
rect 1366 1727 1428 1758
rect 1444 1727 1506 1758
rect 1575 1756 1624 1781
rect 1639 1756 1669 1772
rect 1538 1742 1568 1750
rect 1575 1748 1685 1756
rect 1538 1734 1583 1742
rect 1270 1716 1289 1718
rect 1304 1716 1350 1718
rect 1270 1700 1350 1716
rect 1377 1714 1412 1727
rect 1453 1724 1490 1727
rect 1453 1722 1495 1724
rect 1382 1711 1412 1714
rect 1391 1707 1398 1711
rect 1398 1706 1399 1707
rect 1357 1700 1367 1706
rect 1116 1692 1151 1700
rect 1116 1666 1117 1692
rect 1124 1666 1151 1692
rect 1059 1648 1089 1662
rect 1116 1658 1151 1666
rect 1153 1692 1194 1700
rect 1153 1666 1168 1692
rect 1175 1666 1194 1692
rect 1258 1688 1289 1700
rect 1304 1688 1407 1700
rect 1419 1690 1445 1716
rect 1460 1711 1490 1722
rect 1522 1718 1584 1734
rect 1522 1716 1568 1718
rect 1522 1700 1584 1716
rect 1596 1700 1602 1748
rect 1605 1740 1685 1748
rect 1605 1738 1624 1740
rect 1639 1738 1673 1740
rect 1605 1722 1685 1738
rect 1605 1700 1624 1722
rect 1639 1706 1669 1722
rect 1697 1716 1703 1790
rect 1706 1716 1725 1860
rect 1740 1716 1746 1860
rect 1755 1790 1768 1860
rect 1820 1856 1842 1860
rect 1813 1834 1842 1848
rect 1895 1834 1911 1848
rect 1949 1844 1955 1846
rect 1962 1844 2070 1860
rect 2077 1844 2083 1846
rect 2091 1844 2106 1860
rect 2172 1854 2191 1857
rect 1813 1832 1911 1834
rect 1938 1832 2106 1844
rect 2121 1834 2137 1848
rect 2172 1835 2194 1854
rect 2204 1848 2220 1849
rect 2203 1846 2220 1848
rect 2204 1841 2220 1846
rect 2194 1834 2200 1835
rect 2203 1834 2232 1841
rect 2121 1833 2232 1834
rect 2121 1832 2238 1833
rect 1797 1824 1848 1832
rect 1895 1824 1929 1832
rect 1797 1812 1822 1824
rect 1829 1812 1848 1824
rect 1902 1822 1929 1824
rect 1938 1822 2159 1832
rect 2194 1829 2200 1832
rect 1902 1818 2159 1822
rect 1797 1804 1848 1812
rect 1895 1804 2159 1818
rect 2203 1824 2238 1832
rect 1749 1756 1768 1790
rect 1813 1796 1842 1804
rect 1813 1790 1830 1796
rect 1813 1788 1847 1790
rect 1895 1788 1911 1804
rect 1912 1794 2120 1804
rect 2121 1794 2137 1804
rect 2185 1800 2200 1815
rect 2203 1812 2204 1824
rect 2211 1812 2238 1824
rect 2203 1804 2238 1812
rect 2203 1803 2232 1804
rect 1923 1790 2137 1794
rect 1938 1788 2137 1790
rect 2172 1790 2185 1800
rect 2203 1790 2220 1803
rect 2172 1788 2220 1790
rect 1814 1784 1847 1788
rect 1810 1782 1847 1784
rect 1810 1781 1877 1782
rect 1810 1776 1841 1781
rect 1847 1776 1877 1781
rect 1810 1772 1877 1776
rect 1783 1769 1877 1772
rect 1783 1762 1832 1769
rect 1783 1756 1813 1762
rect 1832 1757 1837 1762
rect 1749 1740 1829 1756
rect 1841 1748 1877 1769
rect 1938 1764 2127 1788
rect 2172 1787 2219 1788
rect 2185 1782 2219 1787
rect 1953 1761 2127 1764
rect 1946 1758 2127 1761
rect 2155 1781 2219 1782
rect 1749 1738 1768 1740
rect 1783 1738 1817 1740
rect 1749 1722 1829 1738
rect 1749 1716 1768 1722
rect 1465 1690 1568 1700
rect 1419 1688 1568 1690
rect 1589 1688 1624 1700
rect 1258 1686 1420 1688
rect 1270 1666 1289 1686
rect 1304 1684 1334 1686
rect 1153 1658 1194 1666
rect 1276 1662 1289 1666
rect 1341 1670 1420 1686
rect 1452 1686 1624 1688
rect 1452 1670 1531 1686
rect 1538 1684 1568 1686
rect 1116 1648 1145 1658
rect 1159 1648 1188 1658
rect 1203 1648 1233 1662
rect 1276 1648 1319 1662
rect 1341 1658 1531 1670
rect 1596 1666 1602 1686
rect 1326 1648 1356 1658
rect 1357 1648 1515 1658
rect 1519 1648 1549 1658
rect 1553 1648 1583 1662
rect 1611 1648 1624 1686
rect 1696 1700 1725 1716
rect 1739 1700 1768 1716
rect 1783 1706 1813 1722
rect 1841 1700 1847 1748
rect 1850 1742 1869 1748
rect 1884 1742 1914 1750
rect 1850 1734 1914 1742
rect 1850 1718 1930 1734
rect 1946 1727 2008 1758
rect 2024 1727 2086 1758
rect 2155 1756 2204 1781
rect 2219 1756 2249 1772
rect 2118 1742 2148 1750
rect 2155 1748 2265 1756
rect 2118 1734 2163 1742
rect 1850 1716 1869 1718
rect 1884 1716 1930 1718
rect 1850 1700 1930 1716
rect 1957 1714 1992 1727
rect 2033 1724 2070 1727
rect 2033 1722 2075 1724
rect 1962 1711 1992 1714
rect 1971 1707 1978 1711
rect 1978 1706 1979 1707
rect 1937 1700 1947 1706
rect 1696 1692 1731 1700
rect 1696 1666 1697 1692
rect 1704 1666 1731 1692
rect 1639 1648 1669 1662
rect 1696 1658 1731 1666
rect 1733 1692 1774 1700
rect 1733 1666 1748 1692
rect 1755 1666 1774 1692
rect 1838 1688 1869 1700
rect 1884 1688 1987 1700
rect 1999 1690 2025 1716
rect 2040 1711 2070 1722
rect 2102 1718 2164 1734
rect 2102 1716 2148 1718
rect 2102 1700 2164 1716
rect 2176 1700 2182 1748
rect 2185 1740 2265 1748
rect 2185 1738 2204 1740
rect 2219 1738 2253 1740
rect 2185 1722 2265 1738
rect 2185 1700 2204 1722
rect 2219 1706 2249 1722
rect 2277 1716 2283 1790
rect 2286 1716 2305 1860
rect 2320 1716 2326 1860
rect 2335 1790 2348 1860
rect 2400 1856 2422 1860
rect 2393 1834 2422 1848
rect 2475 1834 2491 1848
rect 2529 1844 2535 1846
rect 2542 1844 2650 1860
rect 2657 1844 2663 1846
rect 2671 1844 2686 1860
rect 2752 1854 2771 1857
rect 2393 1832 2491 1834
rect 2518 1832 2686 1844
rect 2701 1834 2717 1848
rect 2752 1835 2774 1854
rect 2784 1848 2800 1849
rect 2783 1846 2800 1848
rect 2784 1841 2800 1846
rect 2774 1834 2780 1835
rect 2783 1834 2812 1841
rect 2701 1833 2812 1834
rect 2701 1832 2818 1833
rect 2377 1824 2428 1832
rect 2475 1824 2509 1832
rect 2377 1812 2402 1824
rect 2409 1812 2428 1824
rect 2482 1822 2509 1824
rect 2518 1822 2739 1832
rect 2774 1829 2780 1832
rect 2482 1818 2739 1822
rect 2377 1804 2428 1812
rect 2475 1804 2739 1818
rect 2783 1824 2818 1832
rect 2329 1756 2348 1790
rect 2393 1796 2422 1804
rect 2393 1790 2410 1796
rect 2393 1788 2427 1790
rect 2475 1788 2491 1804
rect 2492 1794 2700 1804
rect 2701 1794 2717 1804
rect 2765 1800 2780 1815
rect 2783 1812 2784 1824
rect 2791 1812 2818 1824
rect 2783 1804 2818 1812
rect 2783 1803 2812 1804
rect 2503 1790 2717 1794
rect 2518 1788 2717 1790
rect 2752 1790 2765 1800
rect 2783 1790 2800 1803
rect 2752 1788 2800 1790
rect 2394 1784 2427 1788
rect 2390 1782 2427 1784
rect 2390 1781 2457 1782
rect 2390 1776 2421 1781
rect 2427 1776 2457 1781
rect 2390 1772 2457 1776
rect 2363 1769 2457 1772
rect 2363 1762 2412 1769
rect 2363 1756 2393 1762
rect 2412 1757 2417 1762
rect 2329 1740 2409 1756
rect 2421 1748 2457 1769
rect 2518 1764 2707 1788
rect 2752 1787 2799 1788
rect 2765 1782 2799 1787
rect 2533 1761 2707 1764
rect 2526 1758 2707 1761
rect 2735 1781 2799 1782
rect 2329 1738 2348 1740
rect 2363 1738 2397 1740
rect 2329 1722 2409 1738
rect 2329 1716 2348 1722
rect 2045 1690 2148 1700
rect 1999 1688 2148 1690
rect 2169 1688 2204 1700
rect 1838 1686 2000 1688
rect 1850 1666 1869 1686
rect 1884 1684 1914 1686
rect 1733 1658 1774 1666
rect 1856 1662 1869 1666
rect 1921 1670 2000 1686
rect 2032 1686 2204 1688
rect 2032 1670 2111 1686
rect 2118 1684 2148 1686
rect 1696 1648 1725 1658
rect 1739 1648 1768 1658
rect 1783 1648 1813 1662
rect 1856 1648 1899 1662
rect 1921 1658 2111 1670
rect 2176 1666 2182 1686
rect 1906 1648 1936 1658
rect 1937 1648 2095 1658
rect 2099 1648 2129 1658
rect 2133 1648 2163 1662
rect 2191 1648 2204 1686
rect 2276 1700 2305 1716
rect 2319 1700 2348 1716
rect 2363 1706 2393 1722
rect 2421 1700 2427 1748
rect 2430 1742 2449 1748
rect 2464 1742 2494 1750
rect 2430 1734 2494 1742
rect 2430 1718 2510 1734
rect 2526 1727 2588 1758
rect 2604 1727 2666 1758
rect 2735 1756 2784 1781
rect 2799 1756 2829 1772
rect 2698 1742 2728 1750
rect 2735 1748 2845 1756
rect 2698 1734 2743 1742
rect 2430 1716 2449 1718
rect 2464 1716 2510 1718
rect 2430 1700 2510 1716
rect 2537 1714 2572 1727
rect 2613 1724 2650 1727
rect 2613 1722 2655 1724
rect 2542 1711 2572 1714
rect 2551 1707 2558 1711
rect 2558 1706 2559 1707
rect 2517 1700 2527 1706
rect 2276 1692 2311 1700
rect 2276 1666 2277 1692
rect 2284 1666 2311 1692
rect 2219 1648 2249 1662
rect 2276 1658 2311 1666
rect 2313 1692 2354 1700
rect 2313 1666 2328 1692
rect 2335 1666 2354 1692
rect 2418 1688 2449 1700
rect 2464 1688 2567 1700
rect 2579 1690 2605 1716
rect 2620 1711 2650 1722
rect 2682 1718 2744 1734
rect 2682 1716 2728 1718
rect 2682 1700 2744 1716
rect 2756 1700 2762 1748
rect 2765 1740 2845 1748
rect 2765 1738 2784 1740
rect 2799 1738 2833 1740
rect 2765 1722 2845 1738
rect 2765 1700 2784 1722
rect 2799 1706 2829 1722
rect 2857 1716 2863 1790
rect 2866 1716 2885 1860
rect 2900 1716 2906 1860
rect 2915 1790 2928 1860
rect 2980 1856 3002 1860
rect 2973 1834 3002 1848
rect 3055 1834 3071 1848
rect 3109 1844 3115 1846
rect 3122 1844 3230 1860
rect 3237 1844 3243 1846
rect 3251 1844 3266 1860
rect 3332 1854 3351 1857
rect 2973 1832 3071 1834
rect 3098 1832 3266 1844
rect 3281 1834 3297 1848
rect 3332 1835 3354 1854
rect 3364 1848 3380 1849
rect 3363 1846 3380 1848
rect 3364 1841 3380 1846
rect 3354 1834 3360 1835
rect 3363 1834 3392 1841
rect 3281 1833 3392 1834
rect 3281 1832 3398 1833
rect 2957 1824 3008 1832
rect 3055 1824 3089 1832
rect 2957 1812 2982 1824
rect 2989 1812 3008 1824
rect 3062 1822 3089 1824
rect 3098 1822 3319 1832
rect 3354 1829 3360 1832
rect 3062 1818 3319 1822
rect 2957 1804 3008 1812
rect 3055 1804 3319 1818
rect 3363 1824 3398 1832
rect 2909 1756 2928 1790
rect 2973 1796 3002 1804
rect 2973 1790 2990 1796
rect 2973 1788 3007 1790
rect 3055 1788 3071 1804
rect 3072 1794 3280 1804
rect 3281 1794 3297 1804
rect 3345 1800 3360 1815
rect 3363 1812 3364 1824
rect 3371 1812 3398 1824
rect 3363 1804 3398 1812
rect 3363 1803 3392 1804
rect 3083 1790 3297 1794
rect 3098 1788 3297 1790
rect 3332 1790 3345 1800
rect 3363 1790 3380 1803
rect 3332 1788 3380 1790
rect 2974 1784 3007 1788
rect 2970 1782 3007 1784
rect 2970 1781 3037 1782
rect 2970 1776 3001 1781
rect 3007 1776 3037 1781
rect 2970 1772 3037 1776
rect 2943 1769 3037 1772
rect 2943 1762 2992 1769
rect 2943 1756 2973 1762
rect 2992 1757 2997 1762
rect 2909 1740 2989 1756
rect 3001 1748 3037 1769
rect 3098 1764 3287 1788
rect 3332 1787 3379 1788
rect 3345 1782 3379 1787
rect 3113 1761 3287 1764
rect 3106 1758 3287 1761
rect 3315 1781 3379 1782
rect 2909 1738 2928 1740
rect 2943 1738 2977 1740
rect 2909 1722 2989 1738
rect 2909 1716 2928 1722
rect 2625 1690 2728 1700
rect 2579 1688 2728 1690
rect 2749 1688 2784 1700
rect 2418 1686 2580 1688
rect 2430 1666 2449 1686
rect 2464 1684 2494 1686
rect 2313 1658 2354 1666
rect 2436 1662 2449 1666
rect 2501 1670 2580 1686
rect 2612 1686 2784 1688
rect 2612 1670 2691 1686
rect 2698 1684 2728 1686
rect 2276 1648 2305 1658
rect 2319 1648 2348 1658
rect 2363 1648 2393 1662
rect 2436 1648 2479 1662
rect 2501 1658 2691 1670
rect 2756 1666 2762 1686
rect 2486 1648 2516 1658
rect 2517 1648 2675 1658
rect 2679 1648 2709 1658
rect 2713 1648 2743 1662
rect 2771 1648 2784 1686
rect 2856 1700 2885 1716
rect 2899 1700 2928 1716
rect 2943 1706 2973 1722
rect 3001 1700 3007 1748
rect 3010 1742 3029 1748
rect 3044 1742 3074 1750
rect 3010 1734 3074 1742
rect 3010 1718 3090 1734
rect 3106 1727 3168 1758
rect 3184 1727 3246 1758
rect 3315 1756 3364 1781
rect 3379 1756 3409 1772
rect 3278 1742 3308 1750
rect 3315 1748 3425 1756
rect 3278 1734 3323 1742
rect 3010 1716 3029 1718
rect 3044 1716 3090 1718
rect 3010 1700 3090 1716
rect 3117 1714 3152 1727
rect 3193 1724 3230 1727
rect 3193 1722 3235 1724
rect 3122 1711 3152 1714
rect 3131 1707 3138 1711
rect 3138 1706 3139 1707
rect 3097 1700 3107 1706
rect 2856 1692 2891 1700
rect 2856 1666 2857 1692
rect 2864 1666 2891 1692
rect 2799 1648 2829 1662
rect 2856 1658 2891 1666
rect 2893 1692 2934 1700
rect 2893 1666 2908 1692
rect 2915 1666 2934 1692
rect 2998 1688 3029 1700
rect 3044 1688 3147 1700
rect 3159 1690 3185 1716
rect 3200 1711 3230 1722
rect 3262 1718 3324 1734
rect 3262 1716 3308 1718
rect 3262 1700 3324 1716
rect 3336 1700 3342 1748
rect 3345 1740 3425 1748
rect 3345 1738 3364 1740
rect 3379 1738 3413 1740
rect 3345 1722 3425 1738
rect 3345 1700 3364 1722
rect 3379 1706 3409 1722
rect 3437 1716 3443 1790
rect 3446 1716 3465 1860
rect 3480 1716 3486 1860
rect 3495 1790 3508 1860
rect 3560 1856 3582 1860
rect 3553 1834 3582 1848
rect 3635 1834 3651 1848
rect 3689 1844 3695 1846
rect 3702 1844 3810 1860
rect 3817 1844 3823 1846
rect 3831 1844 3846 1860
rect 3912 1854 3931 1857
rect 3553 1832 3651 1834
rect 3678 1832 3846 1844
rect 3861 1834 3877 1848
rect 3912 1835 3934 1854
rect 3944 1848 3960 1849
rect 3943 1846 3960 1848
rect 3944 1841 3960 1846
rect 3934 1834 3940 1835
rect 3943 1834 3972 1841
rect 3861 1833 3972 1834
rect 3861 1832 3978 1833
rect 3537 1824 3588 1832
rect 3635 1824 3669 1832
rect 3537 1812 3562 1824
rect 3569 1812 3588 1824
rect 3642 1822 3669 1824
rect 3678 1822 3899 1832
rect 3934 1829 3940 1832
rect 3642 1818 3899 1822
rect 3537 1804 3588 1812
rect 3635 1804 3899 1818
rect 3943 1824 3978 1832
rect 3489 1756 3508 1790
rect 3553 1796 3582 1804
rect 3553 1790 3570 1796
rect 3553 1788 3587 1790
rect 3635 1788 3651 1804
rect 3652 1794 3860 1804
rect 3861 1794 3877 1804
rect 3925 1800 3940 1815
rect 3943 1812 3944 1824
rect 3951 1812 3978 1824
rect 3943 1804 3978 1812
rect 3943 1803 3972 1804
rect 3663 1790 3877 1794
rect 3678 1788 3877 1790
rect 3912 1790 3925 1800
rect 3943 1790 3960 1803
rect 3912 1788 3960 1790
rect 3554 1784 3587 1788
rect 3550 1782 3587 1784
rect 3550 1781 3617 1782
rect 3550 1776 3581 1781
rect 3587 1776 3617 1781
rect 3550 1772 3617 1776
rect 3523 1769 3617 1772
rect 3523 1762 3572 1769
rect 3523 1756 3553 1762
rect 3572 1757 3577 1762
rect 3489 1740 3569 1756
rect 3581 1748 3617 1769
rect 3678 1764 3867 1788
rect 3912 1787 3959 1788
rect 3925 1782 3959 1787
rect 3693 1761 3867 1764
rect 3686 1758 3867 1761
rect 3895 1781 3959 1782
rect 3489 1738 3508 1740
rect 3523 1738 3557 1740
rect 3489 1722 3569 1738
rect 3489 1716 3508 1722
rect 3205 1690 3308 1700
rect 3159 1688 3308 1690
rect 3329 1688 3364 1700
rect 2998 1686 3160 1688
rect 3010 1666 3029 1686
rect 3044 1684 3074 1686
rect 2893 1658 2934 1666
rect 3016 1662 3029 1666
rect 3081 1670 3160 1686
rect 3192 1686 3364 1688
rect 3192 1670 3271 1686
rect 3278 1684 3308 1686
rect 2856 1648 2885 1658
rect 2899 1648 2928 1658
rect 2943 1648 2973 1662
rect 3016 1648 3059 1662
rect 3081 1658 3271 1670
rect 3336 1666 3342 1686
rect 3066 1648 3096 1658
rect 3097 1648 3255 1658
rect 3259 1648 3289 1658
rect 3293 1648 3323 1662
rect 3351 1648 3364 1686
rect 3436 1700 3465 1716
rect 3479 1700 3508 1716
rect 3523 1706 3553 1722
rect 3581 1700 3587 1748
rect 3590 1742 3609 1748
rect 3624 1742 3654 1750
rect 3590 1734 3654 1742
rect 3590 1718 3670 1734
rect 3686 1727 3748 1758
rect 3764 1727 3826 1758
rect 3895 1756 3944 1781
rect 3959 1756 3989 1772
rect 3858 1742 3888 1750
rect 3895 1748 4005 1756
rect 3858 1734 3903 1742
rect 3590 1716 3609 1718
rect 3624 1716 3670 1718
rect 3590 1700 3670 1716
rect 3697 1714 3732 1727
rect 3773 1724 3810 1727
rect 3773 1722 3815 1724
rect 3702 1711 3732 1714
rect 3711 1707 3718 1711
rect 3718 1706 3719 1707
rect 3677 1700 3687 1706
rect 3436 1692 3471 1700
rect 3436 1666 3437 1692
rect 3444 1666 3471 1692
rect 3379 1648 3409 1662
rect 3436 1658 3471 1666
rect 3473 1692 3514 1700
rect 3473 1666 3488 1692
rect 3495 1666 3514 1692
rect 3578 1688 3609 1700
rect 3624 1688 3727 1700
rect 3739 1690 3765 1716
rect 3780 1711 3810 1722
rect 3842 1718 3904 1734
rect 3842 1716 3888 1718
rect 3842 1700 3904 1716
rect 3916 1700 3922 1748
rect 3925 1740 4005 1748
rect 3925 1738 3944 1740
rect 3959 1738 3993 1740
rect 3925 1722 4005 1738
rect 3925 1700 3944 1722
rect 3959 1706 3989 1722
rect 4017 1716 4023 1790
rect 4026 1716 4045 1860
rect 4060 1716 4066 1860
rect 4075 1790 4088 1860
rect 4140 1856 4162 1860
rect 4133 1834 4162 1848
rect 4215 1834 4231 1848
rect 4269 1844 4275 1846
rect 4282 1844 4390 1860
rect 4397 1844 4403 1846
rect 4411 1844 4426 1860
rect 4492 1854 4511 1857
rect 4133 1832 4231 1834
rect 4258 1832 4426 1844
rect 4441 1834 4457 1848
rect 4492 1835 4514 1854
rect 4524 1848 4540 1849
rect 4523 1846 4540 1848
rect 4524 1841 4540 1846
rect 4514 1834 4520 1835
rect 4523 1834 4552 1841
rect 4441 1833 4552 1834
rect 4441 1832 4558 1833
rect 4117 1824 4168 1832
rect 4215 1824 4249 1832
rect 4117 1812 4142 1824
rect 4149 1812 4168 1824
rect 4222 1822 4249 1824
rect 4258 1822 4479 1832
rect 4514 1829 4520 1832
rect 4222 1818 4479 1822
rect 4117 1804 4168 1812
rect 4215 1804 4479 1818
rect 4523 1824 4558 1832
rect 4069 1756 4088 1790
rect 4133 1796 4162 1804
rect 4133 1790 4150 1796
rect 4133 1788 4167 1790
rect 4215 1788 4231 1804
rect 4232 1794 4440 1804
rect 4441 1794 4457 1804
rect 4505 1800 4520 1815
rect 4523 1812 4524 1824
rect 4531 1812 4558 1824
rect 4523 1804 4558 1812
rect 4523 1803 4552 1804
rect 4243 1790 4457 1794
rect 4258 1788 4457 1790
rect 4492 1790 4505 1800
rect 4523 1790 4540 1803
rect 4492 1788 4540 1790
rect 4134 1784 4167 1788
rect 4130 1782 4167 1784
rect 4130 1781 4197 1782
rect 4130 1776 4161 1781
rect 4167 1776 4197 1781
rect 4130 1772 4197 1776
rect 4103 1769 4197 1772
rect 4103 1762 4152 1769
rect 4103 1756 4133 1762
rect 4152 1757 4157 1762
rect 4069 1740 4149 1756
rect 4161 1748 4197 1769
rect 4258 1764 4447 1788
rect 4492 1787 4539 1788
rect 4505 1782 4539 1787
rect 4273 1761 4447 1764
rect 4266 1758 4447 1761
rect 4475 1781 4539 1782
rect 4069 1738 4088 1740
rect 4103 1738 4137 1740
rect 4069 1722 4149 1738
rect 4069 1716 4088 1722
rect 3785 1690 3888 1700
rect 3739 1688 3888 1690
rect 3909 1688 3944 1700
rect 3578 1686 3740 1688
rect 3590 1666 3609 1686
rect 3624 1684 3654 1686
rect 3473 1658 3514 1666
rect 3596 1662 3609 1666
rect 3661 1670 3740 1686
rect 3772 1686 3944 1688
rect 3772 1670 3851 1686
rect 3858 1684 3888 1686
rect 3436 1648 3465 1658
rect 3479 1648 3508 1658
rect 3523 1648 3553 1662
rect 3596 1648 3639 1662
rect 3661 1658 3851 1670
rect 3916 1666 3922 1686
rect 3646 1648 3676 1658
rect 3677 1648 3835 1658
rect 3839 1648 3869 1658
rect 3873 1648 3903 1662
rect 3931 1648 3944 1686
rect 4016 1700 4045 1716
rect 4059 1700 4088 1716
rect 4103 1706 4133 1722
rect 4161 1700 4167 1748
rect 4170 1742 4189 1748
rect 4204 1742 4234 1750
rect 4170 1734 4234 1742
rect 4170 1718 4250 1734
rect 4266 1727 4328 1758
rect 4344 1727 4406 1758
rect 4475 1756 4524 1781
rect 4539 1756 4569 1772
rect 4438 1742 4468 1750
rect 4475 1748 4585 1756
rect 4438 1734 4483 1742
rect 4170 1716 4189 1718
rect 4204 1716 4250 1718
rect 4170 1700 4250 1716
rect 4277 1714 4312 1727
rect 4353 1724 4390 1727
rect 4353 1722 4395 1724
rect 4282 1711 4312 1714
rect 4291 1707 4298 1711
rect 4298 1706 4299 1707
rect 4257 1700 4267 1706
rect 4016 1692 4051 1700
rect 4016 1666 4017 1692
rect 4024 1666 4051 1692
rect 3959 1648 3989 1662
rect 4016 1658 4051 1666
rect 4053 1692 4094 1700
rect 4053 1666 4068 1692
rect 4075 1666 4094 1692
rect 4158 1688 4189 1700
rect 4204 1688 4307 1700
rect 4319 1690 4345 1716
rect 4360 1711 4390 1722
rect 4422 1718 4484 1734
rect 4422 1716 4468 1718
rect 4422 1700 4484 1716
rect 4496 1700 4502 1748
rect 4505 1740 4585 1748
rect 4505 1738 4524 1740
rect 4539 1738 4573 1740
rect 4505 1722 4585 1738
rect 4505 1700 4524 1722
rect 4539 1706 4569 1722
rect 4597 1716 4603 1790
rect 4606 1716 4625 1860
rect 4640 1716 4646 1860
rect 4655 1790 4668 1860
rect 4720 1856 4742 1860
rect 4713 1834 4742 1848
rect 4795 1834 4811 1848
rect 4849 1844 4855 1846
rect 4862 1844 4970 1860
rect 4977 1844 4983 1846
rect 4991 1844 5006 1860
rect 5072 1854 5091 1857
rect 4713 1832 4811 1834
rect 4838 1832 5006 1844
rect 5021 1834 5037 1848
rect 5072 1835 5094 1854
rect 5104 1848 5120 1849
rect 5103 1846 5120 1848
rect 5104 1841 5120 1846
rect 5094 1834 5100 1835
rect 5103 1834 5132 1841
rect 5021 1833 5132 1834
rect 5021 1832 5138 1833
rect 4697 1824 4748 1832
rect 4795 1824 4829 1832
rect 4697 1812 4722 1824
rect 4729 1812 4748 1824
rect 4802 1822 4829 1824
rect 4838 1822 5059 1832
rect 5094 1829 5100 1832
rect 4802 1818 5059 1822
rect 4697 1804 4748 1812
rect 4795 1804 5059 1818
rect 5103 1824 5138 1832
rect 4649 1756 4668 1790
rect 4713 1796 4742 1804
rect 4713 1790 4730 1796
rect 4713 1788 4747 1790
rect 4795 1788 4811 1804
rect 4812 1794 5020 1804
rect 5021 1794 5037 1804
rect 5085 1800 5100 1815
rect 5103 1812 5104 1824
rect 5111 1812 5138 1824
rect 5103 1804 5138 1812
rect 5103 1803 5132 1804
rect 4823 1790 5037 1794
rect 4838 1788 5037 1790
rect 5072 1790 5085 1800
rect 5103 1790 5120 1803
rect 5072 1788 5120 1790
rect 4714 1784 4747 1788
rect 4710 1782 4747 1784
rect 4710 1781 4777 1782
rect 4710 1776 4741 1781
rect 4747 1776 4777 1781
rect 4710 1772 4777 1776
rect 4683 1769 4777 1772
rect 4683 1762 4732 1769
rect 4683 1756 4713 1762
rect 4732 1757 4737 1762
rect 4649 1740 4729 1756
rect 4741 1748 4777 1769
rect 4838 1764 5027 1788
rect 5072 1787 5119 1788
rect 5085 1782 5119 1787
rect 4853 1761 5027 1764
rect 4846 1758 5027 1761
rect 5055 1781 5119 1782
rect 4649 1738 4668 1740
rect 4683 1738 4717 1740
rect 4649 1722 4729 1738
rect 4649 1716 4668 1722
rect 4365 1690 4468 1700
rect 4319 1688 4468 1690
rect 4489 1688 4524 1700
rect 4158 1686 4320 1688
rect 4170 1666 4189 1686
rect 4204 1684 4234 1686
rect 4053 1658 4094 1666
rect 4176 1662 4189 1666
rect 4241 1670 4320 1686
rect 4352 1686 4524 1688
rect 4352 1670 4431 1686
rect 4438 1684 4468 1686
rect 4016 1648 4045 1658
rect 4059 1648 4088 1658
rect 4103 1648 4133 1662
rect 4176 1648 4219 1662
rect 4241 1658 4431 1670
rect 4496 1666 4502 1686
rect 4226 1648 4256 1658
rect 4257 1648 4415 1658
rect 4419 1648 4449 1658
rect 4453 1648 4483 1662
rect 4511 1648 4524 1686
rect 4596 1700 4625 1716
rect 4639 1700 4668 1716
rect 4683 1706 4713 1722
rect 4741 1700 4747 1748
rect 4750 1742 4769 1748
rect 4784 1742 4814 1750
rect 4750 1734 4814 1742
rect 4750 1718 4830 1734
rect 4846 1727 4908 1758
rect 4924 1727 4986 1758
rect 5055 1756 5104 1781
rect 5119 1756 5149 1772
rect 5018 1742 5048 1750
rect 5055 1748 5165 1756
rect 5018 1734 5063 1742
rect 4750 1716 4769 1718
rect 4784 1716 4830 1718
rect 4750 1700 4830 1716
rect 4857 1714 4892 1727
rect 4933 1724 4970 1727
rect 4933 1722 4975 1724
rect 4862 1711 4892 1714
rect 4871 1707 4878 1711
rect 4878 1706 4879 1707
rect 4837 1700 4847 1706
rect 4596 1692 4631 1700
rect 4596 1666 4597 1692
rect 4604 1666 4631 1692
rect 4539 1648 4569 1662
rect 4596 1658 4631 1666
rect 4633 1692 4674 1700
rect 4633 1666 4648 1692
rect 4655 1666 4674 1692
rect 4738 1688 4769 1700
rect 4784 1688 4887 1700
rect 4899 1690 4925 1716
rect 4940 1711 4970 1722
rect 5002 1718 5064 1734
rect 5002 1716 5048 1718
rect 5002 1700 5064 1716
rect 5076 1700 5082 1748
rect 5085 1740 5165 1748
rect 5085 1738 5104 1740
rect 5119 1738 5153 1740
rect 5085 1722 5165 1738
rect 5085 1700 5104 1722
rect 5119 1706 5149 1722
rect 5177 1716 5183 1790
rect 5186 1716 5205 1860
rect 5220 1716 5226 1860
rect 5235 1790 5248 1860
rect 5300 1856 5322 1860
rect 5293 1834 5322 1848
rect 5375 1834 5391 1848
rect 5429 1844 5435 1846
rect 5442 1844 5550 1860
rect 5557 1844 5563 1846
rect 5571 1844 5586 1860
rect 5652 1854 5671 1857
rect 5293 1832 5391 1834
rect 5418 1832 5586 1844
rect 5601 1834 5617 1848
rect 5652 1835 5674 1854
rect 5684 1848 5700 1849
rect 5683 1846 5700 1848
rect 5684 1841 5700 1846
rect 5674 1834 5680 1835
rect 5683 1834 5712 1841
rect 5601 1833 5712 1834
rect 5601 1832 5718 1833
rect 5277 1824 5328 1832
rect 5375 1824 5409 1832
rect 5277 1812 5302 1824
rect 5309 1812 5328 1824
rect 5382 1822 5409 1824
rect 5418 1822 5639 1832
rect 5674 1829 5680 1832
rect 5382 1818 5639 1822
rect 5277 1804 5328 1812
rect 5375 1804 5639 1818
rect 5683 1824 5718 1832
rect 5229 1756 5248 1790
rect 5293 1796 5322 1804
rect 5293 1790 5310 1796
rect 5293 1788 5327 1790
rect 5375 1788 5391 1804
rect 5392 1794 5600 1804
rect 5601 1794 5617 1804
rect 5665 1800 5680 1815
rect 5683 1812 5684 1824
rect 5691 1812 5718 1824
rect 5683 1804 5718 1812
rect 5683 1803 5712 1804
rect 5403 1790 5617 1794
rect 5418 1788 5617 1790
rect 5652 1790 5665 1800
rect 5683 1790 5700 1803
rect 5652 1788 5700 1790
rect 5294 1784 5327 1788
rect 5290 1782 5327 1784
rect 5290 1781 5357 1782
rect 5290 1776 5321 1781
rect 5327 1776 5357 1781
rect 5290 1772 5357 1776
rect 5263 1769 5357 1772
rect 5263 1762 5312 1769
rect 5263 1756 5293 1762
rect 5312 1757 5317 1762
rect 5229 1740 5309 1756
rect 5321 1748 5357 1769
rect 5418 1764 5607 1788
rect 5652 1787 5699 1788
rect 5665 1782 5699 1787
rect 5433 1761 5607 1764
rect 5426 1758 5607 1761
rect 5635 1781 5699 1782
rect 5229 1738 5248 1740
rect 5263 1738 5297 1740
rect 5229 1722 5309 1738
rect 5229 1716 5248 1722
rect 4945 1690 5048 1700
rect 4899 1688 5048 1690
rect 5069 1688 5104 1700
rect 4738 1686 4900 1688
rect 4750 1666 4769 1686
rect 4784 1684 4814 1686
rect 4633 1658 4674 1666
rect 4756 1662 4769 1666
rect 4821 1670 4900 1686
rect 4932 1686 5104 1688
rect 4932 1670 5011 1686
rect 5018 1684 5048 1686
rect 4596 1648 4625 1658
rect 4639 1648 4668 1658
rect 4683 1648 4713 1662
rect 4756 1648 4799 1662
rect 4821 1658 5011 1670
rect 5076 1666 5082 1686
rect 4806 1648 4836 1658
rect 4837 1648 4995 1658
rect 4999 1648 5029 1658
rect 5033 1648 5063 1662
rect 5091 1648 5104 1686
rect 5176 1700 5205 1716
rect 5219 1700 5248 1716
rect 5263 1706 5293 1722
rect 5321 1700 5327 1748
rect 5330 1742 5349 1748
rect 5364 1742 5394 1750
rect 5330 1734 5394 1742
rect 5330 1718 5410 1734
rect 5426 1727 5488 1758
rect 5504 1727 5566 1758
rect 5635 1756 5684 1781
rect 5699 1756 5729 1772
rect 5598 1742 5628 1750
rect 5635 1748 5745 1756
rect 5598 1734 5643 1742
rect 5330 1716 5349 1718
rect 5364 1716 5410 1718
rect 5330 1700 5410 1716
rect 5437 1714 5472 1727
rect 5513 1724 5550 1727
rect 5513 1722 5555 1724
rect 5442 1711 5472 1714
rect 5451 1707 5458 1711
rect 5458 1706 5459 1707
rect 5417 1700 5427 1706
rect 5176 1692 5211 1700
rect 5176 1666 5177 1692
rect 5184 1666 5211 1692
rect 5119 1648 5149 1662
rect 5176 1658 5211 1666
rect 5213 1692 5254 1700
rect 5213 1666 5228 1692
rect 5235 1666 5254 1692
rect 5318 1688 5349 1700
rect 5364 1688 5467 1700
rect 5479 1690 5505 1716
rect 5520 1711 5550 1722
rect 5582 1718 5644 1734
rect 5582 1716 5628 1718
rect 5582 1700 5644 1716
rect 5656 1700 5662 1748
rect 5665 1740 5745 1748
rect 5665 1738 5684 1740
rect 5699 1738 5733 1740
rect 5665 1722 5745 1738
rect 5665 1700 5684 1722
rect 5699 1706 5729 1722
rect 5757 1716 5763 1790
rect 5766 1716 5785 1860
rect 5800 1716 5806 1860
rect 5815 1790 5828 1860
rect 5880 1856 5902 1860
rect 5873 1834 5902 1848
rect 5955 1834 5971 1848
rect 6009 1844 6015 1846
rect 6022 1844 6130 1860
rect 6137 1844 6143 1846
rect 6151 1844 6166 1860
rect 6232 1854 6251 1857
rect 5873 1832 5971 1834
rect 5998 1832 6166 1844
rect 6181 1834 6197 1848
rect 6232 1835 6254 1854
rect 6264 1848 6280 1849
rect 6263 1846 6280 1848
rect 6264 1841 6280 1846
rect 6254 1834 6260 1835
rect 6263 1834 6292 1841
rect 6181 1833 6292 1834
rect 6181 1832 6298 1833
rect 5857 1824 5908 1832
rect 5955 1824 5989 1832
rect 5857 1812 5882 1824
rect 5889 1812 5908 1824
rect 5962 1822 5989 1824
rect 5998 1822 6219 1832
rect 6254 1829 6260 1832
rect 5962 1818 6219 1822
rect 5857 1804 5908 1812
rect 5955 1804 6219 1818
rect 6263 1824 6298 1832
rect 5809 1756 5828 1790
rect 5873 1796 5902 1804
rect 5873 1790 5890 1796
rect 5873 1788 5907 1790
rect 5955 1788 5971 1804
rect 5972 1794 6180 1804
rect 6181 1794 6197 1804
rect 6245 1800 6260 1815
rect 6263 1812 6264 1824
rect 6271 1812 6298 1824
rect 6263 1804 6298 1812
rect 6263 1803 6292 1804
rect 5983 1790 6197 1794
rect 5998 1788 6197 1790
rect 6232 1790 6245 1800
rect 6263 1790 6280 1803
rect 6232 1788 6280 1790
rect 5874 1784 5907 1788
rect 5870 1782 5907 1784
rect 5870 1781 5937 1782
rect 5870 1776 5901 1781
rect 5907 1776 5937 1781
rect 5870 1772 5937 1776
rect 5843 1769 5937 1772
rect 5843 1762 5892 1769
rect 5843 1756 5873 1762
rect 5892 1757 5897 1762
rect 5809 1740 5889 1756
rect 5901 1748 5937 1769
rect 5998 1764 6187 1788
rect 6232 1787 6279 1788
rect 6245 1782 6279 1787
rect 6013 1761 6187 1764
rect 6006 1758 6187 1761
rect 6215 1781 6279 1782
rect 5809 1738 5828 1740
rect 5843 1738 5877 1740
rect 5809 1722 5889 1738
rect 5809 1716 5828 1722
rect 5525 1690 5628 1700
rect 5479 1688 5628 1690
rect 5649 1688 5684 1700
rect 5318 1686 5480 1688
rect 5330 1666 5349 1686
rect 5364 1684 5394 1686
rect 5213 1658 5254 1666
rect 5336 1662 5349 1666
rect 5401 1670 5480 1686
rect 5512 1686 5684 1688
rect 5512 1670 5591 1686
rect 5598 1684 5628 1686
rect 5176 1648 5205 1658
rect 5219 1648 5248 1658
rect 5263 1648 5293 1662
rect 5336 1648 5379 1662
rect 5401 1658 5591 1670
rect 5656 1666 5662 1686
rect 5386 1648 5416 1658
rect 5417 1648 5575 1658
rect 5579 1648 5609 1658
rect 5613 1648 5643 1662
rect 5671 1648 5684 1686
rect 5756 1700 5785 1716
rect 5799 1700 5828 1716
rect 5843 1706 5873 1722
rect 5901 1700 5907 1748
rect 5910 1742 5929 1748
rect 5944 1742 5974 1750
rect 5910 1734 5974 1742
rect 5910 1718 5990 1734
rect 6006 1727 6068 1758
rect 6084 1727 6146 1758
rect 6215 1756 6264 1781
rect 6279 1756 6309 1772
rect 6178 1742 6208 1750
rect 6215 1748 6325 1756
rect 6178 1734 6223 1742
rect 5910 1716 5929 1718
rect 5944 1716 5990 1718
rect 5910 1700 5990 1716
rect 6017 1714 6052 1727
rect 6093 1724 6130 1727
rect 6093 1722 6135 1724
rect 6022 1711 6052 1714
rect 6031 1707 6038 1711
rect 6038 1706 6039 1707
rect 5997 1700 6007 1706
rect 5756 1692 5791 1700
rect 5756 1666 5757 1692
rect 5764 1666 5791 1692
rect 5699 1648 5729 1662
rect 5756 1658 5791 1666
rect 5793 1692 5834 1700
rect 5793 1666 5808 1692
rect 5815 1666 5834 1692
rect 5898 1688 5929 1700
rect 5944 1688 6047 1700
rect 6059 1690 6085 1716
rect 6100 1711 6130 1722
rect 6162 1718 6224 1734
rect 6162 1716 6208 1718
rect 6162 1700 6224 1716
rect 6236 1700 6242 1748
rect 6245 1740 6325 1748
rect 6245 1738 6264 1740
rect 6279 1738 6313 1740
rect 6245 1722 6325 1738
rect 6245 1700 6264 1722
rect 6279 1706 6309 1722
rect 6337 1716 6343 1790
rect 6346 1716 6365 1860
rect 6380 1716 6386 1860
rect 6395 1790 6408 1860
rect 6460 1856 6482 1860
rect 6453 1834 6482 1848
rect 6535 1834 6551 1848
rect 6589 1844 6595 1846
rect 6602 1844 6710 1860
rect 6717 1844 6723 1846
rect 6731 1844 6746 1860
rect 6812 1854 6831 1857
rect 6453 1832 6551 1834
rect 6578 1832 6746 1844
rect 6761 1834 6777 1848
rect 6812 1835 6834 1854
rect 6844 1848 6860 1849
rect 6843 1846 6860 1848
rect 6844 1841 6860 1846
rect 6834 1834 6840 1835
rect 6843 1834 6872 1841
rect 6761 1833 6872 1834
rect 6761 1832 6878 1833
rect 6437 1824 6488 1832
rect 6535 1824 6569 1832
rect 6437 1812 6462 1824
rect 6469 1812 6488 1824
rect 6542 1822 6569 1824
rect 6578 1822 6799 1832
rect 6834 1829 6840 1832
rect 6542 1818 6799 1822
rect 6437 1804 6488 1812
rect 6535 1804 6799 1818
rect 6843 1824 6878 1832
rect 6389 1756 6408 1790
rect 6453 1796 6482 1804
rect 6453 1790 6470 1796
rect 6453 1788 6487 1790
rect 6535 1788 6551 1804
rect 6552 1794 6760 1804
rect 6761 1794 6777 1804
rect 6825 1800 6840 1815
rect 6843 1812 6844 1824
rect 6851 1812 6878 1824
rect 6843 1804 6878 1812
rect 6843 1803 6872 1804
rect 6563 1790 6777 1794
rect 6578 1788 6777 1790
rect 6812 1790 6825 1800
rect 6843 1790 6860 1803
rect 6812 1788 6860 1790
rect 6454 1784 6487 1788
rect 6450 1782 6487 1784
rect 6450 1781 6517 1782
rect 6450 1776 6481 1781
rect 6487 1776 6517 1781
rect 6450 1772 6517 1776
rect 6423 1769 6517 1772
rect 6423 1762 6472 1769
rect 6423 1756 6453 1762
rect 6472 1757 6477 1762
rect 6389 1740 6469 1756
rect 6481 1748 6517 1769
rect 6578 1764 6767 1788
rect 6812 1787 6859 1788
rect 6825 1782 6859 1787
rect 6593 1761 6767 1764
rect 6586 1758 6767 1761
rect 6795 1781 6859 1782
rect 6389 1738 6408 1740
rect 6423 1738 6457 1740
rect 6389 1722 6469 1738
rect 6389 1716 6408 1722
rect 6105 1690 6208 1700
rect 6059 1688 6208 1690
rect 6229 1688 6264 1700
rect 5898 1686 6060 1688
rect 5910 1666 5929 1686
rect 5944 1684 5974 1686
rect 5793 1658 5834 1666
rect 5916 1662 5929 1666
rect 5981 1670 6060 1686
rect 6092 1686 6264 1688
rect 6092 1670 6171 1686
rect 6178 1684 6208 1686
rect 5756 1648 5785 1658
rect 5799 1648 5828 1658
rect 5843 1648 5873 1662
rect 5916 1648 5959 1662
rect 5981 1658 6171 1670
rect 6236 1666 6242 1686
rect 5966 1648 5996 1658
rect 5997 1648 6155 1658
rect 6159 1648 6189 1658
rect 6193 1648 6223 1662
rect 6251 1648 6264 1686
rect 6336 1700 6365 1716
rect 6379 1700 6408 1716
rect 6423 1706 6453 1722
rect 6481 1700 6487 1748
rect 6490 1742 6509 1748
rect 6524 1742 6554 1750
rect 6490 1734 6554 1742
rect 6490 1718 6570 1734
rect 6586 1727 6648 1758
rect 6664 1727 6726 1758
rect 6795 1756 6844 1781
rect 6859 1756 6889 1772
rect 6758 1742 6788 1750
rect 6795 1748 6905 1756
rect 6758 1734 6803 1742
rect 6490 1716 6509 1718
rect 6524 1716 6570 1718
rect 6490 1700 6570 1716
rect 6597 1714 6632 1727
rect 6673 1724 6710 1727
rect 6673 1722 6715 1724
rect 6602 1711 6632 1714
rect 6611 1707 6618 1711
rect 6618 1706 6619 1707
rect 6577 1700 6587 1706
rect 6336 1692 6371 1700
rect 6336 1666 6337 1692
rect 6344 1666 6371 1692
rect 6279 1648 6309 1662
rect 6336 1658 6371 1666
rect 6373 1692 6414 1700
rect 6373 1666 6388 1692
rect 6395 1666 6414 1692
rect 6478 1688 6509 1700
rect 6524 1688 6627 1700
rect 6639 1690 6665 1716
rect 6680 1711 6710 1722
rect 6742 1718 6804 1734
rect 6742 1716 6788 1718
rect 6742 1700 6804 1716
rect 6816 1700 6822 1748
rect 6825 1740 6905 1748
rect 6825 1738 6844 1740
rect 6859 1738 6893 1740
rect 6825 1722 6905 1738
rect 6825 1700 6844 1722
rect 6859 1706 6889 1722
rect 6917 1716 6923 1790
rect 6926 1716 6945 1860
rect 6960 1716 6966 1860
rect 6975 1790 6988 1860
rect 7040 1856 7062 1860
rect 7033 1834 7062 1848
rect 7115 1834 7131 1848
rect 7169 1844 7175 1846
rect 7182 1844 7290 1860
rect 7297 1844 7303 1846
rect 7311 1844 7326 1860
rect 7392 1854 7411 1857
rect 7033 1832 7131 1834
rect 7158 1832 7326 1844
rect 7341 1834 7357 1848
rect 7392 1835 7414 1854
rect 7424 1848 7440 1849
rect 7423 1846 7440 1848
rect 7424 1841 7440 1846
rect 7414 1834 7420 1835
rect 7423 1834 7452 1841
rect 7341 1833 7452 1834
rect 7341 1832 7458 1833
rect 7017 1824 7068 1832
rect 7115 1824 7149 1832
rect 7017 1812 7042 1824
rect 7049 1812 7068 1824
rect 7122 1822 7149 1824
rect 7158 1822 7379 1832
rect 7414 1829 7420 1832
rect 7122 1818 7379 1822
rect 7017 1804 7068 1812
rect 7115 1804 7379 1818
rect 7423 1824 7458 1832
rect 6969 1756 6988 1790
rect 7033 1796 7062 1804
rect 7033 1790 7050 1796
rect 7033 1788 7067 1790
rect 7115 1788 7131 1804
rect 7132 1794 7340 1804
rect 7341 1794 7357 1804
rect 7405 1800 7420 1815
rect 7423 1812 7424 1824
rect 7431 1812 7458 1824
rect 7423 1804 7458 1812
rect 7423 1803 7452 1804
rect 7151 1790 7357 1794
rect 7158 1788 7357 1790
rect 7392 1790 7405 1800
rect 7423 1790 7440 1803
rect 7392 1788 7440 1790
rect 7034 1784 7067 1788
rect 7030 1782 7067 1784
rect 7030 1781 7097 1782
rect 7030 1776 7061 1781
rect 7067 1776 7097 1781
rect 7030 1772 7097 1776
rect 7003 1769 7097 1772
rect 7003 1762 7052 1769
rect 7003 1756 7033 1762
rect 7052 1757 7057 1762
rect 6969 1740 7049 1756
rect 7061 1748 7097 1769
rect 7158 1764 7347 1788
rect 7392 1787 7439 1788
rect 7405 1782 7439 1787
rect 7173 1761 7347 1764
rect 7166 1758 7347 1761
rect 7375 1781 7439 1782
rect 6969 1738 6988 1740
rect 7003 1738 7037 1740
rect 6969 1722 7049 1738
rect 6969 1716 6988 1722
rect 6685 1690 6788 1700
rect 6639 1688 6788 1690
rect 6809 1688 6844 1700
rect 6478 1686 6640 1688
rect 6490 1666 6509 1686
rect 6524 1684 6554 1686
rect 6373 1658 6414 1666
rect 6496 1662 6509 1666
rect 6561 1670 6640 1686
rect 6672 1686 6844 1688
rect 6672 1670 6751 1686
rect 6758 1684 6788 1686
rect 6336 1648 6365 1658
rect 6379 1648 6408 1658
rect 6423 1648 6453 1662
rect 6496 1648 6539 1662
rect 6561 1658 6751 1670
rect 6816 1666 6822 1686
rect 6546 1648 6576 1658
rect 6577 1648 6735 1658
rect 6739 1648 6769 1658
rect 6773 1648 6803 1662
rect 6831 1648 6844 1686
rect 6916 1700 6945 1716
rect 6959 1700 6988 1716
rect 7003 1706 7033 1722
rect 7061 1700 7067 1748
rect 7070 1742 7089 1748
rect 7104 1742 7134 1750
rect 7070 1734 7134 1742
rect 7070 1718 7150 1734
rect 7166 1727 7228 1758
rect 7244 1727 7306 1758
rect 7375 1756 7424 1781
rect 7439 1756 7469 1772
rect 7338 1742 7368 1750
rect 7375 1748 7485 1756
rect 7338 1734 7383 1742
rect 7070 1716 7089 1718
rect 7104 1716 7150 1718
rect 7070 1700 7150 1716
rect 7177 1714 7212 1727
rect 7253 1724 7290 1727
rect 7253 1722 7295 1724
rect 7182 1711 7212 1714
rect 7191 1707 7198 1711
rect 7198 1706 7199 1707
rect 7157 1700 7167 1706
rect 6916 1692 6951 1700
rect 6916 1666 6917 1692
rect 6924 1666 6951 1692
rect 6859 1648 6889 1662
rect 6916 1658 6951 1666
rect 6953 1692 6994 1700
rect 6953 1666 6968 1692
rect 6975 1666 6994 1692
rect 7058 1688 7089 1700
rect 7104 1688 7207 1700
rect 7219 1690 7245 1716
rect 7260 1711 7290 1722
rect 7322 1718 7384 1734
rect 7322 1716 7368 1718
rect 7322 1700 7384 1716
rect 7396 1700 7402 1748
rect 7405 1740 7485 1748
rect 7405 1738 7424 1740
rect 7439 1738 7473 1740
rect 7405 1722 7485 1738
rect 7405 1700 7424 1722
rect 7439 1706 7469 1722
rect 7497 1716 7503 1790
rect 7506 1716 7525 1860
rect 7540 1716 7546 1860
rect 7555 1790 7568 1860
rect 7620 1856 7642 1860
rect 7613 1834 7642 1848
rect 7695 1834 7711 1848
rect 7749 1844 7755 1846
rect 7762 1844 7870 1860
rect 7877 1844 7883 1846
rect 7891 1844 7906 1860
rect 7972 1854 7991 1857
rect 7613 1832 7711 1834
rect 7738 1832 7906 1844
rect 7921 1834 7937 1848
rect 7972 1835 7994 1854
rect 8004 1848 8020 1849
rect 8003 1846 8020 1848
rect 8004 1841 8020 1846
rect 7994 1834 8000 1835
rect 8003 1834 8032 1841
rect 7921 1833 8032 1834
rect 7921 1832 8038 1833
rect 7597 1824 7648 1832
rect 7695 1824 7729 1832
rect 7597 1812 7622 1824
rect 7629 1812 7648 1824
rect 7702 1822 7729 1824
rect 7738 1822 7959 1832
rect 7994 1829 8000 1832
rect 7702 1818 7959 1822
rect 7597 1804 7648 1812
rect 7695 1804 7959 1818
rect 8003 1824 8038 1832
rect 7549 1756 7568 1790
rect 7613 1796 7642 1804
rect 7613 1790 7630 1796
rect 7613 1788 7647 1790
rect 7695 1788 7711 1804
rect 7712 1794 7920 1804
rect 7921 1794 7937 1804
rect 7985 1800 8000 1815
rect 8003 1812 8004 1824
rect 8011 1812 8038 1824
rect 8003 1804 8038 1812
rect 8003 1803 8032 1804
rect 7723 1790 7937 1794
rect 7738 1788 7937 1790
rect 7972 1790 7985 1800
rect 8003 1790 8020 1803
rect 7972 1788 8020 1790
rect 7614 1784 7647 1788
rect 7610 1782 7647 1784
rect 7610 1781 7677 1782
rect 7610 1776 7641 1781
rect 7647 1776 7677 1781
rect 7610 1772 7677 1776
rect 7583 1769 7677 1772
rect 7583 1762 7632 1769
rect 7583 1756 7613 1762
rect 7632 1757 7637 1762
rect 7549 1740 7629 1756
rect 7641 1748 7677 1769
rect 7738 1764 7927 1788
rect 7972 1787 8019 1788
rect 7985 1782 8019 1787
rect 7753 1761 7927 1764
rect 7746 1758 7927 1761
rect 7955 1781 8019 1782
rect 7549 1738 7568 1740
rect 7583 1738 7617 1740
rect 7549 1722 7629 1738
rect 7549 1716 7568 1722
rect 7265 1690 7368 1700
rect 7219 1688 7368 1690
rect 7389 1688 7424 1700
rect 7058 1686 7220 1688
rect 7070 1666 7089 1686
rect 7104 1684 7134 1686
rect 6953 1658 6994 1666
rect 7076 1662 7089 1666
rect 7141 1670 7220 1686
rect 7252 1686 7424 1688
rect 7252 1670 7331 1686
rect 7338 1684 7368 1686
rect 6916 1648 6945 1658
rect 6959 1648 6988 1658
rect 7003 1648 7033 1662
rect 7076 1648 7119 1662
rect 7141 1658 7331 1670
rect 7396 1666 7402 1686
rect 7126 1648 7156 1658
rect 7157 1648 7315 1658
rect 7319 1648 7349 1658
rect 7353 1648 7383 1662
rect 7411 1648 7424 1686
rect 7496 1700 7525 1716
rect 7539 1700 7568 1716
rect 7583 1706 7613 1722
rect 7641 1700 7647 1748
rect 7650 1742 7669 1748
rect 7684 1742 7714 1750
rect 7650 1734 7714 1742
rect 7650 1718 7730 1734
rect 7746 1727 7808 1758
rect 7824 1727 7886 1758
rect 7955 1756 8004 1781
rect 8019 1756 8049 1772
rect 7918 1742 7948 1750
rect 7955 1748 8065 1756
rect 7918 1734 7963 1742
rect 7650 1716 7669 1718
rect 7684 1716 7730 1718
rect 7650 1700 7730 1716
rect 7757 1714 7792 1727
rect 7833 1724 7870 1727
rect 7833 1722 7875 1724
rect 7762 1711 7792 1714
rect 7771 1707 7778 1711
rect 7778 1706 7779 1707
rect 7737 1700 7747 1706
rect 7496 1692 7531 1700
rect 7496 1666 7497 1692
rect 7504 1666 7531 1692
rect 7439 1648 7469 1662
rect 7496 1658 7531 1666
rect 7533 1692 7574 1700
rect 7533 1666 7548 1692
rect 7555 1666 7574 1692
rect 7638 1688 7669 1700
rect 7684 1688 7787 1700
rect 7799 1690 7825 1716
rect 7840 1711 7870 1722
rect 7902 1718 7964 1734
rect 7902 1716 7948 1718
rect 7902 1700 7964 1716
rect 7976 1700 7982 1748
rect 7985 1740 8065 1748
rect 7985 1738 8004 1740
rect 8019 1738 8053 1740
rect 7985 1722 8065 1738
rect 7985 1700 8004 1722
rect 8019 1706 8049 1722
rect 8077 1716 8083 1790
rect 8086 1716 8105 1860
rect 8120 1716 8126 1860
rect 8135 1790 8148 1860
rect 8200 1856 8222 1860
rect 8193 1834 8222 1848
rect 8275 1834 8291 1848
rect 8329 1844 8335 1846
rect 8342 1844 8450 1860
rect 8457 1844 8463 1846
rect 8471 1844 8486 1860
rect 8552 1854 8571 1857
rect 8193 1832 8291 1834
rect 8318 1832 8486 1844
rect 8501 1834 8517 1848
rect 8552 1835 8574 1854
rect 8584 1848 8600 1849
rect 8583 1846 8600 1848
rect 8584 1841 8600 1846
rect 8574 1834 8580 1835
rect 8583 1834 8612 1841
rect 8501 1833 8612 1834
rect 8501 1832 8618 1833
rect 8177 1824 8228 1832
rect 8275 1824 8309 1832
rect 8177 1812 8202 1824
rect 8209 1812 8228 1824
rect 8282 1822 8309 1824
rect 8318 1822 8539 1832
rect 8574 1829 8580 1832
rect 8282 1818 8539 1822
rect 8177 1804 8228 1812
rect 8275 1804 8539 1818
rect 8583 1824 8618 1832
rect 8129 1756 8148 1790
rect 8193 1796 8222 1804
rect 8193 1790 8210 1796
rect 8193 1788 8227 1790
rect 8275 1788 8291 1804
rect 8292 1794 8500 1804
rect 8501 1794 8517 1804
rect 8565 1800 8580 1815
rect 8583 1812 8584 1824
rect 8591 1812 8618 1824
rect 8583 1804 8618 1812
rect 8583 1803 8612 1804
rect 8303 1790 8517 1794
rect 8318 1788 8517 1790
rect 8552 1790 8565 1800
rect 8583 1790 8600 1803
rect 8552 1788 8600 1790
rect 8194 1784 8227 1788
rect 8190 1782 8227 1784
rect 8190 1781 8257 1782
rect 8190 1776 8221 1781
rect 8227 1776 8257 1781
rect 8190 1772 8257 1776
rect 8163 1769 8257 1772
rect 8163 1762 8212 1769
rect 8163 1756 8193 1762
rect 8212 1757 8217 1762
rect 8129 1740 8209 1756
rect 8221 1748 8257 1769
rect 8318 1764 8507 1788
rect 8552 1787 8599 1788
rect 8565 1782 8599 1787
rect 8333 1761 8507 1764
rect 8326 1758 8507 1761
rect 8535 1781 8599 1782
rect 8129 1738 8148 1740
rect 8163 1738 8197 1740
rect 8129 1722 8209 1738
rect 8129 1716 8148 1722
rect 7845 1690 7948 1700
rect 7799 1688 7948 1690
rect 7969 1688 8004 1700
rect 7638 1686 7800 1688
rect 7650 1666 7669 1686
rect 7684 1684 7714 1686
rect 7533 1658 7574 1666
rect 7656 1662 7669 1666
rect 7721 1670 7800 1686
rect 7832 1686 8004 1688
rect 7832 1670 7911 1686
rect 7918 1684 7948 1686
rect 7496 1648 7525 1658
rect 7539 1648 7568 1658
rect 7583 1648 7613 1662
rect 7656 1648 7699 1662
rect 7721 1658 7911 1670
rect 7976 1666 7982 1686
rect 7706 1648 7736 1658
rect 7737 1648 7895 1658
rect 7899 1648 7929 1658
rect 7933 1648 7963 1662
rect 7991 1648 8004 1686
rect 8076 1700 8105 1716
rect 8119 1700 8148 1716
rect 8163 1706 8193 1722
rect 8221 1700 8227 1748
rect 8230 1742 8249 1748
rect 8264 1742 8294 1750
rect 8230 1734 8294 1742
rect 8230 1718 8310 1734
rect 8326 1727 8388 1758
rect 8404 1727 8466 1758
rect 8535 1756 8584 1781
rect 8599 1756 8629 1772
rect 8498 1742 8528 1750
rect 8535 1748 8645 1756
rect 8498 1734 8543 1742
rect 8230 1716 8249 1718
rect 8264 1716 8310 1718
rect 8230 1700 8310 1716
rect 8337 1714 8372 1727
rect 8413 1724 8450 1727
rect 8413 1722 8455 1724
rect 8342 1711 8372 1714
rect 8351 1707 8358 1711
rect 8358 1706 8359 1707
rect 8317 1700 8327 1706
rect 8076 1692 8111 1700
rect 8076 1666 8077 1692
rect 8084 1666 8111 1692
rect 8019 1648 8049 1662
rect 8076 1658 8111 1666
rect 8113 1692 8154 1700
rect 8113 1666 8128 1692
rect 8135 1666 8154 1692
rect 8218 1688 8249 1700
rect 8264 1688 8367 1700
rect 8379 1690 8405 1716
rect 8420 1711 8450 1722
rect 8482 1718 8544 1734
rect 8482 1716 8528 1718
rect 8482 1700 8544 1716
rect 8556 1700 8562 1748
rect 8565 1740 8645 1748
rect 8565 1738 8584 1740
rect 8599 1738 8633 1740
rect 8565 1722 8645 1738
rect 8565 1700 8584 1722
rect 8599 1706 8629 1722
rect 8657 1716 8663 1790
rect 8666 1716 8685 1860
rect 8700 1716 8706 1860
rect 8715 1790 8728 1860
rect 8780 1856 8802 1860
rect 8773 1834 8802 1848
rect 8855 1834 8871 1848
rect 8909 1844 8915 1846
rect 8922 1844 9030 1860
rect 9037 1844 9043 1846
rect 9051 1844 9066 1860
rect 9132 1854 9151 1857
rect 8773 1832 8871 1834
rect 8898 1832 9066 1844
rect 9081 1834 9097 1848
rect 9132 1835 9154 1854
rect 9164 1848 9180 1849
rect 9163 1846 9180 1848
rect 9164 1841 9180 1846
rect 9154 1834 9160 1835
rect 9163 1834 9192 1841
rect 9081 1833 9192 1834
rect 9081 1832 9198 1833
rect 8757 1824 8808 1832
rect 8855 1824 8889 1832
rect 8757 1812 8782 1824
rect 8789 1812 8808 1824
rect 8862 1822 8889 1824
rect 8898 1822 9119 1832
rect 9154 1829 9160 1832
rect 8862 1818 9119 1822
rect 8757 1804 8808 1812
rect 8855 1804 9119 1818
rect 9163 1824 9198 1832
rect 8709 1756 8728 1790
rect 8773 1796 8802 1804
rect 8773 1790 8790 1796
rect 8773 1788 8807 1790
rect 8855 1788 8871 1804
rect 8872 1794 9080 1804
rect 9081 1794 9097 1804
rect 9145 1800 9160 1815
rect 9163 1812 9164 1824
rect 9171 1812 9198 1824
rect 9163 1804 9198 1812
rect 9163 1803 9192 1804
rect 8883 1790 9097 1794
rect 8898 1788 9097 1790
rect 9132 1790 9145 1800
rect 9163 1790 9180 1803
rect 9132 1788 9180 1790
rect 8774 1784 8807 1788
rect 8770 1782 8807 1784
rect 8770 1781 8837 1782
rect 8770 1776 8801 1781
rect 8807 1776 8837 1781
rect 8770 1772 8837 1776
rect 8743 1769 8837 1772
rect 8743 1762 8792 1769
rect 8743 1756 8773 1762
rect 8792 1757 8797 1762
rect 8709 1740 8789 1756
rect 8801 1748 8837 1769
rect 8898 1764 9087 1788
rect 9132 1787 9179 1788
rect 9145 1782 9179 1787
rect 8913 1761 9087 1764
rect 8906 1758 9087 1761
rect 9115 1781 9179 1782
rect 8709 1738 8728 1740
rect 8743 1738 8777 1740
rect 8709 1722 8789 1738
rect 8709 1716 8728 1722
rect 8425 1690 8528 1700
rect 8379 1688 8528 1690
rect 8549 1688 8584 1700
rect 8218 1686 8380 1688
rect 8230 1666 8249 1686
rect 8264 1684 8294 1686
rect 8113 1658 8154 1666
rect 8236 1662 8249 1666
rect 8301 1670 8380 1686
rect 8412 1686 8584 1688
rect 8412 1670 8491 1686
rect 8498 1684 8528 1686
rect 8076 1648 8105 1658
rect 8119 1648 8148 1658
rect 8163 1648 8193 1662
rect 8236 1648 8279 1662
rect 8301 1658 8491 1670
rect 8556 1666 8562 1686
rect 8286 1648 8316 1658
rect 8317 1648 8475 1658
rect 8479 1648 8509 1658
rect 8513 1648 8543 1662
rect 8571 1648 8584 1686
rect 8656 1700 8685 1716
rect 8699 1700 8728 1716
rect 8743 1706 8773 1722
rect 8801 1700 8807 1748
rect 8810 1742 8829 1748
rect 8844 1742 8874 1750
rect 8810 1734 8874 1742
rect 8810 1718 8890 1734
rect 8906 1727 8968 1758
rect 8984 1727 9046 1758
rect 9115 1756 9164 1781
rect 9179 1756 9209 1772
rect 9078 1742 9108 1750
rect 9115 1748 9225 1756
rect 9078 1734 9123 1742
rect 8810 1716 8829 1718
rect 8844 1716 8890 1718
rect 8810 1700 8890 1716
rect 8917 1714 8952 1727
rect 8993 1724 9030 1727
rect 8993 1722 9035 1724
rect 8922 1711 8952 1714
rect 8931 1707 8938 1711
rect 8938 1706 8939 1707
rect 8897 1700 8907 1706
rect 8656 1692 8691 1700
rect 8656 1666 8657 1692
rect 8664 1666 8691 1692
rect 8599 1648 8629 1662
rect 8656 1658 8691 1666
rect 8693 1692 8734 1700
rect 8693 1666 8708 1692
rect 8715 1666 8734 1692
rect 8798 1688 8829 1700
rect 8844 1688 8947 1700
rect 8959 1690 8985 1716
rect 9000 1711 9030 1722
rect 9062 1718 9124 1734
rect 9062 1716 9108 1718
rect 9062 1700 9124 1716
rect 9136 1700 9142 1748
rect 9145 1740 9225 1748
rect 9145 1738 9164 1740
rect 9179 1738 9213 1740
rect 9145 1722 9225 1738
rect 9145 1700 9164 1722
rect 9179 1706 9209 1722
rect 9237 1716 9243 1790
rect 9246 1716 9265 1860
rect 9280 1716 9286 1860
rect 9295 1790 9308 1860
rect 9360 1856 9382 1860
rect 9353 1834 9382 1848
rect 9435 1834 9451 1848
rect 9489 1844 9495 1846
rect 9502 1844 9610 1860
rect 9617 1844 9623 1846
rect 9631 1844 9646 1860
rect 9712 1854 9731 1857
rect 9353 1832 9451 1834
rect 9478 1832 9646 1844
rect 9661 1834 9677 1848
rect 9712 1835 9734 1854
rect 9744 1848 9760 1849
rect 9743 1846 9760 1848
rect 9744 1841 9760 1846
rect 9734 1834 9740 1835
rect 9743 1834 9772 1841
rect 9661 1833 9772 1834
rect 9661 1832 9778 1833
rect 9337 1824 9388 1832
rect 9435 1824 9469 1832
rect 9337 1812 9362 1824
rect 9369 1812 9388 1824
rect 9442 1822 9469 1824
rect 9478 1822 9699 1832
rect 9734 1829 9740 1832
rect 9442 1818 9699 1822
rect 9337 1804 9388 1812
rect 9435 1804 9699 1818
rect 9743 1824 9778 1832
rect 9289 1756 9308 1790
rect 9353 1796 9382 1804
rect 9353 1790 9370 1796
rect 9353 1788 9387 1790
rect 9435 1788 9451 1804
rect 9452 1794 9660 1804
rect 9661 1794 9677 1804
rect 9725 1800 9740 1815
rect 9743 1812 9744 1824
rect 9751 1812 9778 1824
rect 9743 1804 9778 1812
rect 9743 1803 9772 1804
rect 9463 1790 9677 1794
rect 9478 1788 9677 1790
rect 9712 1790 9725 1800
rect 9743 1790 9760 1803
rect 9712 1788 9760 1790
rect 9354 1784 9387 1788
rect 9350 1782 9387 1784
rect 9350 1781 9417 1782
rect 9350 1776 9381 1781
rect 9387 1776 9417 1781
rect 9350 1772 9417 1776
rect 9323 1769 9417 1772
rect 9323 1762 9372 1769
rect 9323 1756 9353 1762
rect 9372 1757 9377 1762
rect 9289 1740 9369 1756
rect 9381 1748 9417 1769
rect 9478 1764 9667 1788
rect 9712 1787 9759 1788
rect 9725 1782 9759 1787
rect 9493 1761 9667 1764
rect 9486 1758 9667 1761
rect 9695 1781 9759 1782
rect 9289 1738 9308 1740
rect 9323 1738 9357 1740
rect 9289 1722 9369 1738
rect 9289 1716 9308 1722
rect 9005 1690 9108 1700
rect 8959 1688 9108 1690
rect 9129 1688 9164 1700
rect 8798 1686 8960 1688
rect 8810 1666 8829 1686
rect 8844 1684 8874 1686
rect 8693 1658 8734 1666
rect 8816 1662 8829 1666
rect 8881 1670 8960 1686
rect 8992 1686 9164 1688
rect 8992 1670 9071 1686
rect 9078 1684 9108 1686
rect 8656 1648 8685 1658
rect 8699 1648 8728 1658
rect 8743 1648 8773 1662
rect 8816 1648 8859 1662
rect 8881 1658 9071 1670
rect 9136 1666 9142 1686
rect 8866 1648 8896 1658
rect 8897 1648 9055 1658
rect 9059 1648 9089 1658
rect 9093 1648 9123 1662
rect 9151 1648 9164 1686
rect 9236 1700 9265 1716
rect 9279 1700 9308 1716
rect 9323 1706 9353 1722
rect 9381 1700 9387 1748
rect 9390 1742 9409 1748
rect 9424 1742 9454 1750
rect 9390 1734 9454 1742
rect 9390 1718 9470 1734
rect 9486 1727 9548 1758
rect 9564 1727 9626 1758
rect 9695 1756 9744 1781
rect 9759 1756 9789 1772
rect 9658 1742 9688 1750
rect 9695 1748 9805 1756
rect 9658 1734 9703 1742
rect 9390 1716 9409 1718
rect 9424 1716 9470 1718
rect 9390 1700 9470 1716
rect 9497 1714 9532 1727
rect 9573 1724 9610 1727
rect 9573 1722 9615 1724
rect 9502 1711 9532 1714
rect 9511 1707 9518 1711
rect 9518 1706 9519 1707
rect 9477 1700 9487 1706
rect 9236 1692 9271 1700
rect 9236 1666 9237 1692
rect 9244 1666 9271 1692
rect 9179 1648 9209 1662
rect 9236 1658 9271 1666
rect 9273 1692 9314 1700
rect 9273 1666 9288 1692
rect 9295 1666 9314 1692
rect 9378 1688 9409 1700
rect 9424 1688 9527 1700
rect 9539 1690 9565 1716
rect 9580 1711 9610 1722
rect 9642 1718 9704 1734
rect 9642 1716 9688 1718
rect 9642 1700 9704 1716
rect 9716 1700 9722 1748
rect 9725 1740 9805 1748
rect 9725 1738 9744 1740
rect 9759 1738 9793 1740
rect 9725 1722 9805 1738
rect 9725 1700 9744 1722
rect 9759 1706 9789 1722
rect 9817 1716 9823 1790
rect 9826 1716 9845 1860
rect 9860 1716 9866 1860
rect 9875 1790 9888 1860
rect 9940 1856 9962 1860
rect 9933 1834 9962 1848
rect 10015 1834 10031 1848
rect 10069 1844 10075 1846
rect 10082 1844 10190 1860
rect 10197 1844 10203 1846
rect 10211 1844 10226 1860
rect 10292 1854 10311 1857
rect 9933 1832 10031 1834
rect 10058 1832 10226 1844
rect 10241 1834 10257 1848
rect 10292 1835 10314 1854
rect 10324 1848 10340 1849
rect 10323 1846 10340 1848
rect 10324 1841 10340 1846
rect 10314 1834 10320 1835
rect 10323 1834 10352 1841
rect 10241 1833 10352 1834
rect 10241 1832 10358 1833
rect 9917 1824 9968 1832
rect 10015 1824 10049 1832
rect 9917 1812 9942 1824
rect 9949 1812 9968 1824
rect 10022 1822 10049 1824
rect 10058 1822 10279 1832
rect 10314 1829 10320 1832
rect 10022 1818 10279 1822
rect 9917 1804 9968 1812
rect 10015 1804 10279 1818
rect 10323 1824 10358 1832
rect 9869 1756 9888 1790
rect 9933 1796 9962 1804
rect 9933 1790 9950 1796
rect 9933 1788 9967 1790
rect 10015 1788 10031 1804
rect 10032 1794 10240 1804
rect 10241 1794 10257 1804
rect 10305 1800 10320 1815
rect 10323 1812 10324 1824
rect 10331 1812 10358 1824
rect 10323 1804 10358 1812
rect 10323 1803 10352 1804
rect 10043 1790 10257 1794
rect 10058 1788 10257 1790
rect 10292 1790 10305 1800
rect 10323 1790 10340 1803
rect 10292 1788 10340 1790
rect 9934 1784 9967 1788
rect 9930 1782 9967 1784
rect 9930 1781 9997 1782
rect 9930 1776 9961 1781
rect 9967 1776 9997 1781
rect 9930 1772 9997 1776
rect 9903 1769 9997 1772
rect 9903 1762 9952 1769
rect 9903 1756 9933 1762
rect 9952 1757 9957 1762
rect 9869 1740 9949 1756
rect 9961 1748 9997 1769
rect 10058 1764 10247 1788
rect 10292 1787 10339 1788
rect 10305 1782 10339 1787
rect 10073 1761 10247 1764
rect 10066 1758 10247 1761
rect 10275 1781 10339 1782
rect 9869 1738 9888 1740
rect 9903 1738 9937 1740
rect 9869 1722 9949 1738
rect 9869 1716 9888 1722
rect 9585 1690 9688 1700
rect 9539 1688 9688 1690
rect 9709 1688 9744 1700
rect 9378 1686 9540 1688
rect 9390 1666 9409 1686
rect 9424 1684 9454 1686
rect 9273 1658 9314 1666
rect 9396 1662 9409 1666
rect 9461 1670 9540 1686
rect 9572 1686 9744 1688
rect 9572 1670 9651 1686
rect 9658 1684 9688 1686
rect 9236 1648 9265 1658
rect 9279 1648 9308 1658
rect 9323 1648 9353 1662
rect 9396 1648 9439 1662
rect 9461 1658 9651 1670
rect 9716 1666 9722 1686
rect 9446 1648 9476 1658
rect 9477 1648 9635 1658
rect 9639 1648 9669 1658
rect 9673 1648 9703 1662
rect 9731 1648 9744 1686
rect 9816 1700 9845 1716
rect 9859 1700 9888 1716
rect 9903 1706 9933 1722
rect 9961 1700 9967 1748
rect 9970 1742 9989 1748
rect 10004 1742 10034 1750
rect 9970 1734 10034 1742
rect 9970 1718 10050 1734
rect 10066 1727 10128 1758
rect 10144 1727 10206 1758
rect 10275 1756 10324 1781
rect 10339 1756 10369 1772
rect 10238 1742 10268 1750
rect 10275 1748 10385 1756
rect 10238 1734 10283 1742
rect 9970 1716 9989 1718
rect 10004 1716 10050 1718
rect 9970 1700 10050 1716
rect 10077 1714 10112 1727
rect 10153 1724 10190 1727
rect 10153 1722 10195 1724
rect 10082 1711 10112 1714
rect 10091 1707 10098 1711
rect 10098 1706 10099 1707
rect 10057 1700 10067 1706
rect 9816 1692 9851 1700
rect 9816 1666 9817 1692
rect 9824 1666 9851 1692
rect 9759 1648 9789 1662
rect 9816 1658 9851 1666
rect 9853 1692 9894 1700
rect 9853 1666 9868 1692
rect 9875 1666 9894 1692
rect 9958 1688 9989 1700
rect 10004 1688 10107 1700
rect 10119 1690 10145 1716
rect 10160 1711 10190 1722
rect 10222 1718 10284 1734
rect 10222 1716 10268 1718
rect 10222 1700 10284 1716
rect 10296 1700 10302 1748
rect 10305 1740 10385 1748
rect 10305 1738 10324 1740
rect 10339 1738 10373 1740
rect 10305 1722 10385 1738
rect 10305 1700 10324 1722
rect 10339 1706 10369 1722
rect 10397 1716 10403 1790
rect 10406 1716 10425 1860
rect 10440 1716 10446 1860
rect 10455 1790 10468 1860
rect 10520 1856 10542 1860
rect 10513 1834 10542 1848
rect 10595 1834 10611 1848
rect 10649 1844 10655 1846
rect 10662 1844 10770 1860
rect 10777 1844 10783 1846
rect 10791 1844 10806 1860
rect 10872 1854 10891 1857
rect 10513 1832 10611 1834
rect 10638 1832 10806 1844
rect 10821 1834 10837 1848
rect 10872 1835 10894 1854
rect 10904 1848 10920 1849
rect 10903 1846 10920 1848
rect 10904 1841 10920 1846
rect 10894 1834 10900 1835
rect 10903 1834 10932 1841
rect 10821 1833 10932 1834
rect 10821 1832 10938 1833
rect 10497 1824 10548 1832
rect 10595 1824 10629 1832
rect 10497 1812 10522 1824
rect 10529 1812 10548 1824
rect 10602 1822 10629 1824
rect 10638 1822 10859 1832
rect 10894 1829 10900 1832
rect 10602 1818 10859 1822
rect 10497 1804 10548 1812
rect 10595 1804 10859 1818
rect 10903 1824 10938 1832
rect 10449 1756 10468 1790
rect 10513 1796 10542 1804
rect 10513 1790 10530 1796
rect 10513 1788 10547 1790
rect 10595 1788 10611 1804
rect 10612 1794 10820 1804
rect 10821 1794 10837 1804
rect 10885 1800 10900 1815
rect 10903 1812 10904 1824
rect 10911 1812 10938 1824
rect 10903 1804 10938 1812
rect 10903 1803 10932 1804
rect 10623 1790 10837 1794
rect 10638 1788 10837 1790
rect 10872 1790 10885 1800
rect 10903 1790 10920 1803
rect 10872 1788 10920 1790
rect 10514 1784 10547 1788
rect 10510 1782 10547 1784
rect 10510 1781 10577 1782
rect 10510 1776 10541 1781
rect 10547 1776 10577 1781
rect 10510 1772 10577 1776
rect 10483 1769 10577 1772
rect 10483 1762 10532 1769
rect 10483 1756 10513 1762
rect 10532 1757 10537 1762
rect 10449 1740 10529 1756
rect 10541 1748 10577 1769
rect 10638 1764 10827 1788
rect 10872 1787 10919 1788
rect 10885 1782 10919 1787
rect 10653 1761 10827 1764
rect 10646 1758 10827 1761
rect 10855 1781 10919 1782
rect 10449 1738 10468 1740
rect 10483 1738 10517 1740
rect 10449 1722 10529 1738
rect 10449 1716 10468 1722
rect 10165 1690 10268 1700
rect 10119 1688 10268 1690
rect 10289 1688 10324 1700
rect 9958 1686 10120 1688
rect 9970 1666 9989 1686
rect 10004 1684 10034 1686
rect 9853 1658 9894 1666
rect 9976 1662 9989 1666
rect 10041 1670 10120 1686
rect 10152 1686 10324 1688
rect 10152 1670 10231 1686
rect 10238 1684 10268 1686
rect 9816 1648 9845 1658
rect 9859 1648 9888 1658
rect 9903 1648 9933 1662
rect 9976 1648 10019 1662
rect 10041 1658 10231 1670
rect 10296 1666 10302 1686
rect 10026 1648 10056 1658
rect 10057 1648 10215 1658
rect 10219 1648 10249 1658
rect 10253 1648 10283 1662
rect 10311 1648 10324 1686
rect 10396 1700 10425 1716
rect 10439 1700 10468 1716
rect 10483 1706 10513 1722
rect 10541 1700 10547 1748
rect 10550 1742 10569 1748
rect 10584 1742 10614 1750
rect 10550 1734 10614 1742
rect 10550 1718 10630 1734
rect 10646 1727 10708 1758
rect 10724 1727 10786 1758
rect 10855 1756 10904 1781
rect 10919 1756 10949 1772
rect 10818 1742 10848 1750
rect 10855 1748 10965 1756
rect 10818 1734 10863 1742
rect 10550 1716 10569 1718
rect 10584 1716 10630 1718
rect 10550 1700 10630 1716
rect 10657 1714 10692 1727
rect 10733 1724 10770 1727
rect 10733 1722 10775 1724
rect 10662 1711 10692 1714
rect 10671 1707 10678 1711
rect 10678 1706 10679 1707
rect 10637 1700 10647 1706
rect 10396 1692 10431 1700
rect 10396 1666 10397 1692
rect 10404 1666 10431 1692
rect 10339 1648 10369 1662
rect 10396 1658 10431 1666
rect 10433 1692 10474 1700
rect 10433 1666 10448 1692
rect 10455 1666 10474 1692
rect 10538 1688 10569 1700
rect 10584 1688 10687 1700
rect 10699 1690 10725 1716
rect 10740 1711 10770 1722
rect 10802 1718 10864 1734
rect 10802 1716 10848 1718
rect 10802 1700 10864 1716
rect 10876 1700 10882 1748
rect 10885 1740 10965 1748
rect 10885 1738 10904 1740
rect 10919 1738 10953 1740
rect 10885 1722 10965 1738
rect 10885 1700 10904 1722
rect 10919 1706 10949 1722
rect 10977 1716 10983 1790
rect 10986 1716 11005 1860
rect 11020 1716 11026 1860
rect 11035 1790 11048 1860
rect 11100 1856 11122 1860
rect 11093 1834 11122 1848
rect 11175 1834 11191 1848
rect 11229 1844 11235 1846
rect 11242 1844 11350 1860
rect 11357 1844 11363 1846
rect 11371 1844 11386 1860
rect 11452 1854 11471 1857
rect 11093 1832 11191 1834
rect 11218 1832 11386 1844
rect 11401 1834 11417 1848
rect 11452 1835 11474 1854
rect 11484 1848 11500 1849
rect 11483 1846 11500 1848
rect 11484 1841 11500 1846
rect 11474 1834 11480 1835
rect 11483 1834 11512 1841
rect 11401 1833 11512 1834
rect 11401 1832 11518 1833
rect 11077 1824 11128 1832
rect 11175 1824 11209 1832
rect 11077 1812 11102 1824
rect 11109 1812 11128 1824
rect 11182 1822 11209 1824
rect 11218 1822 11439 1832
rect 11474 1829 11480 1832
rect 11182 1818 11439 1822
rect 11077 1804 11128 1812
rect 11175 1804 11439 1818
rect 11483 1824 11518 1832
rect 11029 1756 11048 1790
rect 11093 1796 11122 1804
rect 11093 1790 11110 1796
rect 11093 1788 11127 1790
rect 11175 1788 11191 1804
rect 11192 1794 11400 1804
rect 11401 1794 11417 1804
rect 11465 1800 11480 1815
rect 11483 1812 11484 1824
rect 11491 1812 11518 1824
rect 11483 1804 11518 1812
rect 11483 1803 11512 1804
rect 11203 1790 11417 1794
rect 11218 1788 11417 1790
rect 11452 1790 11465 1800
rect 11483 1790 11500 1803
rect 11452 1788 11500 1790
rect 11094 1784 11127 1788
rect 11090 1782 11127 1784
rect 11090 1781 11157 1782
rect 11090 1776 11121 1781
rect 11127 1776 11157 1781
rect 11090 1772 11157 1776
rect 11063 1769 11157 1772
rect 11063 1762 11112 1769
rect 11063 1756 11093 1762
rect 11112 1757 11117 1762
rect 11029 1740 11109 1756
rect 11121 1748 11157 1769
rect 11218 1764 11407 1788
rect 11452 1787 11499 1788
rect 11465 1782 11499 1787
rect 11233 1761 11407 1764
rect 11226 1758 11407 1761
rect 11435 1781 11499 1782
rect 11029 1738 11048 1740
rect 11063 1738 11097 1740
rect 11029 1722 11109 1738
rect 11029 1716 11048 1722
rect 10745 1690 10848 1700
rect 10699 1688 10848 1690
rect 10869 1688 10904 1700
rect 10538 1686 10700 1688
rect 10550 1666 10569 1686
rect 10584 1684 10614 1686
rect 10433 1658 10474 1666
rect 10556 1662 10569 1666
rect 10621 1670 10700 1686
rect 10732 1686 10904 1688
rect 10732 1670 10811 1686
rect 10818 1684 10848 1686
rect 10396 1648 10425 1658
rect 10439 1648 10468 1658
rect 10483 1648 10513 1662
rect 10556 1648 10599 1662
rect 10621 1658 10811 1670
rect 10876 1666 10882 1686
rect 10606 1648 10636 1658
rect 10637 1648 10795 1658
rect 10799 1648 10829 1658
rect 10833 1648 10863 1662
rect 10891 1648 10904 1686
rect 10976 1700 11005 1716
rect 11019 1700 11048 1716
rect 11063 1706 11093 1722
rect 11121 1700 11127 1748
rect 11130 1742 11149 1748
rect 11164 1742 11194 1750
rect 11130 1734 11194 1742
rect 11130 1718 11210 1734
rect 11226 1727 11288 1758
rect 11304 1727 11366 1758
rect 11435 1756 11484 1781
rect 11499 1756 11529 1772
rect 11398 1742 11428 1750
rect 11435 1748 11545 1756
rect 11398 1734 11443 1742
rect 11130 1716 11149 1718
rect 11164 1716 11210 1718
rect 11130 1700 11210 1716
rect 11237 1714 11272 1727
rect 11313 1724 11350 1727
rect 11313 1722 11355 1724
rect 11242 1711 11272 1714
rect 11251 1707 11258 1711
rect 11258 1706 11259 1707
rect 11217 1700 11227 1706
rect 10976 1692 11011 1700
rect 10976 1666 10977 1692
rect 10984 1666 11011 1692
rect 10919 1648 10949 1662
rect 10976 1658 11011 1666
rect 11013 1692 11054 1700
rect 11013 1666 11028 1692
rect 11035 1666 11054 1692
rect 11118 1688 11149 1700
rect 11164 1688 11267 1700
rect 11279 1690 11305 1716
rect 11320 1711 11350 1722
rect 11382 1718 11444 1734
rect 11382 1716 11428 1718
rect 11382 1700 11444 1716
rect 11456 1700 11462 1748
rect 11465 1740 11545 1748
rect 11465 1738 11484 1740
rect 11499 1738 11533 1740
rect 11465 1722 11545 1738
rect 11465 1700 11484 1722
rect 11499 1706 11529 1722
rect 11557 1716 11563 1790
rect 11566 1716 11585 1860
rect 11600 1716 11606 1860
rect 11615 1790 11628 1860
rect 11680 1856 11702 1860
rect 11673 1834 11702 1848
rect 11755 1834 11771 1848
rect 11809 1844 11815 1846
rect 11822 1844 11930 1860
rect 11937 1844 11943 1846
rect 11951 1844 11966 1860
rect 12032 1854 12051 1857
rect 11673 1832 11771 1834
rect 11798 1832 11966 1844
rect 11981 1834 11997 1848
rect 12032 1835 12054 1854
rect 12064 1848 12080 1849
rect 12063 1846 12080 1848
rect 12064 1841 12080 1846
rect 12054 1834 12060 1835
rect 12063 1834 12092 1841
rect 11981 1833 12092 1834
rect 11981 1832 12098 1833
rect 11657 1824 11708 1832
rect 11755 1824 11789 1832
rect 11657 1812 11682 1824
rect 11689 1812 11708 1824
rect 11762 1822 11789 1824
rect 11798 1822 12019 1832
rect 12054 1829 12060 1832
rect 11762 1818 12019 1822
rect 11657 1804 11708 1812
rect 11755 1804 12019 1818
rect 12063 1824 12098 1832
rect 11609 1756 11628 1790
rect 11673 1796 11702 1804
rect 11673 1790 11690 1796
rect 11673 1788 11707 1790
rect 11755 1788 11771 1804
rect 11772 1794 11980 1804
rect 11981 1794 11997 1804
rect 12045 1800 12060 1815
rect 12063 1812 12064 1824
rect 12071 1812 12098 1824
rect 12063 1804 12098 1812
rect 12063 1803 12092 1804
rect 11783 1790 11997 1794
rect 11798 1788 11997 1790
rect 12032 1790 12045 1800
rect 12063 1790 12080 1803
rect 12032 1788 12080 1790
rect 11674 1784 11707 1788
rect 11670 1782 11707 1784
rect 11670 1781 11737 1782
rect 11670 1776 11701 1781
rect 11707 1776 11737 1781
rect 11670 1772 11737 1776
rect 11643 1769 11737 1772
rect 11643 1762 11692 1769
rect 11643 1756 11673 1762
rect 11692 1757 11697 1762
rect 11609 1740 11689 1756
rect 11701 1748 11737 1769
rect 11798 1764 11987 1788
rect 12032 1787 12079 1788
rect 12045 1782 12079 1787
rect 11813 1761 11987 1764
rect 11806 1758 11987 1761
rect 12015 1781 12079 1782
rect 11609 1738 11628 1740
rect 11643 1738 11677 1740
rect 11609 1722 11689 1738
rect 11609 1716 11628 1722
rect 11325 1690 11428 1700
rect 11279 1688 11428 1690
rect 11449 1688 11484 1700
rect 11118 1686 11280 1688
rect 11130 1666 11149 1686
rect 11164 1684 11194 1686
rect 11013 1658 11054 1666
rect 11136 1662 11149 1666
rect 11201 1670 11280 1686
rect 11312 1686 11484 1688
rect 11312 1670 11391 1686
rect 11398 1684 11428 1686
rect 10976 1648 11005 1658
rect 11019 1648 11048 1658
rect 11063 1648 11093 1662
rect 11136 1648 11179 1662
rect 11201 1658 11391 1670
rect 11456 1666 11462 1686
rect 11186 1648 11216 1658
rect 11217 1648 11375 1658
rect 11379 1648 11409 1658
rect 11413 1648 11443 1662
rect 11471 1648 11484 1686
rect 11556 1700 11585 1716
rect 11599 1700 11628 1716
rect 11643 1706 11673 1722
rect 11701 1700 11707 1748
rect 11710 1742 11729 1748
rect 11744 1742 11774 1750
rect 11710 1734 11774 1742
rect 11710 1718 11790 1734
rect 11806 1727 11868 1758
rect 11884 1727 11946 1758
rect 12015 1756 12064 1781
rect 12079 1756 12109 1772
rect 11978 1742 12008 1750
rect 12015 1748 12125 1756
rect 11978 1734 12023 1742
rect 11710 1716 11729 1718
rect 11744 1716 11790 1718
rect 11710 1700 11790 1716
rect 11817 1714 11852 1727
rect 11893 1724 11930 1727
rect 11893 1722 11935 1724
rect 11822 1711 11852 1714
rect 11831 1707 11838 1711
rect 11838 1706 11839 1707
rect 11797 1700 11807 1706
rect 11556 1692 11591 1700
rect 11556 1666 11557 1692
rect 11564 1666 11591 1692
rect 11499 1648 11529 1662
rect 11556 1658 11591 1666
rect 11593 1692 11634 1700
rect 11593 1666 11608 1692
rect 11615 1666 11634 1692
rect 11698 1688 11729 1700
rect 11744 1688 11847 1700
rect 11859 1690 11885 1716
rect 11900 1711 11930 1722
rect 11962 1718 12024 1734
rect 11962 1716 12008 1718
rect 11962 1700 12024 1716
rect 12036 1700 12042 1748
rect 12045 1740 12125 1748
rect 12045 1738 12064 1740
rect 12079 1738 12113 1740
rect 12045 1722 12125 1738
rect 12045 1700 12064 1722
rect 12079 1706 12109 1722
rect 12137 1716 12143 1790
rect 12146 1716 12165 1860
rect 12180 1716 12186 1860
rect 12195 1790 12208 1860
rect 12260 1856 12282 1860
rect 12253 1834 12282 1848
rect 12335 1834 12351 1848
rect 12389 1844 12395 1846
rect 12402 1844 12510 1860
rect 12517 1844 12523 1846
rect 12531 1844 12546 1860
rect 12612 1854 12631 1857
rect 12253 1832 12351 1834
rect 12378 1832 12546 1844
rect 12561 1834 12577 1848
rect 12612 1835 12634 1854
rect 12644 1848 12660 1849
rect 12643 1846 12660 1848
rect 12644 1841 12660 1846
rect 12634 1834 12640 1835
rect 12643 1834 12672 1841
rect 12561 1833 12672 1834
rect 12561 1832 12678 1833
rect 12237 1824 12288 1832
rect 12335 1824 12369 1832
rect 12237 1812 12262 1824
rect 12269 1812 12288 1824
rect 12342 1822 12369 1824
rect 12378 1822 12599 1832
rect 12634 1829 12640 1832
rect 12342 1818 12599 1822
rect 12237 1804 12288 1812
rect 12335 1804 12599 1818
rect 12643 1824 12678 1832
rect 12189 1756 12208 1790
rect 12253 1796 12282 1804
rect 12253 1790 12270 1796
rect 12253 1788 12287 1790
rect 12335 1788 12351 1804
rect 12352 1794 12560 1804
rect 12561 1794 12577 1804
rect 12625 1800 12640 1815
rect 12643 1812 12644 1824
rect 12651 1812 12678 1824
rect 12643 1804 12678 1812
rect 12643 1803 12672 1804
rect 12363 1790 12577 1794
rect 12378 1788 12577 1790
rect 12612 1790 12625 1800
rect 12643 1790 12660 1803
rect 12612 1788 12660 1790
rect 12254 1784 12287 1788
rect 12250 1782 12287 1784
rect 12250 1781 12317 1782
rect 12250 1776 12281 1781
rect 12287 1776 12317 1781
rect 12250 1772 12317 1776
rect 12223 1769 12317 1772
rect 12223 1762 12272 1769
rect 12223 1756 12253 1762
rect 12272 1757 12277 1762
rect 12189 1740 12269 1756
rect 12281 1748 12317 1769
rect 12378 1764 12567 1788
rect 12612 1787 12659 1788
rect 12625 1782 12659 1787
rect 12393 1761 12567 1764
rect 12386 1758 12567 1761
rect 12595 1781 12659 1782
rect 12189 1738 12208 1740
rect 12223 1738 12257 1740
rect 12189 1722 12269 1738
rect 12189 1716 12208 1722
rect 11905 1690 12008 1700
rect 11859 1688 12008 1690
rect 12029 1688 12064 1700
rect 11698 1686 11860 1688
rect 11710 1666 11729 1686
rect 11744 1684 11774 1686
rect 11593 1658 11634 1666
rect 11716 1662 11729 1666
rect 11781 1670 11860 1686
rect 11892 1686 12064 1688
rect 11892 1670 11971 1686
rect 11978 1684 12008 1686
rect 11556 1648 11585 1658
rect 11599 1648 11628 1658
rect 11643 1648 11673 1662
rect 11716 1648 11759 1662
rect 11781 1658 11971 1670
rect 12036 1666 12042 1686
rect 11766 1648 11796 1658
rect 11797 1648 11955 1658
rect 11959 1648 11989 1658
rect 11993 1648 12023 1662
rect 12051 1648 12064 1686
rect 12136 1700 12165 1716
rect 12179 1700 12208 1716
rect 12223 1706 12253 1722
rect 12281 1700 12287 1748
rect 12290 1742 12309 1748
rect 12324 1742 12354 1750
rect 12290 1734 12354 1742
rect 12290 1718 12370 1734
rect 12386 1727 12448 1758
rect 12464 1727 12526 1758
rect 12595 1756 12644 1781
rect 12659 1756 12689 1772
rect 12558 1742 12588 1750
rect 12595 1748 12705 1756
rect 12558 1734 12603 1742
rect 12290 1716 12309 1718
rect 12324 1716 12370 1718
rect 12290 1700 12370 1716
rect 12397 1714 12432 1727
rect 12473 1724 12510 1727
rect 12473 1722 12515 1724
rect 12402 1711 12432 1714
rect 12411 1707 12418 1711
rect 12418 1706 12419 1707
rect 12377 1700 12387 1706
rect 12136 1692 12171 1700
rect 12136 1666 12137 1692
rect 12144 1666 12171 1692
rect 12079 1648 12109 1662
rect 12136 1658 12171 1666
rect 12173 1692 12214 1700
rect 12173 1666 12188 1692
rect 12195 1666 12214 1692
rect 12278 1688 12309 1700
rect 12324 1688 12427 1700
rect 12439 1690 12465 1716
rect 12480 1711 12510 1722
rect 12542 1718 12604 1734
rect 12542 1716 12588 1718
rect 12542 1700 12604 1716
rect 12616 1700 12622 1748
rect 12625 1740 12705 1748
rect 12625 1738 12644 1740
rect 12659 1738 12693 1740
rect 12625 1722 12705 1738
rect 12625 1700 12644 1722
rect 12659 1706 12689 1722
rect 12717 1716 12723 1790
rect 12726 1716 12745 1860
rect 12760 1716 12766 1860
rect 12775 1790 12788 1860
rect 12840 1856 12862 1860
rect 12833 1834 12862 1848
rect 12915 1834 12931 1848
rect 12969 1844 12975 1846
rect 12982 1844 13090 1860
rect 13097 1844 13103 1846
rect 13111 1844 13126 1860
rect 13192 1854 13211 1857
rect 12833 1832 12931 1834
rect 12958 1832 13126 1844
rect 13141 1834 13157 1848
rect 13192 1835 13214 1854
rect 13224 1848 13240 1849
rect 13223 1846 13240 1848
rect 13224 1841 13240 1846
rect 13214 1834 13220 1835
rect 13223 1834 13252 1841
rect 13141 1833 13252 1834
rect 13141 1832 13258 1833
rect 12817 1824 12868 1832
rect 12915 1824 12949 1832
rect 12817 1812 12842 1824
rect 12849 1812 12868 1824
rect 12922 1822 12949 1824
rect 12958 1822 13179 1832
rect 13214 1829 13220 1832
rect 12922 1818 13179 1822
rect 12817 1804 12868 1812
rect 12915 1804 13179 1818
rect 13223 1824 13258 1832
rect 12769 1756 12788 1790
rect 12833 1796 12862 1804
rect 12833 1790 12850 1796
rect 12833 1788 12867 1790
rect 12915 1788 12931 1804
rect 12932 1794 13140 1804
rect 13141 1794 13157 1804
rect 13205 1800 13220 1815
rect 13223 1812 13224 1824
rect 13231 1812 13258 1824
rect 13223 1804 13258 1812
rect 13223 1803 13252 1804
rect 12943 1790 13157 1794
rect 12958 1788 13157 1790
rect 13192 1790 13205 1800
rect 13223 1790 13240 1803
rect 13192 1788 13240 1790
rect 12834 1784 12867 1788
rect 12830 1782 12867 1784
rect 12830 1781 12897 1782
rect 12830 1776 12861 1781
rect 12867 1776 12897 1781
rect 12830 1772 12897 1776
rect 12803 1769 12897 1772
rect 12803 1762 12852 1769
rect 12803 1756 12833 1762
rect 12852 1757 12857 1762
rect 12769 1740 12849 1756
rect 12861 1748 12897 1769
rect 12958 1764 13147 1788
rect 13192 1787 13239 1788
rect 13205 1782 13239 1787
rect 12973 1761 13147 1764
rect 12966 1758 13147 1761
rect 13175 1781 13239 1782
rect 12769 1738 12788 1740
rect 12803 1738 12837 1740
rect 12769 1722 12849 1738
rect 12769 1716 12788 1722
rect 12485 1690 12588 1700
rect 12439 1688 12588 1690
rect 12609 1688 12644 1700
rect 12278 1686 12440 1688
rect 12290 1666 12309 1686
rect 12324 1684 12354 1686
rect 12173 1658 12214 1666
rect 12296 1662 12309 1666
rect 12361 1670 12440 1686
rect 12472 1686 12644 1688
rect 12472 1670 12551 1686
rect 12558 1684 12588 1686
rect 12136 1648 12165 1658
rect 12179 1648 12208 1658
rect 12223 1648 12253 1662
rect 12296 1648 12339 1662
rect 12361 1658 12551 1670
rect 12616 1666 12622 1686
rect 12346 1648 12376 1658
rect 12377 1648 12535 1658
rect 12539 1648 12569 1658
rect 12573 1648 12603 1662
rect 12631 1648 12644 1686
rect 12716 1700 12745 1716
rect 12759 1700 12788 1716
rect 12803 1706 12833 1722
rect 12861 1700 12867 1748
rect 12870 1742 12889 1748
rect 12904 1742 12934 1750
rect 12870 1734 12934 1742
rect 12870 1718 12950 1734
rect 12966 1727 13028 1758
rect 13044 1727 13106 1758
rect 13175 1756 13224 1781
rect 13239 1756 13269 1772
rect 13138 1742 13168 1750
rect 13175 1748 13285 1756
rect 13138 1734 13183 1742
rect 12870 1716 12889 1718
rect 12904 1716 12950 1718
rect 12870 1700 12950 1716
rect 12977 1714 13012 1727
rect 13053 1724 13090 1727
rect 13053 1722 13095 1724
rect 12982 1711 13012 1714
rect 12991 1707 12998 1711
rect 12998 1706 12999 1707
rect 12957 1700 12967 1706
rect 12716 1692 12751 1700
rect 12716 1666 12717 1692
rect 12724 1666 12751 1692
rect 12659 1648 12689 1662
rect 12716 1658 12751 1666
rect 12753 1692 12794 1700
rect 12753 1666 12768 1692
rect 12775 1666 12794 1692
rect 12858 1688 12889 1700
rect 12904 1688 13007 1700
rect 13019 1690 13045 1716
rect 13060 1711 13090 1722
rect 13122 1718 13184 1734
rect 13122 1716 13168 1718
rect 13122 1700 13184 1716
rect 13196 1700 13202 1748
rect 13205 1740 13285 1748
rect 13205 1738 13224 1740
rect 13239 1738 13273 1740
rect 13205 1722 13285 1738
rect 13205 1700 13224 1722
rect 13239 1706 13269 1722
rect 13297 1716 13303 1790
rect 13306 1716 13325 1860
rect 13340 1716 13346 1860
rect 13355 1790 13368 1860
rect 13420 1856 13442 1860
rect 13413 1834 13442 1848
rect 13495 1834 13511 1848
rect 13549 1844 13555 1846
rect 13562 1844 13670 1860
rect 13677 1844 13683 1846
rect 13691 1844 13706 1860
rect 13772 1854 13791 1857
rect 13413 1832 13511 1834
rect 13538 1832 13706 1844
rect 13721 1834 13737 1848
rect 13772 1835 13794 1854
rect 13804 1848 13820 1849
rect 13803 1846 13820 1848
rect 13804 1841 13820 1846
rect 13794 1834 13800 1835
rect 13803 1834 13832 1841
rect 13721 1833 13832 1834
rect 13721 1832 13838 1833
rect 13397 1824 13448 1832
rect 13495 1824 13529 1832
rect 13397 1812 13422 1824
rect 13429 1812 13448 1824
rect 13502 1822 13529 1824
rect 13538 1822 13759 1832
rect 13794 1829 13800 1832
rect 13502 1818 13759 1822
rect 13397 1804 13448 1812
rect 13495 1804 13759 1818
rect 13803 1824 13838 1832
rect 13349 1756 13368 1790
rect 13413 1796 13442 1804
rect 13413 1790 13430 1796
rect 13413 1788 13447 1790
rect 13495 1788 13511 1804
rect 13512 1794 13720 1804
rect 13721 1794 13737 1804
rect 13785 1800 13800 1815
rect 13803 1812 13804 1824
rect 13811 1812 13838 1824
rect 13803 1804 13838 1812
rect 13803 1803 13832 1804
rect 13523 1790 13737 1794
rect 13538 1788 13737 1790
rect 13772 1790 13785 1800
rect 13803 1790 13820 1803
rect 13772 1788 13820 1790
rect 13414 1784 13447 1788
rect 13410 1782 13447 1784
rect 13410 1781 13477 1782
rect 13410 1776 13441 1781
rect 13447 1776 13477 1781
rect 13410 1772 13477 1776
rect 13383 1769 13477 1772
rect 13383 1762 13432 1769
rect 13383 1756 13413 1762
rect 13432 1757 13437 1762
rect 13349 1740 13429 1756
rect 13441 1748 13477 1769
rect 13538 1764 13727 1788
rect 13772 1787 13819 1788
rect 13785 1782 13819 1787
rect 13553 1761 13727 1764
rect 13546 1758 13727 1761
rect 13755 1781 13819 1782
rect 13349 1738 13368 1740
rect 13383 1738 13417 1740
rect 13349 1722 13429 1738
rect 13349 1716 13368 1722
rect 13065 1690 13168 1700
rect 13019 1688 13168 1690
rect 13189 1688 13224 1700
rect 12858 1686 13020 1688
rect 12870 1666 12889 1686
rect 12904 1684 12934 1686
rect 12753 1658 12794 1666
rect 12876 1662 12889 1666
rect 12941 1670 13020 1686
rect 13052 1686 13224 1688
rect 13052 1670 13131 1686
rect 13138 1684 13168 1686
rect 12716 1648 12745 1658
rect 12759 1648 12788 1658
rect 12803 1648 12833 1662
rect 12876 1648 12919 1662
rect 12941 1658 13131 1670
rect 13196 1666 13202 1686
rect 12926 1648 12956 1658
rect 12957 1648 13115 1658
rect 13119 1648 13149 1658
rect 13153 1648 13183 1662
rect 13211 1648 13224 1686
rect 13296 1700 13325 1716
rect 13339 1700 13368 1716
rect 13383 1706 13413 1722
rect 13441 1700 13447 1748
rect 13450 1742 13469 1748
rect 13484 1742 13514 1750
rect 13450 1734 13514 1742
rect 13450 1718 13530 1734
rect 13546 1727 13608 1758
rect 13624 1727 13686 1758
rect 13755 1756 13804 1781
rect 13819 1756 13849 1772
rect 13718 1742 13748 1750
rect 13755 1748 13865 1756
rect 13718 1734 13763 1742
rect 13450 1716 13469 1718
rect 13484 1716 13530 1718
rect 13450 1700 13530 1716
rect 13557 1714 13592 1727
rect 13633 1724 13670 1727
rect 13633 1722 13675 1724
rect 13562 1711 13592 1714
rect 13571 1707 13578 1711
rect 13578 1706 13579 1707
rect 13537 1700 13547 1706
rect 13296 1692 13331 1700
rect 13296 1666 13297 1692
rect 13304 1666 13331 1692
rect 13239 1648 13269 1662
rect 13296 1658 13331 1666
rect 13333 1692 13374 1700
rect 13333 1666 13348 1692
rect 13355 1666 13374 1692
rect 13438 1688 13469 1700
rect 13484 1688 13587 1700
rect 13599 1690 13625 1716
rect 13640 1711 13670 1722
rect 13702 1718 13764 1734
rect 13702 1716 13748 1718
rect 13702 1700 13764 1716
rect 13776 1700 13782 1748
rect 13785 1740 13865 1748
rect 13785 1738 13804 1740
rect 13819 1738 13853 1740
rect 13785 1722 13865 1738
rect 13785 1700 13804 1722
rect 13819 1706 13849 1722
rect 13877 1716 13883 1790
rect 13886 1716 13905 1860
rect 13920 1716 13926 1860
rect 13935 1790 13948 1860
rect 14000 1856 14022 1860
rect 13993 1834 14022 1848
rect 14075 1834 14091 1848
rect 14129 1844 14135 1846
rect 14142 1844 14250 1860
rect 14257 1844 14263 1846
rect 14271 1844 14286 1860
rect 14352 1854 14371 1857
rect 13993 1832 14091 1834
rect 14118 1832 14286 1844
rect 14301 1834 14317 1848
rect 14352 1835 14374 1854
rect 14384 1848 14400 1849
rect 14383 1846 14400 1848
rect 14384 1841 14400 1846
rect 14374 1834 14380 1835
rect 14383 1834 14412 1841
rect 14301 1833 14412 1834
rect 14301 1832 14418 1833
rect 13977 1824 14028 1832
rect 14075 1824 14109 1832
rect 13977 1812 14002 1824
rect 14009 1812 14028 1824
rect 14082 1822 14109 1824
rect 14118 1822 14339 1832
rect 14374 1829 14380 1832
rect 14082 1818 14339 1822
rect 13977 1804 14028 1812
rect 14075 1804 14339 1818
rect 14383 1824 14418 1832
rect 13929 1756 13948 1790
rect 13993 1796 14022 1804
rect 13993 1790 14010 1796
rect 13993 1788 14027 1790
rect 14075 1788 14091 1804
rect 14092 1794 14300 1804
rect 14301 1794 14317 1804
rect 14365 1800 14380 1815
rect 14383 1812 14384 1824
rect 14391 1812 14418 1824
rect 14383 1804 14418 1812
rect 14383 1803 14412 1804
rect 14103 1790 14317 1794
rect 14118 1788 14317 1790
rect 14352 1790 14365 1800
rect 14383 1790 14400 1803
rect 14352 1788 14400 1790
rect 13994 1784 14027 1788
rect 13990 1782 14027 1784
rect 13990 1781 14057 1782
rect 13990 1776 14021 1781
rect 14027 1776 14057 1781
rect 13990 1772 14057 1776
rect 13963 1769 14057 1772
rect 13963 1762 14012 1769
rect 13963 1756 13993 1762
rect 14012 1757 14017 1762
rect 13929 1740 14009 1756
rect 14021 1748 14057 1769
rect 14118 1764 14307 1788
rect 14352 1787 14399 1788
rect 14365 1782 14399 1787
rect 14133 1761 14307 1764
rect 14126 1758 14307 1761
rect 14335 1781 14399 1782
rect 13929 1738 13948 1740
rect 13963 1738 13997 1740
rect 13929 1722 14009 1738
rect 13929 1716 13948 1722
rect 13645 1690 13748 1700
rect 13599 1688 13748 1690
rect 13769 1688 13804 1700
rect 13438 1686 13600 1688
rect 13450 1666 13469 1686
rect 13484 1684 13514 1686
rect 13333 1658 13374 1666
rect 13456 1662 13469 1666
rect 13521 1670 13600 1686
rect 13632 1686 13804 1688
rect 13632 1670 13711 1686
rect 13718 1684 13748 1686
rect 13296 1648 13325 1658
rect 13339 1648 13368 1658
rect 13383 1648 13413 1662
rect 13456 1648 13499 1662
rect 13521 1658 13711 1670
rect 13776 1666 13782 1686
rect 13506 1648 13536 1658
rect 13537 1648 13695 1658
rect 13699 1648 13729 1658
rect 13733 1648 13763 1662
rect 13791 1648 13804 1686
rect 13876 1700 13905 1716
rect 13919 1700 13948 1716
rect 13963 1706 13993 1722
rect 14021 1700 14027 1748
rect 14030 1742 14049 1748
rect 14064 1742 14094 1750
rect 14030 1734 14094 1742
rect 14030 1718 14110 1734
rect 14126 1727 14188 1758
rect 14204 1727 14266 1758
rect 14335 1756 14384 1781
rect 14399 1756 14429 1772
rect 14298 1742 14328 1750
rect 14335 1748 14445 1756
rect 14298 1734 14343 1742
rect 14030 1716 14049 1718
rect 14064 1716 14110 1718
rect 14030 1700 14110 1716
rect 14137 1714 14172 1727
rect 14213 1724 14250 1727
rect 14213 1722 14255 1724
rect 14142 1711 14172 1714
rect 14151 1707 14158 1711
rect 14158 1706 14159 1707
rect 14117 1700 14127 1706
rect 13876 1692 13911 1700
rect 13876 1666 13877 1692
rect 13884 1666 13911 1692
rect 13819 1648 13849 1662
rect 13876 1658 13911 1666
rect 13913 1692 13954 1700
rect 13913 1666 13928 1692
rect 13935 1666 13954 1692
rect 14018 1688 14049 1700
rect 14064 1688 14167 1700
rect 14179 1690 14205 1716
rect 14220 1711 14250 1722
rect 14282 1718 14344 1734
rect 14282 1716 14328 1718
rect 14282 1700 14344 1716
rect 14356 1700 14362 1748
rect 14365 1740 14445 1748
rect 14365 1738 14384 1740
rect 14399 1738 14433 1740
rect 14365 1722 14445 1738
rect 14365 1700 14384 1722
rect 14399 1706 14429 1722
rect 14457 1716 14463 1790
rect 14466 1716 14485 1860
rect 14500 1716 14506 1860
rect 14515 1790 14528 1860
rect 14580 1856 14602 1860
rect 14573 1834 14602 1848
rect 14655 1834 14671 1848
rect 14709 1844 14715 1846
rect 14722 1844 14830 1860
rect 14837 1844 14843 1846
rect 14851 1844 14866 1860
rect 14932 1854 14951 1857
rect 14573 1832 14671 1834
rect 14698 1832 14866 1844
rect 14881 1834 14897 1848
rect 14932 1835 14954 1854
rect 14964 1848 14980 1849
rect 14963 1846 14980 1848
rect 14964 1841 14980 1846
rect 14954 1834 14960 1835
rect 14963 1834 14992 1841
rect 14881 1833 14992 1834
rect 14881 1832 14998 1833
rect 14557 1824 14608 1832
rect 14655 1824 14689 1832
rect 14557 1812 14582 1824
rect 14589 1812 14608 1824
rect 14662 1822 14689 1824
rect 14698 1822 14919 1832
rect 14954 1829 14960 1832
rect 14662 1818 14919 1822
rect 14557 1804 14608 1812
rect 14655 1804 14919 1818
rect 14963 1824 14998 1832
rect 14509 1756 14528 1790
rect 14573 1796 14602 1804
rect 14573 1790 14590 1796
rect 14573 1788 14607 1790
rect 14655 1788 14671 1804
rect 14672 1794 14880 1804
rect 14881 1794 14897 1804
rect 14945 1800 14960 1815
rect 14963 1812 14964 1824
rect 14971 1812 14998 1824
rect 14963 1804 14998 1812
rect 14963 1803 14992 1804
rect 14683 1790 14897 1794
rect 14698 1788 14897 1790
rect 14932 1790 14945 1800
rect 14963 1790 14980 1803
rect 14932 1788 14980 1790
rect 14574 1784 14607 1788
rect 14570 1782 14607 1784
rect 14570 1781 14637 1782
rect 14570 1776 14601 1781
rect 14607 1776 14637 1781
rect 14570 1772 14637 1776
rect 14543 1769 14637 1772
rect 14543 1762 14592 1769
rect 14543 1756 14573 1762
rect 14592 1757 14597 1762
rect 14509 1740 14589 1756
rect 14601 1748 14637 1769
rect 14698 1764 14887 1788
rect 14932 1787 14979 1788
rect 14945 1782 14979 1787
rect 14713 1761 14887 1764
rect 14706 1758 14887 1761
rect 14915 1781 14979 1782
rect 14509 1738 14528 1740
rect 14543 1738 14577 1740
rect 14509 1722 14589 1738
rect 14509 1716 14528 1722
rect 14225 1690 14328 1700
rect 14179 1688 14328 1690
rect 14349 1688 14384 1700
rect 14018 1686 14180 1688
rect 14030 1666 14049 1686
rect 14064 1684 14094 1686
rect 13913 1658 13954 1666
rect 14036 1662 14049 1666
rect 14101 1670 14180 1686
rect 14212 1686 14384 1688
rect 14212 1670 14291 1686
rect 14298 1684 14328 1686
rect 13876 1648 13905 1658
rect 13919 1648 13948 1658
rect 13963 1648 13993 1662
rect 14036 1648 14079 1662
rect 14101 1658 14291 1670
rect 14356 1666 14362 1686
rect 14086 1648 14116 1658
rect 14117 1648 14275 1658
rect 14279 1648 14309 1658
rect 14313 1648 14343 1662
rect 14371 1648 14384 1686
rect 14456 1700 14485 1716
rect 14499 1700 14528 1716
rect 14543 1706 14573 1722
rect 14601 1700 14607 1748
rect 14610 1742 14629 1748
rect 14644 1742 14674 1750
rect 14610 1734 14674 1742
rect 14610 1718 14690 1734
rect 14706 1727 14768 1758
rect 14784 1727 14846 1758
rect 14915 1756 14964 1781
rect 14979 1756 15009 1772
rect 14878 1742 14908 1750
rect 14915 1748 15025 1756
rect 14878 1734 14923 1742
rect 14610 1716 14629 1718
rect 14644 1716 14690 1718
rect 14610 1700 14690 1716
rect 14717 1714 14752 1727
rect 14793 1724 14830 1727
rect 14793 1722 14835 1724
rect 14722 1711 14752 1714
rect 14731 1707 14738 1711
rect 14738 1706 14739 1707
rect 14697 1700 14707 1706
rect 14456 1692 14491 1700
rect 14456 1666 14457 1692
rect 14464 1666 14491 1692
rect 14399 1648 14429 1662
rect 14456 1658 14491 1666
rect 14493 1692 14534 1700
rect 14493 1666 14508 1692
rect 14515 1666 14534 1692
rect 14598 1688 14629 1700
rect 14644 1688 14747 1700
rect 14759 1690 14785 1716
rect 14800 1711 14830 1722
rect 14862 1718 14924 1734
rect 14862 1716 14908 1718
rect 14862 1700 14924 1716
rect 14936 1700 14942 1748
rect 14945 1740 15025 1748
rect 14945 1738 14964 1740
rect 14979 1738 15013 1740
rect 14945 1722 15025 1738
rect 14945 1700 14964 1722
rect 14979 1706 15009 1722
rect 15037 1716 15043 1790
rect 15046 1716 15065 1860
rect 15080 1716 15086 1860
rect 15095 1790 15108 1860
rect 15160 1856 15182 1860
rect 15153 1834 15182 1848
rect 15235 1834 15251 1848
rect 15289 1844 15295 1846
rect 15302 1844 15410 1860
rect 15417 1844 15423 1846
rect 15431 1844 15446 1860
rect 15512 1854 15531 1857
rect 15153 1832 15251 1834
rect 15278 1832 15446 1844
rect 15461 1834 15477 1848
rect 15512 1835 15534 1854
rect 15544 1848 15560 1849
rect 15543 1846 15560 1848
rect 15544 1841 15560 1846
rect 15534 1834 15540 1835
rect 15543 1834 15572 1841
rect 15461 1833 15572 1834
rect 15461 1832 15578 1833
rect 15137 1824 15188 1832
rect 15235 1824 15269 1832
rect 15137 1812 15162 1824
rect 15169 1812 15188 1824
rect 15242 1822 15269 1824
rect 15278 1822 15499 1832
rect 15534 1829 15540 1832
rect 15242 1818 15499 1822
rect 15137 1804 15188 1812
rect 15235 1804 15499 1818
rect 15543 1824 15578 1832
rect 15089 1756 15108 1790
rect 15153 1796 15182 1804
rect 15153 1790 15170 1796
rect 15153 1788 15187 1790
rect 15235 1788 15251 1804
rect 15252 1794 15460 1804
rect 15461 1794 15477 1804
rect 15525 1800 15540 1815
rect 15543 1812 15544 1824
rect 15551 1812 15578 1824
rect 15543 1804 15578 1812
rect 15543 1803 15572 1804
rect 15263 1790 15477 1794
rect 15278 1788 15477 1790
rect 15512 1790 15525 1800
rect 15543 1790 15560 1803
rect 15512 1788 15560 1790
rect 15154 1784 15187 1788
rect 15150 1782 15187 1784
rect 15150 1781 15217 1782
rect 15150 1776 15181 1781
rect 15187 1776 15217 1781
rect 15150 1772 15217 1776
rect 15123 1769 15217 1772
rect 15123 1762 15172 1769
rect 15123 1756 15153 1762
rect 15172 1757 15177 1762
rect 15089 1740 15169 1756
rect 15181 1748 15217 1769
rect 15278 1764 15467 1788
rect 15512 1787 15559 1788
rect 15525 1782 15559 1787
rect 15293 1761 15467 1764
rect 15286 1758 15467 1761
rect 15495 1781 15559 1782
rect 15089 1738 15108 1740
rect 15123 1738 15157 1740
rect 15089 1722 15169 1738
rect 15089 1716 15108 1722
rect 14805 1690 14908 1700
rect 14759 1688 14908 1690
rect 14929 1688 14964 1700
rect 14598 1686 14760 1688
rect 14610 1666 14629 1686
rect 14644 1684 14674 1686
rect 14493 1658 14534 1666
rect 14616 1662 14629 1666
rect 14681 1670 14760 1686
rect 14792 1686 14964 1688
rect 14792 1670 14871 1686
rect 14878 1684 14908 1686
rect 14456 1648 14485 1658
rect 14499 1648 14528 1658
rect 14543 1648 14573 1662
rect 14616 1648 14659 1662
rect 14681 1658 14871 1670
rect 14936 1666 14942 1686
rect 14666 1648 14696 1658
rect 14697 1648 14855 1658
rect 14859 1648 14889 1658
rect 14893 1648 14923 1662
rect 14951 1648 14964 1686
rect 15036 1700 15065 1716
rect 15079 1700 15108 1716
rect 15123 1706 15153 1722
rect 15181 1700 15187 1748
rect 15190 1742 15209 1748
rect 15224 1742 15254 1750
rect 15190 1734 15254 1742
rect 15190 1718 15270 1734
rect 15286 1727 15348 1758
rect 15364 1727 15426 1758
rect 15495 1756 15544 1781
rect 15559 1756 15589 1772
rect 15458 1742 15488 1750
rect 15495 1748 15605 1756
rect 15458 1734 15503 1742
rect 15190 1716 15209 1718
rect 15224 1716 15270 1718
rect 15190 1700 15270 1716
rect 15297 1714 15332 1727
rect 15373 1724 15410 1727
rect 15373 1722 15415 1724
rect 15302 1711 15332 1714
rect 15311 1707 15318 1711
rect 15318 1706 15319 1707
rect 15277 1700 15287 1706
rect 15036 1692 15071 1700
rect 15036 1666 15037 1692
rect 15044 1666 15071 1692
rect 14979 1648 15009 1662
rect 15036 1658 15071 1666
rect 15073 1692 15114 1700
rect 15073 1666 15088 1692
rect 15095 1666 15114 1692
rect 15178 1688 15209 1700
rect 15224 1688 15327 1700
rect 15339 1690 15365 1716
rect 15380 1711 15410 1722
rect 15442 1718 15504 1734
rect 15442 1716 15488 1718
rect 15442 1700 15504 1716
rect 15516 1700 15522 1748
rect 15525 1740 15605 1748
rect 15525 1738 15544 1740
rect 15559 1738 15593 1740
rect 15525 1722 15605 1738
rect 15525 1700 15544 1722
rect 15559 1706 15589 1722
rect 15617 1716 15623 1790
rect 15626 1716 15645 1860
rect 15660 1716 15666 1860
rect 15675 1790 15688 1860
rect 15740 1856 15762 1860
rect 15733 1834 15762 1848
rect 15815 1834 15831 1848
rect 15869 1844 15875 1846
rect 15882 1844 15990 1860
rect 15997 1844 16003 1846
rect 16011 1844 16026 1860
rect 16092 1854 16111 1857
rect 15733 1832 15831 1834
rect 15858 1832 16026 1844
rect 16041 1834 16057 1848
rect 16092 1835 16114 1854
rect 16124 1848 16140 1849
rect 16123 1846 16140 1848
rect 16124 1841 16140 1846
rect 16114 1834 16120 1835
rect 16123 1834 16152 1841
rect 16041 1833 16152 1834
rect 16041 1832 16158 1833
rect 15717 1824 15768 1832
rect 15815 1824 15849 1832
rect 15717 1812 15742 1824
rect 15749 1812 15768 1824
rect 15822 1822 15849 1824
rect 15858 1822 16079 1832
rect 16114 1829 16120 1832
rect 15822 1818 16079 1822
rect 15717 1804 15768 1812
rect 15815 1804 16079 1818
rect 16123 1824 16158 1832
rect 15669 1756 15688 1790
rect 15733 1796 15762 1804
rect 15733 1790 15750 1796
rect 15733 1788 15767 1790
rect 15815 1788 15831 1804
rect 15832 1794 16040 1804
rect 16041 1794 16057 1804
rect 16105 1800 16120 1815
rect 16123 1812 16124 1824
rect 16131 1812 16158 1824
rect 16123 1804 16158 1812
rect 16123 1803 16152 1804
rect 15843 1790 16057 1794
rect 15858 1788 16057 1790
rect 16092 1790 16105 1800
rect 16123 1790 16140 1803
rect 16092 1788 16140 1790
rect 15734 1784 15767 1788
rect 15730 1782 15767 1784
rect 15730 1781 15797 1782
rect 15730 1776 15761 1781
rect 15767 1776 15797 1781
rect 15730 1772 15797 1776
rect 15703 1769 15797 1772
rect 15703 1762 15752 1769
rect 15703 1756 15733 1762
rect 15752 1757 15757 1762
rect 15669 1740 15749 1756
rect 15761 1748 15797 1769
rect 15858 1764 16047 1788
rect 16092 1787 16139 1788
rect 16105 1782 16139 1787
rect 15873 1761 16047 1764
rect 15866 1758 16047 1761
rect 16075 1781 16139 1782
rect 15669 1738 15688 1740
rect 15703 1738 15737 1740
rect 15669 1722 15749 1738
rect 15669 1716 15688 1722
rect 15385 1690 15488 1700
rect 15339 1688 15488 1690
rect 15509 1688 15544 1700
rect 15178 1686 15340 1688
rect 15190 1666 15209 1686
rect 15224 1684 15254 1686
rect 15073 1658 15114 1666
rect 15196 1662 15209 1666
rect 15261 1670 15340 1686
rect 15372 1686 15544 1688
rect 15372 1670 15451 1686
rect 15458 1684 15488 1686
rect 15036 1648 15065 1658
rect 15079 1648 15108 1658
rect 15123 1648 15153 1662
rect 15196 1648 15239 1662
rect 15261 1658 15451 1670
rect 15516 1666 15522 1686
rect 15246 1648 15276 1658
rect 15277 1648 15435 1658
rect 15439 1648 15469 1658
rect 15473 1648 15503 1662
rect 15531 1648 15544 1686
rect 15616 1700 15645 1716
rect 15659 1700 15688 1716
rect 15703 1706 15733 1722
rect 15761 1700 15767 1748
rect 15770 1742 15789 1748
rect 15804 1742 15834 1750
rect 15770 1734 15834 1742
rect 15770 1718 15850 1734
rect 15866 1727 15928 1758
rect 15944 1727 16006 1758
rect 16075 1756 16124 1781
rect 16139 1756 16169 1772
rect 16038 1742 16068 1750
rect 16075 1748 16185 1756
rect 16038 1734 16083 1742
rect 15770 1716 15789 1718
rect 15804 1716 15850 1718
rect 15770 1700 15850 1716
rect 15877 1714 15912 1727
rect 15953 1724 15990 1727
rect 15953 1722 15995 1724
rect 15882 1711 15912 1714
rect 15891 1707 15898 1711
rect 15898 1706 15899 1707
rect 15857 1700 15867 1706
rect 15616 1692 15651 1700
rect 15616 1666 15617 1692
rect 15624 1666 15651 1692
rect 15559 1648 15589 1662
rect 15616 1658 15651 1666
rect 15653 1692 15694 1700
rect 15653 1666 15668 1692
rect 15675 1666 15694 1692
rect 15758 1688 15789 1700
rect 15804 1688 15907 1700
rect 15919 1690 15945 1716
rect 15960 1711 15990 1722
rect 16022 1718 16084 1734
rect 16022 1716 16068 1718
rect 16022 1700 16084 1716
rect 16096 1700 16102 1748
rect 16105 1740 16185 1748
rect 16105 1738 16124 1740
rect 16139 1738 16173 1740
rect 16105 1722 16185 1738
rect 16105 1700 16124 1722
rect 16139 1706 16169 1722
rect 16197 1716 16203 1790
rect 16206 1716 16225 1860
rect 16240 1716 16246 1860
rect 16255 1790 16268 1860
rect 16320 1856 16342 1860
rect 16313 1834 16342 1848
rect 16395 1834 16411 1848
rect 16449 1844 16455 1846
rect 16462 1844 16570 1860
rect 16577 1844 16583 1846
rect 16591 1844 16606 1860
rect 16672 1854 16691 1857
rect 16313 1832 16411 1834
rect 16438 1832 16606 1844
rect 16621 1834 16637 1848
rect 16672 1835 16694 1854
rect 16704 1848 16720 1849
rect 16703 1846 16720 1848
rect 16704 1841 16720 1846
rect 16694 1834 16700 1835
rect 16703 1834 16732 1841
rect 16621 1833 16732 1834
rect 16621 1832 16738 1833
rect 16297 1824 16348 1832
rect 16395 1824 16429 1832
rect 16297 1812 16322 1824
rect 16329 1812 16348 1824
rect 16402 1822 16429 1824
rect 16438 1822 16659 1832
rect 16694 1829 16700 1832
rect 16402 1818 16659 1822
rect 16297 1804 16348 1812
rect 16395 1804 16659 1818
rect 16703 1824 16738 1832
rect 16249 1756 16268 1790
rect 16313 1796 16342 1804
rect 16313 1790 16330 1796
rect 16313 1788 16347 1790
rect 16395 1788 16411 1804
rect 16412 1794 16620 1804
rect 16621 1794 16637 1804
rect 16685 1800 16700 1815
rect 16703 1812 16704 1824
rect 16711 1812 16738 1824
rect 16703 1804 16738 1812
rect 16703 1803 16732 1804
rect 16423 1790 16637 1794
rect 16438 1788 16637 1790
rect 16672 1790 16685 1800
rect 16703 1790 16720 1803
rect 16672 1788 16720 1790
rect 16314 1784 16347 1788
rect 16310 1782 16347 1784
rect 16310 1781 16377 1782
rect 16310 1776 16341 1781
rect 16347 1776 16377 1781
rect 16310 1772 16377 1776
rect 16283 1769 16377 1772
rect 16283 1762 16332 1769
rect 16283 1756 16313 1762
rect 16332 1757 16337 1762
rect 16249 1740 16329 1756
rect 16341 1748 16377 1769
rect 16438 1764 16627 1788
rect 16672 1787 16719 1788
rect 16685 1782 16719 1787
rect 16453 1761 16627 1764
rect 16446 1758 16627 1761
rect 16655 1781 16719 1782
rect 16249 1738 16268 1740
rect 16283 1738 16317 1740
rect 16249 1722 16329 1738
rect 16249 1716 16268 1722
rect 15965 1690 16068 1700
rect 15919 1688 16068 1690
rect 16089 1688 16124 1700
rect 15758 1686 15920 1688
rect 15770 1666 15789 1686
rect 15804 1684 15834 1686
rect 15653 1658 15694 1666
rect 15776 1662 15789 1666
rect 15841 1670 15920 1686
rect 15952 1686 16124 1688
rect 15952 1670 16031 1686
rect 16038 1684 16068 1686
rect 15616 1648 15645 1658
rect 15659 1648 15688 1658
rect 15703 1648 15733 1662
rect 15776 1648 15819 1662
rect 15841 1658 16031 1670
rect 16096 1666 16102 1686
rect 15826 1648 15856 1658
rect 15857 1648 16015 1658
rect 16019 1648 16049 1658
rect 16053 1648 16083 1662
rect 16111 1648 16124 1686
rect 16196 1700 16225 1716
rect 16239 1700 16268 1716
rect 16283 1706 16313 1722
rect 16341 1700 16347 1748
rect 16350 1742 16369 1748
rect 16384 1742 16414 1750
rect 16350 1734 16414 1742
rect 16350 1718 16430 1734
rect 16446 1727 16508 1758
rect 16524 1727 16586 1758
rect 16655 1756 16704 1781
rect 16719 1756 16749 1772
rect 16618 1742 16648 1750
rect 16655 1748 16765 1756
rect 16618 1734 16663 1742
rect 16350 1716 16369 1718
rect 16384 1716 16430 1718
rect 16350 1700 16430 1716
rect 16457 1714 16492 1727
rect 16533 1724 16570 1727
rect 16533 1722 16575 1724
rect 16462 1711 16492 1714
rect 16471 1707 16478 1711
rect 16478 1706 16479 1707
rect 16437 1700 16447 1706
rect 16196 1692 16231 1700
rect 16196 1666 16197 1692
rect 16204 1666 16231 1692
rect 16139 1648 16169 1662
rect 16196 1658 16231 1666
rect 16233 1692 16274 1700
rect 16233 1666 16248 1692
rect 16255 1666 16274 1692
rect 16338 1688 16369 1700
rect 16384 1688 16487 1700
rect 16499 1690 16525 1716
rect 16540 1711 16570 1722
rect 16602 1718 16664 1734
rect 16602 1716 16648 1718
rect 16602 1700 16664 1716
rect 16676 1700 16682 1748
rect 16685 1740 16765 1748
rect 16685 1738 16704 1740
rect 16719 1738 16753 1740
rect 16685 1722 16765 1738
rect 16685 1700 16704 1722
rect 16719 1706 16749 1722
rect 16777 1716 16783 1790
rect 16786 1716 16805 1860
rect 16820 1716 16826 1860
rect 16835 1790 16848 1860
rect 16900 1856 16922 1860
rect 16893 1834 16922 1848
rect 16975 1834 16991 1848
rect 17029 1844 17035 1846
rect 17042 1844 17150 1860
rect 17157 1844 17163 1846
rect 17171 1844 17186 1860
rect 17252 1854 17271 1857
rect 16893 1832 16991 1834
rect 17018 1832 17186 1844
rect 17201 1834 17217 1848
rect 17252 1835 17274 1854
rect 17284 1848 17300 1849
rect 17283 1846 17300 1848
rect 17284 1841 17300 1846
rect 17274 1834 17280 1835
rect 17283 1834 17312 1841
rect 17201 1833 17312 1834
rect 17201 1832 17318 1833
rect 16877 1824 16928 1832
rect 16975 1824 17009 1832
rect 16877 1812 16902 1824
rect 16909 1812 16928 1824
rect 16982 1822 17009 1824
rect 17018 1822 17239 1832
rect 17274 1829 17280 1832
rect 16982 1818 17239 1822
rect 16877 1804 16928 1812
rect 16975 1804 17239 1818
rect 17283 1824 17318 1832
rect 16829 1756 16848 1790
rect 16893 1796 16922 1804
rect 16893 1790 16910 1796
rect 16893 1788 16927 1790
rect 16975 1788 16991 1804
rect 16992 1794 17200 1804
rect 17201 1794 17217 1804
rect 17265 1800 17280 1815
rect 17283 1812 17284 1824
rect 17291 1812 17318 1824
rect 17283 1804 17318 1812
rect 17283 1803 17312 1804
rect 17003 1790 17217 1794
rect 17018 1788 17217 1790
rect 17252 1790 17265 1800
rect 17283 1790 17300 1803
rect 17252 1788 17300 1790
rect 16894 1784 16927 1788
rect 16890 1782 16927 1784
rect 16890 1781 16957 1782
rect 16890 1776 16921 1781
rect 16927 1776 16957 1781
rect 16890 1772 16957 1776
rect 16863 1769 16957 1772
rect 16863 1762 16912 1769
rect 16863 1756 16893 1762
rect 16912 1757 16917 1762
rect 16829 1740 16909 1756
rect 16921 1748 16957 1769
rect 17018 1764 17207 1788
rect 17252 1787 17299 1788
rect 17265 1782 17299 1787
rect 17033 1761 17207 1764
rect 17026 1758 17207 1761
rect 17235 1781 17299 1782
rect 16829 1738 16848 1740
rect 16863 1738 16897 1740
rect 16829 1722 16909 1738
rect 16829 1716 16848 1722
rect 16545 1690 16648 1700
rect 16499 1688 16648 1690
rect 16669 1688 16704 1700
rect 16338 1686 16500 1688
rect 16350 1666 16369 1686
rect 16384 1684 16414 1686
rect 16233 1658 16274 1666
rect 16356 1662 16369 1666
rect 16421 1670 16500 1686
rect 16532 1686 16704 1688
rect 16532 1670 16611 1686
rect 16618 1684 16648 1686
rect 16196 1648 16225 1658
rect 16239 1648 16268 1658
rect 16283 1648 16313 1662
rect 16356 1648 16399 1662
rect 16421 1658 16611 1670
rect 16676 1666 16682 1686
rect 16406 1648 16436 1658
rect 16437 1648 16595 1658
rect 16599 1648 16629 1658
rect 16633 1648 16663 1662
rect 16691 1648 16704 1686
rect 16776 1700 16805 1716
rect 16819 1700 16848 1716
rect 16863 1706 16893 1722
rect 16921 1700 16927 1748
rect 16930 1742 16949 1748
rect 16964 1742 16994 1750
rect 16930 1734 16994 1742
rect 16930 1718 17010 1734
rect 17026 1727 17088 1758
rect 17104 1727 17166 1758
rect 17235 1756 17284 1781
rect 17299 1756 17329 1772
rect 17198 1742 17228 1750
rect 17235 1748 17345 1756
rect 17198 1734 17243 1742
rect 16930 1716 16949 1718
rect 16964 1716 17010 1718
rect 16930 1700 17010 1716
rect 17037 1714 17072 1727
rect 17113 1724 17150 1727
rect 17113 1722 17155 1724
rect 17042 1711 17072 1714
rect 17051 1707 17058 1711
rect 17058 1706 17059 1707
rect 17017 1700 17027 1706
rect 16776 1692 16811 1700
rect 16776 1666 16777 1692
rect 16784 1666 16811 1692
rect 16719 1648 16749 1662
rect 16776 1658 16811 1666
rect 16813 1692 16854 1700
rect 16813 1666 16828 1692
rect 16835 1666 16854 1692
rect 16918 1688 16949 1700
rect 16964 1688 17067 1700
rect 17079 1690 17105 1716
rect 17120 1711 17150 1722
rect 17182 1718 17244 1734
rect 17182 1716 17228 1718
rect 17182 1700 17244 1716
rect 17256 1700 17262 1748
rect 17265 1740 17345 1748
rect 17265 1738 17284 1740
rect 17299 1738 17333 1740
rect 17265 1722 17345 1738
rect 17265 1700 17284 1722
rect 17299 1706 17329 1722
rect 17357 1716 17363 1790
rect 17366 1716 17385 1860
rect 17400 1716 17406 1860
rect 17415 1790 17428 1860
rect 17480 1856 17502 1860
rect 17473 1834 17502 1848
rect 17555 1834 17571 1848
rect 17609 1844 17615 1846
rect 17622 1844 17730 1860
rect 17737 1844 17743 1846
rect 17751 1844 17766 1860
rect 17832 1854 17851 1857
rect 17473 1832 17571 1834
rect 17598 1832 17766 1844
rect 17781 1834 17797 1848
rect 17832 1835 17854 1854
rect 17864 1848 17880 1849
rect 17863 1846 17880 1848
rect 17864 1841 17880 1846
rect 17854 1834 17860 1835
rect 17863 1834 17892 1841
rect 17781 1833 17892 1834
rect 17781 1832 17898 1833
rect 17457 1824 17508 1832
rect 17555 1824 17589 1832
rect 17457 1812 17482 1824
rect 17489 1812 17508 1824
rect 17562 1822 17589 1824
rect 17598 1822 17819 1832
rect 17854 1829 17860 1832
rect 17562 1818 17819 1822
rect 17457 1804 17508 1812
rect 17555 1804 17819 1818
rect 17863 1824 17898 1832
rect 17409 1756 17428 1790
rect 17473 1796 17502 1804
rect 17473 1790 17490 1796
rect 17473 1788 17507 1790
rect 17555 1788 17571 1804
rect 17572 1794 17780 1804
rect 17781 1794 17797 1804
rect 17845 1800 17860 1815
rect 17863 1812 17864 1824
rect 17871 1812 17898 1824
rect 17863 1804 17898 1812
rect 17863 1803 17892 1804
rect 17583 1790 17797 1794
rect 17598 1788 17797 1790
rect 17832 1790 17845 1800
rect 17863 1790 17880 1803
rect 17832 1788 17880 1790
rect 17474 1784 17507 1788
rect 17470 1782 17507 1784
rect 17470 1781 17537 1782
rect 17470 1776 17501 1781
rect 17507 1776 17537 1781
rect 17470 1772 17537 1776
rect 17443 1769 17537 1772
rect 17443 1762 17492 1769
rect 17443 1756 17473 1762
rect 17492 1757 17497 1762
rect 17409 1740 17489 1756
rect 17501 1748 17537 1769
rect 17598 1764 17787 1788
rect 17832 1787 17879 1788
rect 17845 1782 17879 1787
rect 17613 1761 17787 1764
rect 17606 1758 17787 1761
rect 17815 1781 17879 1782
rect 17409 1738 17428 1740
rect 17443 1738 17477 1740
rect 17409 1722 17489 1738
rect 17409 1716 17428 1722
rect 17125 1690 17228 1700
rect 17079 1688 17228 1690
rect 17249 1688 17284 1700
rect 16918 1686 17080 1688
rect 16930 1666 16949 1686
rect 16964 1684 16994 1686
rect 16813 1658 16854 1666
rect 16936 1662 16949 1666
rect 17001 1670 17080 1686
rect 17112 1686 17284 1688
rect 17112 1670 17191 1686
rect 17198 1684 17228 1686
rect 16776 1648 16805 1658
rect 16819 1648 16848 1658
rect 16863 1648 16893 1662
rect 16936 1648 16979 1662
rect 17001 1658 17191 1670
rect 17256 1666 17262 1686
rect 16986 1648 17016 1658
rect 17017 1648 17175 1658
rect 17179 1648 17209 1658
rect 17213 1648 17243 1662
rect 17271 1648 17284 1686
rect 17356 1700 17385 1716
rect 17399 1700 17428 1716
rect 17443 1706 17473 1722
rect 17501 1700 17507 1748
rect 17510 1742 17529 1748
rect 17544 1742 17574 1750
rect 17510 1734 17574 1742
rect 17510 1718 17590 1734
rect 17606 1727 17668 1758
rect 17684 1727 17746 1758
rect 17815 1756 17864 1781
rect 17879 1756 17909 1772
rect 17778 1742 17808 1750
rect 17815 1748 17925 1756
rect 17778 1734 17823 1742
rect 17510 1716 17529 1718
rect 17544 1716 17590 1718
rect 17510 1700 17590 1716
rect 17617 1714 17652 1727
rect 17693 1724 17730 1727
rect 17693 1722 17735 1724
rect 17622 1711 17652 1714
rect 17631 1707 17638 1711
rect 17638 1706 17639 1707
rect 17597 1700 17607 1706
rect 17356 1692 17391 1700
rect 17356 1666 17357 1692
rect 17364 1666 17391 1692
rect 17299 1648 17329 1662
rect 17356 1658 17391 1666
rect 17393 1692 17434 1700
rect 17393 1666 17408 1692
rect 17415 1666 17434 1692
rect 17498 1688 17529 1700
rect 17544 1688 17647 1700
rect 17659 1690 17685 1716
rect 17700 1711 17730 1722
rect 17762 1718 17824 1734
rect 17762 1716 17808 1718
rect 17762 1700 17824 1716
rect 17836 1700 17842 1748
rect 17845 1740 17925 1748
rect 17845 1738 17864 1740
rect 17879 1738 17913 1740
rect 17845 1722 17925 1738
rect 17845 1700 17864 1722
rect 17879 1706 17909 1722
rect 17937 1716 17943 1790
rect 17946 1716 17965 1860
rect 17980 1716 17986 1860
rect 17995 1790 18008 1860
rect 18060 1856 18082 1860
rect 18053 1834 18082 1848
rect 18135 1834 18151 1848
rect 18189 1844 18195 1846
rect 18202 1844 18310 1860
rect 18317 1844 18323 1846
rect 18331 1844 18346 1860
rect 18412 1854 18431 1857
rect 18053 1832 18151 1834
rect 18178 1832 18346 1844
rect 18361 1834 18377 1848
rect 18412 1835 18434 1854
rect 18444 1848 18460 1849
rect 18443 1846 18460 1848
rect 18444 1841 18460 1846
rect 18434 1834 18440 1835
rect 18443 1834 18472 1841
rect 18361 1833 18472 1834
rect 18361 1832 18478 1833
rect 18037 1824 18088 1832
rect 18135 1824 18169 1832
rect 18037 1812 18062 1824
rect 18069 1812 18088 1824
rect 18142 1822 18169 1824
rect 18178 1822 18399 1832
rect 18434 1829 18440 1832
rect 18142 1818 18399 1822
rect 18037 1804 18088 1812
rect 18135 1804 18399 1818
rect 18443 1824 18478 1832
rect 17989 1756 18008 1790
rect 18053 1796 18082 1804
rect 18053 1790 18070 1796
rect 18053 1788 18087 1790
rect 18135 1788 18151 1804
rect 18152 1794 18360 1804
rect 18361 1794 18377 1804
rect 18425 1800 18440 1815
rect 18443 1812 18444 1824
rect 18451 1812 18478 1824
rect 18443 1804 18478 1812
rect 18443 1803 18472 1804
rect 18163 1790 18377 1794
rect 18178 1788 18377 1790
rect 18412 1790 18425 1800
rect 18443 1790 18460 1803
rect 18412 1788 18460 1790
rect 18054 1784 18087 1788
rect 18050 1782 18087 1784
rect 18050 1781 18117 1782
rect 18050 1776 18081 1781
rect 18087 1776 18117 1781
rect 18050 1772 18117 1776
rect 18023 1769 18117 1772
rect 18023 1762 18072 1769
rect 18023 1756 18053 1762
rect 18072 1757 18077 1762
rect 17989 1740 18069 1756
rect 18081 1748 18117 1769
rect 18178 1764 18367 1788
rect 18412 1787 18459 1788
rect 18425 1782 18459 1787
rect 18193 1761 18367 1764
rect 18186 1758 18367 1761
rect 18395 1781 18459 1782
rect 17989 1738 18008 1740
rect 18023 1738 18057 1740
rect 17989 1722 18069 1738
rect 17989 1716 18008 1722
rect 17705 1690 17808 1700
rect 17659 1688 17808 1690
rect 17829 1688 17864 1700
rect 17498 1686 17660 1688
rect 17510 1666 17529 1686
rect 17544 1684 17574 1686
rect 17393 1658 17434 1666
rect 17516 1662 17529 1666
rect 17581 1670 17660 1686
rect 17692 1686 17864 1688
rect 17692 1670 17771 1686
rect 17778 1684 17808 1686
rect 17356 1648 17385 1658
rect 17399 1648 17428 1658
rect 17443 1648 17473 1662
rect 17516 1648 17559 1662
rect 17581 1658 17771 1670
rect 17836 1666 17842 1686
rect 17566 1648 17596 1658
rect 17597 1648 17755 1658
rect 17759 1648 17789 1658
rect 17793 1648 17823 1662
rect 17851 1648 17864 1686
rect 17936 1700 17965 1716
rect 17979 1700 18008 1716
rect 18023 1706 18053 1722
rect 18081 1700 18087 1748
rect 18090 1742 18109 1748
rect 18124 1742 18154 1750
rect 18090 1734 18154 1742
rect 18090 1718 18170 1734
rect 18186 1727 18248 1758
rect 18264 1727 18326 1758
rect 18395 1756 18444 1781
rect 18459 1756 18489 1772
rect 18358 1742 18388 1750
rect 18395 1748 18505 1756
rect 18358 1734 18403 1742
rect 18090 1716 18109 1718
rect 18124 1716 18170 1718
rect 18090 1700 18170 1716
rect 18197 1714 18232 1727
rect 18273 1724 18310 1727
rect 18273 1722 18315 1724
rect 18202 1711 18232 1714
rect 18211 1707 18218 1711
rect 18218 1706 18219 1707
rect 18177 1700 18187 1706
rect 17936 1692 17971 1700
rect 17936 1666 17937 1692
rect 17944 1666 17971 1692
rect 17879 1648 17909 1662
rect 17936 1658 17971 1666
rect 17973 1692 18014 1700
rect 17973 1666 17988 1692
rect 17995 1666 18014 1692
rect 18078 1688 18109 1700
rect 18124 1688 18227 1700
rect 18239 1690 18265 1716
rect 18280 1711 18310 1722
rect 18342 1718 18404 1734
rect 18342 1716 18388 1718
rect 18342 1700 18404 1716
rect 18416 1700 18422 1748
rect 18425 1740 18505 1748
rect 18425 1738 18444 1740
rect 18459 1738 18493 1740
rect 18425 1722 18505 1738
rect 18425 1700 18444 1722
rect 18459 1706 18489 1722
rect 18517 1716 18523 1790
rect 18532 1716 18545 1860
rect 18285 1690 18388 1700
rect 18239 1688 18388 1690
rect 18409 1688 18444 1700
rect 18078 1686 18240 1688
rect 18090 1666 18109 1686
rect 18124 1684 18154 1686
rect 17973 1658 18014 1666
rect 18096 1662 18109 1666
rect 18161 1670 18240 1686
rect 18272 1686 18444 1688
rect 18272 1670 18351 1686
rect 18358 1684 18388 1686
rect 17936 1648 17965 1658
rect 17979 1648 18008 1658
rect 18023 1648 18053 1662
rect 18096 1648 18139 1662
rect 18161 1658 18351 1670
rect 18416 1666 18422 1686
rect 18146 1648 18176 1658
rect 18177 1648 18335 1658
rect 18339 1648 18369 1658
rect 18373 1648 18403 1662
rect 18431 1648 18444 1686
rect 18516 1700 18545 1716
rect 18516 1692 18551 1700
rect 18516 1666 18517 1692
rect 18524 1666 18551 1692
rect 18459 1648 18489 1662
rect 18516 1658 18551 1666
rect 18516 1648 18545 1658
rect -1 1642 18545 1648
rect 0 1634 18545 1642
rect 15 1604 28 1634
rect 43 1620 73 1634
rect 116 1620 159 1634
rect 166 1620 386 1634
rect 393 1620 423 1634
rect 83 1606 98 1618
rect 117 1606 130 1620
rect 198 1616 351 1620
rect 80 1604 102 1606
rect 180 1604 372 1616
rect 451 1604 464 1634
rect 479 1620 509 1634
rect 546 1604 565 1634
rect 580 1604 586 1634
rect 595 1604 608 1634
rect 623 1620 653 1634
rect 696 1620 739 1634
rect 746 1620 966 1634
rect 973 1620 1003 1634
rect 663 1606 678 1618
rect 697 1606 710 1620
rect 778 1616 931 1620
rect 660 1604 682 1606
rect 760 1604 952 1616
rect 1031 1604 1044 1634
rect 1059 1620 1089 1634
rect 1126 1604 1145 1634
rect 1160 1604 1166 1634
rect 1175 1604 1188 1634
rect 1203 1620 1233 1634
rect 1276 1620 1319 1634
rect 1326 1620 1546 1634
rect 1553 1620 1583 1634
rect 1243 1606 1258 1618
rect 1277 1606 1290 1620
rect 1358 1616 1511 1620
rect 1240 1604 1262 1606
rect 1340 1604 1532 1616
rect 1611 1604 1624 1634
rect 1639 1620 1669 1634
rect 1706 1604 1725 1634
rect 1740 1604 1746 1634
rect 1755 1604 1768 1634
rect 1783 1620 1813 1634
rect 1856 1620 1899 1634
rect 1906 1620 2126 1634
rect 2133 1620 2163 1634
rect 1823 1606 1838 1618
rect 1857 1606 1870 1620
rect 1938 1616 2091 1620
rect 1820 1604 1842 1606
rect 1920 1604 2112 1616
rect 2191 1604 2204 1634
rect 2219 1620 2249 1634
rect 2286 1604 2305 1634
rect 2320 1604 2326 1634
rect 2335 1604 2348 1634
rect 2363 1620 2393 1634
rect 2436 1620 2479 1634
rect 2486 1620 2706 1634
rect 2713 1620 2743 1634
rect 2403 1606 2418 1618
rect 2437 1606 2450 1620
rect 2518 1616 2671 1620
rect 2400 1604 2422 1606
rect 2500 1604 2692 1616
rect 2771 1604 2784 1634
rect 2799 1620 2829 1634
rect 2866 1604 2885 1634
rect 2900 1604 2906 1634
rect 2915 1604 2928 1634
rect 2943 1620 2973 1634
rect 3016 1620 3059 1634
rect 3066 1620 3286 1634
rect 3293 1620 3323 1634
rect 2983 1606 2998 1618
rect 3017 1606 3030 1620
rect 3098 1616 3251 1620
rect 2980 1604 3002 1606
rect 3080 1604 3272 1616
rect 3351 1604 3364 1634
rect 3379 1620 3409 1634
rect 3446 1604 3465 1634
rect 3480 1604 3486 1634
rect 3495 1604 3508 1634
rect 3523 1620 3553 1634
rect 3596 1620 3639 1634
rect 3646 1620 3866 1634
rect 3873 1620 3903 1634
rect 3563 1606 3578 1618
rect 3597 1606 3610 1620
rect 3678 1616 3831 1620
rect 3560 1604 3582 1606
rect 3660 1604 3852 1616
rect 3931 1604 3944 1634
rect 3959 1620 3989 1634
rect 4026 1604 4045 1634
rect 4060 1604 4066 1634
rect 4075 1604 4088 1634
rect 4103 1620 4133 1634
rect 4176 1620 4219 1634
rect 4226 1620 4446 1634
rect 4453 1620 4483 1634
rect 4143 1606 4158 1618
rect 4177 1606 4190 1620
rect 4258 1616 4411 1620
rect 4140 1604 4162 1606
rect 4240 1604 4432 1616
rect 4511 1604 4524 1634
rect 4539 1620 4569 1634
rect 4606 1604 4625 1634
rect 4640 1604 4646 1634
rect 4655 1604 4668 1634
rect 4683 1620 4713 1634
rect 4756 1620 4799 1634
rect 4806 1620 5026 1634
rect 5033 1620 5063 1634
rect 4723 1606 4738 1618
rect 4757 1606 4770 1620
rect 4838 1616 4991 1620
rect 4720 1604 4742 1606
rect 4820 1604 5012 1616
rect 5091 1604 5104 1634
rect 5119 1620 5149 1634
rect 5186 1604 5205 1634
rect 5220 1604 5226 1634
rect 5235 1604 5248 1634
rect 5263 1620 5293 1634
rect 5336 1620 5379 1634
rect 5386 1620 5606 1634
rect 5613 1620 5643 1634
rect 5303 1606 5318 1618
rect 5337 1606 5350 1620
rect 5418 1616 5571 1620
rect 5300 1604 5322 1606
rect 5400 1604 5592 1616
rect 5671 1604 5684 1634
rect 5699 1620 5729 1634
rect 5766 1604 5785 1634
rect 5800 1604 5806 1634
rect 5815 1604 5828 1634
rect 5843 1620 5873 1634
rect 5916 1620 5959 1634
rect 5966 1620 6186 1634
rect 6193 1620 6223 1634
rect 5883 1606 5898 1618
rect 5917 1606 5930 1620
rect 5998 1616 6151 1620
rect 5880 1604 5902 1606
rect 5980 1604 6172 1616
rect 6251 1604 6264 1634
rect 6279 1620 6309 1634
rect 6346 1604 6365 1634
rect 6380 1604 6386 1634
rect 6395 1604 6408 1634
rect 6423 1620 6453 1634
rect 6496 1620 6539 1634
rect 6546 1620 6766 1634
rect 6773 1620 6803 1634
rect 6463 1606 6478 1618
rect 6497 1606 6510 1620
rect 6578 1616 6731 1620
rect 6460 1604 6482 1606
rect 6560 1604 6752 1616
rect 6831 1604 6844 1634
rect 6859 1620 6889 1634
rect 6926 1604 6945 1634
rect 6960 1604 6966 1634
rect 6975 1604 6988 1634
rect 7003 1620 7033 1634
rect 7076 1620 7119 1634
rect 7126 1620 7346 1634
rect 7353 1620 7383 1634
rect 7043 1606 7058 1618
rect 7077 1606 7090 1620
rect 7158 1616 7311 1620
rect 7040 1604 7062 1606
rect 7140 1604 7332 1616
rect 7411 1604 7424 1634
rect 7439 1620 7469 1634
rect 7506 1604 7525 1634
rect 7540 1604 7546 1634
rect 7555 1604 7568 1634
rect 7583 1620 7613 1634
rect 7656 1620 7699 1634
rect 7706 1620 7926 1634
rect 7933 1620 7963 1634
rect 7623 1606 7638 1618
rect 7657 1606 7670 1620
rect 7738 1616 7891 1620
rect 7620 1604 7642 1606
rect 7720 1604 7912 1616
rect 7991 1604 8004 1634
rect 8019 1620 8049 1634
rect 8086 1604 8105 1634
rect 8120 1604 8126 1634
rect 8135 1604 8148 1634
rect 8163 1620 8193 1634
rect 8236 1620 8279 1634
rect 8286 1620 8506 1634
rect 8513 1620 8543 1634
rect 8203 1606 8218 1618
rect 8237 1606 8250 1620
rect 8318 1616 8471 1620
rect 8200 1604 8222 1606
rect 8300 1604 8492 1616
rect 8571 1604 8584 1634
rect 8599 1620 8629 1634
rect 8666 1604 8685 1634
rect 8700 1604 8706 1634
rect 8715 1604 8728 1634
rect 8743 1620 8773 1634
rect 8816 1620 8859 1634
rect 8866 1620 9086 1634
rect 9093 1620 9123 1634
rect 8783 1606 8798 1618
rect 8817 1606 8830 1620
rect 8898 1616 9051 1620
rect 8780 1604 8802 1606
rect 8880 1604 9072 1616
rect 9151 1604 9164 1634
rect 9179 1620 9209 1634
rect 9246 1604 9265 1634
rect 9280 1604 9286 1634
rect 9295 1604 9308 1634
rect 9323 1620 9353 1634
rect 9396 1620 9439 1634
rect 9446 1620 9666 1634
rect 9673 1620 9703 1634
rect 9363 1606 9378 1618
rect 9397 1606 9410 1620
rect 9478 1616 9631 1620
rect 9360 1604 9382 1606
rect 9460 1604 9652 1616
rect 9731 1604 9744 1634
rect 9759 1620 9789 1634
rect 9826 1604 9845 1634
rect 9860 1604 9866 1634
rect 9875 1604 9888 1634
rect 9903 1620 9933 1634
rect 9976 1620 10019 1634
rect 10026 1620 10246 1634
rect 10253 1620 10283 1634
rect 9943 1606 9958 1618
rect 9977 1606 9990 1620
rect 10058 1616 10211 1620
rect 9940 1604 9962 1606
rect 10040 1604 10232 1616
rect 10311 1604 10324 1634
rect 10339 1620 10369 1634
rect 10406 1604 10425 1634
rect 10440 1604 10446 1634
rect 10455 1604 10468 1634
rect 10483 1620 10513 1634
rect 10556 1620 10599 1634
rect 10606 1620 10826 1634
rect 10833 1620 10863 1634
rect 10523 1606 10538 1618
rect 10557 1606 10570 1620
rect 10638 1616 10791 1620
rect 10520 1604 10542 1606
rect 10620 1604 10812 1616
rect 10891 1604 10904 1634
rect 10919 1620 10949 1634
rect 10986 1604 11005 1634
rect 11020 1604 11026 1634
rect 11035 1604 11048 1634
rect 11063 1620 11093 1634
rect 11136 1620 11179 1634
rect 11186 1620 11406 1634
rect 11413 1620 11443 1634
rect 11103 1606 11118 1618
rect 11137 1606 11150 1620
rect 11218 1616 11371 1620
rect 11100 1604 11122 1606
rect 11200 1604 11392 1616
rect 11471 1604 11484 1634
rect 11499 1620 11529 1634
rect 11566 1604 11585 1634
rect 11600 1604 11606 1634
rect 11615 1604 11628 1634
rect 11643 1620 11673 1634
rect 11716 1620 11759 1634
rect 11766 1620 11986 1634
rect 11993 1620 12023 1634
rect 11683 1606 11698 1618
rect 11717 1606 11730 1620
rect 11798 1616 11951 1620
rect 11680 1604 11702 1606
rect 11780 1604 11972 1616
rect 12051 1604 12064 1634
rect 12079 1620 12109 1634
rect 12146 1604 12165 1634
rect 12180 1604 12186 1634
rect 12195 1604 12208 1634
rect 12223 1620 12253 1634
rect 12296 1620 12339 1634
rect 12346 1620 12566 1634
rect 12573 1620 12603 1634
rect 12263 1606 12278 1618
rect 12297 1606 12310 1620
rect 12378 1616 12531 1620
rect 12260 1604 12282 1606
rect 12360 1604 12552 1616
rect 12631 1604 12644 1634
rect 12659 1620 12689 1634
rect 12726 1604 12745 1634
rect 12760 1604 12766 1634
rect 12775 1604 12788 1634
rect 12803 1620 12833 1634
rect 12876 1620 12919 1634
rect 12926 1620 13146 1634
rect 13153 1620 13183 1634
rect 12843 1606 12858 1618
rect 12877 1606 12890 1620
rect 12958 1616 13111 1620
rect 12840 1604 12862 1606
rect 12940 1604 13132 1616
rect 13211 1604 13224 1634
rect 13239 1620 13269 1634
rect 13306 1604 13325 1634
rect 13340 1604 13346 1634
rect 13355 1604 13368 1634
rect 13383 1620 13413 1634
rect 13456 1620 13499 1634
rect 13506 1620 13726 1634
rect 13733 1620 13763 1634
rect 13423 1606 13438 1618
rect 13457 1606 13470 1620
rect 13538 1616 13691 1620
rect 13420 1604 13442 1606
rect 13520 1604 13712 1616
rect 13791 1604 13804 1634
rect 13819 1620 13849 1634
rect 13886 1604 13905 1634
rect 13920 1604 13926 1634
rect 13935 1604 13948 1634
rect 13963 1620 13993 1634
rect 14036 1620 14079 1634
rect 14086 1620 14306 1634
rect 14313 1620 14343 1634
rect 14003 1606 14018 1618
rect 14037 1606 14050 1620
rect 14118 1616 14271 1620
rect 14000 1604 14022 1606
rect 14100 1604 14292 1616
rect 14371 1604 14384 1634
rect 14399 1620 14429 1634
rect 14466 1604 14485 1634
rect 14500 1604 14506 1634
rect 14515 1604 14528 1634
rect 14543 1620 14573 1634
rect 14616 1620 14659 1634
rect 14666 1620 14886 1634
rect 14893 1620 14923 1634
rect 14583 1606 14598 1618
rect 14617 1606 14630 1620
rect 14698 1616 14851 1620
rect 14580 1604 14602 1606
rect 14680 1604 14872 1616
rect 14951 1604 14964 1634
rect 14979 1620 15009 1634
rect 15046 1604 15065 1634
rect 15080 1604 15086 1634
rect 15095 1604 15108 1634
rect 15123 1620 15153 1634
rect 15196 1620 15239 1634
rect 15246 1620 15466 1634
rect 15473 1620 15503 1634
rect 15163 1606 15178 1618
rect 15197 1606 15210 1620
rect 15278 1616 15431 1620
rect 15160 1604 15182 1606
rect 15260 1604 15452 1616
rect 15531 1604 15544 1634
rect 15559 1620 15589 1634
rect 15626 1604 15645 1634
rect 15660 1604 15666 1634
rect 15675 1604 15688 1634
rect 15703 1620 15733 1634
rect 15776 1620 15819 1634
rect 15826 1620 16046 1634
rect 16053 1620 16083 1634
rect 15743 1606 15758 1618
rect 15777 1606 15790 1620
rect 15858 1616 16011 1620
rect 15740 1604 15762 1606
rect 15840 1604 16032 1616
rect 16111 1604 16124 1634
rect 16139 1620 16169 1634
rect 16206 1604 16225 1634
rect 16240 1604 16246 1634
rect 16255 1604 16268 1634
rect 16283 1620 16313 1634
rect 16356 1620 16399 1634
rect 16406 1620 16626 1634
rect 16633 1620 16663 1634
rect 16323 1606 16338 1618
rect 16357 1606 16370 1620
rect 16438 1616 16591 1620
rect 16320 1604 16342 1606
rect 16420 1604 16612 1616
rect 16691 1604 16704 1634
rect 16719 1620 16749 1634
rect 16786 1604 16805 1634
rect 16820 1604 16826 1634
rect 16835 1604 16848 1634
rect 16863 1620 16893 1634
rect 16936 1620 16979 1634
rect 16986 1620 17206 1634
rect 17213 1620 17243 1634
rect 16903 1606 16918 1618
rect 16937 1606 16950 1620
rect 17018 1616 17171 1620
rect 16900 1604 16922 1606
rect 17000 1604 17192 1616
rect 17271 1604 17284 1634
rect 17299 1620 17329 1634
rect 17366 1604 17385 1634
rect 17400 1604 17406 1634
rect 17415 1604 17428 1634
rect 17443 1620 17473 1634
rect 17516 1620 17559 1634
rect 17566 1620 17786 1634
rect 17793 1620 17823 1634
rect 17483 1606 17498 1618
rect 17517 1606 17530 1620
rect 17598 1616 17751 1620
rect 17480 1604 17502 1606
rect 17580 1604 17772 1616
rect 17851 1604 17864 1634
rect 17879 1620 17909 1634
rect 17946 1604 17965 1634
rect 17980 1604 17986 1634
rect 17995 1604 18008 1634
rect 18023 1620 18053 1634
rect 18096 1620 18139 1634
rect 18146 1620 18366 1634
rect 18373 1620 18403 1634
rect 18063 1606 18078 1618
rect 18097 1606 18110 1620
rect 18178 1616 18331 1620
rect 18060 1604 18082 1606
rect 18160 1604 18352 1616
rect 18431 1604 18444 1634
rect 18459 1620 18489 1634
rect 18532 1604 18545 1634
rect 0 1590 18545 1604
rect 15 1520 28 1590
rect 80 1586 102 1590
rect 73 1564 102 1578
rect 155 1564 171 1578
rect 209 1574 215 1576
rect 222 1574 330 1590
rect 337 1574 343 1576
rect 351 1574 366 1590
rect 432 1584 451 1587
rect 73 1562 171 1564
rect 198 1562 366 1574
rect 381 1564 397 1578
rect 432 1565 454 1584
rect 464 1578 480 1579
rect 463 1576 480 1578
rect 464 1571 480 1576
rect 454 1564 460 1565
rect 463 1564 492 1571
rect 381 1563 492 1564
rect 381 1562 498 1563
rect 57 1554 108 1562
rect 155 1554 189 1562
rect 57 1542 82 1554
rect 89 1542 108 1554
rect 162 1552 189 1554
rect 198 1552 419 1562
rect 454 1559 460 1562
rect 162 1548 419 1552
rect 57 1534 108 1542
rect 155 1534 419 1548
rect 463 1554 498 1562
rect 9 1486 28 1520
rect 73 1526 102 1534
rect 73 1520 90 1526
rect 73 1518 107 1520
rect 155 1518 171 1534
rect 172 1524 380 1534
rect 381 1524 397 1534
rect 445 1530 460 1545
rect 463 1542 464 1554
rect 471 1542 498 1554
rect 463 1534 498 1542
rect 463 1533 492 1534
rect 183 1520 397 1524
rect 198 1518 397 1520
rect 432 1520 445 1530
rect 463 1520 480 1533
rect 432 1518 480 1520
rect 74 1514 107 1518
rect 70 1512 107 1514
rect 70 1511 137 1512
rect 70 1506 101 1511
rect 107 1506 137 1511
rect 70 1502 137 1506
rect 43 1499 137 1502
rect 43 1492 92 1499
rect 43 1486 73 1492
rect 92 1487 97 1492
rect 9 1470 89 1486
rect 101 1478 137 1499
rect 198 1494 387 1518
rect 432 1517 479 1518
rect 445 1512 479 1517
rect 213 1491 387 1494
rect 206 1488 387 1491
rect 415 1511 479 1512
rect 9 1468 28 1470
rect 43 1468 77 1470
rect 9 1452 89 1468
rect 9 1446 28 1452
rect -1 1430 28 1446
rect 43 1436 73 1452
rect 101 1430 107 1478
rect 110 1472 129 1478
rect 144 1472 174 1480
rect 110 1464 174 1472
rect 110 1448 190 1464
rect 206 1457 268 1488
rect 284 1457 346 1488
rect 415 1486 464 1511
rect 479 1486 509 1502
rect 378 1472 408 1480
rect 415 1478 525 1486
rect 378 1464 423 1472
rect 110 1446 129 1448
rect 144 1446 190 1448
rect 110 1430 190 1446
rect 217 1444 252 1457
rect 293 1454 330 1457
rect 293 1452 335 1454
rect 222 1441 252 1444
rect 231 1437 238 1441
rect 238 1436 239 1437
rect 197 1430 207 1436
rect -7 1422 34 1430
rect -7 1396 8 1422
rect 15 1396 34 1422
rect 98 1418 129 1430
rect 144 1418 247 1430
rect 259 1420 285 1446
rect 300 1441 330 1452
rect 362 1448 424 1464
rect 362 1446 408 1448
rect 362 1430 424 1446
rect 436 1430 442 1478
rect 445 1470 525 1478
rect 445 1468 464 1470
rect 479 1468 513 1470
rect 445 1452 525 1468
rect 445 1430 464 1452
rect 479 1436 509 1452
rect 537 1446 543 1520
rect 546 1446 565 1590
rect 580 1446 586 1590
rect 595 1520 608 1590
rect 660 1586 682 1590
rect 653 1564 682 1578
rect 735 1564 751 1578
rect 789 1574 795 1576
rect 802 1574 910 1590
rect 917 1574 923 1576
rect 931 1574 946 1590
rect 1012 1584 1031 1587
rect 653 1562 751 1564
rect 778 1562 946 1574
rect 961 1564 977 1578
rect 1012 1565 1034 1584
rect 1044 1578 1060 1579
rect 1043 1576 1060 1578
rect 1044 1571 1060 1576
rect 1034 1564 1040 1565
rect 1043 1564 1072 1571
rect 961 1563 1072 1564
rect 961 1562 1078 1563
rect 637 1554 688 1562
rect 735 1554 769 1562
rect 637 1542 662 1554
rect 669 1542 688 1554
rect 742 1552 769 1554
rect 778 1552 999 1562
rect 1034 1559 1040 1562
rect 742 1548 999 1552
rect 637 1534 688 1542
rect 735 1534 999 1548
rect 1043 1554 1078 1562
rect 589 1486 608 1520
rect 653 1526 682 1534
rect 653 1520 670 1526
rect 653 1518 687 1520
rect 735 1518 751 1534
rect 752 1524 960 1534
rect 961 1524 977 1534
rect 1025 1530 1040 1545
rect 1043 1542 1044 1554
rect 1051 1542 1078 1554
rect 1043 1534 1078 1542
rect 1043 1533 1072 1534
rect 763 1520 977 1524
rect 778 1518 977 1520
rect 1012 1520 1025 1530
rect 1043 1520 1060 1533
rect 1012 1518 1060 1520
rect 654 1514 687 1518
rect 650 1512 687 1514
rect 650 1511 717 1512
rect 650 1506 681 1511
rect 687 1506 717 1511
rect 650 1502 717 1506
rect 623 1499 717 1502
rect 623 1492 672 1499
rect 623 1486 653 1492
rect 672 1487 677 1492
rect 589 1470 669 1486
rect 681 1478 717 1499
rect 778 1494 967 1518
rect 1012 1517 1059 1518
rect 1025 1512 1059 1517
rect 793 1491 967 1494
rect 786 1488 967 1491
rect 995 1511 1059 1512
rect 589 1468 608 1470
rect 623 1468 657 1470
rect 589 1452 669 1468
rect 589 1446 608 1452
rect 305 1420 408 1430
rect 259 1418 408 1420
rect 429 1418 464 1430
rect 98 1416 260 1418
rect 110 1396 129 1416
rect 144 1414 174 1416
rect -7 1388 34 1396
rect 116 1392 129 1396
rect 181 1400 260 1416
rect 292 1416 464 1418
rect 292 1400 371 1416
rect 378 1414 408 1416
rect -1 1378 28 1388
rect 43 1378 73 1392
rect 116 1378 159 1392
rect 181 1388 371 1400
rect 436 1396 442 1416
rect 166 1378 196 1388
rect 197 1378 355 1388
rect 359 1378 389 1388
rect 393 1378 423 1392
rect 451 1378 464 1416
rect 536 1430 565 1446
rect 579 1430 608 1446
rect 623 1436 653 1452
rect 681 1430 687 1478
rect 690 1472 709 1478
rect 724 1472 754 1480
rect 690 1464 754 1472
rect 690 1448 770 1464
rect 786 1457 848 1488
rect 864 1457 926 1488
rect 995 1486 1044 1511
rect 1059 1486 1089 1502
rect 958 1472 988 1480
rect 995 1478 1105 1486
rect 958 1464 1003 1472
rect 690 1446 709 1448
rect 724 1446 770 1448
rect 690 1430 770 1446
rect 797 1444 832 1457
rect 873 1454 910 1457
rect 873 1452 915 1454
rect 802 1441 832 1444
rect 811 1437 818 1441
rect 818 1436 819 1437
rect 777 1430 787 1436
rect 536 1422 571 1430
rect 536 1396 537 1422
rect 544 1396 571 1422
rect 479 1378 509 1392
rect 536 1388 571 1396
rect 573 1422 614 1430
rect 573 1396 588 1422
rect 595 1396 614 1422
rect 678 1418 709 1430
rect 724 1418 827 1430
rect 839 1420 865 1446
rect 880 1441 910 1452
rect 942 1448 1004 1464
rect 942 1446 988 1448
rect 942 1430 1004 1446
rect 1016 1430 1022 1478
rect 1025 1470 1105 1478
rect 1025 1468 1044 1470
rect 1059 1468 1093 1470
rect 1025 1452 1105 1468
rect 1025 1430 1044 1452
rect 1059 1436 1089 1452
rect 1117 1446 1123 1520
rect 1126 1446 1145 1590
rect 1160 1446 1166 1590
rect 1175 1520 1188 1590
rect 1240 1586 1262 1590
rect 1233 1564 1262 1578
rect 1315 1564 1331 1578
rect 1369 1574 1375 1576
rect 1382 1574 1490 1590
rect 1497 1574 1503 1576
rect 1511 1574 1526 1590
rect 1592 1584 1611 1587
rect 1233 1562 1331 1564
rect 1358 1562 1526 1574
rect 1541 1564 1557 1578
rect 1592 1565 1614 1584
rect 1624 1578 1640 1579
rect 1623 1576 1640 1578
rect 1624 1571 1640 1576
rect 1614 1564 1620 1565
rect 1623 1564 1652 1571
rect 1541 1563 1652 1564
rect 1541 1562 1658 1563
rect 1217 1554 1268 1562
rect 1315 1554 1349 1562
rect 1217 1542 1242 1554
rect 1249 1542 1268 1554
rect 1322 1552 1349 1554
rect 1358 1552 1579 1562
rect 1614 1559 1620 1562
rect 1322 1548 1579 1552
rect 1217 1534 1268 1542
rect 1315 1534 1579 1548
rect 1623 1554 1658 1562
rect 1169 1486 1188 1520
rect 1233 1526 1262 1534
rect 1233 1520 1250 1526
rect 1233 1518 1267 1520
rect 1315 1518 1331 1534
rect 1332 1524 1540 1534
rect 1541 1524 1557 1534
rect 1605 1530 1620 1545
rect 1623 1542 1624 1554
rect 1631 1542 1658 1554
rect 1623 1534 1658 1542
rect 1623 1533 1652 1534
rect 1343 1520 1557 1524
rect 1358 1518 1557 1520
rect 1592 1520 1605 1530
rect 1623 1520 1640 1533
rect 1592 1518 1640 1520
rect 1234 1514 1267 1518
rect 1230 1512 1267 1514
rect 1230 1511 1297 1512
rect 1230 1506 1261 1511
rect 1267 1506 1297 1511
rect 1230 1502 1297 1506
rect 1203 1499 1297 1502
rect 1203 1492 1252 1499
rect 1203 1486 1233 1492
rect 1252 1487 1257 1492
rect 1169 1470 1249 1486
rect 1261 1478 1297 1499
rect 1358 1494 1547 1518
rect 1592 1517 1639 1518
rect 1605 1512 1639 1517
rect 1373 1491 1547 1494
rect 1366 1488 1547 1491
rect 1575 1511 1639 1512
rect 1169 1468 1188 1470
rect 1203 1468 1237 1470
rect 1169 1452 1249 1468
rect 1169 1446 1188 1452
rect 885 1420 988 1430
rect 839 1418 988 1420
rect 1009 1418 1044 1430
rect 678 1416 840 1418
rect 690 1396 709 1416
rect 724 1414 754 1416
rect 573 1388 614 1396
rect 696 1392 709 1396
rect 761 1400 840 1416
rect 872 1416 1044 1418
rect 872 1400 951 1416
rect 958 1414 988 1416
rect 536 1378 565 1388
rect 579 1378 608 1388
rect 623 1378 653 1392
rect 696 1378 739 1392
rect 761 1388 951 1400
rect 1016 1396 1022 1416
rect 746 1378 776 1388
rect 777 1378 935 1388
rect 939 1378 969 1388
rect 973 1378 1003 1392
rect 1031 1378 1044 1416
rect 1116 1430 1145 1446
rect 1159 1430 1188 1446
rect 1203 1436 1233 1452
rect 1261 1430 1267 1478
rect 1270 1472 1289 1478
rect 1304 1472 1334 1480
rect 1270 1464 1334 1472
rect 1270 1448 1350 1464
rect 1366 1457 1428 1488
rect 1444 1457 1506 1488
rect 1575 1486 1624 1511
rect 1639 1486 1669 1502
rect 1538 1472 1568 1480
rect 1575 1478 1685 1486
rect 1538 1464 1583 1472
rect 1270 1446 1289 1448
rect 1304 1446 1350 1448
rect 1270 1430 1350 1446
rect 1377 1444 1412 1457
rect 1453 1454 1490 1457
rect 1453 1452 1495 1454
rect 1382 1441 1412 1444
rect 1391 1437 1398 1441
rect 1398 1436 1399 1437
rect 1357 1430 1367 1436
rect 1116 1422 1151 1430
rect 1116 1396 1117 1422
rect 1124 1396 1151 1422
rect 1059 1378 1089 1392
rect 1116 1388 1151 1396
rect 1153 1422 1194 1430
rect 1153 1396 1168 1422
rect 1175 1396 1194 1422
rect 1258 1418 1289 1430
rect 1304 1418 1407 1430
rect 1419 1420 1445 1446
rect 1460 1441 1490 1452
rect 1522 1448 1584 1464
rect 1522 1446 1568 1448
rect 1522 1430 1584 1446
rect 1596 1430 1602 1478
rect 1605 1470 1685 1478
rect 1605 1468 1624 1470
rect 1639 1468 1673 1470
rect 1605 1452 1685 1468
rect 1605 1430 1624 1452
rect 1639 1436 1669 1452
rect 1697 1446 1703 1520
rect 1706 1446 1725 1590
rect 1740 1446 1746 1590
rect 1755 1520 1768 1590
rect 1820 1586 1842 1590
rect 1813 1564 1842 1578
rect 1895 1564 1911 1578
rect 1949 1574 1955 1576
rect 1962 1574 2070 1590
rect 2077 1574 2083 1576
rect 2091 1574 2106 1590
rect 2172 1584 2191 1587
rect 1813 1562 1911 1564
rect 1938 1562 2106 1574
rect 2121 1564 2137 1578
rect 2172 1565 2194 1584
rect 2204 1578 2220 1579
rect 2203 1576 2220 1578
rect 2204 1571 2220 1576
rect 2194 1564 2200 1565
rect 2203 1564 2232 1571
rect 2121 1563 2232 1564
rect 2121 1562 2238 1563
rect 1797 1554 1848 1562
rect 1895 1554 1929 1562
rect 1797 1542 1822 1554
rect 1829 1542 1848 1554
rect 1902 1552 1929 1554
rect 1938 1552 2159 1562
rect 2194 1559 2200 1562
rect 1902 1548 2159 1552
rect 1797 1534 1848 1542
rect 1895 1534 2159 1548
rect 2203 1554 2238 1562
rect 1749 1486 1768 1520
rect 1813 1526 1842 1534
rect 1813 1520 1830 1526
rect 1813 1518 1847 1520
rect 1895 1518 1911 1534
rect 1912 1524 2120 1534
rect 2121 1524 2137 1534
rect 2185 1530 2200 1545
rect 2203 1542 2204 1554
rect 2211 1542 2238 1554
rect 2203 1534 2238 1542
rect 2203 1533 2232 1534
rect 1923 1520 2137 1524
rect 1938 1518 2137 1520
rect 2172 1520 2185 1530
rect 2203 1520 2220 1533
rect 2172 1518 2220 1520
rect 1814 1514 1847 1518
rect 1810 1512 1847 1514
rect 1810 1511 1877 1512
rect 1810 1506 1841 1511
rect 1847 1506 1877 1511
rect 1810 1502 1877 1506
rect 1783 1499 1877 1502
rect 1783 1492 1832 1499
rect 1783 1486 1813 1492
rect 1832 1487 1837 1492
rect 1749 1470 1829 1486
rect 1841 1478 1877 1499
rect 1938 1494 2127 1518
rect 2172 1517 2219 1518
rect 2185 1512 2219 1517
rect 1953 1491 2127 1494
rect 1946 1488 2127 1491
rect 2155 1511 2219 1512
rect 1749 1468 1768 1470
rect 1783 1468 1817 1470
rect 1749 1452 1829 1468
rect 1749 1446 1768 1452
rect 1465 1420 1568 1430
rect 1419 1418 1568 1420
rect 1589 1418 1624 1430
rect 1258 1416 1420 1418
rect 1270 1396 1289 1416
rect 1304 1414 1334 1416
rect 1153 1388 1194 1396
rect 1276 1392 1289 1396
rect 1341 1400 1420 1416
rect 1452 1416 1624 1418
rect 1452 1400 1531 1416
rect 1538 1414 1568 1416
rect 1116 1378 1145 1388
rect 1159 1378 1188 1388
rect 1203 1378 1233 1392
rect 1276 1378 1319 1392
rect 1341 1388 1531 1400
rect 1596 1396 1602 1416
rect 1326 1378 1356 1388
rect 1357 1378 1515 1388
rect 1519 1378 1549 1388
rect 1553 1378 1583 1392
rect 1611 1378 1624 1416
rect 1696 1430 1725 1446
rect 1739 1430 1768 1446
rect 1783 1436 1813 1452
rect 1841 1430 1847 1478
rect 1850 1472 1869 1478
rect 1884 1472 1914 1480
rect 1850 1464 1914 1472
rect 1850 1448 1930 1464
rect 1946 1457 2008 1488
rect 2024 1457 2086 1488
rect 2155 1486 2204 1511
rect 2219 1486 2249 1502
rect 2118 1472 2148 1480
rect 2155 1478 2265 1486
rect 2118 1464 2163 1472
rect 1850 1446 1869 1448
rect 1884 1446 1930 1448
rect 1850 1430 1930 1446
rect 1957 1444 1992 1457
rect 2033 1454 2070 1457
rect 2033 1452 2075 1454
rect 1962 1441 1992 1444
rect 1971 1437 1978 1441
rect 1978 1436 1979 1437
rect 1937 1430 1947 1436
rect 1696 1422 1731 1430
rect 1696 1396 1697 1422
rect 1704 1396 1731 1422
rect 1639 1378 1669 1392
rect 1696 1388 1731 1396
rect 1733 1422 1774 1430
rect 1733 1396 1748 1422
rect 1755 1396 1774 1422
rect 1838 1418 1869 1430
rect 1884 1418 1987 1430
rect 1999 1420 2025 1446
rect 2040 1441 2070 1452
rect 2102 1448 2164 1464
rect 2102 1446 2148 1448
rect 2102 1430 2164 1446
rect 2176 1430 2182 1478
rect 2185 1470 2265 1478
rect 2185 1468 2204 1470
rect 2219 1468 2253 1470
rect 2185 1452 2265 1468
rect 2185 1430 2204 1452
rect 2219 1436 2249 1452
rect 2277 1446 2283 1520
rect 2286 1446 2305 1590
rect 2320 1446 2326 1590
rect 2335 1520 2348 1590
rect 2400 1586 2422 1590
rect 2393 1564 2422 1578
rect 2475 1564 2491 1578
rect 2529 1574 2535 1576
rect 2542 1574 2650 1590
rect 2657 1574 2663 1576
rect 2671 1574 2686 1590
rect 2752 1584 2771 1587
rect 2393 1562 2491 1564
rect 2518 1562 2686 1574
rect 2701 1564 2717 1578
rect 2752 1565 2774 1584
rect 2784 1578 2800 1579
rect 2783 1576 2800 1578
rect 2784 1571 2800 1576
rect 2774 1564 2780 1565
rect 2783 1564 2812 1571
rect 2701 1563 2812 1564
rect 2701 1562 2818 1563
rect 2377 1554 2428 1562
rect 2475 1554 2509 1562
rect 2377 1542 2402 1554
rect 2409 1542 2428 1554
rect 2482 1552 2509 1554
rect 2518 1552 2739 1562
rect 2774 1559 2780 1562
rect 2482 1548 2739 1552
rect 2377 1534 2428 1542
rect 2475 1534 2739 1548
rect 2783 1554 2818 1562
rect 2329 1486 2348 1520
rect 2393 1526 2422 1534
rect 2393 1520 2410 1526
rect 2393 1518 2427 1520
rect 2475 1518 2491 1534
rect 2492 1524 2700 1534
rect 2701 1524 2717 1534
rect 2765 1530 2780 1545
rect 2783 1542 2784 1554
rect 2791 1542 2818 1554
rect 2783 1534 2818 1542
rect 2783 1533 2812 1534
rect 2503 1520 2717 1524
rect 2518 1518 2717 1520
rect 2752 1520 2765 1530
rect 2783 1520 2800 1533
rect 2752 1518 2800 1520
rect 2394 1514 2427 1518
rect 2390 1512 2427 1514
rect 2390 1511 2457 1512
rect 2390 1506 2421 1511
rect 2427 1506 2457 1511
rect 2390 1502 2457 1506
rect 2363 1499 2457 1502
rect 2363 1492 2412 1499
rect 2363 1486 2393 1492
rect 2412 1487 2417 1492
rect 2329 1470 2409 1486
rect 2421 1478 2457 1499
rect 2518 1494 2707 1518
rect 2752 1517 2799 1518
rect 2765 1512 2799 1517
rect 2533 1491 2707 1494
rect 2526 1488 2707 1491
rect 2735 1511 2799 1512
rect 2329 1468 2348 1470
rect 2363 1468 2397 1470
rect 2329 1452 2409 1468
rect 2329 1446 2348 1452
rect 2045 1420 2148 1430
rect 1999 1418 2148 1420
rect 2169 1418 2204 1430
rect 1838 1416 2000 1418
rect 1850 1396 1869 1416
rect 1884 1414 1914 1416
rect 1733 1388 1774 1396
rect 1856 1392 1869 1396
rect 1921 1400 2000 1416
rect 2032 1416 2204 1418
rect 2032 1400 2111 1416
rect 2118 1414 2148 1416
rect 1696 1378 1725 1388
rect 1739 1378 1768 1388
rect 1783 1378 1813 1392
rect 1856 1378 1899 1392
rect 1921 1388 2111 1400
rect 2176 1396 2182 1416
rect 1906 1378 1936 1388
rect 1937 1378 2095 1388
rect 2099 1378 2129 1388
rect 2133 1378 2163 1392
rect 2191 1378 2204 1416
rect 2276 1430 2305 1446
rect 2319 1430 2348 1446
rect 2363 1436 2393 1452
rect 2421 1430 2427 1478
rect 2430 1472 2449 1478
rect 2464 1472 2494 1480
rect 2430 1464 2494 1472
rect 2430 1448 2510 1464
rect 2526 1457 2588 1488
rect 2604 1457 2666 1488
rect 2735 1486 2784 1511
rect 2799 1486 2829 1502
rect 2698 1472 2728 1480
rect 2735 1478 2845 1486
rect 2698 1464 2743 1472
rect 2430 1446 2449 1448
rect 2464 1446 2510 1448
rect 2430 1430 2510 1446
rect 2537 1444 2572 1457
rect 2613 1454 2650 1457
rect 2613 1452 2655 1454
rect 2542 1441 2572 1444
rect 2551 1437 2558 1441
rect 2558 1436 2559 1437
rect 2517 1430 2527 1436
rect 2276 1422 2311 1430
rect 2276 1396 2277 1422
rect 2284 1396 2311 1422
rect 2219 1378 2249 1392
rect 2276 1388 2311 1396
rect 2313 1422 2354 1430
rect 2313 1396 2328 1422
rect 2335 1396 2354 1422
rect 2418 1418 2449 1430
rect 2464 1418 2567 1430
rect 2579 1420 2605 1446
rect 2620 1441 2650 1452
rect 2682 1448 2744 1464
rect 2682 1446 2728 1448
rect 2682 1430 2744 1446
rect 2756 1430 2762 1478
rect 2765 1470 2845 1478
rect 2765 1468 2784 1470
rect 2799 1468 2833 1470
rect 2765 1452 2845 1468
rect 2765 1430 2784 1452
rect 2799 1436 2829 1452
rect 2857 1446 2863 1520
rect 2866 1446 2885 1590
rect 2900 1446 2906 1590
rect 2915 1520 2928 1590
rect 2980 1586 3002 1590
rect 2973 1564 3002 1578
rect 3055 1564 3071 1578
rect 3109 1574 3115 1576
rect 3122 1574 3230 1590
rect 3237 1574 3243 1576
rect 3251 1574 3266 1590
rect 3332 1584 3351 1587
rect 2973 1562 3071 1564
rect 3098 1562 3266 1574
rect 3281 1564 3297 1578
rect 3332 1565 3354 1584
rect 3364 1578 3380 1579
rect 3363 1576 3380 1578
rect 3364 1571 3380 1576
rect 3354 1564 3360 1565
rect 3363 1564 3392 1571
rect 3281 1563 3392 1564
rect 3281 1562 3398 1563
rect 2957 1554 3008 1562
rect 3055 1554 3089 1562
rect 2957 1542 2982 1554
rect 2989 1542 3008 1554
rect 3062 1552 3089 1554
rect 3098 1552 3319 1562
rect 3354 1559 3360 1562
rect 3062 1548 3319 1552
rect 2957 1534 3008 1542
rect 3055 1534 3319 1548
rect 3363 1554 3398 1562
rect 2909 1486 2928 1520
rect 2973 1526 3002 1534
rect 2973 1520 2990 1526
rect 2973 1518 3007 1520
rect 3055 1518 3071 1534
rect 3072 1524 3280 1534
rect 3281 1524 3297 1534
rect 3345 1530 3360 1545
rect 3363 1542 3364 1554
rect 3371 1542 3398 1554
rect 3363 1534 3398 1542
rect 3363 1533 3392 1534
rect 3083 1520 3297 1524
rect 3098 1518 3297 1520
rect 3332 1520 3345 1530
rect 3363 1520 3380 1533
rect 3332 1518 3380 1520
rect 2974 1514 3007 1518
rect 2970 1512 3007 1514
rect 2970 1511 3037 1512
rect 2970 1506 3001 1511
rect 3007 1506 3037 1511
rect 2970 1502 3037 1506
rect 2943 1499 3037 1502
rect 2943 1492 2992 1499
rect 2943 1486 2973 1492
rect 2992 1487 2997 1492
rect 2909 1470 2989 1486
rect 3001 1478 3037 1499
rect 3098 1494 3287 1518
rect 3332 1517 3379 1518
rect 3345 1512 3379 1517
rect 3113 1491 3287 1494
rect 3106 1488 3287 1491
rect 3315 1511 3379 1512
rect 2909 1468 2928 1470
rect 2943 1468 2977 1470
rect 2909 1452 2989 1468
rect 2909 1446 2928 1452
rect 2625 1420 2728 1430
rect 2579 1418 2728 1420
rect 2749 1418 2784 1430
rect 2418 1416 2580 1418
rect 2430 1396 2449 1416
rect 2464 1414 2494 1416
rect 2313 1388 2354 1396
rect 2436 1392 2449 1396
rect 2501 1400 2580 1416
rect 2612 1416 2784 1418
rect 2612 1400 2691 1416
rect 2698 1414 2728 1416
rect 2276 1378 2305 1388
rect 2319 1378 2348 1388
rect 2363 1378 2393 1392
rect 2436 1378 2479 1392
rect 2501 1388 2691 1400
rect 2756 1396 2762 1416
rect 2486 1378 2516 1388
rect 2517 1378 2675 1388
rect 2679 1378 2709 1388
rect 2713 1378 2743 1392
rect 2771 1378 2784 1416
rect 2856 1430 2885 1446
rect 2899 1430 2928 1446
rect 2943 1436 2973 1452
rect 3001 1430 3007 1478
rect 3010 1472 3029 1478
rect 3044 1472 3074 1480
rect 3010 1464 3074 1472
rect 3010 1448 3090 1464
rect 3106 1457 3168 1488
rect 3184 1457 3246 1488
rect 3315 1486 3364 1511
rect 3379 1486 3409 1502
rect 3278 1472 3308 1480
rect 3315 1478 3425 1486
rect 3278 1464 3323 1472
rect 3010 1446 3029 1448
rect 3044 1446 3090 1448
rect 3010 1430 3090 1446
rect 3117 1444 3152 1457
rect 3193 1454 3230 1457
rect 3193 1452 3235 1454
rect 3122 1441 3152 1444
rect 3131 1437 3138 1441
rect 3138 1436 3139 1437
rect 3097 1430 3107 1436
rect 2856 1422 2891 1430
rect 2856 1396 2857 1422
rect 2864 1396 2891 1422
rect 2799 1378 2829 1392
rect 2856 1388 2891 1396
rect 2893 1422 2934 1430
rect 2893 1396 2908 1422
rect 2915 1396 2934 1422
rect 2998 1418 3029 1430
rect 3044 1418 3147 1430
rect 3159 1420 3185 1446
rect 3200 1441 3230 1452
rect 3262 1448 3324 1464
rect 3262 1446 3308 1448
rect 3262 1430 3324 1446
rect 3336 1430 3342 1478
rect 3345 1470 3425 1478
rect 3345 1468 3364 1470
rect 3379 1468 3413 1470
rect 3345 1452 3425 1468
rect 3345 1430 3364 1452
rect 3379 1436 3409 1452
rect 3437 1446 3443 1520
rect 3446 1446 3465 1590
rect 3480 1446 3486 1590
rect 3495 1520 3508 1590
rect 3560 1586 3582 1590
rect 3553 1564 3582 1578
rect 3635 1564 3651 1578
rect 3689 1574 3695 1576
rect 3702 1574 3810 1590
rect 3817 1574 3823 1576
rect 3831 1574 3846 1590
rect 3912 1584 3931 1587
rect 3553 1562 3651 1564
rect 3678 1562 3846 1574
rect 3861 1564 3877 1578
rect 3912 1565 3934 1584
rect 3944 1578 3960 1579
rect 3943 1576 3960 1578
rect 3944 1571 3960 1576
rect 3934 1564 3940 1565
rect 3943 1564 3972 1571
rect 3861 1563 3972 1564
rect 3861 1562 3978 1563
rect 3537 1554 3588 1562
rect 3635 1554 3669 1562
rect 3537 1542 3562 1554
rect 3569 1542 3588 1554
rect 3642 1552 3669 1554
rect 3678 1552 3899 1562
rect 3934 1559 3940 1562
rect 3642 1548 3899 1552
rect 3537 1534 3588 1542
rect 3635 1534 3899 1548
rect 3943 1554 3978 1562
rect 3489 1486 3508 1520
rect 3553 1526 3582 1534
rect 3553 1520 3570 1526
rect 3553 1518 3587 1520
rect 3635 1518 3651 1534
rect 3652 1524 3860 1534
rect 3861 1524 3877 1534
rect 3925 1530 3940 1545
rect 3943 1542 3944 1554
rect 3951 1542 3978 1554
rect 3943 1534 3978 1542
rect 3943 1533 3972 1534
rect 3663 1520 3877 1524
rect 3678 1518 3877 1520
rect 3912 1520 3925 1530
rect 3943 1520 3960 1533
rect 3912 1518 3960 1520
rect 3554 1514 3587 1518
rect 3550 1512 3587 1514
rect 3550 1511 3617 1512
rect 3550 1506 3581 1511
rect 3587 1506 3617 1511
rect 3550 1502 3617 1506
rect 3523 1499 3617 1502
rect 3523 1492 3572 1499
rect 3523 1486 3553 1492
rect 3572 1487 3577 1492
rect 3489 1470 3569 1486
rect 3581 1478 3617 1499
rect 3678 1494 3867 1518
rect 3912 1517 3959 1518
rect 3925 1512 3959 1517
rect 3693 1491 3867 1494
rect 3686 1488 3867 1491
rect 3895 1511 3959 1512
rect 3489 1468 3508 1470
rect 3523 1468 3557 1470
rect 3489 1452 3569 1468
rect 3489 1446 3508 1452
rect 3205 1420 3308 1430
rect 3159 1418 3308 1420
rect 3329 1418 3364 1430
rect 2998 1416 3160 1418
rect 3010 1396 3029 1416
rect 3044 1414 3074 1416
rect 2893 1388 2934 1396
rect 3016 1392 3029 1396
rect 3081 1400 3160 1416
rect 3192 1416 3364 1418
rect 3192 1400 3271 1416
rect 3278 1414 3308 1416
rect 2856 1378 2885 1388
rect 2899 1378 2928 1388
rect 2943 1378 2973 1392
rect 3016 1378 3059 1392
rect 3081 1388 3271 1400
rect 3336 1396 3342 1416
rect 3066 1378 3096 1388
rect 3097 1378 3255 1388
rect 3259 1378 3289 1388
rect 3293 1378 3323 1392
rect 3351 1378 3364 1416
rect 3436 1430 3465 1446
rect 3479 1430 3508 1446
rect 3523 1436 3553 1452
rect 3581 1430 3587 1478
rect 3590 1472 3609 1478
rect 3624 1472 3654 1480
rect 3590 1464 3654 1472
rect 3590 1448 3670 1464
rect 3686 1457 3748 1488
rect 3764 1457 3826 1488
rect 3895 1486 3944 1511
rect 3959 1486 3989 1502
rect 3858 1472 3888 1480
rect 3895 1478 4005 1486
rect 3858 1464 3903 1472
rect 3590 1446 3609 1448
rect 3624 1446 3670 1448
rect 3590 1430 3670 1446
rect 3697 1444 3732 1457
rect 3773 1454 3810 1457
rect 3773 1452 3815 1454
rect 3702 1441 3732 1444
rect 3711 1437 3718 1441
rect 3718 1436 3719 1437
rect 3677 1430 3687 1436
rect 3436 1422 3471 1430
rect 3436 1396 3437 1422
rect 3444 1396 3471 1422
rect 3379 1378 3409 1392
rect 3436 1388 3471 1396
rect 3473 1422 3514 1430
rect 3473 1396 3488 1422
rect 3495 1396 3514 1422
rect 3578 1418 3609 1430
rect 3624 1418 3727 1430
rect 3739 1420 3765 1446
rect 3780 1441 3810 1452
rect 3842 1448 3904 1464
rect 3842 1446 3888 1448
rect 3842 1430 3904 1446
rect 3916 1430 3922 1478
rect 3925 1470 4005 1478
rect 3925 1468 3944 1470
rect 3959 1468 3993 1470
rect 3925 1452 4005 1468
rect 3925 1430 3944 1452
rect 3959 1436 3989 1452
rect 4017 1446 4023 1520
rect 4026 1446 4045 1590
rect 4060 1446 4066 1590
rect 4075 1520 4088 1590
rect 4140 1586 4162 1590
rect 4133 1564 4162 1578
rect 4215 1564 4231 1578
rect 4269 1574 4275 1576
rect 4282 1574 4390 1590
rect 4397 1574 4403 1576
rect 4411 1574 4426 1590
rect 4492 1584 4511 1587
rect 4133 1562 4231 1564
rect 4258 1562 4426 1574
rect 4441 1564 4457 1578
rect 4492 1565 4514 1584
rect 4524 1578 4540 1579
rect 4523 1576 4540 1578
rect 4524 1571 4540 1576
rect 4514 1564 4520 1565
rect 4523 1564 4552 1571
rect 4441 1563 4552 1564
rect 4441 1562 4558 1563
rect 4117 1554 4168 1562
rect 4215 1554 4249 1562
rect 4117 1542 4142 1554
rect 4149 1542 4168 1554
rect 4222 1552 4249 1554
rect 4258 1552 4479 1562
rect 4514 1559 4520 1562
rect 4222 1548 4479 1552
rect 4117 1534 4168 1542
rect 4215 1534 4479 1548
rect 4523 1554 4558 1562
rect 4069 1486 4088 1520
rect 4133 1526 4162 1534
rect 4133 1520 4150 1526
rect 4133 1518 4167 1520
rect 4215 1518 4231 1534
rect 4232 1524 4440 1534
rect 4441 1524 4457 1534
rect 4505 1530 4520 1545
rect 4523 1542 4524 1554
rect 4531 1542 4558 1554
rect 4523 1534 4558 1542
rect 4523 1533 4552 1534
rect 4243 1520 4457 1524
rect 4258 1518 4457 1520
rect 4492 1520 4505 1530
rect 4523 1520 4540 1533
rect 4492 1518 4540 1520
rect 4134 1514 4167 1518
rect 4130 1512 4167 1514
rect 4130 1511 4197 1512
rect 4130 1506 4161 1511
rect 4167 1506 4197 1511
rect 4130 1502 4197 1506
rect 4103 1499 4197 1502
rect 4103 1492 4152 1499
rect 4103 1486 4133 1492
rect 4152 1487 4157 1492
rect 4069 1470 4149 1486
rect 4161 1478 4197 1499
rect 4258 1494 4447 1518
rect 4492 1517 4539 1518
rect 4505 1512 4539 1517
rect 4273 1491 4447 1494
rect 4266 1488 4447 1491
rect 4475 1511 4539 1512
rect 4069 1468 4088 1470
rect 4103 1468 4137 1470
rect 4069 1452 4149 1468
rect 4069 1446 4088 1452
rect 3785 1420 3888 1430
rect 3739 1418 3888 1420
rect 3909 1418 3944 1430
rect 3578 1416 3740 1418
rect 3590 1396 3609 1416
rect 3624 1414 3654 1416
rect 3473 1388 3514 1396
rect 3596 1392 3609 1396
rect 3661 1400 3740 1416
rect 3772 1416 3944 1418
rect 3772 1400 3851 1416
rect 3858 1414 3888 1416
rect 3436 1378 3465 1388
rect 3479 1378 3508 1388
rect 3523 1378 3553 1392
rect 3596 1378 3639 1392
rect 3661 1388 3851 1400
rect 3916 1396 3922 1416
rect 3646 1378 3676 1388
rect 3677 1378 3835 1388
rect 3839 1378 3869 1388
rect 3873 1378 3903 1392
rect 3931 1378 3944 1416
rect 4016 1430 4045 1446
rect 4059 1430 4088 1446
rect 4103 1436 4133 1452
rect 4161 1430 4167 1478
rect 4170 1472 4189 1478
rect 4204 1472 4234 1480
rect 4170 1464 4234 1472
rect 4170 1448 4250 1464
rect 4266 1457 4328 1488
rect 4344 1457 4406 1488
rect 4475 1486 4524 1511
rect 4539 1486 4569 1502
rect 4438 1472 4468 1480
rect 4475 1478 4585 1486
rect 4438 1464 4483 1472
rect 4170 1446 4189 1448
rect 4204 1446 4250 1448
rect 4170 1430 4250 1446
rect 4277 1444 4312 1457
rect 4353 1454 4390 1457
rect 4353 1452 4395 1454
rect 4282 1441 4312 1444
rect 4291 1437 4298 1441
rect 4298 1436 4299 1437
rect 4257 1430 4267 1436
rect 4016 1422 4051 1430
rect 4016 1396 4017 1422
rect 4024 1396 4051 1422
rect 3959 1378 3989 1392
rect 4016 1388 4051 1396
rect 4053 1422 4094 1430
rect 4053 1396 4068 1422
rect 4075 1396 4094 1422
rect 4158 1418 4189 1430
rect 4204 1418 4307 1430
rect 4319 1420 4345 1446
rect 4360 1441 4390 1452
rect 4422 1448 4484 1464
rect 4422 1446 4468 1448
rect 4422 1430 4484 1446
rect 4496 1430 4502 1478
rect 4505 1470 4585 1478
rect 4505 1468 4524 1470
rect 4539 1468 4573 1470
rect 4505 1452 4585 1468
rect 4505 1430 4524 1452
rect 4539 1436 4569 1452
rect 4597 1446 4603 1520
rect 4606 1446 4625 1590
rect 4640 1446 4646 1590
rect 4655 1520 4668 1590
rect 4720 1586 4742 1590
rect 4713 1564 4742 1578
rect 4795 1564 4811 1578
rect 4849 1574 4855 1576
rect 4862 1574 4970 1590
rect 4977 1574 4983 1576
rect 4991 1574 5006 1590
rect 5072 1584 5091 1587
rect 4713 1562 4811 1564
rect 4838 1562 5006 1574
rect 5021 1564 5037 1578
rect 5072 1565 5094 1584
rect 5104 1578 5120 1579
rect 5103 1576 5120 1578
rect 5104 1571 5120 1576
rect 5094 1564 5100 1565
rect 5103 1564 5132 1571
rect 5021 1563 5132 1564
rect 5021 1562 5138 1563
rect 4697 1554 4748 1562
rect 4795 1554 4829 1562
rect 4697 1542 4722 1554
rect 4729 1542 4748 1554
rect 4802 1552 4829 1554
rect 4838 1552 5059 1562
rect 5094 1559 5100 1562
rect 4802 1548 5059 1552
rect 4697 1534 4748 1542
rect 4795 1534 5059 1548
rect 5103 1554 5138 1562
rect 4649 1486 4668 1520
rect 4713 1526 4742 1534
rect 4713 1520 4730 1526
rect 4713 1518 4747 1520
rect 4795 1518 4811 1534
rect 4812 1524 5020 1534
rect 5021 1524 5037 1534
rect 5085 1530 5100 1545
rect 5103 1542 5104 1554
rect 5111 1542 5138 1554
rect 5103 1534 5138 1542
rect 5103 1533 5132 1534
rect 4823 1520 5037 1524
rect 4838 1518 5037 1520
rect 5072 1520 5085 1530
rect 5103 1520 5120 1533
rect 5072 1518 5120 1520
rect 4714 1514 4747 1518
rect 4710 1512 4747 1514
rect 4710 1511 4777 1512
rect 4710 1506 4741 1511
rect 4747 1506 4777 1511
rect 4710 1502 4777 1506
rect 4683 1499 4777 1502
rect 4683 1492 4732 1499
rect 4683 1486 4713 1492
rect 4732 1487 4737 1492
rect 4649 1470 4729 1486
rect 4741 1478 4777 1499
rect 4838 1494 5027 1518
rect 5072 1517 5119 1518
rect 5085 1512 5119 1517
rect 4853 1491 5027 1494
rect 4846 1488 5027 1491
rect 5055 1511 5119 1512
rect 4649 1468 4668 1470
rect 4683 1468 4717 1470
rect 4649 1452 4729 1468
rect 4649 1446 4668 1452
rect 4365 1420 4468 1430
rect 4319 1418 4468 1420
rect 4489 1418 4524 1430
rect 4158 1416 4320 1418
rect 4170 1396 4189 1416
rect 4204 1414 4234 1416
rect 4053 1388 4094 1396
rect 4176 1392 4189 1396
rect 4241 1400 4320 1416
rect 4352 1416 4524 1418
rect 4352 1400 4431 1416
rect 4438 1414 4468 1416
rect 4016 1378 4045 1388
rect 4059 1378 4088 1388
rect 4103 1378 4133 1392
rect 4176 1378 4219 1392
rect 4241 1388 4431 1400
rect 4496 1396 4502 1416
rect 4226 1378 4256 1388
rect 4257 1378 4415 1388
rect 4419 1378 4449 1388
rect 4453 1378 4483 1392
rect 4511 1378 4524 1416
rect 4596 1430 4625 1446
rect 4639 1430 4668 1446
rect 4683 1436 4713 1452
rect 4741 1430 4747 1478
rect 4750 1472 4769 1478
rect 4784 1472 4814 1480
rect 4750 1464 4814 1472
rect 4750 1448 4830 1464
rect 4846 1457 4908 1488
rect 4924 1457 4986 1488
rect 5055 1486 5104 1511
rect 5119 1486 5149 1502
rect 5018 1472 5048 1480
rect 5055 1478 5165 1486
rect 5018 1464 5063 1472
rect 4750 1446 4769 1448
rect 4784 1446 4830 1448
rect 4750 1430 4830 1446
rect 4857 1444 4892 1457
rect 4933 1454 4970 1457
rect 4933 1452 4975 1454
rect 4862 1441 4892 1444
rect 4871 1437 4878 1441
rect 4878 1436 4879 1437
rect 4837 1430 4847 1436
rect 4596 1422 4631 1430
rect 4596 1396 4597 1422
rect 4604 1396 4631 1422
rect 4539 1378 4569 1392
rect 4596 1388 4631 1396
rect 4633 1422 4674 1430
rect 4633 1396 4648 1422
rect 4655 1396 4674 1422
rect 4738 1418 4769 1430
rect 4784 1418 4887 1430
rect 4899 1420 4925 1446
rect 4940 1441 4970 1452
rect 5002 1448 5064 1464
rect 5002 1446 5048 1448
rect 5002 1430 5064 1446
rect 5076 1430 5082 1478
rect 5085 1470 5165 1478
rect 5085 1468 5104 1470
rect 5119 1468 5153 1470
rect 5085 1452 5165 1468
rect 5085 1430 5104 1452
rect 5119 1436 5149 1452
rect 5177 1446 5183 1520
rect 5186 1446 5205 1590
rect 5220 1446 5226 1590
rect 5235 1520 5248 1590
rect 5300 1586 5322 1590
rect 5293 1564 5322 1578
rect 5375 1564 5391 1578
rect 5429 1574 5435 1576
rect 5442 1574 5550 1590
rect 5557 1574 5563 1576
rect 5571 1574 5586 1590
rect 5652 1584 5671 1587
rect 5293 1562 5391 1564
rect 5418 1562 5586 1574
rect 5601 1564 5617 1578
rect 5652 1565 5674 1584
rect 5684 1578 5700 1579
rect 5683 1576 5700 1578
rect 5684 1571 5700 1576
rect 5674 1564 5680 1565
rect 5683 1564 5712 1571
rect 5601 1563 5712 1564
rect 5601 1562 5718 1563
rect 5277 1554 5328 1562
rect 5375 1554 5409 1562
rect 5277 1542 5302 1554
rect 5309 1542 5328 1554
rect 5382 1552 5409 1554
rect 5418 1552 5639 1562
rect 5674 1559 5680 1562
rect 5382 1548 5639 1552
rect 5277 1534 5328 1542
rect 5375 1534 5639 1548
rect 5683 1554 5718 1562
rect 5229 1486 5248 1520
rect 5293 1526 5322 1534
rect 5293 1520 5310 1526
rect 5293 1518 5327 1520
rect 5375 1518 5391 1534
rect 5392 1524 5600 1534
rect 5601 1524 5617 1534
rect 5665 1530 5680 1545
rect 5683 1542 5684 1554
rect 5691 1542 5718 1554
rect 5683 1534 5718 1542
rect 5683 1533 5712 1534
rect 5403 1520 5617 1524
rect 5418 1518 5617 1520
rect 5652 1520 5665 1530
rect 5683 1520 5700 1533
rect 5652 1518 5700 1520
rect 5294 1514 5327 1518
rect 5290 1512 5327 1514
rect 5290 1511 5357 1512
rect 5290 1506 5321 1511
rect 5327 1506 5357 1511
rect 5290 1502 5357 1506
rect 5263 1499 5357 1502
rect 5263 1492 5312 1499
rect 5263 1486 5293 1492
rect 5312 1487 5317 1492
rect 5229 1470 5309 1486
rect 5321 1478 5357 1499
rect 5418 1494 5607 1518
rect 5652 1517 5699 1518
rect 5665 1512 5699 1517
rect 5433 1491 5607 1494
rect 5426 1488 5607 1491
rect 5635 1511 5699 1512
rect 5229 1468 5248 1470
rect 5263 1468 5297 1470
rect 5229 1452 5309 1468
rect 5229 1446 5248 1452
rect 4945 1420 5048 1430
rect 4899 1418 5048 1420
rect 5069 1418 5104 1430
rect 4738 1416 4900 1418
rect 4750 1396 4769 1416
rect 4784 1414 4814 1416
rect 4633 1388 4674 1396
rect 4756 1392 4769 1396
rect 4821 1400 4900 1416
rect 4932 1416 5104 1418
rect 4932 1400 5011 1416
rect 5018 1414 5048 1416
rect 4596 1378 4625 1388
rect 4639 1378 4668 1388
rect 4683 1378 4713 1392
rect 4756 1378 4799 1392
rect 4821 1388 5011 1400
rect 5076 1396 5082 1416
rect 4806 1378 4836 1388
rect 4837 1378 4995 1388
rect 4999 1378 5029 1388
rect 5033 1378 5063 1392
rect 5091 1378 5104 1416
rect 5176 1430 5205 1446
rect 5219 1430 5248 1446
rect 5263 1436 5293 1452
rect 5321 1430 5327 1478
rect 5330 1472 5349 1478
rect 5364 1472 5394 1480
rect 5330 1464 5394 1472
rect 5330 1448 5410 1464
rect 5426 1457 5488 1488
rect 5504 1457 5566 1488
rect 5635 1486 5684 1511
rect 5699 1486 5729 1502
rect 5598 1472 5628 1480
rect 5635 1478 5745 1486
rect 5598 1464 5643 1472
rect 5330 1446 5349 1448
rect 5364 1446 5410 1448
rect 5330 1430 5410 1446
rect 5437 1444 5472 1457
rect 5513 1454 5550 1457
rect 5513 1452 5555 1454
rect 5442 1441 5472 1444
rect 5451 1437 5458 1441
rect 5458 1436 5459 1437
rect 5417 1430 5427 1436
rect 5176 1422 5211 1430
rect 5176 1396 5177 1422
rect 5184 1396 5211 1422
rect 5119 1378 5149 1392
rect 5176 1388 5211 1396
rect 5213 1422 5254 1430
rect 5213 1396 5228 1422
rect 5235 1396 5254 1422
rect 5318 1418 5349 1430
rect 5364 1418 5467 1430
rect 5479 1420 5505 1446
rect 5520 1441 5550 1452
rect 5582 1448 5644 1464
rect 5582 1446 5628 1448
rect 5582 1430 5644 1446
rect 5656 1430 5662 1478
rect 5665 1470 5745 1478
rect 5665 1468 5684 1470
rect 5699 1468 5733 1470
rect 5665 1452 5745 1468
rect 5665 1430 5684 1452
rect 5699 1436 5729 1452
rect 5757 1446 5763 1520
rect 5766 1446 5785 1590
rect 5800 1446 5806 1590
rect 5815 1520 5828 1590
rect 5880 1586 5902 1590
rect 5873 1564 5902 1578
rect 5955 1564 5971 1578
rect 6009 1574 6015 1576
rect 6022 1574 6130 1590
rect 6137 1574 6143 1576
rect 6151 1574 6166 1590
rect 6232 1584 6251 1587
rect 5873 1562 5971 1564
rect 5998 1562 6166 1574
rect 6181 1564 6197 1578
rect 6232 1565 6254 1584
rect 6264 1578 6280 1579
rect 6263 1576 6280 1578
rect 6264 1571 6280 1576
rect 6254 1564 6260 1565
rect 6263 1564 6292 1571
rect 6181 1563 6292 1564
rect 6181 1562 6298 1563
rect 5857 1554 5908 1562
rect 5955 1554 5989 1562
rect 5857 1542 5882 1554
rect 5889 1542 5908 1554
rect 5962 1552 5989 1554
rect 5998 1552 6219 1562
rect 6254 1559 6260 1562
rect 5962 1548 6219 1552
rect 5857 1534 5908 1542
rect 5955 1534 6219 1548
rect 6263 1554 6298 1562
rect 5809 1486 5828 1520
rect 5873 1526 5902 1534
rect 5873 1520 5890 1526
rect 5873 1518 5907 1520
rect 5955 1518 5971 1534
rect 5972 1524 6180 1534
rect 6181 1524 6197 1534
rect 6245 1530 6260 1545
rect 6263 1542 6264 1554
rect 6271 1542 6298 1554
rect 6263 1534 6298 1542
rect 6263 1533 6292 1534
rect 5983 1520 6197 1524
rect 5998 1518 6197 1520
rect 6232 1520 6245 1530
rect 6263 1520 6280 1533
rect 6232 1518 6280 1520
rect 5874 1514 5907 1518
rect 5870 1512 5907 1514
rect 5870 1511 5937 1512
rect 5870 1506 5901 1511
rect 5907 1506 5937 1511
rect 5870 1502 5937 1506
rect 5843 1499 5937 1502
rect 5843 1492 5892 1499
rect 5843 1486 5873 1492
rect 5892 1487 5897 1492
rect 5809 1470 5889 1486
rect 5901 1478 5937 1499
rect 5998 1494 6187 1518
rect 6232 1517 6279 1518
rect 6245 1512 6279 1517
rect 6013 1491 6187 1494
rect 6006 1488 6187 1491
rect 6215 1511 6279 1512
rect 5809 1468 5828 1470
rect 5843 1468 5877 1470
rect 5809 1452 5889 1468
rect 5809 1446 5828 1452
rect 5525 1420 5628 1430
rect 5479 1418 5628 1420
rect 5649 1418 5684 1430
rect 5318 1416 5480 1418
rect 5330 1396 5349 1416
rect 5364 1414 5394 1416
rect 5213 1388 5254 1396
rect 5336 1392 5349 1396
rect 5401 1400 5480 1416
rect 5512 1416 5684 1418
rect 5512 1400 5591 1416
rect 5598 1414 5628 1416
rect 5176 1378 5205 1388
rect 5219 1378 5248 1388
rect 5263 1378 5293 1392
rect 5336 1378 5379 1392
rect 5401 1388 5591 1400
rect 5656 1396 5662 1416
rect 5386 1378 5416 1388
rect 5417 1378 5575 1388
rect 5579 1378 5609 1388
rect 5613 1378 5643 1392
rect 5671 1378 5684 1416
rect 5756 1430 5785 1446
rect 5799 1430 5828 1446
rect 5843 1436 5873 1452
rect 5901 1430 5907 1478
rect 5910 1472 5929 1478
rect 5944 1472 5974 1480
rect 5910 1464 5974 1472
rect 5910 1448 5990 1464
rect 6006 1457 6068 1488
rect 6084 1457 6146 1488
rect 6215 1486 6264 1511
rect 6279 1486 6309 1502
rect 6178 1472 6208 1480
rect 6215 1478 6325 1486
rect 6178 1464 6223 1472
rect 5910 1446 5929 1448
rect 5944 1446 5990 1448
rect 5910 1430 5990 1446
rect 6017 1444 6052 1457
rect 6093 1454 6130 1457
rect 6093 1452 6135 1454
rect 6022 1441 6052 1444
rect 6031 1437 6038 1441
rect 6038 1436 6039 1437
rect 5997 1430 6007 1436
rect 5756 1422 5791 1430
rect 5756 1396 5757 1422
rect 5764 1396 5791 1422
rect 5699 1378 5729 1392
rect 5756 1388 5791 1396
rect 5793 1422 5834 1430
rect 5793 1396 5808 1422
rect 5815 1396 5834 1422
rect 5898 1418 5929 1430
rect 5944 1418 6047 1430
rect 6059 1420 6085 1446
rect 6100 1441 6130 1452
rect 6162 1448 6224 1464
rect 6162 1446 6208 1448
rect 6162 1430 6224 1446
rect 6236 1430 6242 1478
rect 6245 1470 6325 1478
rect 6245 1468 6264 1470
rect 6279 1468 6313 1470
rect 6245 1452 6325 1468
rect 6245 1430 6264 1452
rect 6279 1436 6309 1452
rect 6337 1446 6343 1520
rect 6346 1446 6365 1590
rect 6380 1446 6386 1590
rect 6395 1520 6408 1590
rect 6460 1586 6482 1590
rect 6453 1564 6482 1578
rect 6535 1564 6551 1578
rect 6589 1574 6595 1576
rect 6602 1574 6710 1590
rect 6717 1574 6723 1576
rect 6731 1574 6746 1590
rect 6812 1584 6831 1587
rect 6453 1562 6551 1564
rect 6578 1562 6746 1574
rect 6761 1564 6777 1578
rect 6812 1565 6834 1584
rect 6844 1578 6860 1579
rect 6843 1576 6860 1578
rect 6844 1571 6860 1576
rect 6834 1564 6840 1565
rect 6843 1564 6872 1571
rect 6761 1563 6872 1564
rect 6761 1562 6878 1563
rect 6437 1554 6488 1562
rect 6535 1554 6569 1562
rect 6437 1542 6462 1554
rect 6469 1542 6488 1554
rect 6542 1552 6569 1554
rect 6578 1552 6799 1562
rect 6834 1559 6840 1562
rect 6542 1548 6799 1552
rect 6437 1534 6488 1542
rect 6535 1534 6799 1548
rect 6843 1554 6878 1562
rect 6389 1486 6408 1520
rect 6453 1526 6482 1534
rect 6453 1520 6470 1526
rect 6453 1518 6487 1520
rect 6535 1518 6551 1534
rect 6552 1524 6760 1534
rect 6761 1524 6777 1534
rect 6825 1530 6840 1545
rect 6843 1542 6844 1554
rect 6851 1542 6878 1554
rect 6843 1534 6878 1542
rect 6843 1533 6872 1534
rect 6563 1520 6777 1524
rect 6578 1518 6777 1520
rect 6812 1520 6825 1530
rect 6843 1520 6860 1533
rect 6812 1518 6860 1520
rect 6454 1514 6487 1518
rect 6450 1512 6487 1514
rect 6450 1511 6517 1512
rect 6450 1506 6481 1511
rect 6487 1506 6517 1511
rect 6450 1502 6517 1506
rect 6423 1499 6517 1502
rect 6423 1492 6472 1499
rect 6423 1486 6453 1492
rect 6472 1487 6477 1492
rect 6389 1470 6469 1486
rect 6481 1478 6517 1499
rect 6578 1494 6767 1518
rect 6812 1517 6859 1518
rect 6825 1512 6859 1517
rect 6593 1491 6767 1494
rect 6586 1488 6767 1491
rect 6795 1511 6859 1512
rect 6389 1468 6408 1470
rect 6423 1468 6457 1470
rect 6389 1452 6469 1468
rect 6389 1446 6408 1452
rect 6105 1420 6208 1430
rect 6059 1418 6208 1420
rect 6229 1418 6264 1430
rect 5898 1416 6060 1418
rect 5910 1396 5929 1416
rect 5944 1414 5974 1416
rect 5793 1388 5834 1396
rect 5916 1392 5929 1396
rect 5981 1400 6060 1416
rect 6092 1416 6264 1418
rect 6092 1400 6171 1416
rect 6178 1414 6208 1416
rect 5756 1378 5785 1388
rect 5799 1378 5828 1388
rect 5843 1378 5873 1392
rect 5916 1378 5959 1392
rect 5981 1388 6171 1400
rect 6236 1396 6242 1416
rect 5966 1378 5996 1388
rect 5997 1378 6155 1388
rect 6159 1378 6189 1388
rect 6193 1378 6223 1392
rect 6251 1378 6264 1416
rect 6336 1430 6365 1446
rect 6379 1430 6408 1446
rect 6423 1436 6453 1452
rect 6481 1430 6487 1478
rect 6490 1472 6509 1478
rect 6524 1472 6554 1480
rect 6490 1464 6554 1472
rect 6490 1448 6570 1464
rect 6586 1457 6648 1488
rect 6664 1457 6726 1488
rect 6795 1486 6844 1511
rect 6859 1486 6889 1502
rect 6758 1472 6788 1480
rect 6795 1478 6905 1486
rect 6758 1464 6803 1472
rect 6490 1446 6509 1448
rect 6524 1446 6570 1448
rect 6490 1430 6570 1446
rect 6597 1444 6632 1457
rect 6673 1454 6710 1457
rect 6673 1452 6715 1454
rect 6602 1441 6632 1444
rect 6611 1437 6618 1441
rect 6618 1436 6619 1437
rect 6577 1430 6587 1436
rect 6336 1422 6371 1430
rect 6336 1396 6337 1422
rect 6344 1396 6371 1422
rect 6279 1378 6309 1392
rect 6336 1388 6371 1396
rect 6373 1422 6414 1430
rect 6373 1396 6388 1422
rect 6395 1396 6414 1422
rect 6478 1418 6509 1430
rect 6524 1418 6627 1430
rect 6639 1420 6665 1446
rect 6680 1441 6710 1452
rect 6742 1448 6804 1464
rect 6742 1446 6788 1448
rect 6742 1430 6804 1446
rect 6816 1430 6822 1478
rect 6825 1470 6905 1478
rect 6825 1468 6844 1470
rect 6859 1468 6893 1470
rect 6825 1452 6905 1468
rect 6825 1430 6844 1452
rect 6859 1436 6889 1452
rect 6917 1446 6923 1520
rect 6926 1446 6945 1590
rect 6960 1446 6966 1590
rect 6975 1520 6988 1590
rect 7040 1586 7062 1590
rect 7033 1564 7062 1578
rect 7115 1564 7131 1578
rect 7169 1574 7175 1576
rect 7182 1574 7290 1590
rect 7297 1574 7303 1576
rect 7311 1574 7326 1590
rect 7392 1584 7411 1587
rect 7033 1562 7131 1564
rect 7158 1562 7326 1574
rect 7341 1564 7357 1578
rect 7392 1565 7414 1584
rect 7424 1578 7440 1579
rect 7423 1576 7440 1578
rect 7424 1571 7440 1576
rect 7414 1564 7420 1565
rect 7423 1564 7452 1571
rect 7341 1563 7452 1564
rect 7341 1562 7458 1563
rect 7017 1554 7068 1562
rect 7115 1554 7149 1562
rect 7017 1542 7042 1554
rect 7049 1542 7068 1554
rect 7122 1552 7149 1554
rect 7158 1552 7379 1562
rect 7414 1559 7420 1562
rect 7122 1548 7379 1552
rect 7017 1534 7068 1542
rect 7115 1534 7379 1548
rect 7423 1554 7458 1562
rect 6969 1486 6988 1520
rect 7033 1526 7062 1534
rect 7033 1520 7050 1526
rect 7033 1518 7067 1520
rect 7115 1518 7131 1534
rect 7132 1524 7340 1534
rect 7341 1524 7357 1534
rect 7405 1530 7420 1545
rect 7423 1542 7424 1554
rect 7431 1542 7458 1554
rect 7423 1534 7458 1542
rect 7423 1533 7452 1534
rect 7151 1520 7357 1524
rect 7158 1518 7357 1520
rect 7392 1520 7405 1530
rect 7423 1520 7440 1533
rect 7392 1518 7440 1520
rect 7034 1514 7067 1518
rect 7030 1512 7067 1514
rect 7030 1511 7097 1512
rect 7030 1506 7061 1511
rect 7067 1506 7097 1511
rect 7030 1502 7097 1506
rect 7003 1499 7097 1502
rect 7003 1492 7052 1499
rect 7003 1486 7033 1492
rect 7052 1487 7057 1492
rect 6969 1470 7049 1486
rect 7061 1478 7097 1499
rect 7158 1494 7347 1518
rect 7392 1517 7439 1518
rect 7405 1512 7439 1517
rect 7173 1491 7347 1494
rect 7166 1488 7347 1491
rect 7375 1511 7439 1512
rect 6969 1468 6988 1470
rect 7003 1468 7037 1470
rect 6969 1452 7049 1468
rect 6969 1446 6988 1452
rect 6685 1420 6788 1430
rect 6639 1418 6788 1420
rect 6809 1418 6844 1430
rect 6478 1416 6640 1418
rect 6490 1396 6509 1416
rect 6524 1414 6554 1416
rect 6373 1388 6414 1396
rect 6496 1392 6509 1396
rect 6561 1400 6640 1416
rect 6672 1416 6844 1418
rect 6672 1400 6751 1416
rect 6758 1414 6788 1416
rect 6336 1378 6365 1388
rect 6379 1378 6408 1388
rect 6423 1378 6453 1392
rect 6496 1378 6539 1392
rect 6561 1388 6751 1400
rect 6816 1396 6822 1416
rect 6546 1378 6576 1388
rect 6577 1378 6735 1388
rect 6739 1378 6769 1388
rect 6773 1378 6803 1392
rect 6831 1378 6844 1416
rect 6916 1430 6945 1446
rect 6959 1430 6988 1446
rect 7003 1436 7033 1452
rect 7061 1430 7067 1478
rect 7070 1472 7089 1478
rect 7104 1472 7134 1480
rect 7070 1464 7134 1472
rect 7070 1448 7150 1464
rect 7166 1457 7228 1488
rect 7244 1457 7306 1488
rect 7375 1486 7424 1511
rect 7439 1486 7469 1502
rect 7338 1472 7368 1480
rect 7375 1478 7485 1486
rect 7338 1464 7383 1472
rect 7070 1446 7089 1448
rect 7104 1446 7150 1448
rect 7070 1430 7150 1446
rect 7177 1444 7212 1457
rect 7253 1454 7290 1457
rect 7253 1452 7295 1454
rect 7182 1441 7212 1444
rect 7191 1437 7198 1441
rect 7198 1436 7199 1437
rect 7157 1430 7167 1436
rect 6916 1422 6951 1430
rect 6916 1396 6917 1422
rect 6924 1396 6951 1422
rect 6859 1378 6889 1392
rect 6916 1388 6951 1396
rect 6953 1422 6994 1430
rect 6953 1396 6968 1422
rect 6975 1396 6994 1422
rect 7058 1418 7089 1430
rect 7104 1418 7207 1430
rect 7219 1420 7245 1446
rect 7260 1441 7290 1452
rect 7322 1448 7384 1464
rect 7322 1446 7368 1448
rect 7322 1430 7384 1446
rect 7396 1430 7402 1478
rect 7405 1470 7485 1478
rect 7405 1468 7424 1470
rect 7439 1468 7473 1470
rect 7405 1452 7485 1468
rect 7405 1430 7424 1452
rect 7439 1436 7469 1452
rect 7497 1446 7503 1520
rect 7506 1446 7525 1590
rect 7540 1446 7546 1590
rect 7555 1520 7568 1590
rect 7620 1586 7642 1590
rect 7613 1564 7642 1578
rect 7695 1564 7711 1578
rect 7749 1574 7755 1576
rect 7762 1574 7870 1590
rect 7877 1574 7883 1576
rect 7891 1574 7906 1590
rect 7972 1584 7991 1587
rect 7613 1562 7711 1564
rect 7738 1562 7906 1574
rect 7921 1564 7937 1578
rect 7972 1565 7994 1584
rect 8004 1578 8020 1579
rect 8003 1576 8020 1578
rect 8004 1571 8020 1576
rect 7994 1564 8000 1565
rect 8003 1564 8032 1571
rect 7921 1563 8032 1564
rect 7921 1562 8038 1563
rect 7597 1554 7648 1562
rect 7695 1554 7729 1562
rect 7597 1542 7622 1554
rect 7629 1542 7648 1554
rect 7702 1552 7729 1554
rect 7738 1552 7959 1562
rect 7994 1559 8000 1562
rect 7702 1548 7959 1552
rect 7597 1534 7648 1542
rect 7695 1534 7959 1548
rect 8003 1554 8038 1562
rect 7549 1486 7568 1520
rect 7613 1526 7642 1534
rect 7613 1520 7630 1526
rect 7613 1518 7647 1520
rect 7695 1518 7711 1534
rect 7712 1524 7920 1534
rect 7921 1524 7937 1534
rect 7985 1530 8000 1545
rect 8003 1542 8004 1554
rect 8011 1542 8038 1554
rect 8003 1534 8038 1542
rect 8003 1533 8032 1534
rect 7723 1520 7937 1524
rect 7738 1518 7937 1520
rect 7972 1520 7985 1530
rect 8003 1520 8020 1533
rect 7972 1518 8020 1520
rect 7614 1514 7647 1518
rect 7610 1512 7647 1514
rect 7610 1511 7677 1512
rect 7610 1506 7641 1511
rect 7647 1506 7677 1511
rect 7610 1502 7677 1506
rect 7583 1499 7677 1502
rect 7583 1492 7632 1499
rect 7583 1486 7613 1492
rect 7632 1487 7637 1492
rect 7549 1470 7629 1486
rect 7641 1478 7677 1499
rect 7738 1494 7927 1518
rect 7972 1517 8019 1518
rect 7985 1512 8019 1517
rect 7753 1491 7927 1494
rect 7746 1488 7927 1491
rect 7955 1511 8019 1512
rect 7549 1468 7568 1470
rect 7583 1468 7617 1470
rect 7549 1452 7629 1468
rect 7549 1446 7568 1452
rect 7265 1420 7368 1430
rect 7219 1418 7368 1420
rect 7389 1418 7424 1430
rect 7058 1416 7220 1418
rect 7070 1396 7089 1416
rect 7104 1414 7134 1416
rect 6953 1388 6994 1396
rect 7076 1392 7089 1396
rect 7141 1400 7220 1416
rect 7252 1416 7424 1418
rect 7252 1400 7331 1416
rect 7338 1414 7368 1416
rect 6916 1378 6945 1388
rect 6959 1378 6988 1388
rect 7003 1378 7033 1392
rect 7076 1378 7119 1392
rect 7141 1388 7331 1400
rect 7396 1396 7402 1416
rect 7126 1378 7156 1388
rect 7157 1378 7315 1388
rect 7319 1378 7349 1388
rect 7353 1378 7383 1392
rect 7411 1378 7424 1416
rect 7496 1430 7525 1446
rect 7539 1430 7568 1446
rect 7583 1436 7613 1452
rect 7641 1430 7647 1478
rect 7650 1472 7669 1478
rect 7684 1472 7714 1480
rect 7650 1464 7714 1472
rect 7650 1448 7730 1464
rect 7746 1457 7808 1488
rect 7824 1457 7886 1488
rect 7955 1486 8004 1511
rect 8019 1486 8049 1502
rect 7918 1472 7948 1480
rect 7955 1478 8065 1486
rect 7918 1464 7963 1472
rect 7650 1446 7669 1448
rect 7684 1446 7730 1448
rect 7650 1430 7730 1446
rect 7757 1444 7792 1457
rect 7833 1454 7870 1457
rect 7833 1452 7875 1454
rect 7762 1441 7792 1444
rect 7771 1437 7778 1441
rect 7778 1436 7779 1437
rect 7737 1430 7747 1436
rect 7496 1422 7531 1430
rect 7496 1396 7497 1422
rect 7504 1396 7531 1422
rect 7439 1378 7469 1392
rect 7496 1388 7531 1396
rect 7533 1422 7574 1430
rect 7533 1396 7548 1422
rect 7555 1396 7574 1422
rect 7638 1418 7669 1430
rect 7684 1418 7787 1430
rect 7799 1420 7825 1446
rect 7840 1441 7870 1452
rect 7902 1448 7964 1464
rect 7902 1446 7948 1448
rect 7902 1430 7964 1446
rect 7976 1430 7982 1478
rect 7985 1470 8065 1478
rect 7985 1468 8004 1470
rect 8019 1468 8053 1470
rect 7985 1452 8065 1468
rect 7985 1430 8004 1452
rect 8019 1436 8049 1452
rect 8077 1446 8083 1520
rect 8086 1446 8105 1590
rect 8120 1446 8126 1590
rect 8135 1520 8148 1590
rect 8200 1586 8222 1590
rect 8193 1564 8222 1578
rect 8275 1564 8291 1578
rect 8329 1574 8335 1576
rect 8342 1574 8450 1590
rect 8457 1574 8463 1576
rect 8471 1574 8486 1590
rect 8552 1584 8571 1587
rect 8193 1562 8291 1564
rect 8318 1562 8486 1574
rect 8501 1564 8517 1578
rect 8552 1565 8574 1584
rect 8584 1578 8600 1579
rect 8583 1576 8600 1578
rect 8584 1571 8600 1576
rect 8574 1564 8580 1565
rect 8583 1564 8612 1571
rect 8501 1563 8612 1564
rect 8501 1562 8618 1563
rect 8177 1554 8228 1562
rect 8275 1554 8309 1562
rect 8177 1542 8202 1554
rect 8209 1542 8228 1554
rect 8282 1552 8309 1554
rect 8318 1552 8539 1562
rect 8574 1559 8580 1562
rect 8282 1548 8539 1552
rect 8177 1534 8228 1542
rect 8275 1534 8539 1548
rect 8583 1554 8618 1562
rect 8129 1486 8148 1520
rect 8193 1526 8222 1534
rect 8193 1520 8210 1526
rect 8193 1518 8227 1520
rect 8275 1518 8291 1534
rect 8292 1524 8500 1534
rect 8501 1524 8517 1534
rect 8565 1530 8580 1545
rect 8583 1542 8584 1554
rect 8591 1542 8618 1554
rect 8583 1534 8618 1542
rect 8583 1533 8612 1534
rect 8303 1520 8517 1524
rect 8318 1518 8517 1520
rect 8552 1520 8565 1530
rect 8583 1520 8600 1533
rect 8552 1518 8600 1520
rect 8194 1514 8227 1518
rect 8190 1512 8227 1514
rect 8190 1511 8257 1512
rect 8190 1506 8221 1511
rect 8227 1506 8257 1511
rect 8190 1502 8257 1506
rect 8163 1499 8257 1502
rect 8163 1492 8212 1499
rect 8163 1486 8193 1492
rect 8212 1487 8217 1492
rect 8129 1470 8209 1486
rect 8221 1478 8257 1499
rect 8318 1494 8507 1518
rect 8552 1517 8599 1518
rect 8565 1512 8599 1517
rect 8333 1491 8507 1494
rect 8326 1488 8507 1491
rect 8535 1511 8599 1512
rect 8129 1468 8148 1470
rect 8163 1468 8197 1470
rect 8129 1452 8209 1468
rect 8129 1446 8148 1452
rect 7845 1420 7948 1430
rect 7799 1418 7948 1420
rect 7969 1418 8004 1430
rect 7638 1416 7800 1418
rect 7650 1396 7669 1416
rect 7684 1414 7714 1416
rect 7533 1388 7574 1396
rect 7656 1392 7669 1396
rect 7721 1400 7800 1416
rect 7832 1416 8004 1418
rect 7832 1400 7911 1416
rect 7918 1414 7948 1416
rect 7496 1378 7525 1388
rect 7539 1378 7568 1388
rect 7583 1378 7613 1392
rect 7656 1378 7699 1392
rect 7721 1388 7911 1400
rect 7976 1396 7982 1416
rect 7706 1378 7736 1388
rect 7737 1378 7895 1388
rect 7899 1378 7929 1388
rect 7933 1378 7963 1392
rect 7991 1378 8004 1416
rect 8076 1430 8105 1446
rect 8119 1430 8148 1446
rect 8163 1436 8193 1452
rect 8221 1430 8227 1478
rect 8230 1472 8249 1478
rect 8264 1472 8294 1480
rect 8230 1464 8294 1472
rect 8230 1448 8310 1464
rect 8326 1457 8388 1488
rect 8404 1457 8466 1488
rect 8535 1486 8584 1511
rect 8599 1486 8629 1502
rect 8498 1472 8528 1480
rect 8535 1478 8645 1486
rect 8498 1464 8543 1472
rect 8230 1446 8249 1448
rect 8264 1446 8310 1448
rect 8230 1430 8310 1446
rect 8337 1444 8372 1457
rect 8413 1454 8450 1457
rect 8413 1452 8455 1454
rect 8342 1441 8372 1444
rect 8351 1437 8358 1441
rect 8358 1436 8359 1437
rect 8317 1430 8327 1436
rect 8076 1422 8111 1430
rect 8076 1396 8077 1422
rect 8084 1396 8111 1422
rect 8019 1378 8049 1392
rect 8076 1388 8111 1396
rect 8113 1422 8154 1430
rect 8113 1396 8128 1422
rect 8135 1396 8154 1422
rect 8218 1418 8249 1430
rect 8264 1418 8367 1430
rect 8379 1420 8405 1446
rect 8420 1441 8450 1452
rect 8482 1448 8544 1464
rect 8482 1446 8528 1448
rect 8482 1430 8544 1446
rect 8556 1430 8562 1478
rect 8565 1470 8645 1478
rect 8565 1468 8584 1470
rect 8599 1468 8633 1470
rect 8565 1452 8645 1468
rect 8565 1430 8584 1452
rect 8599 1436 8629 1452
rect 8657 1446 8663 1520
rect 8666 1446 8685 1590
rect 8700 1446 8706 1590
rect 8715 1520 8728 1590
rect 8780 1586 8802 1590
rect 8773 1564 8802 1578
rect 8855 1564 8871 1578
rect 8909 1574 8915 1576
rect 8922 1574 9030 1590
rect 9037 1574 9043 1576
rect 9051 1574 9066 1590
rect 9132 1584 9151 1587
rect 8773 1562 8871 1564
rect 8898 1562 9066 1574
rect 9081 1564 9097 1578
rect 9132 1565 9154 1584
rect 9164 1578 9180 1579
rect 9163 1576 9180 1578
rect 9164 1571 9180 1576
rect 9154 1564 9160 1565
rect 9163 1564 9192 1571
rect 9081 1563 9192 1564
rect 9081 1562 9198 1563
rect 8757 1554 8808 1562
rect 8855 1554 8889 1562
rect 8757 1542 8782 1554
rect 8789 1542 8808 1554
rect 8862 1552 8889 1554
rect 8898 1552 9119 1562
rect 9154 1559 9160 1562
rect 8862 1548 9119 1552
rect 8757 1534 8808 1542
rect 8855 1534 9119 1548
rect 9163 1554 9198 1562
rect 8709 1486 8728 1520
rect 8773 1526 8802 1534
rect 8773 1520 8790 1526
rect 8773 1518 8807 1520
rect 8855 1518 8871 1534
rect 8872 1524 9080 1534
rect 9081 1524 9097 1534
rect 9145 1530 9160 1545
rect 9163 1542 9164 1554
rect 9171 1542 9198 1554
rect 9163 1534 9198 1542
rect 9163 1533 9192 1534
rect 8883 1520 9097 1524
rect 8898 1518 9097 1520
rect 9132 1520 9145 1530
rect 9163 1520 9180 1533
rect 9132 1518 9180 1520
rect 8774 1514 8807 1518
rect 8770 1512 8807 1514
rect 8770 1511 8837 1512
rect 8770 1506 8801 1511
rect 8807 1506 8837 1511
rect 8770 1502 8837 1506
rect 8743 1499 8837 1502
rect 8743 1492 8792 1499
rect 8743 1486 8773 1492
rect 8792 1487 8797 1492
rect 8709 1470 8789 1486
rect 8801 1478 8837 1499
rect 8898 1494 9087 1518
rect 9132 1517 9179 1518
rect 9145 1512 9179 1517
rect 8913 1491 9087 1494
rect 8906 1488 9087 1491
rect 9115 1511 9179 1512
rect 8709 1468 8728 1470
rect 8743 1468 8777 1470
rect 8709 1452 8789 1468
rect 8709 1446 8728 1452
rect 8425 1420 8528 1430
rect 8379 1418 8528 1420
rect 8549 1418 8584 1430
rect 8218 1416 8380 1418
rect 8230 1396 8249 1416
rect 8264 1414 8294 1416
rect 8113 1388 8154 1396
rect 8236 1392 8249 1396
rect 8301 1400 8380 1416
rect 8412 1416 8584 1418
rect 8412 1400 8491 1416
rect 8498 1414 8528 1416
rect 8076 1378 8105 1388
rect 8119 1378 8148 1388
rect 8163 1378 8193 1392
rect 8236 1378 8279 1392
rect 8301 1388 8491 1400
rect 8556 1396 8562 1416
rect 8286 1378 8316 1388
rect 8317 1378 8475 1388
rect 8479 1378 8509 1388
rect 8513 1378 8543 1392
rect 8571 1378 8584 1416
rect 8656 1430 8685 1446
rect 8699 1430 8728 1446
rect 8743 1436 8773 1452
rect 8801 1430 8807 1478
rect 8810 1472 8829 1478
rect 8844 1472 8874 1480
rect 8810 1464 8874 1472
rect 8810 1448 8890 1464
rect 8906 1457 8968 1488
rect 8984 1457 9046 1488
rect 9115 1486 9164 1511
rect 9179 1486 9209 1502
rect 9078 1472 9108 1480
rect 9115 1478 9225 1486
rect 9078 1464 9123 1472
rect 8810 1446 8829 1448
rect 8844 1446 8890 1448
rect 8810 1430 8890 1446
rect 8917 1444 8952 1457
rect 8993 1454 9030 1457
rect 8993 1452 9035 1454
rect 8922 1441 8952 1444
rect 8931 1437 8938 1441
rect 8938 1436 8939 1437
rect 8897 1430 8907 1436
rect 8656 1422 8691 1430
rect 8656 1396 8657 1422
rect 8664 1396 8691 1422
rect 8599 1378 8629 1392
rect 8656 1388 8691 1396
rect 8693 1422 8734 1430
rect 8693 1396 8708 1422
rect 8715 1396 8734 1422
rect 8798 1418 8829 1430
rect 8844 1418 8947 1430
rect 8959 1420 8985 1446
rect 9000 1441 9030 1452
rect 9062 1448 9124 1464
rect 9062 1446 9108 1448
rect 9062 1430 9124 1446
rect 9136 1430 9142 1478
rect 9145 1470 9225 1478
rect 9145 1468 9164 1470
rect 9179 1468 9213 1470
rect 9145 1452 9225 1468
rect 9145 1430 9164 1452
rect 9179 1436 9209 1452
rect 9237 1446 9243 1520
rect 9246 1446 9265 1590
rect 9280 1446 9286 1590
rect 9295 1520 9308 1590
rect 9360 1586 9382 1590
rect 9353 1564 9382 1578
rect 9435 1564 9451 1578
rect 9489 1574 9495 1576
rect 9502 1574 9610 1590
rect 9617 1574 9623 1576
rect 9631 1574 9646 1590
rect 9712 1584 9731 1587
rect 9353 1562 9451 1564
rect 9478 1562 9646 1574
rect 9661 1564 9677 1578
rect 9712 1565 9734 1584
rect 9744 1578 9760 1579
rect 9743 1576 9760 1578
rect 9744 1571 9760 1576
rect 9734 1564 9740 1565
rect 9743 1564 9772 1571
rect 9661 1563 9772 1564
rect 9661 1562 9778 1563
rect 9337 1554 9388 1562
rect 9435 1554 9469 1562
rect 9337 1542 9362 1554
rect 9369 1542 9388 1554
rect 9442 1552 9469 1554
rect 9478 1552 9699 1562
rect 9734 1559 9740 1562
rect 9442 1548 9699 1552
rect 9337 1534 9388 1542
rect 9435 1534 9699 1548
rect 9743 1554 9778 1562
rect 9289 1486 9308 1520
rect 9353 1526 9382 1534
rect 9353 1520 9370 1526
rect 9353 1518 9387 1520
rect 9435 1518 9451 1534
rect 9452 1524 9660 1534
rect 9661 1524 9677 1534
rect 9725 1530 9740 1545
rect 9743 1542 9744 1554
rect 9751 1542 9778 1554
rect 9743 1534 9778 1542
rect 9743 1533 9772 1534
rect 9463 1520 9677 1524
rect 9478 1518 9677 1520
rect 9712 1520 9725 1530
rect 9743 1520 9760 1533
rect 9712 1518 9760 1520
rect 9354 1514 9387 1518
rect 9350 1512 9387 1514
rect 9350 1511 9417 1512
rect 9350 1506 9381 1511
rect 9387 1506 9417 1511
rect 9350 1502 9417 1506
rect 9323 1499 9417 1502
rect 9323 1492 9372 1499
rect 9323 1486 9353 1492
rect 9372 1487 9377 1492
rect 9289 1470 9369 1486
rect 9381 1478 9417 1499
rect 9478 1494 9667 1518
rect 9712 1517 9759 1518
rect 9725 1512 9759 1517
rect 9493 1491 9667 1494
rect 9486 1488 9667 1491
rect 9695 1511 9759 1512
rect 9289 1468 9308 1470
rect 9323 1468 9357 1470
rect 9289 1452 9369 1468
rect 9289 1446 9308 1452
rect 9005 1420 9108 1430
rect 8959 1418 9108 1420
rect 9129 1418 9164 1430
rect 8798 1416 8960 1418
rect 8810 1396 8829 1416
rect 8844 1414 8874 1416
rect 8693 1388 8734 1396
rect 8816 1392 8829 1396
rect 8881 1400 8960 1416
rect 8992 1416 9164 1418
rect 8992 1400 9071 1416
rect 9078 1414 9108 1416
rect 8656 1378 8685 1388
rect 8699 1378 8728 1388
rect 8743 1378 8773 1392
rect 8816 1378 8859 1392
rect 8881 1388 9071 1400
rect 9136 1396 9142 1416
rect 8866 1378 8896 1388
rect 8897 1378 9055 1388
rect 9059 1378 9089 1388
rect 9093 1378 9123 1392
rect 9151 1378 9164 1416
rect 9236 1430 9265 1446
rect 9279 1430 9308 1446
rect 9323 1436 9353 1452
rect 9381 1430 9387 1478
rect 9390 1472 9409 1478
rect 9424 1472 9454 1480
rect 9390 1464 9454 1472
rect 9390 1448 9470 1464
rect 9486 1457 9548 1488
rect 9564 1457 9626 1488
rect 9695 1486 9744 1511
rect 9759 1486 9789 1502
rect 9658 1472 9688 1480
rect 9695 1478 9805 1486
rect 9658 1464 9703 1472
rect 9390 1446 9409 1448
rect 9424 1446 9470 1448
rect 9390 1430 9470 1446
rect 9497 1444 9532 1457
rect 9573 1454 9610 1457
rect 9573 1452 9615 1454
rect 9502 1441 9532 1444
rect 9511 1437 9518 1441
rect 9518 1436 9519 1437
rect 9477 1430 9487 1436
rect 9236 1422 9271 1430
rect 9236 1396 9237 1422
rect 9244 1396 9271 1422
rect 9179 1378 9209 1392
rect 9236 1388 9271 1396
rect 9273 1422 9314 1430
rect 9273 1396 9288 1422
rect 9295 1396 9314 1422
rect 9378 1418 9409 1430
rect 9424 1418 9527 1430
rect 9539 1420 9565 1446
rect 9580 1441 9610 1452
rect 9642 1448 9704 1464
rect 9642 1446 9688 1448
rect 9642 1430 9704 1446
rect 9716 1430 9722 1478
rect 9725 1470 9805 1478
rect 9725 1468 9744 1470
rect 9759 1468 9793 1470
rect 9725 1452 9805 1468
rect 9725 1430 9744 1452
rect 9759 1436 9789 1452
rect 9817 1446 9823 1520
rect 9826 1446 9845 1590
rect 9860 1446 9866 1590
rect 9875 1520 9888 1590
rect 9940 1586 9962 1590
rect 9933 1564 9962 1578
rect 10015 1564 10031 1578
rect 10069 1574 10075 1576
rect 10082 1574 10190 1590
rect 10197 1574 10203 1576
rect 10211 1574 10226 1590
rect 10292 1584 10311 1587
rect 9933 1562 10031 1564
rect 10058 1562 10226 1574
rect 10241 1564 10257 1578
rect 10292 1565 10314 1584
rect 10324 1578 10340 1579
rect 10323 1576 10340 1578
rect 10324 1571 10340 1576
rect 10314 1564 10320 1565
rect 10323 1564 10352 1571
rect 10241 1563 10352 1564
rect 10241 1562 10358 1563
rect 9917 1554 9968 1562
rect 10015 1554 10049 1562
rect 9917 1542 9942 1554
rect 9949 1542 9968 1554
rect 10022 1552 10049 1554
rect 10058 1552 10279 1562
rect 10314 1559 10320 1562
rect 10022 1548 10279 1552
rect 9917 1534 9968 1542
rect 10015 1534 10279 1548
rect 10323 1554 10358 1562
rect 9869 1486 9888 1520
rect 9933 1526 9962 1534
rect 9933 1520 9950 1526
rect 9933 1518 9967 1520
rect 10015 1518 10031 1534
rect 10032 1524 10240 1534
rect 10241 1524 10257 1534
rect 10305 1530 10320 1545
rect 10323 1542 10324 1554
rect 10331 1542 10358 1554
rect 10323 1534 10358 1542
rect 10323 1533 10352 1534
rect 10043 1520 10257 1524
rect 10058 1518 10257 1520
rect 10292 1520 10305 1530
rect 10323 1520 10340 1533
rect 10292 1518 10340 1520
rect 9934 1514 9967 1518
rect 9930 1512 9967 1514
rect 9930 1511 9997 1512
rect 9930 1506 9961 1511
rect 9967 1506 9997 1511
rect 9930 1502 9997 1506
rect 9903 1499 9997 1502
rect 9903 1492 9952 1499
rect 9903 1486 9933 1492
rect 9952 1487 9957 1492
rect 9869 1470 9949 1486
rect 9961 1478 9997 1499
rect 10058 1494 10247 1518
rect 10292 1517 10339 1518
rect 10305 1512 10339 1517
rect 10073 1491 10247 1494
rect 10066 1488 10247 1491
rect 10275 1511 10339 1512
rect 9869 1468 9888 1470
rect 9903 1468 9937 1470
rect 9869 1452 9949 1468
rect 9869 1446 9888 1452
rect 9585 1420 9688 1430
rect 9539 1418 9688 1420
rect 9709 1418 9744 1430
rect 9378 1416 9540 1418
rect 9390 1396 9409 1416
rect 9424 1414 9454 1416
rect 9273 1388 9314 1396
rect 9396 1392 9409 1396
rect 9461 1400 9540 1416
rect 9572 1416 9744 1418
rect 9572 1400 9651 1416
rect 9658 1414 9688 1416
rect 9236 1378 9265 1388
rect 9279 1378 9308 1388
rect 9323 1378 9353 1392
rect 9396 1378 9439 1392
rect 9461 1388 9651 1400
rect 9716 1396 9722 1416
rect 9446 1378 9476 1388
rect 9477 1378 9635 1388
rect 9639 1378 9669 1388
rect 9673 1378 9703 1392
rect 9731 1378 9744 1416
rect 9816 1430 9845 1446
rect 9859 1430 9888 1446
rect 9903 1436 9933 1452
rect 9961 1430 9967 1478
rect 9970 1472 9989 1478
rect 10004 1472 10034 1480
rect 9970 1464 10034 1472
rect 9970 1448 10050 1464
rect 10066 1457 10128 1488
rect 10144 1457 10206 1488
rect 10275 1486 10324 1511
rect 10339 1486 10369 1502
rect 10238 1472 10268 1480
rect 10275 1478 10385 1486
rect 10238 1464 10283 1472
rect 9970 1446 9989 1448
rect 10004 1446 10050 1448
rect 9970 1430 10050 1446
rect 10077 1444 10112 1457
rect 10153 1454 10190 1457
rect 10153 1452 10195 1454
rect 10082 1441 10112 1444
rect 10091 1437 10098 1441
rect 10098 1436 10099 1437
rect 10057 1430 10067 1436
rect 9816 1422 9851 1430
rect 9816 1396 9817 1422
rect 9824 1396 9851 1422
rect 9759 1378 9789 1392
rect 9816 1388 9851 1396
rect 9853 1422 9894 1430
rect 9853 1396 9868 1422
rect 9875 1396 9894 1422
rect 9958 1418 9989 1430
rect 10004 1418 10107 1430
rect 10119 1420 10145 1446
rect 10160 1441 10190 1452
rect 10222 1448 10284 1464
rect 10222 1446 10268 1448
rect 10222 1430 10284 1446
rect 10296 1430 10302 1478
rect 10305 1470 10385 1478
rect 10305 1468 10324 1470
rect 10339 1468 10373 1470
rect 10305 1452 10385 1468
rect 10305 1430 10324 1452
rect 10339 1436 10369 1452
rect 10397 1446 10403 1520
rect 10406 1446 10425 1590
rect 10440 1446 10446 1590
rect 10455 1520 10468 1590
rect 10520 1586 10542 1590
rect 10513 1564 10542 1578
rect 10595 1564 10611 1578
rect 10649 1574 10655 1576
rect 10662 1574 10770 1590
rect 10777 1574 10783 1576
rect 10791 1574 10806 1590
rect 10872 1584 10891 1587
rect 10513 1562 10611 1564
rect 10638 1562 10806 1574
rect 10821 1564 10837 1578
rect 10872 1565 10894 1584
rect 10904 1578 10920 1579
rect 10903 1576 10920 1578
rect 10904 1571 10920 1576
rect 10894 1564 10900 1565
rect 10903 1564 10932 1571
rect 10821 1563 10932 1564
rect 10821 1562 10938 1563
rect 10497 1554 10548 1562
rect 10595 1554 10629 1562
rect 10497 1542 10522 1554
rect 10529 1542 10548 1554
rect 10602 1552 10629 1554
rect 10638 1552 10859 1562
rect 10894 1559 10900 1562
rect 10602 1548 10859 1552
rect 10497 1534 10548 1542
rect 10595 1534 10859 1548
rect 10903 1554 10938 1562
rect 10449 1486 10468 1520
rect 10513 1526 10542 1534
rect 10513 1520 10530 1526
rect 10513 1518 10547 1520
rect 10595 1518 10611 1534
rect 10612 1524 10820 1534
rect 10821 1524 10837 1534
rect 10885 1530 10900 1545
rect 10903 1542 10904 1554
rect 10911 1542 10938 1554
rect 10903 1534 10938 1542
rect 10903 1533 10932 1534
rect 10623 1520 10837 1524
rect 10638 1518 10837 1520
rect 10872 1520 10885 1530
rect 10903 1520 10920 1533
rect 10872 1518 10920 1520
rect 10514 1514 10547 1518
rect 10510 1512 10547 1514
rect 10510 1511 10577 1512
rect 10510 1506 10541 1511
rect 10547 1506 10577 1511
rect 10510 1502 10577 1506
rect 10483 1499 10577 1502
rect 10483 1492 10532 1499
rect 10483 1486 10513 1492
rect 10532 1487 10537 1492
rect 10449 1470 10529 1486
rect 10541 1478 10577 1499
rect 10638 1494 10827 1518
rect 10872 1517 10919 1518
rect 10885 1512 10919 1517
rect 10653 1491 10827 1494
rect 10646 1488 10827 1491
rect 10855 1511 10919 1512
rect 10449 1468 10468 1470
rect 10483 1468 10517 1470
rect 10449 1452 10529 1468
rect 10449 1446 10468 1452
rect 10165 1420 10268 1430
rect 10119 1418 10268 1420
rect 10289 1418 10324 1430
rect 9958 1416 10120 1418
rect 9970 1396 9989 1416
rect 10004 1414 10034 1416
rect 9853 1388 9894 1396
rect 9976 1392 9989 1396
rect 10041 1400 10120 1416
rect 10152 1416 10324 1418
rect 10152 1400 10231 1416
rect 10238 1414 10268 1416
rect 9816 1378 9845 1388
rect 9859 1378 9888 1388
rect 9903 1378 9933 1392
rect 9976 1378 10019 1392
rect 10041 1388 10231 1400
rect 10296 1396 10302 1416
rect 10026 1378 10056 1388
rect 10057 1378 10215 1388
rect 10219 1378 10249 1388
rect 10253 1378 10283 1392
rect 10311 1378 10324 1416
rect 10396 1430 10425 1446
rect 10439 1430 10468 1446
rect 10483 1436 10513 1452
rect 10541 1430 10547 1478
rect 10550 1472 10569 1478
rect 10584 1472 10614 1480
rect 10550 1464 10614 1472
rect 10550 1448 10630 1464
rect 10646 1457 10708 1488
rect 10724 1457 10786 1488
rect 10855 1486 10904 1511
rect 10919 1486 10949 1502
rect 10818 1472 10848 1480
rect 10855 1478 10965 1486
rect 10818 1464 10863 1472
rect 10550 1446 10569 1448
rect 10584 1446 10630 1448
rect 10550 1430 10630 1446
rect 10657 1444 10692 1457
rect 10733 1454 10770 1457
rect 10733 1452 10775 1454
rect 10662 1441 10692 1444
rect 10671 1437 10678 1441
rect 10678 1436 10679 1437
rect 10637 1430 10647 1436
rect 10396 1422 10431 1430
rect 10396 1396 10397 1422
rect 10404 1396 10431 1422
rect 10339 1378 10369 1392
rect 10396 1388 10431 1396
rect 10433 1422 10474 1430
rect 10433 1396 10448 1422
rect 10455 1396 10474 1422
rect 10538 1418 10569 1430
rect 10584 1418 10687 1430
rect 10699 1420 10725 1446
rect 10740 1441 10770 1452
rect 10802 1448 10864 1464
rect 10802 1446 10848 1448
rect 10802 1430 10864 1446
rect 10876 1430 10882 1478
rect 10885 1470 10965 1478
rect 10885 1468 10904 1470
rect 10919 1468 10953 1470
rect 10885 1452 10965 1468
rect 10885 1430 10904 1452
rect 10919 1436 10949 1452
rect 10977 1446 10983 1520
rect 10986 1446 11005 1590
rect 11020 1446 11026 1590
rect 11035 1520 11048 1590
rect 11100 1586 11122 1590
rect 11093 1564 11122 1578
rect 11175 1564 11191 1578
rect 11229 1574 11235 1576
rect 11242 1574 11350 1590
rect 11357 1574 11363 1576
rect 11371 1574 11386 1590
rect 11452 1584 11471 1587
rect 11093 1562 11191 1564
rect 11218 1562 11386 1574
rect 11401 1564 11417 1578
rect 11452 1565 11474 1584
rect 11484 1578 11500 1579
rect 11483 1576 11500 1578
rect 11484 1571 11500 1576
rect 11474 1564 11480 1565
rect 11483 1564 11512 1571
rect 11401 1563 11512 1564
rect 11401 1562 11518 1563
rect 11077 1554 11128 1562
rect 11175 1554 11209 1562
rect 11077 1542 11102 1554
rect 11109 1542 11128 1554
rect 11182 1552 11209 1554
rect 11218 1552 11439 1562
rect 11474 1559 11480 1562
rect 11182 1548 11439 1552
rect 11077 1534 11128 1542
rect 11175 1534 11439 1548
rect 11483 1554 11518 1562
rect 11029 1486 11048 1520
rect 11093 1526 11122 1534
rect 11093 1520 11110 1526
rect 11093 1518 11127 1520
rect 11175 1518 11191 1534
rect 11192 1524 11400 1534
rect 11401 1524 11417 1534
rect 11465 1530 11480 1545
rect 11483 1542 11484 1554
rect 11491 1542 11518 1554
rect 11483 1534 11518 1542
rect 11483 1533 11512 1534
rect 11203 1520 11417 1524
rect 11218 1518 11417 1520
rect 11452 1520 11465 1530
rect 11483 1520 11500 1533
rect 11452 1518 11500 1520
rect 11094 1514 11127 1518
rect 11090 1512 11127 1514
rect 11090 1511 11157 1512
rect 11090 1506 11121 1511
rect 11127 1506 11157 1511
rect 11090 1502 11157 1506
rect 11063 1499 11157 1502
rect 11063 1492 11112 1499
rect 11063 1486 11093 1492
rect 11112 1487 11117 1492
rect 11029 1470 11109 1486
rect 11121 1478 11157 1499
rect 11218 1494 11407 1518
rect 11452 1517 11499 1518
rect 11465 1512 11499 1517
rect 11233 1491 11407 1494
rect 11226 1488 11407 1491
rect 11435 1511 11499 1512
rect 11029 1468 11048 1470
rect 11063 1468 11097 1470
rect 11029 1452 11109 1468
rect 11029 1446 11048 1452
rect 10745 1420 10848 1430
rect 10699 1418 10848 1420
rect 10869 1418 10904 1430
rect 10538 1416 10700 1418
rect 10550 1396 10569 1416
rect 10584 1414 10614 1416
rect 10433 1388 10474 1396
rect 10556 1392 10569 1396
rect 10621 1400 10700 1416
rect 10732 1416 10904 1418
rect 10732 1400 10811 1416
rect 10818 1414 10848 1416
rect 10396 1378 10425 1388
rect 10439 1378 10468 1388
rect 10483 1378 10513 1392
rect 10556 1378 10599 1392
rect 10621 1388 10811 1400
rect 10876 1396 10882 1416
rect 10606 1378 10636 1388
rect 10637 1378 10795 1388
rect 10799 1378 10829 1388
rect 10833 1378 10863 1392
rect 10891 1378 10904 1416
rect 10976 1430 11005 1446
rect 11019 1430 11048 1446
rect 11063 1436 11093 1452
rect 11121 1430 11127 1478
rect 11130 1472 11149 1478
rect 11164 1472 11194 1480
rect 11130 1464 11194 1472
rect 11130 1448 11210 1464
rect 11226 1457 11288 1488
rect 11304 1457 11366 1488
rect 11435 1486 11484 1511
rect 11499 1486 11529 1502
rect 11398 1472 11428 1480
rect 11435 1478 11545 1486
rect 11398 1464 11443 1472
rect 11130 1446 11149 1448
rect 11164 1446 11210 1448
rect 11130 1430 11210 1446
rect 11237 1444 11272 1457
rect 11313 1454 11350 1457
rect 11313 1452 11355 1454
rect 11242 1441 11272 1444
rect 11251 1437 11258 1441
rect 11258 1436 11259 1437
rect 11217 1430 11227 1436
rect 10976 1422 11011 1430
rect 10976 1396 10977 1422
rect 10984 1396 11011 1422
rect 10919 1378 10949 1392
rect 10976 1388 11011 1396
rect 11013 1422 11054 1430
rect 11013 1396 11028 1422
rect 11035 1396 11054 1422
rect 11118 1418 11149 1430
rect 11164 1418 11267 1430
rect 11279 1420 11305 1446
rect 11320 1441 11350 1452
rect 11382 1448 11444 1464
rect 11382 1446 11428 1448
rect 11382 1430 11444 1446
rect 11456 1430 11462 1478
rect 11465 1470 11545 1478
rect 11465 1468 11484 1470
rect 11499 1468 11533 1470
rect 11465 1452 11545 1468
rect 11465 1430 11484 1452
rect 11499 1436 11529 1452
rect 11557 1446 11563 1520
rect 11566 1446 11585 1590
rect 11600 1446 11606 1590
rect 11615 1520 11628 1590
rect 11680 1586 11702 1590
rect 11673 1564 11702 1578
rect 11755 1564 11771 1578
rect 11809 1574 11815 1576
rect 11822 1574 11930 1590
rect 11937 1574 11943 1576
rect 11951 1574 11966 1590
rect 12032 1584 12051 1587
rect 11673 1562 11771 1564
rect 11798 1562 11966 1574
rect 11981 1564 11997 1578
rect 12032 1565 12054 1584
rect 12064 1578 12080 1579
rect 12063 1576 12080 1578
rect 12064 1571 12080 1576
rect 12054 1564 12060 1565
rect 12063 1564 12092 1571
rect 11981 1563 12092 1564
rect 11981 1562 12098 1563
rect 11657 1554 11708 1562
rect 11755 1554 11789 1562
rect 11657 1542 11682 1554
rect 11689 1542 11708 1554
rect 11762 1552 11789 1554
rect 11798 1552 12019 1562
rect 12054 1559 12060 1562
rect 11762 1548 12019 1552
rect 11657 1534 11708 1542
rect 11755 1534 12019 1548
rect 12063 1554 12098 1562
rect 11609 1486 11628 1520
rect 11673 1526 11702 1534
rect 11673 1520 11690 1526
rect 11673 1518 11707 1520
rect 11755 1518 11771 1534
rect 11772 1524 11980 1534
rect 11981 1524 11997 1534
rect 12045 1530 12060 1545
rect 12063 1542 12064 1554
rect 12071 1542 12098 1554
rect 12063 1534 12098 1542
rect 12063 1533 12092 1534
rect 11783 1520 11997 1524
rect 11798 1518 11997 1520
rect 12032 1520 12045 1530
rect 12063 1520 12080 1533
rect 12032 1518 12080 1520
rect 11674 1514 11707 1518
rect 11670 1512 11707 1514
rect 11670 1511 11737 1512
rect 11670 1506 11701 1511
rect 11707 1506 11737 1511
rect 11670 1502 11737 1506
rect 11643 1499 11737 1502
rect 11643 1492 11692 1499
rect 11643 1486 11673 1492
rect 11692 1487 11697 1492
rect 11609 1470 11689 1486
rect 11701 1478 11737 1499
rect 11798 1494 11987 1518
rect 12032 1517 12079 1518
rect 12045 1512 12079 1517
rect 11813 1491 11987 1494
rect 11806 1488 11987 1491
rect 12015 1511 12079 1512
rect 11609 1468 11628 1470
rect 11643 1468 11677 1470
rect 11609 1452 11689 1468
rect 11609 1446 11628 1452
rect 11325 1420 11428 1430
rect 11279 1418 11428 1420
rect 11449 1418 11484 1430
rect 11118 1416 11280 1418
rect 11130 1396 11149 1416
rect 11164 1414 11194 1416
rect 11013 1388 11054 1396
rect 11136 1392 11149 1396
rect 11201 1400 11280 1416
rect 11312 1416 11484 1418
rect 11312 1400 11391 1416
rect 11398 1414 11428 1416
rect 10976 1378 11005 1388
rect 11019 1378 11048 1388
rect 11063 1378 11093 1392
rect 11136 1378 11179 1392
rect 11201 1388 11391 1400
rect 11456 1396 11462 1416
rect 11186 1378 11216 1388
rect 11217 1378 11375 1388
rect 11379 1378 11409 1388
rect 11413 1378 11443 1392
rect 11471 1378 11484 1416
rect 11556 1430 11585 1446
rect 11599 1430 11628 1446
rect 11643 1436 11673 1452
rect 11701 1430 11707 1478
rect 11710 1472 11729 1478
rect 11744 1472 11774 1480
rect 11710 1464 11774 1472
rect 11710 1448 11790 1464
rect 11806 1457 11868 1488
rect 11884 1457 11946 1488
rect 12015 1486 12064 1511
rect 12079 1486 12109 1502
rect 11978 1472 12008 1480
rect 12015 1478 12125 1486
rect 11978 1464 12023 1472
rect 11710 1446 11729 1448
rect 11744 1446 11790 1448
rect 11710 1430 11790 1446
rect 11817 1444 11852 1457
rect 11893 1454 11930 1457
rect 11893 1452 11935 1454
rect 11822 1441 11852 1444
rect 11831 1437 11838 1441
rect 11838 1436 11839 1437
rect 11797 1430 11807 1436
rect 11556 1422 11591 1430
rect 11556 1396 11557 1422
rect 11564 1396 11591 1422
rect 11499 1378 11529 1392
rect 11556 1388 11591 1396
rect 11593 1422 11634 1430
rect 11593 1396 11608 1422
rect 11615 1396 11634 1422
rect 11698 1418 11729 1430
rect 11744 1418 11847 1430
rect 11859 1420 11885 1446
rect 11900 1441 11930 1452
rect 11962 1448 12024 1464
rect 11962 1446 12008 1448
rect 11962 1430 12024 1446
rect 12036 1430 12042 1478
rect 12045 1470 12125 1478
rect 12045 1468 12064 1470
rect 12079 1468 12113 1470
rect 12045 1452 12125 1468
rect 12045 1430 12064 1452
rect 12079 1436 12109 1452
rect 12137 1446 12143 1520
rect 12146 1446 12165 1590
rect 12180 1446 12186 1590
rect 12195 1520 12208 1590
rect 12260 1586 12282 1590
rect 12253 1564 12282 1578
rect 12335 1564 12351 1578
rect 12389 1574 12395 1576
rect 12402 1574 12510 1590
rect 12517 1574 12523 1576
rect 12531 1574 12546 1590
rect 12612 1584 12631 1587
rect 12253 1562 12351 1564
rect 12378 1562 12546 1574
rect 12561 1564 12577 1578
rect 12612 1565 12634 1584
rect 12644 1578 12660 1579
rect 12643 1576 12660 1578
rect 12644 1571 12660 1576
rect 12634 1564 12640 1565
rect 12643 1564 12672 1571
rect 12561 1563 12672 1564
rect 12561 1562 12678 1563
rect 12237 1554 12288 1562
rect 12335 1554 12369 1562
rect 12237 1542 12262 1554
rect 12269 1542 12288 1554
rect 12342 1552 12369 1554
rect 12378 1552 12599 1562
rect 12634 1559 12640 1562
rect 12342 1548 12599 1552
rect 12237 1534 12288 1542
rect 12335 1534 12599 1548
rect 12643 1554 12678 1562
rect 12189 1486 12208 1520
rect 12253 1526 12282 1534
rect 12253 1520 12270 1526
rect 12253 1518 12287 1520
rect 12335 1518 12351 1534
rect 12352 1524 12560 1534
rect 12561 1524 12577 1534
rect 12625 1530 12640 1545
rect 12643 1542 12644 1554
rect 12651 1542 12678 1554
rect 12643 1534 12678 1542
rect 12643 1533 12672 1534
rect 12363 1520 12577 1524
rect 12378 1518 12577 1520
rect 12612 1520 12625 1530
rect 12643 1520 12660 1533
rect 12612 1518 12660 1520
rect 12254 1514 12287 1518
rect 12250 1512 12287 1514
rect 12250 1511 12317 1512
rect 12250 1506 12281 1511
rect 12287 1506 12317 1511
rect 12250 1502 12317 1506
rect 12223 1499 12317 1502
rect 12223 1492 12272 1499
rect 12223 1486 12253 1492
rect 12272 1487 12277 1492
rect 12189 1470 12269 1486
rect 12281 1478 12317 1499
rect 12378 1494 12567 1518
rect 12612 1517 12659 1518
rect 12625 1512 12659 1517
rect 12393 1491 12567 1494
rect 12386 1488 12567 1491
rect 12595 1511 12659 1512
rect 12189 1468 12208 1470
rect 12223 1468 12257 1470
rect 12189 1452 12269 1468
rect 12189 1446 12208 1452
rect 11905 1420 12008 1430
rect 11859 1418 12008 1420
rect 12029 1418 12064 1430
rect 11698 1416 11860 1418
rect 11710 1396 11729 1416
rect 11744 1414 11774 1416
rect 11593 1388 11634 1396
rect 11716 1392 11729 1396
rect 11781 1400 11860 1416
rect 11892 1416 12064 1418
rect 11892 1400 11971 1416
rect 11978 1414 12008 1416
rect 11556 1378 11585 1388
rect 11599 1378 11628 1388
rect 11643 1378 11673 1392
rect 11716 1378 11759 1392
rect 11781 1388 11971 1400
rect 12036 1396 12042 1416
rect 11766 1378 11796 1388
rect 11797 1378 11955 1388
rect 11959 1378 11989 1388
rect 11993 1378 12023 1392
rect 12051 1378 12064 1416
rect 12136 1430 12165 1446
rect 12179 1430 12208 1446
rect 12223 1436 12253 1452
rect 12281 1430 12287 1478
rect 12290 1472 12309 1478
rect 12324 1472 12354 1480
rect 12290 1464 12354 1472
rect 12290 1448 12370 1464
rect 12386 1457 12448 1488
rect 12464 1457 12526 1488
rect 12595 1486 12644 1511
rect 12659 1486 12689 1502
rect 12558 1472 12588 1480
rect 12595 1478 12705 1486
rect 12558 1464 12603 1472
rect 12290 1446 12309 1448
rect 12324 1446 12370 1448
rect 12290 1430 12370 1446
rect 12397 1444 12432 1457
rect 12473 1454 12510 1457
rect 12473 1452 12515 1454
rect 12402 1441 12432 1444
rect 12411 1437 12418 1441
rect 12418 1436 12419 1437
rect 12377 1430 12387 1436
rect 12136 1422 12171 1430
rect 12136 1396 12137 1422
rect 12144 1396 12171 1422
rect 12079 1378 12109 1392
rect 12136 1388 12171 1396
rect 12173 1422 12214 1430
rect 12173 1396 12188 1422
rect 12195 1396 12214 1422
rect 12278 1418 12309 1430
rect 12324 1418 12427 1430
rect 12439 1420 12465 1446
rect 12480 1441 12510 1452
rect 12542 1448 12604 1464
rect 12542 1446 12588 1448
rect 12542 1430 12604 1446
rect 12616 1430 12622 1478
rect 12625 1470 12705 1478
rect 12625 1468 12644 1470
rect 12659 1468 12693 1470
rect 12625 1452 12705 1468
rect 12625 1430 12644 1452
rect 12659 1436 12689 1452
rect 12717 1446 12723 1520
rect 12726 1446 12745 1590
rect 12760 1446 12766 1590
rect 12775 1520 12788 1590
rect 12840 1586 12862 1590
rect 12833 1564 12862 1578
rect 12915 1564 12931 1578
rect 12969 1574 12975 1576
rect 12982 1574 13090 1590
rect 13097 1574 13103 1576
rect 13111 1574 13126 1590
rect 13192 1584 13211 1587
rect 12833 1562 12931 1564
rect 12958 1562 13126 1574
rect 13141 1564 13157 1578
rect 13192 1565 13214 1584
rect 13224 1578 13240 1579
rect 13223 1576 13240 1578
rect 13224 1571 13240 1576
rect 13214 1564 13220 1565
rect 13223 1564 13252 1571
rect 13141 1563 13252 1564
rect 13141 1562 13258 1563
rect 12817 1554 12868 1562
rect 12915 1554 12949 1562
rect 12817 1542 12842 1554
rect 12849 1542 12868 1554
rect 12922 1552 12949 1554
rect 12958 1552 13179 1562
rect 13214 1559 13220 1562
rect 12922 1548 13179 1552
rect 12817 1534 12868 1542
rect 12915 1534 13179 1548
rect 13223 1554 13258 1562
rect 12769 1486 12788 1520
rect 12833 1526 12862 1534
rect 12833 1520 12850 1526
rect 12833 1518 12867 1520
rect 12915 1518 12931 1534
rect 12932 1524 13140 1534
rect 13141 1524 13157 1534
rect 13205 1530 13220 1545
rect 13223 1542 13224 1554
rect 13231 1542 13258 1554
rect 13223 1534 13258 1542
rect 13223 1533 13252 1534
rect 12943 1520 13157 1524
rect 12958 1518 13157 1520
rect 13192 1520 13205 1530
rect 13223 1520 13240 1533
rect 13192 1518 13240 1520
rect 12834 1514 12867 1518
rect 12830 1512 12867 1514
rect 12830 1511 12897 1512
rect 12830 1506 12861 1511
rect 12867 1506 12897 1511
rect 12830 1502 12897 1506
rect 12803 1499 12897 1502
rect 12803 1492 12852 1499
rect 12803 1486 12833 1492
rect 12852 1487 12857 1492
rect 12769 1470 12849 1486
rect 12861 1478 12897 1499
rect 12958 1494 13147 1518
rect 13192 1517 13239 1518
rect 13205 1512 13239 1517
rect 12973 1491 13147 1494
rect 12966 1488 13147 1491
rect 13175 1511 13239 1512
rect 12769 1468 12788 1470
rect 12803 1468 12837 1470
rect 12769 1452 12849 1468
rect 12769 1446 12788 1452
rect 12485 1420 12588 1430
rect 12439 1418 12588 1420
rect 12609 1418 12644 1430
rect 12278 1416 12440 1418
rect 12290 1396 12309 1416
rect 12324 1414 12354 1416
rect 12173 1388 12214 1396
rect 12296 1392 12309 1396
rect 12361 1400 12440 1416
rect 12472 1416 12644 1418
rect 12472 1400 12551 1416
rect 12558 1414 12588 1416
rect 12136 1378 12165 1388
rect 12179 1378 12208 1388
rect 12223 1378 12253 1392
rect 12296 1378 12339 1392
rect 12361 1388 12551 1400
rect 12616 1396 12622 1416
rect 12346 1378 12376 1388
rect 12377 1378 12535 1388
rect 12539 1378 12569 1388
rect 12573 1378 12603 1392
rect 12631 1378 12644 1416
rect 12716 1430 12745 1446
rect 12759 1430 12788 1446
rect 12803 1436 12833 1452
rect 12861 1430 12867 1478
rect 12870 1472 12889 1478
rect 12904 1472 12934 1480
rect 12870 1464 12934 1472
rect 12870 1448 12950 1464
rect 12966 1457 13028 1488
rect 13044 1457 13106 1488
rect 13175 1486 13224 1511
rect 13239 1486 13269 1502
rect 13138 1472 13168 1480
rect 13175 1478 13285 1486
rect 13138 1464 13183 1472
rect 12870 1446 12889 1448
rect 12904 1446 12950 1448
rect 12870 1430 12950 1446
rect 12977 1444 13012 1457
rect 13053 1454 13090 1457
rect 13053 1452 13095 1454
rect 12982 1441 13012 1444
rect 12991 1437 12998 1441
rect 12998 1436 12999 1437
rect 12957 1430 12967 1436
rect 12716 1422 12751 1430
rect 12716 1396 12717 1422
rect 12724 1396 12751 1422
rect 12659 1378 12689 1392
rect 12716 1388 12751 1396
rect 12753 1422 12794 1430
rect 12753 1396 12768 1422
rect 12775 1396 12794 1422
rect 12858 1418 12889 1430
rect 12904 1418 13007 1430
rect 13019 1420 13045 1446
rect 13060 1441 13090 1452
rect 13122 1448 13184 1464
rect 13122 1446 13168 1448
rect 13122 1430 13184 1446
rect 13196 1430 13202 1478
rect 13205 1470 13285 1478
rect 13205 1468 13224 1470
rect 13239 1468 13273 1470
rect 13205 1452 13285 1468
rect 13205 1430 13224 1452
rect 13239 1436 13269 1452
rect 13297 1446 13303 1520
rect 13306 1446 13325 1590
rect 13340 1446 13346 1590
rect 13355 1520 13368 1590
rect 13420 1586 13442 1590
rect 13413 1564 13442 1578
rect 13495 1564 13511 1578
rect 13549 1574 13555 1576
rect 13562 1574 13670 1590
rect 13677 1574 13683 1576
rect 13691 1574 13706 1590
rect 13772 1584 13791 1587
rect 13413 1562 13511 1564
rect 13538 1562 13706 1574
rect 13721 1564 13737 1578
rect 13772 1565 13794 1584
rect 13804 1578 13820 1579
rect 13803 1576 13820 1578
rect 13804 1571 13820 1576
rect 13794 1564 13800 1565
rect 13803 1564 13832 1571
rect 13721 1563 13832 1564
rect 13721 1562 13838 1563
rect 13397 1554 13448 1562
rect 13495 1554 13529 1562
rect 13397 1542 13422 1554
rect 13429 1542 13448 1554
rect 13502 1552 13529 1554
rect 13538 1552 13759 1562
rect 13794 1559 13800 1562
rect 13502 1548 13759 1552
rect 13397 1534 13448 1542
rect 13495 1534 13759 1548
rect 13803 1554 13838 1562
rect 13349 1486 13368 1520
rect 13413 1526 13442 1534
rect 13413 1520 13430 1526
rect 13413 1518 13447 1520
rect 13495 1518 13511 1534
rect 13512 1524 13720 1534
rect 13721 1524 13737 1534
rect 13785 1530 13800 1545
rect 13803 1542 13804 1554
rect 13811 1542 13838 1554
rect 13803 1534 13838 1542
rect 13803 1533 13832 1534
rect 13523 1520 13737 1524
rect 13538 1518 13737 1520
rect 13772 1520 13785 1530
rect 13803 1520 13820 1533
rect 13772 1518 13820 1520
rect 13414 1514 13447 1518
rect 13410 1512 13447 1514
rect 13410 1511 13477 1512
rect 13410 1506 13441 1511
rect 13447 1506 13477 1511
rect 13410 1502 13477 1506
rect 13383 1499 13477 1502
rect 13383 1492 13432 1499
rect 13383 1486 13413 1492
rect 13432 1487 13437 1492
rect 13349 1470 13429 1486
rect 13441 1478 13477 1499
rect 13538 1494 13727 1518
rect 13772 1517 13819 1518
rect 13785 1512 13819 1517
rect 13553 1491 13727 1494
rect 13546 1488 13727 1491
rect 13755 1511 13819 1512
rect 13349 1468 13368 1470
rect 13383 1468 13417 1470
rect 13349 1452 13429 1468
rect 13349 1446 13368 1452
rect 13065 1420 13168 1430
rect 13019 1418 13168 1420
rect 13189 1418 13224 1430
rect 12858 1416 13020 1418
rect 12870 1396 12889 1416
rect 12904 1414 12934 1416
rect 12753 1388 12794 1396
rect 12876 1392 12889 1396
rect 12941 1400 13020 1416
rect 13052 1416 13224 1418
rect 13052 1400 13131 1416
rect 13138 1414 13168 1416
rect 12716 1378 12745 1388
rect 12759 1378 12788 1388
rect 12803 1378 12833 1392
rect 12876 1378 12919 1392
rect 12941 1388 13131 1400
rect 13196 1396 13202 1416
rect 12926 1378 12956 1388
rect 12957 1378 13115 1388
rect 13119 1378 13149 1388
rect 13153 1378 13183 1392
rect 13211 1378 13224 1416
rect 13296 1430 13325 1446
rect 13339 1430 13368 1446
rect 13383 1436 13413 1452
rect 13441 1430 13447 1478
rect 13450 1472 13469 1478
rect 13484 1472 13514 1480
rect 13450 1464 13514 1472
rect 13450 1448 13530 1464
rect 13546 1457 13608 1488
rect 13624 1457 13686 1488
rect 13755 1486 13804 1511
rect 13819 1486 13849 1502
rect 13718 1472 13748 1480
rect 13755 1478 13865 1486
rect 13718 1464 13763 1472
rect 13450 1446 13469 1448
rect 13484 1446 13530 1448
rect 13450 1430 13530 1446
rect 13557 1444 13592 1457
rect 13633 1454 13670 1457
rect 13633 1452 13675 1454
rect 13562 1441 13592 1444
rect 13571 1437 13578 1441
rect 13578 1436 13579 1437
rect 13537 1430 13547 1436
rect 13296 1422 13331 1430
rect 13296 1396 13297 1422
rect 13304 1396 13331 1422
rect 13239 1378 13269 1392
rect 13296 1388 13331 1396
rect 13333 1422 13374 1430
rect 13333 1396 13348 1422
rect 13355 1396 13374 1422
rect 13438 1418 13469 1430
rect 13484 1418 13587 1430
rect 13599 1420 13625 1446
rect 13640 1441 13670 1452
rect 13702 1448 13764 1464
rect 13702 1446 13748 1448
rect 13702 1430 13764 1446
rect 13776 1430 13782 1478
rect 13785 1470 13865 1478
rect 13785 1468 13804 1470
rect 13819 1468 13853 1470
rect 13785 1452 13865 1468
rect 13785 1430 13804 1452
rect 13819 1436 13849 1452
rect 13877 1446 13883 1520
rect 13886 1446 13905 1590
rect 13920 1446 13926 1590
rect 13935 1520 13948 1590
rect 14000 1586 14022 1590
rect 13993 1564 14022 1578
rect 14075 1564 14091 1578
rect 14129 1574 14135 1576
rect 14142 1574 14250 1590
rect 14257 1574 14263 1576
rect 14271 1574 14286 1590
rect 14352 1584 14371 1587
rect 13993 1562 14091 1564
rect 14118 1562 14286 1574
rect 14301 1564 14317 1578
rect 14352 1565 14374 1584
rect 14384 1578 14400 1579
rect 14383 1576 14400 1578
rect 14384 1571 14400 1576
rect 14374 1564 14380 1565
rect 14383 1564 14412 1571
rect 14301 1563 14412 1564
rect 14301 1562 14418 1563
rect 13977 1554 14028 1562
rect 14075 1554 14109 1562
rect 13977 1542 14002 1554
rect 14009 1542 14028 1554
rect 14082 1552 14109 1554
rect 14118 1552 14339 1562
rect 14374 1559 14380 1562
rect 14082 1548 14339 1552
rect 13977 1534 14028 1542
rect 14075 1534 14339 1548
rect 14383 1554 14418 1562
rect 13929 1486 13948 1520
rect 13993 1526 14022 1534
rect 13993 1520 14010 1526
rect 13993 1518 14027 1520
rect 14075 1518 14091 1534
rect 14092 1524 14300 1534
rect 14301 1524 14317 1534
rect 14365 1530 14380 1545
rect 14383 1542 14384 1554
rect 14391 1542 14418 1554
rect 14383 1534 14418 1542
rect 14383 1533 14412 1534
rect 14103 1520 14317 1524
rect 14118 1518 14317 1520
rect 14352 1520 14365 1530
rect 14383 1520 14400 1533
rect 14352 1518 14400 1520
rect 13994 1514 14027 1518
rect 13990 1512 14027 1514
rect 13990 1511 14057 1512
rect 13990 1506 14021 1511
rect 14027 1506 14057 1511
rect 13990 1502 14057 1506
rect 13963 1499 14057 1502
rect 13963 1492 14012 1499
rect 13963 1486 13993 1492
rect 14012 1487 14017 1492
rect 13929 1470 14009 1486
rect 14021 1478 14057 1499
rect 14118 1494 14307 1518
rect 14352 1517 14399 1518
rect 14365 1512 14399 1517
rect 14133 1491 14307 1494
rect 14126 1488 14307 1491
rect 14335 1511 14399 1512
rect 13929 1468 13948 1470
rect 13963 1468 13997 1470
rect 13929 1452 14009 1468
rect 13929 1446 13948 1452
rect 13645 1420 13748 1430
rect 13599 1418 13748 1420
rect 13769 1418 13804 1430
rect 13438 1416 13600 1418
rect 13450 1396 13469 1416
rect 13484 1414 13514 1416
rect 13333 1388 13374 1396
rect 13456 1392 13469 1396
rect 13521 1400 13600 1416
rect 13632 1416 13804 1418
rect 13632 1400 13711 1416
rect 13718 1414 13748 1416
rect 13296 1378 13325 1388
rect 13339 1378 13368 1388
rect 13383 1378 13413 1392
rect 13456 1378 13499 1392
rect 13521 1388 13711 1400
rect 13776 1396 13782 1416
rect 13506 1378 13536 1388
rect 13537 1378 13695 1388
rect 13699 1378 13729 1388
rect 13733 1378 13763 1392
rect 13791 1378 13804 1416
rect 13876 1430 13905 1446
rect 13919 1430 13948 1446
rect 13963 1436 13993 1452
rect 14021 1430 14027 1478
rect 14030 1472 14049 1478
rect 14064 1472 14094 1480
rect 14030 1464 14094 1472
rect 14030 1448 14110 1464
rect 14126 1457 14188 1488
rect 14204 1457 14266 1488
rect 14335 1486 14384 1511
rect 14399 1486 14429 1502
rect 14298 1472 14328 1480
rect 14335 1478 14445 1486
rect 14298 1464 14343 1472
rect 14030 1446 14049 1448
rect 14064 1446 14110 1448
rect 14030 1430 14110 1446
rect 14137 1444 14172 1457
rect 14213 1454 14250 1457
rect 14213 1452 14255 1454
rect 14142 1441 14172 1444
rect 14151 1437 14158 1441
rect 14158 1436 14159 1437
rect 14117 1430 14127 1436
rect 13876 1422 13911 1430
rect 13876 1396 13877 1422
rect 13884 1396 13911 1422
rect 13819 1378 13849 1392
rect 13876 1388 13911 1396
rect 13913 1422 13954 1430
rect 13913 1396 13928 1422
rect 13935 1396 13954 1422
rect 14018 1418 14049 1430
rect 14064 1418 14167 1430
rect 14179 1420 14205 1446
rect 14220 1441 14250 1452
rect 14282 1448 14344 1464
rect 14282 1446 14328 1448
rect 14282 1430 14344 1446
rect 14356 1430 14362 1478
rect 14365 1470 14445 1478
rect 14365 1468 14384 1470
rect 14399 1468 14433 1470
rect 14365 1452 14445 1468
rect 14365 1430 14384 1452
rect 14399 1436 14429 1452
rect 14457 1446 14463 1520
rect 14466 1446 14485 1590
rect 14500 1446 14506 1590
rect 14515 1520 14528 1590
rect 14580 1586 14602 1590
rect 14573 1564 14602 1578
rect 14655 1564 14671 1578
rect 14709 1574 14715 1576
rect 14722 1574 14830 1590
rect 14837 1574 14843 1576
rect 14851 1574 14866 1590
rect 14932 1584 14951 1587
rect 14573 1562 14671 1564
rect 14698 1562 14866 1574
rect 14881 1564 14897 1578
rect 14932 1565 14954 1584
rect 14964 1578 14980 1579
rect 14963 1576 14980 1578
rect 14964 1571 14980 1576
rect 14954 1564 14960 1565
rect 14963 1564 14992 1571
rect 14881 1563 14992 1564
rect 14881 1562 14998 1563
rect 14557 1554 14608 1562
rect 14655 1554 14689 1562
rect 14557 1542 14582 1554
rect 14589 1542 14608 1554
rect 14662 1552 14689 1554
rect 14698 1552 14919 1562
rect 14954 1559 14960 1562
rect 14662 1548 14919 1552
rect 14557 1534 14608 1542
rect 14655 1534 14919 1548
rect 14963 1554 14998 1562
rect 14509 1486 14528 1520
rect 14573 1526 14602 1534
rect 14573 1520 14590 1526
rect 14573 1518 14607 1520
rect 14655 1518 14671 1534
rect 14672 1524 14880 1534
rect 14881 1524 14897 1534
rect 14945 1530 14960 1545
rect 14963 1542 14964 1554
rect 14971 1542 14998 1554
rect 14963 1534 14998 1542
rect 14963 1533 14992 1534
rect 14683 1520 14897 1524
rect 14698 1518 14897 1520
rect 14932 1520 14945 1530
rect 14963 1520 14980 1533
rect 14932 1518 14980 1520
rect 14574 1514 14607 1518
rect 14570 1512 14607 1514
rect 14570 1511 14637 1512
rect 14570 1506 14601 1511
rect 14607 1506 14637 1511
rect 14570 1502 14637 1506
rect 14543 1499 14637 1502
rect 14543 1492 14592 1499
rect 14543 1486 14573 1492
rect 14592 1487 14597 1492
rect 14509 1470 14589 1486
rect 14601 1478 14637 1499
rect 14698 1494 14887 1518
rect 14932 1517 14979 1518
rect 14945 1512 14979 1517
rect 14713 1491 14887 1494
rect 14706 1488 14887 1491
rect 14915 1511 14979 1512
rect 14509 1468 14528 1470
rect 14543 1468 14577 1470
rect 14509 1452 14589 1468
rect 14509 1446 14528 1452
rect 14225 1420 14328 1430
rect 14179 1418 14328 1420
rect 14349 1418 14384 1430
rect 14018 1416 14180 1418
rect 14030 1396 14049 1416
rect 14064 1414 14094 1416
rect 13913 1388 13954 1396
rect 14036 1392 14049 1396
rect 14101 1400 14180 1416
rect 14212 1416 14384 1418
rect 14212 1400 14291 1416
rect 14298 1414 14328 1416
rect 13876 1378 13905 1388
rect 13919 1378 13948 1388
rect 13963 1378 13993 1392
rect 14036 1378 14079 1392
rect 14101 1388 14291 1400
rect 14356 1396 14362 1416
rect 14086 1378 14116 1388
rect 14117 1378 14275 1388
rect 14279 1378 14309 1388
rect 14313 1378 14343 1392
rect 14371 1378 14384 1416
rect 14456 1430 14485 1446
rect 14499 1430 14528 1446
rect 14543 1436 14573 1452
rect 14601 1430 14607 1478
rect 14610 1472 14629 1478
rect 14644 1472 14674 1480
rect 14610 1464 14674 1472
rect 14610 1448 14690 1464
rect 14706 1457 14768 1488
rect 14784 1457 14846 1488
rect 14915 1486 14964 1511
rect 14979 1486 15009 1502
rect 14878 1472 14908 1480
rect 14915 1478 15025 1486
rect 14878 1464 14923 1472
rect 14610 1446 14629 1448
rect 14644 1446 14690 1448
rect 14610 1430 14690 1446
rect 14717 1444 14752 1457
rect 14793 1454 14830 1457
rect 14793 1452 14835 1454
rect 14722 1441 14752 1444
rect 14731 1437 14738 1441
rect 14738 1436 14739 1437
rect 14697 1430 14707 1436
rect 14456 1422 14491 1430
rect 14456 1396 14457 1422
rect 14464 1396 14491 1422
rect 14399 1378 14429 1392
rect 14456 1388 14491 1396
rect 14493 1422 14534 1430
rect 14493 1396 14508 1422
rect 14515 1396 14534 1422
rect 14598 1418 14629 1430
rect 14644 1418 14747 1430
rect 14759 1420 14785 1446
rect 14800 1441 14830 1452
rect 14862 1448 14924 1464
rect 14862 1446 14908 1448
rect 14862 1430 14924 1446
rect 14936 1430 14942 1478
rect 14945 1470 15025 1478
rect 14945 1468 14964 1470
rect 14979 1468 15013 1470
rect 14945 1452 15025 1468
rect 14945 1430 14964 1452
rect 14979 1436 15009 1452
rect 15037 1446 15043 1520
rect 15046 1446 15065 1590
rect 15080 1446 15086 1590
rect 15095 1520 15108 1590
rect 15160 1586 15182 1590
rect 15153 1564 15182 1578
rect 15235 1564 15251 1578
rect 15289 1574 15295 1576
rect 15302 1574 15410 1590
rect 15417 1574 15423 1576
rect 15431 1574 15446 1590
rect 15512 1584 15531 1587
rect 15153 1562 15251 1564
rect 15278 1562 15446 1574
rect 15461 1564 15477 1578
rect 15512 1565 15534 1584
rect 15544 1578 15560 1579
rect 15543 1576 15560 1578
rect 15544 1571 15560 1576
rect 15534 1564 15540 1565
rect 15543 1564 15572 1571
rect 15461 1563 15572 1564
rect 15461 1562 15578 1563
rect 15137 1554 15188 1562
rect 15235 1554 15269 1562
rect 15137 1542 15162 1554
rect 15169 1542 15188 1554
rect 15242 1552 15269 1554
rect 15278 1552 15499 1562
rect 15534 1559 15540 1562
rect 15242 1548 15499 1552
rect 15137 1534 15188 1542
rect 15235 1534 15499 1548
rect 15543 1554 15578 1562
rect 15089 1486 15108 1520
rect 15153 1526 15182 1534
rect 15153 1520 15170 1526
rect 15153 1518 15187 1520
rect 15235 1518 15251 1534
rect 15252 1524 15460 1534
rect 15461 1524 15477 1534
rect 15525 1530 15540 1545
rect 15543 1542 15544 1554
rect 15551 1542 15578 1554
rect 15543 1534 15578 1542
rect 15543 1533 15572 1534
rect 15263 1520 15477 1524
rect 15278 1518 15477 1520
rect 15512 1520 15525 1530
rect 15543 1520 15560 1533
rect 15512 1518 15560 1520
rect 15154 1514 15187 1518
rect 15150 1512 15187 1514
rect 15150 1511 15217 1512
rect 15150 1506 15181 1511
rect 15187 1506 15217 1511
rect 15150 1502 15217 1506
rect 15123 1499 15217 1502
rect 15123 1492 15172 1499
rect 15123 1486 15153 1492
rect 15172 1487 15177 1492
rect 15089 1470 15169 1486
rect 15181 1478 15217 1499
rect 15278 1494 15467 1518
rect 15512 1517 15559 1518
rect 15525 1512 15559 1517
rect 15293 1491 15467 1494
rect 15286 1488 15467 1491
rect 15495 1511 15559 1512
rect 15089 1468 15108 1470
rect 15123 1468 15157 1470
rect 15089 1452 15169 1468
rect 15089 1446 15108 1452
rect 14805 1420 14908 1430
rect 14759 1418 14908 1420
rect 14929 1418 14964 1430
rect 14598 1416 14760 1418
rect 14610 1396 14629 1416
rect 14644 1414 14674 1416
rect 14493 1388 14534 1396
rect 14616 1392 14629 1396
rect 14681 1400 14760 1416
rect 14792 1416 14964 1418
rect 14792 1400 14871 1416
rect 14878 1414 14908 1416
rect 14456 1378 14485 1388
rect 14499 1378 14528 1388
rect 14543 1378 14573 1392
rect 14616 1378 14659 1392
rect 14681 1388 14871 1400
rect 14936 1396 14942 1416
rect 14666 1378 14696 1388
rect 14697 1378 14855 1388
rect 14859 1378 14889 1388
rect 14893 1378 14923 1392
rect 14951 1378 14964 1416
rect 15036 1430 15065 1446
rect 15079 1430 15108 1446
rect 15123 1436 15153 1452
rect 15181 1430 15187 1478
rect 15190 1472 15209 1478
rect 15224 1472 15254 1480
rect 15190 1464 15254 1472
rect 15190 1448 15270 1464
rect 15286 1457 15348 1488
rect 15364 1457 15426 1488
rect 15495 1486 15544 1511
rect 15559 1486 15589 1502
rect 15458 1472 15488 1480
rect 15495 1478 15605 1486
rect 15458 1464 15503 1472
rect 15190 1446 15209 1448
rect 15224 1446 15270 1448
rect 15190 1430 15270 1446
rect 15297 1444 15332 1457
rect 15373 1454 15410 1457
rect 15373 1452 15415 1454
rect 15302 1441 15332 1444
rect 15311 1437 15318 1441
rect 15318 1436 15319 1437
rect 15277 1430 15287 1436
rect 15036 1422 15071 1430
rect 15036 1396 15037 1422
rect 15044 1396 15071 1422
rect 14979 1378 15009 1392
rect 15036 1388 15071 1396
rect 15073 1422 15114 1430
rect 15073 1396 15088 1422
rect 15095 1396 15114 1422
rect 15178 1418 15209 1430
rect 15224 1418 15327 1430
rect 15339 1420 15365 1446
rect 15380 1441 15410 1452
rect 15442 1448 15504 1464
rect 15442 1446 15488 1448
rect 15442 1430 15504 1446
rect 15516 1430 15522 1478
rect 15525 1470 15605 1478
rect 15525 1468 15544 1470
rect 15559 1468 15593 1470
rect 15525 1452 15605 1468
rect 15525 1430 15544 1452
rect 15559 1436 15589 1452
rect 15617 1446 15623 1520
rect 15626 1446 15645 1590
rect 15660 1446 15666 1590
rect 15675 1520 15688 1590
rect 15740 1586 15762 1590
rect 15733 1564 15762 1578
rect 15815 1564 15831 1578
rect 15869 1574 15875 1576
rect 15882 1574 15990 1590
rect 15997 1574 16003 1576
rect 16011 1574 16026 1590
rect 16092 1584 16111 1587
rect 15733 1562 15831 1564
rect 15858 1562 16026 1574
rect 16041 1564 16057 1578
rect 16092 1565 16114 1584
rect 16124 1578 16140 1579
rect 16123 1576 16140 1578
rect 16124 1571 16140 1576
rect 16114 1564 16120 1565
rect 16123 1564 16152 1571
rect 16041 1563 16152 1564
rect 16041 1562 16158 1563
rect 15717 1554 15768 1562
rect 15815 1554 15849 1562
rect 15717 1542 15742 1554
rect 15749 1542 15768 1554
rect 15822 1552 15849 1554
rect 15858 1552 16079 1562
rect 16114 1559 16120 1562
rect 15822 1548 16079 1552
rect 15717 1534 15768 1542
rect 15815 1534 16079 1548
rect 16123 1554 16158 1562
rect 15669 1486 15688 1520
rect 15733 1526 15762 1534
rect 15733 1520 15750 1526
rect 15733 1518 15767 1520
rect 15815 1518 15831 1534
rect 15832 1524 16040 1534
rect 16041 1524 16057 1534
rect 16105 1530 16120 1545
rect 16123 1542 16124 1554
rect 16131 1542 16158 1554
rect 16123 1534 16158 1542
rect 16123 1533 16152 1534
rect 15843 1520 16057 1524
rect 15858 1518 16057 1520
rect 16092 1520 16105 1530
rect 16123 1520 16140 1533
rect 16092 1518 16140 1520
rect 15734 1514 15767 1518
rect 15730 1512 15767 1514
rect 15730 1511 15797 1512
rect 15730 1506 15761 1511
rect 15767 1506 15797 1511
rect 15730 1502 15797 1506
rect 15703 1499 15797 1502
rect 15703 1492 15752 1499
rect 15703 1486 15733 1492
rect 15752 1487 15757 1492
rect 15669 1470 15749 1486
rect 15761 1478 15797 1499
rect 15858 1494 16047 1518
rect 16092 1517 16139 1518
rect 16105 1512 16139 1517
rect 15873 1491 16047 1494
rect 15866 1488 16047 1491
rect 16075 1511 16139 1512
rect 15669 1468 15688 1470
rect 15703 1468 15737 1470
rect 15669 1452 15749 1468
rect 15669 1446 15688 1452
rect 15385 1420 15488 1430
rect 15339 1418 15488 1420
rect 15509 1418 15544 1430
rect 15178 1416 15340 1418
rect 15190 1396 15209 1416
rect 15224 1414 15254 1416
rect 15073 1388 15114 1396
rect 15196 1392 15209 1396
rect 15261 1400 15340 1416
rect 15372 1416 15544 1418
rect 15372 1400 15451 1416
rect 15458 1414 15488 1416
rect 15036 1378 15065 1388
rect 15079 1378 15108 1388
rect 15123 1378 15153 1392
rect 15196 1378 15239 1392
rect 15261 1388 15451 1400
rect 15516 1396 15522 1416
rect 15246 1378 15276 1388
rect 15277 1378 15435 1388
rect 15439 1378 15469 1388
rect 15473 1378 15503 1392
rect 15531 1378 15544 1416
rect 15616 1430 15645 1446
rect 15659 1430 15688 1446
rect 15703 1436 15733 1452
rect 15761 1430 15767 1478
rect 15770 1472 15789 1478
rect 15804 1472 15834 1480
rect 15770 1464 15834 1472
rect 15770 1448 15850 1464
rect 15866 1457 15928 1488
rect 15944 1457 16006 1488
rect 16075 1486 16124 1511
rect 16139 1486 16169 1502
rect 16038 1472 16068 1480
rect 16075 1478 16185 1486
rect 16038 1464 16083 1472
rect 15770 1446 15789 1448
rect 15804 1446 15850 1448
rect 15770 1430 15850 1446
rect 15877 1444 15912 1457
rect 15953 1454 15990 1457
rect 15953 1452 15995 1454
rect 15882 1441 15912 1444
rect 15891 1437 15898 1441
rect 15898 1436 15899 1437
rect 15857 1430 15867 1436
rect 15616 1422 15651 1430
rect 15616 1396 15617 1422
rect 15624 1396 15651 1422
rect 15559 1378 15589 1392
rect 15616 1388 15651 1396
rect 15653 1422 15694 1430
rect 15653 1396 15668 1422
rect 15675 1396 15694 1422
rect 15758 1418 15789 1430
rect 15804 1418 15907 1430
rect 15919 1420 15945 1446
rect 15960 1441 15990 1452
rect 16022 1448 16084 1464
rect 16022 1446 16068 1448
rect 16022 1430 16084 1446
rect 16096 1430 16102 1478
rect 16105 1470 16185 1478
rect 16105 1468 16124 1470
rect 16139 1468 16173 1470
rect 16105 1452 16185 1468
rect 16105 1430 16124 1452
rect 16139 1436 16169 1452
rect 16197 1446 16203 1520
rect 16206 1446 16225 1590
rect 16240 1446 16246 1590
rect 16255 1520 16268 1590
rect 16320 1586 16342 1590
rect 16313 1564 16342 1578
rect 16395 1564 16411 1578
rect 16449 1574 16455 1576
rect 16462 1574 16570 1590
rect 16577 1574 16583 1576
rect 16591 1574 16606 1590
rect 16672 1584 16691 1587
rect 16313 1562 16411 1564
rect 16438 1562 16606 1574
rect 16621 1564 16637 1578
rect 16672 1565 16694 1584
rect 16704 1578 16720 1579
rect 16703 1576 16720 1578
rect 16704 1571 16720 1576
rect 16694 1564 16700 1565
rect 16703 1564 16732 1571
rect 16621 1563 16732 1564
rect 16621 1562 16738 1563
rect 16297 1554 16348 1562
rect 16395 1554 16429 1562
rect 16297 1542 16322 1554
rect 16329 1542 16348 1554
rect 16402 1552 16429 1554
rect 16438 1552 16659 1562
rect 16694 1559 16700 1562
rect 16402 1548 16659 1552
rect 16297 1534 16348 1542
rect 16395 1534 16659 1548
rect 16703 1554 16738 1562
rect 16249 1486 16268 1520
rect 16313 1526 16342 1534
rect 16313 1520 16330 1526
rect 16313 1518 16347 1520
rect 16395 1518 16411 1534
rect 16412 1524 16620 1534
rect 16621 1524 16637 1534
rect 16685 1530 16700 1545
rect 16703 1542 16704 1554
rect 16711 1542 16738 1554
rect 16703 1534 16738 1542
rect 16703 1533 16732 1534
rect 16423 1520 16637 1524
rect 16438 1518 16637 1520
rect 16672 1520 16685 1530
rect 16703 1520 16720 1533
rect 16672 1518 16720 1520
rect 16314 1514 16347 1518
rect 16310 1512 16347 1514
rect 16310 1511 16377 1512
rect 16310 1506 16341 1511
rect 16347 1506 16377 1511
rect 16310 1502 16377 1506
rect 16283 1499 16377 1502
rect 16283 1492 16332 1499
rect 16283 1486 16313 1492
rect 16332 1487 16337 1492
rect 16249 1470 16329 1486
rect 16341 1478 16377 1499
rect 16438 1494 16627 1518
rect 16672 1517 16719 1518
rect 16685 1512 16719 1517
rect 16453 1491 16627 1494
rect 16446 1488 16627 1491
rect 16655 1511 16719 1512
rect 16249 1468 16268 1470
rect 16283 1468 16317 1470
rect 16249 1452 16329 1468
rect 16249 1446 16268 1452
rect 15965 1420 16068 1430
rect 15919 1418 16068 1420
rect 16089 1418 16124 1430
rect 15758 1416 15920 1418
rect 15770 1396 15789 1416
rect 15804 1414 15834 1416
rect 15653 1388 15694 1396
rect 15776 1392 15789 1396
rect 15841 1400 15920 1416
rect 15952 1416 16124 1418
rect 15952 1400 16031 1416
rect 16038 1414 16068 1416
rect 15616 1378 15645 1388
rect 15659 1378 15688 1388
rect 15703 1378 15733 1392
rect 15776 1378 15819 1392
rect 15841 1388 16031 1400
rect 16096 1396 16102 1416
rect 15826 1378 15856 1388
rect 15857 1378 16015 1388
rect 16019 1378 16049 1388
rect 16053 1378 16083 1392
rect 16111 1378 16124 1416
rect 16196 1430 16225 1446
rect 16239 1430 16268 1446
rect 16283 1436 16313 1452
rect 16341 1430 16347 1478
rect 16350 1472 16369 1478
rect 16384 1472 16414 1480
rect 16350 1464 16414 1472
rect 16350 1448 16430 1464
rect 16446 1457 16508 1488
rect 16524 1457 16586 1488
rect 16655 1486 16704 1511
rect 16719 1486 16749 1502
rect 16618 1472 16648 1480
rect 16655 1478 16765 1486
rect 16618 1464 16663 1472
rect 16350 1446 16369 1448
rect 16384 1446 16430 1448
rect 16350 1430 16430 1446
rect 16457 1444 16492 1457
rect 16533 1454 16570 1457
rect 16533 1452 16575 1454
rect 16462 1441 16492 1444
rect 16471 1437 16478 1441
rect 16478 1436 16479 1437
rect 16437 1430 16447 1436
rect 16196 1422 16231 1430
rect 16196 1396 16197 1422
rect 16204 1396 16231 1422
rect 16139 1378 16169 1392
rect 16196 1388 16231 1396
rect 16233 1422 16274 1430
rect 16233 1396 16248 1422
rect 16255 1396 16274 1422
rect 16338 1418 16369 1430
rect 16384 1418 16487 1430
rect 16499 1420 16525 1446
rect 16540 1441 16570 1452
rect 16602 1448 16664 1464
rect 16602 1446 16648 1448
rect 16602 1430 16664 1446
rect 16676 1430 16682 1478
rect 16685 1470 16765 1478
rect 16685 1468 16704 1470
rect 16719 1468 16753 1470
rect 16685 1452 16765 1468
rect 16685 1430 16704 1452
rect 16719 1436 16749 1452
rect 16777 1446 16783 1520
rect 16786 1446 16805 1590
rect 16820 1446 16826 1590
rect 16835 1520 16848 1590
rect 16900 1586 16922 1590
rect 16893 1564 16922 1578
rect 16975 1564 16991 1578
rect 17029 1574 17035 1576
rect 17042 1574 17150 1590
rect 17157 1574 17163 1576
rect 17171 1574 17186 1590
rect 17252 1584 17271 1587
rect 16893 1562 16991 1564
rect 17018 1562 17186 1574
rect 17201 1564 17217 1578
rect 17252 1565 17274 1584
rect 17284 1578 17300 1579
rect 17283 1576 17300 1578
rect 17284 1571 17300 1576
rect 17274 1564 17280 1565
rect 17283 1564 17312 1571
rect 17201 1563 17312 1564
rect 17201 1562 17318 1563
rect 16877 1554 16928 1562
rect 16975 1554 17009 1562
rect 16877 1542 16902 1554
rect 16909 1542 16928 1554
rect 16982 1552 17009 1554
rect 17018 1552 17239 1562
rect 17274 1559 17280 1562
rect 16982 1548 17239 1552
rect 16877 1534 16928 1542
rect 16975 1534 17239 1548
rect 17283 1554 17318 1562
rect 16829 1486 16848 1520
rect 16893 1526 16922 1534
rect 16893 1520 16910 1526
rect 16893 1518 16927 1520
rect 16975 1518 16991 1534
rect 16992 1524 17200 1534
rect 17201 1524 17217 1534
rect 17265 1530 17280 1545
rect 17283 1542 17284 1554
rect 17291 1542 17318 1554
rect 17283 1534 17318 1542
rect 17283 1533 17312 1534
rect 17003 1520 17217 1524
rect 17018 1518 17217 1520
rect 17252 1520 17265 1530
rect 17283 1520 17300 1533
rect 17252 1518 17300 1520
rect 16894 1514 16927 1518
rect 16890 1512 16927 1514
rect 16890 1511 16957 1512
rect 16890 1506 16921 1511
rect 16927 1506 16957 1511
rect 16890 1502 16957 1506
rect 16863 1499 16957 1502
rect 16863 1492 16912 1499
rect 16863 1486 16893 1492
rect 16912 1487 16917 1492
rect 16829 1470 16909 1486
rect 16921 1478 16957 1499
rect 17018 1494 17207 1518
rect 17252 1517 17299 1518
rect 17265 1512 17299 1517
rect 17033 1491 17207 1494
rect 17026 1488 17207 1491
rect 17235 1511 17299 1512
rect 16829 1468 16848 1470
rect 16863 1468 16897 1470
rect 16829 1452 16909 1468
rect 16829 1446 16848 1452
rect 16545 1420 16648 1430
rect 16499 1418 16648 1420
rect 16669 1418 16704 1430
rect 16338 1416 16500 1418
rect 16350 1396 16369 1416
rect 16384 1414 16414 1416
rect 16233 1388 16274 1396
rect 16356 1392 16369 1396
rect 16421 1400 16500 1416
rect 16532 1416 16704 1418
rect 16532 1400 16611 1416
rect 16618 1414 16648 1416
rect 16196 1378 16225 1388
rect 16239 1378 16268 1388
rect 16283 1378 16313 1392
rect 16356 1378 16399 1392
rect 16421 1388 16611 1400
rect 16676 1396 16682 1416
rect 16406 1378 16436 1388
rect 16437 1378 16595 1388
rect 16599 1378 16629 1388
rect 16633 1378 16663 1392
rect 16691 1378 16704 1416
rect 16776 1430 16805 1446
rect 16819 1430 16848 1446
rect 16863 1436 16893 1452
rect 16921 1430 16927 1478
rect 16930 1472 16949 1478
rect 16964 1472 16994 1480
rect 16930 1464 16994 1472
rect 16930 1448 17010 1464
rect 17026 1457 17088 1488
rect 17104 1457 17166 1488
rect 17235 1486 17284 1511
rect 17299 1486 17329 1502
rect 17198 1472 17228 1480
rect 17235 1478 17345 1486
rect 17198 1464 17243 1472
rect 16930 1446 16949 1448
rect 16964 1446 17010 1448
rect 16930 1430 17010 1446
rect 17037 1444 17072 1457
rect 17113 1454 17150 1457
rect 17113 1452 17155 1454
rect 17042 1441 17072 1444
rect 17051 1437 17058 1441
rect 17058 1436 17059 1437
rect 17017 1430 17027 1436
rect 16776 1422 16811 1430
rect 16776 1396 16777 1422
rect 16784 1396 16811 1422
rect 16719 1378 16749 1392
rect 16776 1388 16811 1396
rect 16813 1422 16854 1430
rect 16813 1396 16828 1422
rect 16835 1396 16854 1422
rect 16918 1418 16949 1430
rect 16964 1418 17067 1430
rect 17079 1420 17105 1446
rect 17120 1441 17150 1452
rect 17182 1448 17244 1464
rect 17182 1446 17228 1448
rect 17182 1430 17244 1446
rect 17256 1430 17262 1478
rect 17265 1470 17345 1478
rect 17265 1468 17284 1470
rect 17299 1468 17333 1470
rect 17265 1452 17345 1468
rect 17265 1430 17284 1452
rect 17299 1436 17329 1452
rect 17357 1446 17363 1520
rect 17366 1446 17385 1590
rect 17400 1446 17406 1590
rect 17415 1520 17428 1590
rect 17480 1586 17502 1590
rect 17473 1564 17502 1578
rect 17555 1564 17571 1578
rect 17609 1574 17615 1576
rect 17622 1574 17730 1590
rect 17737 1574 17743 1576
rect 17751 1574 17766 1590
rect 17832 1584 17851 1587
rect 17473 1562 17571 1564
rect 17598 1562 17766 1574
rect 17781 1564 17797 1578
rect 17832 1565 17854 1584
rect 17864 1578 17880 1579
rect 17863 1576 17880 1578
rect 17864 1571 17880 1576
rect 17854 1564 17860 1565
rect 17863 1564 17892 1571
rect 17781 1563 17892 1564
rect 17781 1562 17898 1563
rect 17457 1554 17508 1562
rect 17555 1554 17589 1562
rect 17457 1542 17482 1554
rect 17489 1542 17508 1554
rect 17562 1552 17589 1554
rect 17598 1552 17819 1562
rect 17854 1559 17860 1562
rect 17562 1548 17819 1552
rect 17457 1534 17508 1542
rect 17555 1534 17819 1548
rect 17863 1554 17898 1562
rect 17409 1486 17428 1520
rect 17473 1526 17502 1534
rect 17473 1520 17490 1526
rect 17473 1518 17507 1520
rect 17555 1518 17571 1534
rect 17572 1524 17780 1534
rect 17781 1524 17797 1534
rect 17845 1530 17860 1545
rect 17863 1542 17864 1554
rect 17871 1542 17898 1554
rect 17863 1534 17898 1542
rect 17863 1533 17892 1534
rect 17583 1520 17797 1524
rect 17598 1518 17797 1520
rect 17832 1520 17845 1530
rect 17863 1520 17880 1533
rect 17832 1518 17880 1520
rect 17474 1514 17507 1518
rect 17470 1512 17507 1514
rect 17470 1511 17537 1512
rect 17470 1506 17501 1511
rect 17507 1506 17537 1511
rect 17470 1502 17537 1506
rect 17443 1499 17537 1502
rect 17443 1492 17492 1499
rect 17443 1486 17473 1492
rect 17492 1487 17497 1492
rect 17409 1470 17489 1486
rect 17501 1478 17537 1499
rect 17598 1494 17787 1518
rect 17832 1517 17879 1518
rect 17845 1512 17879 1517
rect 17613 1491 17787 1494
rect 17606 1488 17787 1491
rect 17815 1511 17879 1512
rect 17409 1468 17428 1470
rect 17443 1468 17477 1470
rect 17409 1452 17489 1468
rect 17409 1446 17428 1452
rect 17125 1420 17228 1430
rect 17079 1418 17228 1420
rect 17249 1418 17284 1430
rect 16918 1416 17080 1418
rect 16930 1396 16949 1416
rect 16964 1414 16994 1416
rect 16813 1388 16854 1396
rect 16936 1392 16949 1396
rect 17001 1400 17080 1416
rect 17112 1416 17284 1418
rect 17112 1400 17191 1416
rect 17198 1414 17228 1416
rect 16776 1378 16805 1388
rect 16819 1378 16848 1388
rect 16863 1378 16893 1392
rect 16936 1378 16979 1392
rect 17001 1388 17191 1400
rect 17256 1396 17262 1416
rect 16986 1378 17016 1388
rect 17017 1378 17175 1388
rect 17179 1378 17209 1388
rect 17213 1378 17243 1392
rect 17271 1378 17284 1416
rect 17356 1430 17385 1446
rect 17399 1430 17428 1446
rect 17443 1436 17473 1452
rect 17501 1430 17507 1478
rect 17510 1472 17529 1478
rect 17544 1472 17574 1480
rect 17510 1464 17574 1472
rect 17510 1448 17590 1464
rect 17606 1457 17668 1488
rect 17684 1457 17746 1488
rect 17815 1486 17864 1511
rect 17879 1486 17909 1502
rect 17778 1472 17808 1480
rect 17815 1478 17925 1486
rect 17778 1464 17823 1472
rect 17510 1446 17529 1448
rect 17544 1446 17590 1448
rect 17510 1430 17590 1446
rect 17617 1444 17652 1457
rect 17693 1454 17730 1457
rect 17693 1452 17735 1454
rect 17622 1441 17652 1444
rect 17631 1437 17638 1441
rect 17638 1436 17639 1437
rect 17597 1430 17607 1436
rect 17356 1422 17391 1430
rect 17356 1396 17357 1422
rect 17364 1396 17391 1422
rect 17299 1378 17329 1392
rect 17356 1388 17391 1396
rect 17393 1422 17434 1430
rect 17393 1396 17408 1422
rect 17415 1396 17434 1422
rect 17498 1418 17529 1430
rect 17544 1418 17647 1430
rect 17659 1420 17685 1446
rect 17700 1441 17730 1452
rect 17762 1448 17824 1464
rect 17762 1446 17808 1448
rect 17762 1430 17824 1446
rect 17836 1430 17842 1478
rect 17845 1470 17925 1478
rect 17845 1468 17864 1470
rect 17879 1468 17913 1470
rect 17845 1452 17925 1468
rect 17845 1430 17864 1452
rect 17879 1436 17909 1452
rect 17937 1446 17943 1520
rect 17946 1446 17965 1590
rect 17980 1446 17986 1590
rect 17995 1520 18008 1590
rect 18060 1586 18082 1590
rect 18053 1564 18082 1578
rect 18135 1564 18151 1578
rect 18189 1574 18195 1576
rect 18202 1574 18310 1590
rect 18317 1574 18323 1576
rect 18331 1574 18346 1590
rect 18412 1584 18431 1587
rect 18053 1562 18151 1564
rect 18178 1562 18346 1574
rect 18361 1564 18377 1578
rect 18412 1565 18434 1584
rect 18444 1578 18460 1579
rect 18443 1576 18460 1578
rect 18444 1571 18460 1576
rect 18434 1564 18440 1565
rect 18443 1564 18472 1571
rect 18361 1563 18472 1564
rect 18361 1562 18478 1563
rect 18037 1554 18088 1562
rect 18135 1554 18169 1562
rect 18037 1542 18062 1554
rect 18069 1542 18088 1554
rect 18142 1552 18169 1554
rect 18178 1552 18399 1562
rect 18434 1559 18440 1562
rect 18142 1548 18399 1552
rect 18037 1534 18088 1542
rect 18135 1534 18399 1548
rect 18443 1554 18478 1562
rect 17989 1486 18008 1520
rect 18053 1526 18082 1534
rect 18053 1520 18070 1526
rect 18053 1518 18087 1520
rect 18135 1518 18151 1534
rect 18152 1524 18360 1534
rect 18361 1524 18377 1534
rect 18425 1530 18440 1545
rect 18443 1542 18444 1554
rect 18451 1542 18478 1554
rect 18443 1534 18478 1542
rect 18443 1533 18472 1534
rect 18163 1520 18377 1524
rect 18178 1518 18377 1520
rect 18412 1520 18425 1530
rect 18443 1520 18460 1533
rect 18412 1518 18460 1520
rect 18054 1514 18087 1518
rect 18050 1512 18087 1514
rect 18050 1511 18117 1512
rect 18050 1506 18081 1511
rect 18087 1506 18117 1511
rect 18050 1502 18117 1506
rect 18023 1499 18117 1502
rect 18023 1492 18072 1499
rect 18023 1486 18053 1492
rect 18072 1487 18077 1492
rect 17989 1470 18069 1486
rect 18081 1478 18117 1499
rect 18178 1494 18367 1518
rect 18412 1517 18459 1518
rect 18425 1512 18459 1517
rect 18193 1491 18367 1494
rect 18186 1488 18367 1491
rect 18395 1511 18459 1512
rect 17989 1468 18008 1470
rect 18023 1468 18057 1470
rect 17989 1452 18069 1468
rect 17989 1446 18008 1452
rect 17705 1420 17808 1430
rect 17659 1418 17808 1420
rect 17829 1418 17864 1430
rect 17498 1416 17660 1418
rect 17510 1396 17529 1416
rect 17544 1414 17574 1416
rect 17393 1388 17434 1396
rect 17516 1392 17529 1396
rect 17581 1400 17660 1416
rect 17692 1416 17864 1418
rect 17692 1400 17771 1416
rect 17778 1414 17808 1416
rect 17356 1378 17385 1388
rect 17399 1378 17428 1388
rect 17443 1378 17473 1392
rect 17516 1378 17559 1392
rect 17581 1388 17771 1400
rect 17836 1396 17842 1416
rect 17566 1378 17596 1388
rect 17597 1378 17755 1388
rect 17759 1378 17789 1388
rect 17793 1378 17823 1392
rect 17851 1378 17864 1416
rect 17936 1430 17965 1446
rect 17979 1430 18008 1446
rect 18023 1436 18053 1452
rect 18081 1430 18087 1478
rect 18090 1472 18109 1478
rect 18124 1472 18154 1480
rect 18090 1464 18154 1472
rect 18090 1448 18170 1464
rect 18186 1457 18248 1488
rect 18264 1457 18326 1488
rect 18395 1486 18444 1511
rect 18459 1486 18489 1502
rect 18358 1472 18388 1480
rect 18395 1478 18505 1486
rect 18358 1464 18403 1472
rect 18090 1446 18109 1448
rect 18124 1446 18170 1448
rect 18090 1430 18170 1446
rect 18197 1444 18232 1457
rect 18273 1454 18310 1457
rect 18273 1452 18315 1454
rect 18202 1441 18232 1444
rect 18211 1437 18218 1441
rect 18218 1436 18219 1437
rect 18177 1430 18187 1436
rect 17936 1422 17971 1430
rect 17936 1396 17937 1422
rect 17944 1396 17971 1422
rect 17879 1378 17909 1392
rect 17936 1388 17971 1396
rect 17973 1422 18014 1430
rect 17973 1396 17988 1422
rect 17995 1396 18014 1422
rect 18078 1418 18109 1430
rect 18124 1418 18227 1430
rect 18239 1420 18265 1446
rect 18280 1441 18310 1452
rect 18342 1448 18404 1464
rect 18342 1446 18388 1448
rect 18342 1430 18404 1446
rect 18416 1430 18422 1478
rect 18425 1470 18505 1478
rect 18425 1468 18444 1470
rect 18459 1468 18493 1470
rect 18425 1452 18505 1468
rect 18425 1430 18444 1452
rect 18459 1436 18489 1452
rect 18517 1446 18523 1520
rect 18532 1446 18545 1590
rect 18285 1420 18388 1430
rect 18239 1418 18388 1420
rect 18409 1418 18444 1430
rect 18078 1416 18240 1418
rect 18090 1396 18109 1416
rect 18124 1414 18154 1416
rect 17973 1388 18014 1396
rect 18096 1392 18109 1396
rect 18161 1400 18240 1416
rect 18272 1416 18444 1418
rect 18272 1400 18351 1416
rect 18358 1414 18388 1416
rect 17936 1378 17965 1388
rect 17979 1378 18008 1388
rect 18023 1378 18053 1392
rect 18096 1378 18139 1392
rect 18161 1388 18351 1400
rect 18416 1396 18422 1416
rect 18146 1378 18176 1388
rect 18177 1378 18335 1388
rect 18339 1378 18369 1388
rect 18373 1378 18403 1392
rect 18431 1378 18444 1416
rect 18516 1430 18545 1446
rect 18516 1422 18551 1430
rect 18516 1396 18517 1422
rect 18524 1396 18551 1422
rect 18459 1378 18489 1392
rect 18516 1388 18551 1396
rect 18516 1378 18545 1388
rect -1 1372 18545 1378
rect 0 1364 18545 1372
rect 15 1334 28 1364
rect 43 1350 73 1364
rect 116 1350 159 1364
rect 166 1350 386 1364
rect 393 1350 423 1364
rect 83 1336 98 1348
rect 117 1336 130 1350
rect 198 1346 351 1350
rect 80 1334 102 1336
rect 180 1334 372 1346
rect 451 1334 464 1364
rect 479 1350 509 1364
rect 546 1334 565 1364
rect 580 1334 586 1364
rect 595 1334 608 1364
rect 623 1350 653 1364
rect 696 1350 739 1364
rect 746 1350 966 1364
rect 973 1350 1003 1364
rect 663 1336 678 1348
rect 697 1336 710 1350
rect 778 1346 931 1350
rect 660 1334 682 1336
rect 760 1334 952 1346
rect 1031 1334 1044 1364
rect 1059 1350 1089 1364
rect 1126 1334 1145 1364
rect 1160 1334 1166 1364
rect 1175 1334 1188 1364
rect 1203 1350 1233 1364
rect 1276 1350 1319 1364
rect 1326 1350 1546 1364
rect 1553 1350 1583 1364
rect 1243 1336 1258 1348
rect 1277 1336 1290 1350
rect 1358 1346 1511 1350
rect 1240 1334 1262 1336
rect 1340 1334 1532 1346
rect 1611 1334 1624 1364
rect 1639 1350 1669 1364
rect 1706 1334 1725 1364
rect 1740 1334 1746 1364
rect 1755 1334 1768 1364
rect 1783 1350 1813 1364
rect 1856 1350 1899 1364
rect 1906 1350 2126 1364
rect 2133 1350 2163 1364
rect 1823 1336 1838 1348
rect 1857 1336 1870 1350
rect 1938 1346 2091 1350
rect 1820 1334 1842 1336
rect 1920 1334 2112 1346
rect 2191 1334 2204 1364
rect 2219 1350 2249 1364
rect 2286 1334 2305 1364
rect 2320 1334 2326 1364
rect 2335 1334 2348 1364
rect 2363 1350 2393 1364
rect 2436 1350 2479 1364
rect 2486 1350 2706 1364
rect 2713 1350 2743 1364
rect 2403 1336 2418 1348
rect 2437 1336 2450 1350
rect 2518 1346 2671 1350
rect 2400 1334 2422 1336
rect 2500 1334 2692 1346
rect 2771 1334 2784 1364
rect 2799 1350 2829 1364
rect 2866 1334 2885 1364
rect 2900 1334 2906 1364
rect 2915 1334 2928 1364
rect 2943 1350 2973 1364
rect 3016 1350 3059 1364
rect 3066 1350 3286 1364
rect 3293 1350 3323 1364
rect 2983 1336 2998 1348
rect 3017 1336 3030 1350
rect 3098 1346 3251 1350
rect 2980 1334 3002 1336
rect 3080 1334 3272 1346
rect 3351 1334 3364 1364
rect 3379 1350 3409 1364
rect 3446 1334 3465 1364
rect 3480 1334 3486 1364
rect 3495 1334 3508 1364
rect 3523 1350 3553 1364
rect 3596 1350 3639 1364
rect 3646 1350 3866 1364
rect 3873 1350 3903 1364
rect 3563 1336 3578 1348
rect 3597 1336 3610 1350
rect 3678 1346 3831 1350
rect 3560 1334 3582 1336
rect 3660 1334 3852 1346
rect 3931 1334 3944 1364
rect 3959 1350 3989 1364
rect 4026 1334 4045 1364
rect 4060 1334 4066 1364
rect 4075 1334 4088 1364
rect 4103 1350 4133 1364
rect 4176 1350 4219 1364
rect 4226 1350 4446 1364
rect 4453 1350 4483 1364
rect 4143 1336 4158 1348
rect 4177 1336 4190 1350
rect 4258 1346 4411 1350
rect 4140 1334 4162 1336
rect 4240 1334 4432 1346
rect 4511 1334 4524 1364
rect 4539 1350 4569 1364
rect 4606 1334 4625 1364
rect 4640 1334 4646 1364
rect 4655 1334 4668 1364
rect 4683 1350 4713 1364
rect 4756 1350 4799 1364
rect 4806 1350 5026 1364
rect 5033 1350 5063 1364
rect 4723 1336 4738 1348
rect 4757 1336 4770 1350
rect 4838 1346 4991 1350
rect 4720 1334 4742 1336
rect 4820 1334 5012 1346
rect 5091 1334 5104 1364
rect 5119 1350 5149 1364
rect 5186 1334 5205 1364
rect 5220 1334 5226 1364
rect 5235 1334 5248 1364
rect 5263 1350 5293 1364
rect 5336 1350 5379 1364
rect 5386 1350 5606 1364
rect 5613 1350 5643 1364
rect 5303 1336 5318 1348
rect 5337 1336 5350 1350
rect 5418 1346 5571 1350
rect 5300 1334 5322 1336
rect 5400 1334 5592 1346
rect 5671 1334 5684 1364
rect 5699 1350 5729 1364
rect 5766 1334 5785 1364
rect 5800 1334 5806 1364
rect 5815 1334 5828 1364
rect 5843 1350 5873 1364
rect 5916 1350 5959 1364
rect 5966 1350 6186 1364
rect 6193 1350 6223 1364
rect 5883 1336 5898 1348
rect 5917 1336 5930 1350
rect 5998 1346 6151 1350
rect 5880 1334 5902 1336
rect 5980 1334 6172 1346
rect 6251 1334 6264 1364
rect 6279 1350 6309 1364
rect 6346 1334 6365 1364
rect 6380 1334 6386 1364
rect 6395 1334 6408 1364
rect 6423 1350 6453 1364
rect 6496 1350 6539 1364
rect 6546 1350 6766 1364
rect 6773 1350 6803 1364
rect 6463 1336 6478 1348
rect 6497 1336 6510 1350
rect 6578 1346 6731 1350
rect 6460 1334 6482 1336
rect 6560 1334 6752 1346
rect 6831 1334 6844 1364
rect 6859 1350 6889 1364
rect 6926 1334 6945 1364
rect 6960 1334 6966 1364
rect 6975 1334 6988 1364
rect 7003 1350 7033 1364
rect 7076 1350 7119 1364
rect 7126 1350 7346 1364
rect 7353 1350 7383 1364
rect 7043 1336 7058 1348
rect 7077 1336 7090 1350
rect 7158 1346 7311 1350
rect 7040 1334 7062 1336
rect 7140 1334 7332 1346
rect 7411 1334 7424 1364
rect 7439 1350 7469 1364
rect 7506 1334 7525 1364
rect 7540 1334 7546 1364
rect 7555 1334 7568 1364
rect 7583 1350 7613 1364
rect 7656 1350 7699 1364
rect 7706 1350 7926 1364
rect 7933 1350 7963 1364
rect 7623 1336 7638 1348
rect 7657 1336 7670 1350
rect 7738 1346 7891 1350
rect 7620 1334 7642 1336
rect 7720 1334 7912 1346
rect 7991 1334 8004 1364
rect 8019 1350 8049 1364
rect 8086 1334 8105 1364
rect 8120 1334 8126 1364
rect 8135 1334 8148 1364
rect 8163 1350 8193 1364
rect 8236 1350 8279 1364
rect 8286 1350 8506 1364
rect 8513 1350 8543 1364
rect 8203 1336 8218 1348
rect 8237 1336 8250 1350
rect 8318 1346 8471 1350
rect 8200 1334 8222 1336
rect 8300 1334 8492 1346
rect 8571 1334 8584 1364
rect 8599 1350 8629 1364
rect 8666 1334 8685 1364
rect 8700 1334 8706 1364
rect 8715 1334 8728 1364
rect 8743 1350 8773 1364
rect 8816 1350 8859 1364
rect 8866 1350 9086 1364
rect 9093 1350 9123 1364
rect 8783 1336 8798 1348
rect 8817 1336 8830 1350
rect 8898 1346 9051 1350
rect 8780 1334 8802 1336
rect 8880 1334 9072 1346
rect 9151 1334 9164 1364
rect 9179 1350 9209 1364
rect 9246 1334 9265 1364
rect 9280 1334 9286 1364
rect 9295 1334 9308 1364
rect 9323 1350 9353 1364
rect 9396 1350 9439 1364
rect 9446 1350 9666 1364
rect 9673 1350 9703 1364
rect 9363 1336 9378 1348
rect 9397 1336 9410 1350
rect 9478 1346 9631 1350
rect 9360 1334 9382 1336
rect 9460 1334 9652 1346
rect 9731 1334 9744 1364
rect 9759 1350 9789 1364
rect 9826 1334 9845 1364
rect 9860 1334 9866 1364
rect 9875 1334 9888 1364
rect 9903 1350 9933 1364
rect 9976 1350 10019 1364
rect 10026 1350 10246 1364
rect 10253 1350 10283 1364
rect 9943 1336 9958 1348
rect 9977 1336 9990 1350
rect 10058 1346 10211 1350
rect 9940 1334 9962 1336
rect 10040 1334 10232 1346
rect 10311 1334 10324 1364
rect 10339 1350 10369 1364
rect 10406 1334 10425 1364
rect 10440 1334 10446 1364
rect 10455 1334 10468 1364
rect 10483 1350 10513 1364
rect 10556 1350 10599 1364
rect 10606 1350 10826 1364
rect 10833 1350 10863 1364
rect 10523 1336 10538 1348
rect 10557 1336 10570 1350
rect 10638 1346 10791 1350
rect 10520 1334 10542 1336
rect 10620 1334 10812 1346
rect 10891 1334 10904 1364
rect 10919 1350 10949 1364
rect 10986 1334 11005 1364
rect 11020 1334 11026 1364
rect 11035 1334 11048 1364
rect 11063 1350 11093 1364
rect 11136 1350 11179 1364
rect 11186 1350 11406 1364
rect 11413 1350 11443 1364
rect 11103 1336 11118 1348
rect 11137 1336 11150 1350
rect 11218 1346 11371 1350
rect 11100 1334 11122 1336
rect 11200 1334 11392 1346
rect 11471 1334 11484 1364
rect 11499 1350 11529 1364
rect 11566 1334 11585 1364
rect 11600 1334 11606 1364
rect 11615 1334 11628 1364
rect 11643 1350 11673 1364
rect 11716 1350 11759 1364
rect 11766 1350 11986 1364
rect 11993 1350 12023 1364
rect 11683 1336 11698 1348
rect 11717 1336 11730 1350
rect 11798 1346 11951 1350
rect 11680 1334 11702 1336
rect 11780 1334 11972 1346
rect 12051 1334 12064 1364
rect 12079 1350 12109 1364
rect 12146 1334 12165 1364
rect 12180 1334 12186 1364
rect 12195 1334 12208 1364
rect 12223 1350 12253 1364
rect 12296 1350 12339 1364
rect 12346 1350 12566 1364
rect 12573 1350 12603 1364
rect 12263 1336 12278 1348
rect 12297 1336 12310 1350
rect 12378 1346 12531 1350
rect 12260 1334 12282 1336
rect 12360 1334 12552 1346
rect 12631 1334 12644 1364
rect 12659 1350 12689 1364
rect 12726 1334 12745 1364
rect 12760 1334 12766 1364
rect 12775 1334 12788 1364
rect 12803 1350 12833 1364
rect 12876 1350 12919 1364
rect 12926 1350 13146 1364
rect 13153 1350 13183 1364
rect 12843 1336 12858 1348
rect 12877 1336 12890 1350
rect 12958 1346 13111 1350
rect 12840 1334 12862 1336
rect 12940 1334 13132 1346
rect 13211 1334 13224 1364
rect 13239 1350 13269 1364
rect 13306 1334 13325 1364
rect 13340 1334 13346 1364
rect 13355 1334 13368 1364
rect 13383 1350 13413 1364
rect 13456 1350 13499 1364
rect 13506 1350 13726 1364
rect 13733 1350 13763 1364
rect 13423 1336 13438 1348
rect 13457 1336 13470 1350
rect 13538 1346 13691 1350
rect 13420 1334 13442 1336
rect 13520 1334 13712 1346
rect 13791 1334 13804 1364
rect 13819 1350 13849 1364
rect 13886 1334 13905 1364
rect 13920 1334 13926 1364
rect 13935 1334 13948 1364
rect 13963 1350 13993 1364
rect 14036 1350 14079 1364
rect 14086 1350 14306 1364
rect 14313 1350 14343 1364
rect 14003 1336 14018 1348
rect 14037 1336 14050 1350
rect 14118 1346 14271 1350
rect 14000 1334 14022 1336
rect 14100 1334 14292 1346
rect 14371 1334 14384 1364
rect 14399 1350 14429 1364
rect 14466 1334 14485 1364
rect 14500 1334 14506 1364
rect 14515 1334 14528 1364
rect 14543 1350 14573 1364
rect 14616 1350 14659 1364
rect 14666 1350 14886 1364
rect 14893 1350 14923 1364
rect 14583 1336 14598 1348
rect 14617 1336 14630 1350
rect 14698 1346 14851 1350
rect 14580 1334 14602 1336
rect 14680 1334 14872 1346
rect 14951 1334 14964 1364
rect 14979 1350 15009 1364
rect 15046 1334 15065 1364
rect 15080 1334 15086 1364
rect 15095 1334 15108 1364
rect 15123 1350 15153 1364
rect 15196 1350 15239 1364
rect 15246 1350 15466 1364
rect 15473 1350 15503 1364
rect 15163 1336 15178 1348
rect 15197 1336 15210 1350
rect 15278 1346 15431 1350
rect 15160 1334 15182 1336
rect 15260 1334 15452 1346
rect 15531 1334 15544 1364
rect 15559 1350 15589 1364
rect 15626 1334 15645 1364
rect 15660 1334 15666 1364
rect 15675 1334 15688 1364
rect 15703 1350 15733 1364
rect 15776 1350 15819 1364
rect 15826 1350 16046 1364
rect 16053 1350 16083 1364
rect 15743 1336 15758 1348
rect 15777 1336 15790 1350
rect 15858 1346 16011 1350
rect 15740 1334 15762 1336
rect 15840 1334 16032 1346
rect 16111 1334 16124 1364
rect 16139 1350 16169 1364
rect 16206 1334 16225 1364
rect 16240 1334 16246 1364
rect 16255 1334 16268 1364
rect 16283 1350 16313 1364
rect 16356 1350 16399 1364
rect 16406 1350 16626 1364
rect 16633 1350 16663 1364
rect 16323 1336 16338 1348
rect 16357 1336 16370 1350
rect 16438 1346 16591 1350
rect 16320 1334 16342 1336
rect 16420 1334 16612 1346
rect 16691 1334 16704 1364
rect 16719 1350 16749 1364
rect 16786 1334 16805 1364
rect 16820 1334 16826 1364
rect 16835 1334 16848 1364
rect 16863 1350 16893 1364
rect 16936 1350 16979 1364
rect 16986 1350 17206 1364
rect 17213 1350 17243 1364
rect 16903 1336 16918 1348
rect 16937 1336 16950 1350
rect 17018 1346 17171 1350
rect 16900 1334 16922 1336
rect 17000 1334 17192 1346
rect 17271 1334 17284 1364
rect 17299 1350 17329 1364
rect 17366 1334 17385 1364
rect 17400 1334 17406 1364
rect 17415 1334 17428 1364
rect 17443 1350 17473 1364
rect 17516 1350 17559 1364
rect 17566 1350 17786 1364
rect 17793 1350 17823 1364
rect 17483 1336 17498 1348
rect 17517 1336 17530 1350
rect 17598 1346 17751 1350
rect 17480 1334 17502 1336
rect 17580 1334 17772 1346
rect 17851 1334 17864 1364
rect 17879 1350 17909 1364
rect 17946 1334 17965 1364
rect 17980 1334 17986 1364
rect 17995 1334 18008 1364
rect 18023 1350 18053 1364
rect 18096 1350 18139 1364
rect 18146 1350 18366 1364
rect 18373 1350 18403 1364
rect 18063 1336 18078 1348
rect 18097 1336 18110 1350
rect 18178 1346 18331 1350
rect 18060 1334 18082 1336
rect 18160 1334 18352 1346
rect 18431 1334 18444 1364
rect 18459 1350 18489 1364
rect 18532 1334 18545 1364
rect 0 1320 18545 1334
rect 15 1250 28 1320
rect 80 1316 102 1320
rect 73 1294 102 1308
rect 155 1294 171 1308
rect 209 1304 215 1306
rect 222 1304 330 1320
rect 337 1304 343 1306
rect 351 1304 366 1320
rect 432 1314 451 1317
rect 73 1292 171 1294
rect 198 1292 366 1304
rect 381 1294 397 1308
rect 432 1295 454 1314
rect 464 1308 480 1309
rect 463 1306 480 1308
rect 464 1301 480 1306
rect 454 1294 460 1295
rect 463 1294 492 1301
rect 381 1293 492 1294
rect 381 1292 498 1293
rect 57 1284 108 1292
rect 155 1284 189 1292
rect 57 1272 82 1284
rect 89 1272 108 1284
rect 162 1282 189 1284
rect 198 1282 419 1292
rect 454 1289 460 1292
rect 162 1278 419 1282
rect 57 1264 108 1272
rect 155 1264 419 1278
rect 463 1284 498 1292
rect 9 1216 28 1250
rect 73 1256 102 1264
rect 73 1250 90 1256
rect 73 1248 107 1250
rect 155 1248 171 1264
rect 172 1254 380 1264
rect 381 1254 397 1264
rect 445 1260 460 1275
rect 463 1272 464 1284
rect 471 1272 498 1284
rect 463 1264 498 1272
rect 463 1263 492 1264
rect 183 1250 397 1254
rect 198 1248 397 1250
rect 432 1250 445 1260
rect 463 1250 480 1263
rect 432 1248 480 1250
rect 74 1244 107 1248
rect 70 1242 107 1244
rect 70 1241 137 1242
rect 70 1236 101 1241
rect 107 1236 137 1241
rect 70 1232 137 1236
rect 43 1229 137 1232
rect 43 1222 92 1229
rect 43 1216 73 1222
rect 92 1217 97 1222
rect 9 1200 89 1216
rect 101 1208 137 1229
rect 198 1224 387 1248
rect 432 1247 479 1248
rect 445 1242 479 1247
rect 213 1221 387 1224
rect 206 1218 387 1221
rect 415 1241 479 1242
rect 9 1198 28 1200
rect 43 1198 77 1200
rect 9 1182 89 1198
rect 9 1176 28 1182
rect -1 1160 28 1176
rect 43 1166 73 1182
rect 101 1160 107 1208
rect 110 1202 129 1208
rect 144 1202 174 1210
rect 110 1194 174 1202
rect 110 1178 190 1194
rect 206 1187 268 1218
rect 284 1187 346 1218
rect 415 1216 464 1241
rect 479 1216 509 1232
rect 378 1202 408 1210
rect 415 1208 525 1216
rect 378 1194 423 1202
rect 110 1176 129 1178
rect 144 1176 190 1178
rect 110 1160 190 1176
rect 217 1174 252 1187
rect 293 1184 330 1187
rect 293 1182 335 1184
rect 222 1171 252 1174
rect 231 1167 238 1171
rect 238 1166 239 1167
rect 197 1160 207 1166
rect -7 1152 34 1160
rect -7 1126 8 1152
rect 15 1126 34 1152
rect 98 1148 129 1160
rect 144 1148 247 1160
rect 259 1150 285 1176
rect 300 1171 330 1182
rect 362 1178 424 1194
rect 362 1176 408 1178
rect 362 1160 424 1176
rect 436 1160 442 1208
rect 445 1200 525 1208
rect 445 1198 464 1200
rect 479 1198 513 1200
rect 445 1182 525 1198
rect 445 1160 464 1182
rect 479 1166 509 1182
rect 537 1176 543 1250
rect 546 1176 565 1320
rect 580 1176 586 1320
rect 595 1250 608 1320
rect 660 1316 682 1320
rect 653 1294 682 1308
rect 735 1294 751 1308
rect 789 1304 795 1306
rect 802 1304 910 1320
rect 917 1304 923 1306
rect 931 1304 946 1320
rect 1012 1314 1031 1317
rect 653 1292 751 1294
rect 778 1292 946 1304
rect 961 1294 977 1308
rect 1012 1295 1034 1314
rect 1044 1308 1060 1309
rect 1043 1306 1060 1308
rect 1044 1301 1060 1306
rect 1034 1294 1040 1295
rect 1043 1294 1072 1301
rect 961 1293 1072 1294
rect 961 1292 1078 1293
rect 637 1284 688 1292
rect 735 1284 769 1292
rect 637 1272 662 1284
rect 669 1272 688 1284
rect 742 1282 769 1284
rect 778 1282 999 1292
rect 1034 1289 1040 1292
rect 742 1278 999 1282
rect 637 1264 688 1272
rect 735 1264 999 1278
rect 1043 1284 1078 1292
rect 589 1216 608 1250
rect 653 1256 682 1264
rect 653 1250 670 1256
rect 653 1248 687 1250
rect 735 1248 751 1264
rect 752 1254 960 1264
rect 961 1254 977 1264
rect 1025 1260 1040 1275
rect 1043 1272 1044 1284
rect 1051 1272 1078 1284
rect 1043 1264 1078 1272
rect 1043 1263 1072 1264
rect 763 1250 977 1254
rect 778 1248 977 1250
rect 1012 1250 1025 1260
rect 1043 1250 1060 1263
rect 1012 1248 1060 1250
rect 654 1244 687 1248
rect 650 1242 687 1244
rect 650 1241 717 1242
rect 650 1236 681 1241
rect 687 1236 717 1241
rect 650 1232 717 1236
rect 623 1229 717 1232
rect 623 1222 672 1229
rect 623 1216 653 1222
rect 672 1217 677 1222
rect 589 1200 669 1216
rect 681 1208 717 1229
rect 778 1224 967 1248
rect 1012 1247 1059 1248
rect 1025 1242 1059 1247
rect 793 1221 967 1224
rect 786 1218 967 1221
rect 995 1241 1059 1242
rect 589 1198 608 1200
rect 623 1198 657 1200
rect 589 1182 669 1198
rect 589 1176 608 1182
rect 305 1150 408 1160
rect 259 1148 408 1150
rect 429 1148 464 1160
rect 98 1146 260 1148
rect 110 1126 129 1146
rect 144 1144 174 1146
rect -7 1118 34 1126
rect 116 1122 129 1126
rect 181 1130 260 1146
rect 292 1146 464 1148
rect 292 1130 371 1146
rect 378 1144 408 1146
rect -1 1108 28 1118
rect 43 1108 73 1122
rect 116 1108 159 1122
rect 181 1118 371 1130
rect 436 1126 442 1146
rect 166 1108 196 1118
rect 197 1108 355 1118
rect 359 1108 389 1118
rect 393 1108 423 1122
rect 451 1108 464 1146
rect 536 1160 565 1176
rect 579 1160 608 1176
rect 623 1166 653 1182
rect 681 1160 687 1208
rect 690 1202 709 1208
rect 724 1202 754 1210
rect 690 1194 754 1202
rect 690 1178 770 1194
rect 786 1187 848 1218
rect 864 1187 926 1218
rect 995 1216 1044 1241
rect 1059 1216 1089 1232
rect 958 1202 988 1210
rect 995 1208 1105 1216
rect 958 1194 1003 1202
rect 690 1176 709 1178
rect 724 1176 770 1178
rect 690 1160 770 1176
rect 797 1174 832 1187
rect 873 1184 910 1187
rect 873 1182 915 1184
rect 802 1171 832 1174
rect 811 1167 818 1171
rect 818 1166 819 1167
rect 777 1160 787 1166
rect 536 1152 571 1160
rect 536 1126 537 1152
rect 544 1126 571 1152
rect 479 1108 509 1122
rect 536 1118 571 1126
rect 573 1152 614 1160
rect 573 1126 588 1152
rect 595 1126 614 1152
rect 678 1148 709 1160
rect 724 1148 827 1160
rect 839 1150 865 1176
rect 880 1171 910 1182
rect 942 1178 1004 1194
rect 942 1176 988 1178
rect 942 1160 1004 1176
rect 1016 1160 1022 1208
rect 1025 1200 1105 1208
rect 1025 1198 1044 1200
rect 1059 1198 1093 1200
rect 1025 1182 1105 1198
rect 1025 1160 1044 1182
rect 1059 1166 1089 1182
rect 1117 1176 1123 1250
rect 1126 1176 1145 1320
rect 1160 1176 1166 1320
rect 1175 1250 1188 1320
rect 1240 1316 1262 1320
rect 1233 1294 1262 1308
rect 1315 1294 1331 1308
rect 1369 1304 1375 1306
rect 1382 1304 1490 1320
rect 1497 1304 1503 1306
rect 1511 1304 1526 1320
rect 1592 1314 1611 1317
rect 1233 1292 1331 1294
rect 1358 1292 1526 1304
rect 1541 1294 1557 1308
rect 1592 1295 1614 1314
rect 1624 1308 1640 1309
rect 1623 1306 1640 1308
rect 1624 1301 1640 1306
rect 1614 1294 1620 1295
rect 1623 1294 1652 1301
rect 1541 1293 1652 1294
rect 1541 1292 1658 1293
rect 1217 1284 1268 1292
rect 1315 1284 1349 1292
rect 1217 1272 1242 1284
rect 1249 1272 1268 1284
rect 1322 1282 1349 1284
rect 1358 1282 1579 1292
rect 1614 1289 1620 1292
rect 1322 1278 1579 1282
rect 1217 1264 1268 1272
rect 1315 1264 1579 1278
rect 1623 1284 1658 1292
rect 1169 1216 1188 1250
rect 1233 1256 1262 1264
rect 1233 1250 1250 1256
rect 1233 1248 1267 1250
rect 1315 1248 1331 1264
rect 1332 1254 1540 1264
rect 1541 1254 1557 1264
rect 1605 1260 1620 1275
rect 1623 1272 1624 1284
rect 1631 1272 1658 1284
rect 1623 1264 1658 1272
rect 1623 1263 1652 1264
rect 1343 1250 1557 1254
rect 1358 1248 1557 1250
rect 1592 1250 1605 1260
rect 1623 1250 1640 1263
rect 1592 1248 1640 1250
rect 1234 1244 1267 1248
rect 1230 1242 1267 1244
rect 1230 1241 1297 1242
rect 1230 1236 1261 1241
rect 1267 1236 1297 1241
rect 1230 1232 1297 1236
rect 1203 1229 1297 1232
rect 1203 1222 1252 1229
rect 1203 1216 1233 1222
rect 1252 1217 1257 1222
rect 1169 1200 1249 1216
rect 1261 1208 1297 1229
rect 1358 1224 1547 1248
rect 1592 1247 1639 1248
rect 1605 1242 1639 1247
rect 1373 1221 1547 1224
rect 1366 1218 1547 1221
rect 1575 1241 1639 1242
rect 1169 1198 1188 1200
rect 1203 1198 1237 1200
rect 1169 1182 1249 1198
rect 1169 1176 1188 1182
rect 885 1150 988 1160
rect 839 1148 988 1150
rect 1009 1148 1044 1160
rect 678 1146 840 1148
rect 690 1126 709 1146
rect 724 1144 754 1146
rect 573 1118 614 1126
rect 696 1122 709 1126
rect 761 1130 840 1146
rect 872 1146 1044 1148
rect 872 1130 951 1146
rect 958 1144 988 1146
rect 536 1108 565 1118
rect 579 1108 608 1118
rect 623 1108 653 1122
rect 696 1108 739 1122
rect 761 1118 951 1130
rect 1016 1126 1022 1146
rect 746 1108 776 1118
rect 777 1108 935 1118
rect 939 1108 969 1118
rect 973 1108 1003 1122
rect 1031 1108 1044 1146
rect 1116 1160 1145 1176
rect 1159 1160 1188 1176
rect 1203 1166 1233 1182
rect 1261 1160 1267 1208
rect 1270 1202 1289 1208
rect 1304 1202 1334 1210
rect 1270 1194 1334 1202
rect 1270 1178 1350 1194
rect 1366 1187 1428 1218
rect 1444 1187 1506 1218
rect 1575 1216 1624 1241
rect 1639 1216 1669 1232
rect 1538 1202 1568 1210
rect 1575 1208 1685 1216
rect 1538 1194 1583 1202
rect 1270 1176 1289 1178
rect 1304 1176 1350 1178
rect 1270 1160 1350 1176
rect 1377 1174 1412 1187
rect 1453 1184 1490 1187
rect 1453 1182 1495 1184
rect 1382 1171 1412 1174
rect 1391 1167 1398 1171
rect 1398 1166 1399 1167
rect 1357 1160 1367 1166
rect 1116 1152 1151 1160
rect 1116 1126 1117 1152
rect 1124 1126 1151 1152
rect 1059 1108 1089 1122
rect 1116 1118 1151 1126
rect 1153 1152 1194 1160
rect 1153 1126 1168 1152
rect 1175 1126 1194 1152
rect 1258 1148 1289 1160
rect 1304 1148 1407 1160
rect 1419 1150 1445 1176
rect 1460 1171 1490 1182
rect 1522 1178 1584 1194
rect 1522 1176 1568 1178
rect 1522 1160 1584 1176
rect 1596 1160 1602 1208
rect 1605 1200 1685 1208
rect 1605 1198 1624 1200
rect 1639 1198 1673 1200
rect 1605 1182 1685 1198
rect 1605 1160 1624 1182
rect 1639 1166 1669 1182
rect 1697 1176 1703 1250
rect 1706 1176 1725 1320
rect 1740 1176 1746 1320
rect 1755 1250 1768 1320
rect 1820 1316 1842 1320
rect 1813 1294 1842 1308
rect 1895 1294 1911 1308
rect 1949 1304 1955 1306
rect 1962 1304 2070 1320
rect 2077 1304 2083 1306
rect 2091 1304 2106 1320
rect 2172 1314 2191 1317
rect 1813 1292 1911 1294
rect 1938 1292 2106 1304
rect 2121 1294 2137 1308
rect 2172 1295 2194 1314
rect 2204 1308 2220 1309
rect 2203 1306 2220 1308
rect 2204 1301 2220 1306
rect 2194 1294 2200 1295
rect 2203 1294 2232 1301
rect 2121 1293 2232 1294
rect 2121 1292 2238 1293
rect 1797 1284 1848 1292
rect 1895 1284 1929 1292
rect 1797 1272 1822 1284
rect 1829 1272 1848 1284
rect 1902 1282 1929 1284
rect 1938 1282 2159 1292
rect 2194 1289 2200 1292
rect 1902 1278 2159 1282
rect 1797 1264 1848 1272
rect 1895 1264 2159 1278
rect 2203 1284 2238 1292
rect 1749 1216 1768 1250
rect 1813 1256 1842 1264
rect 1813 1250 1830 1256
rect 1813 1248 1847 1250
rect 1895 1248 1911 1264
rect 1912 1254 2120 1264
rect 2121 1254 2137 1264
rect 2185 1260 2200 1275
rect 2203 1272 2204 1284
rect 2211 1272 2238 1284
rect 2203 1264 2238 1272
rect 2203 1263 2232 1264
rect 1923 1250 2137 1254
rect 1938 1248 2137 1250
rect 2172 1250 2185 1260
rect 2203 1250 2220 1263
rect 2172 1248 2220 1250
rect 1814 1244 1847 1248
rect 1810 1242 1847 1244
rect 1810 1241 1877 1242
rect 1810 1236 1841 1241
rect 1847 1236 1877 1241
rect 1810 1232 1877 1236
rect 1783 1229 1877 1232
rect 1783 1222 1832 1229
rect 1783 1216 1813 1222
rect 1832 1217 1837 1222
rect 1749 1200 1829 1216
rect 1841 1208 1877 1229
rect 1938 1224 2127 1248
rect 2172 1247 2219 1248
rect 2185 1242 2219 1247
rect 1953 1221 2127 1224
rect 1946 1218 2127 1221
rect 2155 1241 2219 1242
rect 1749 1198 1768 1200
rect 1783 1198 1817 1200
rect 1749 1182 1829 1198
rect 1749 1176 1768 1182
rect 1465 1150 1568 1160
rect 1419 1148 1568 1150
rect 1589 1148 1624 1160
rect 1258 1146 1420 1148
rect 1270 1126 1289 1146
rect 1304 1144 1334 1146
rect 1153 1118 1194 1126
rect 1276 1122 1289 1126
rect 1341 1130 1420 1146
rect 1452 1146 1624 1148
rect 1452 1130 1531 1146
rect 1538 1144 1568 1146
rect 1116 1108 1145 1118
rect 1159 1108 1188 1118
rect 1203 1108 1233 1122
rect 1276 1108 1319 1122
rect 1341 1118 1531 1130
rect 1596 1126 1602 1146
rect 1326 1108 1356 1118
rect 1357 1108 1515 1118
rect 1519 1108 1549 1118
rect 1553 1108 1583 1122
rect 1611 1108 1624 1146
rect 1696 1160 1725 1176
rect 1739 1160 1768 1176
rect 1783 1166 1813 1182
rect 1841 1160 1847 1208
rect 1850 1202 1869 1208
rect 1884 1202 1914 1210
rect 1850 1194 1914 1202
rect 1850 1178 1930 1194
rect 1946 1187 2008 1218
rect 2024 1187 2086 1218
rect 2155 1216 2204 1241
rect 2219 1216 2249 1232
rect 2118 1202 2148 1210
rect 2155 1208 2265 1216
rect 2118 1194 2163 1202
rect 1850 1176 1869 1178
rect 1884 1176 1930 1178
rect 1850 1160 1930 1176
rect 1957 1174 1992 1187
rect 2033 1184 2070 1187
rect 2033 1182 2075 1184
rect 1962 1171 1992 1174
rect 1971 1167 1978 1171
rect 1978 1166 1979 1167
rect 1937 1160 1947 1166
rect 1696 1152 1731 1160
rect 1696 1126 1697 1152
rect 1704 1126 1731 1152
rect 1639 1108 1669 1122
rect 1696 1118 1731 1126
rect 1733 1152 1774 1160
rect 1733 1126 1748 1152
rect 1755 1126 1774 1152
rect 1838 1148 1869 1160
rect 1884 1148 1987 1160
rect 1999 1150 2025 1176
rect 2040 1171 2070 1182
rect 2102 1178 2164 1194
rect 2102 1176 2148 1178
rect 2102 1160 2164 1176
rect 2176 1160 2182 1208
rect 2185 1200 2265 1208
rect 2185 1198 2204 1200
rect 2219 1198 2253 1200
rect 2185 1182 2265 1198
rect 2185 1160 2204 1182
rect 2219 1166 2249 1182
rect 2277 1176 2283 1250
rect 2286 1176 2305 1320
rect 2320 1176 2326 1320
rect 2335 1250 2348 1320
rect 2400 1316 2422 1320
rect 2393 1294 2422 1308
rect 2475 1294 2491 1308
rect 2529 1304 2535 1306
rect 2542 1304 2650 1320
rect 2657 1304 2663 1306
rect 2671 1304 2686 1320
rect 2752 1314 2771 1317
rect 2393 1292 2491 1294
rect 2518 1292 2686 1304
rect 2701 1294 2717 1308
rect 2752 1295 2774 1314
rect 2784 1308 2800 1309
rect 2783 1306 2800 1308
rect 2784 1301 2800 1306
rect 2774 1294 2780 1295
rect 2783 1294 2812 1301
rect 2701 1293 2812 1294
rect 2701 1292 2818 1293
rect 2377 1284 2428 1292
rect 2475 1284 2509 1292
rect 2377 1272 2402 1284
rect 2409 1272 2428 1284
rect 2482 1282 2509 1284
rect 2518 1282 2739 1292
rect 2774 1289 2780 1292
rect 2482 1278 2739 1282
rect 2377 1264 2428 1272
rect 2475 1264 2739 1278
rect 2783 1284 2818 1292
rect 2329 1216 2348 1250
rect 2393 1256 2422 1264
rect 2393 1250 2410 1256
rect 2393 1248 2427 1250
rect 2475 1248 2491 1264
rect 2492 1254 2700 1264
rect 2701 1254 2717 1264
rect 2765 1260 2780 1275
rect 2783 1272 2784 1284
rect 2791 1272 2818 1284
rect 2783 1264 2818 1272
rect 2783 1263 2812 1264
rect 2503 1250 2717 1254
rect 2518 1248 2717 1250
rect 2752 1250 2765 1260
rect 2783 1250 2800 1263
rect 2752 1248 2800 1250
rect 2394 1244 2427 1248
rect 2390 1242 2427 1244
rect 2390 1241 2457 1242
rect 2390 1236 2421 1241
rect 2427 1236 2457 1241
rect 2390 1232 2457 1236
rect 2363 1229 2457 1232
rect 2363 1222 2412 1229
rect 2363 1216 2393 1222
rect 2412 1217 2417 1222
rect 2329 1200 2409 1216
rect 2421 1208 2457 1229
rect 2518 1224 2707 1248
rect 2752 1247 2799 1248
rect 2765 1242 2799 1247
rect 2533 1221 2707 1224
rect 2526 1218 2707 1221
rect 2735 1241 2799 1242
rect 2329 1198 2348 1200
rect 2363 1198 2397 1200
rect 2329 1182 2409 1198
rect 2329 1176 2348 1182
rect 2045 1150 2148 1160
rect 1999 1148 2148 1150
rect 2169 1148 2204 1160
rect 1838 1146 2000 1148
rect 1850 1126 1869 1146
rect 1884 1144 1914 1146
rect 1733 1118 1774 1126
rect 1856 1122 1869 1126
rect 1921 1130 2000 1146
rect 2032 1146 2204 1148
rect 2032 1130 2111 1146
rect 2118 1144 2148 1146
rect 1696 1108 1725 1118
rect 1739 1108 1768 1118
rect 1783 1108 1813 1122
rect 1856 1108 1899 1122
rect 1921 1118 2111 1130
rect 2176 1126 2182 1146
rect 1906 1108 1936 1118
rect 1937 1108 2095 1118
rect 2099 1108 2129 1118
rect 2133 1108 2163 1122
rect 2191 1108 2204 1146
rect 2276 1160 2305 1176
rect 2319 1160 2348 1176
rect 2363 1166 2393 1182
rect 2421 1160 2427 1208
rect 2430 1202 2449 1208
rect 2464 1202 2494 1210
rect 2430 1194 2494 1202
rect 2430 1178 2510 1194
rect 2526 1187 2588 1218
rect 2604 1187 2666 1218
rect 2735 1216 2784 1241
rect 2799 1216 2829 1232
rect 2698 1202 2728 1210
rect 2735 1208 2845 1216
rect 2698 1194 2743 1202
rect 2430 1176 2449 1178
rect 2464 1176 2510 1178
rect 2430 1160 2510 1176
rect 2537 1174 2572 1187
rect 2613 1184 2650 1187
rect 2613 1182 2655 1184
rect 2542 1171 2572 1174
rect 2551 1167 2558 1171
rect 2558 1166 2559 1167
rect 2517 1160 2527 1166
rect 2276 1152 2311 1160
rect 2276 1126 2277 1152
rect 2284 1126 2311 1152
rect 2219 1108 2249 1122
rect 2276 1118 2311 1126
rect 2313 1152 2354 1160
rect 2313 1126 2328 1152
rect 2335 1126 2354 1152
rect 2418 1148 2449 1160
rect 2464 1148 2567 1160
rect 2579 1150 2605 1176
rect 2620 1171 2650 1182
rect 2682 1178 2744 1194
rect 2682 1176 2728 1178
rect 2682 1160 2744 1176
rect 2756 1160 2762 1208
rect 2765 1200 2845 1208
rect 2765 1198 2784 1200
rect 2799 1198 2833 1200
rect 2765 1182 2845 1198
rect 2765 1160 2784 1182
rect 2799 1166 2829 1182
rect 2857 1176 2863 1250
rect 2866 1176 2885 1320
rect 2900 1176 2906 1320
rect 2915 1250 2928 1320
rect 2980 1316 3002 1320
rect 2973 1294 3002 1308
rect 3055 1294 3071 1308
rect 3109 1304 3115 1306
rect 3122 1304 3230 1320
rect 3237 1304 3243 1306
rect 3251 1304 3266 1320
rect 3332 1314 3351 1317
rect 2973 1292 3071 1294
rect 3098 1292 3266 1304
rect 3281 1294 3297 1308
rect 3332 1295 3354 1314
rect 3364 1308 3380 1309
rect 3363 1306 3380 1308
rect 3364 1301 3380 1306
rect 3354 1294 3360 1295
rect 3363 1294 3392 1301
rect 3281 1293 3392 1294
rect 3281 1292 3398 1293
rect 2957 1284 3008 1292
rect 3055 1284 3089 1292
rect 2957 1272 2982 1284
rect 2989 1272 3008 1284
rect 3062 1282 3089 1284
rect 3098 1282 3319 1292
rect 3354 1289 3360 1292
rect 3062 1278 3319 1282
rect 2957 1264 3008 1272
rect 3055 1264 3319 1278
rect 3363 1284 3398 1292
rect 2909 1216 2928 1250
rect 2973 1256 3002 1264
rect 2973 1250 2990 1256
rect 2973 1248 3007 1250
rect 3055 1248 3071 1264
rect 3072 1254 3280 1264
rect 3281 1254 3297 1264
rect 3345 1260 3360 1275
rect 3363 1272 3364 1284
rect 3371 1272 3398 1284
rect 3363 1264 3398 1272
rect 3363 1263 3392 1264
rect 3083 1250 3297 1254
rect 3098 1248 3297 1250
rect 3332 1250 3345 1260
rect 3363 1250 3380 1263
rect 3332 1248 3380 1250
rect 2974 1244 3007 1248
rect 2970 1242 3007 1244
rect 2970 1241 3037 1242
rect 2970 1236 3001 1241
rect 3007 1236 3037 1241
rect 2970 1232 3037 1236
rect 2943 1229 3037 1232
rect 2943 1222 2992 1229
rect 2943 1216 2973 1222
rect 2992 1217 2997 1222
rect 2909 1200 2989 1216
rect 3001 1208 3037 1229
rect 3098 1224 3287 1248
rect 3332 1247 3379 1248
rect 3345 1242 3379 1247
rect 3113 1221 3287 1224
rect 3106 1218 3287 1221
rect 3315 1241 3379 1242
rect 2909 1198 2928 1200
rect 2943 1198 2977 1200
rect 2909 1182 2989 1198
rect 2909 1176 2928 1182
rect 2625 1150 2728 1160
rect 2579 1148 2728 1150
rect 2749 1148 2784 1160
rect 2418 1146 2580 1148
rect 2430 1126 2449 1146
rect 2464 1144 2494 1146
rect 2313 1118 2354 1126
rect 2436 1122 2449 1126
rect 2501 1130 2580 1146
rect 2612 1146 2784 1148
rect 2612 1130 2691 1146
rect 2698 1144 2728 1146
rect 2276 1108 2305 1118
rect 2319 1108 2348 1118
rect 2363 1108 2393 1122
rect 2436 1108 2479 1122
rect 2501 1118 2691 1130
rect 2756 1126 2762 1146
rect 2486 1108 2516 1118
rect 2517 1108 2675 1118
rect 2679 1108 2709 1118
rect 2713 1108 2743 1122
rect 2771 1108 2784 1146
rect 2856 1160 2885 1176
rect 2899 1160 2928 1176
rect 2943 1166 2973 1182
rect 3001 1160 3007 1208
rect 3010 1202 3029 1208
rect 3044 1202 3074 1210
rect 3010 1194 3074 1202
rect 3010 1178 3090 1194
rect 3106 1187 3168 1218
rect 3184 1187 3246 1218
rect 3315 1216 3364 1241
rect 3379 1216 3409 1232
rect 3278 1202 3308 1210
rect 3315 1208 3425 1216
rect 3278 1194 3323 1202
rect 3010 1176 3029 1178
rect 3044 1176 3090 1178
rect 3010 1160 3090 1176
rect 3117 1174 3152 1187
rect 3193 1184 3230 1187
rect 3193 1182 3235 1184
rect 3122 1171 3152 1174
rect 3131 1167 3138 1171
rect 3138 1166 3139 1167
rect 3097 1160 3107 1166
rect 2856 1152 2891 1160
rect 2856 1126 2857 1152
rect 2864 1126 2891 1152
rect 2799 1108 2829 1122
rect 2856 1118 2891 1126
rect 2893 1152 2934 1160
rect 2893 1126 2908 1152
rect 2915 1126 2934 1152
rect 2998 1148 3029 1160
rect 3044 1148 3147 1160
rect 3159 1150 3185 1176
rect 3200 1171 3230 1182
rect 3262 1178 3324 1194
rect 3262 1176 3308 1178
rect 3262 1160 3324 1176
rect 3336 1160 3342 1208
rect 3345 1200 3425 1208
rect 3345 1198 3364 1200
rect 3379 1198 3413 1200
rect 3345 1182 3425 1198
rect 3345 1160 3364 1182
rect 3379 1166 3409 1182
rect 3437 1176 3443 1250
rect 3446 1176 3465 1320
rect 3480 1176 3486 1320
rect 3495 1250 3508 1320
rect 3560 1316 3582 1320
rect 3553 1294 3582 1308
rect 3635 1294 3651 1308
rect 3689 1304 3695 1306
rect 3702 1304 3810 1320
rect 3817 1304 3823 1306
rect 3831 1304 3846 1320
rect 3912 1314 3931 1317
rect 3553 1292 3651 1294
rect 3678 1292 3846 1304
rect 3861 1294 3877 1308
rect 3912 1295 3934 1314
rect 3944 1308 3960 1309
rect 3943 1306 3960 1308
rect 3944 1301 3960 1306
rect 3934 1294 3940 1295
rect 3943 1294 3972 1301
rect 3861 1293 3972 1294
rect 3861 1292 3978 1293
rect 3537 1284 3588 1292
rect 3635 1284 3669 1292
rect 3537 1272 3562 1284
rect 3569 1272 3588 1284
rect 3642 1282 3669 1284
rect 3678 1282 3899 1292
rect 3934 1289 3940 1292
rect 3642 1278 3899 1282
rect 3537 1264 3588 1272
rect 3635 1264 3899 1278
rect 3943 1284 3978 1292
rect 3489 1216 3508 1250
rect 3553 1256 3582 1264
rect 3553 1250 3570 1256
rect 3553 1248 3587 1250
rect 3635 1248 3651 1264
rect 3652 1254 3860 1264
rect 3861 1254 3877 1264
rect 3925 1260 3940 1275
rect 3943 1272 3944 1284
rect 3951 1272 3978 1284
rect 3943 1264 3978 1272
rect 3943 1263 3972 1264
rect 3663 1250 3877 1254
rect 3678 1248 3877 1250
rect 3912 1250 3925 1260
rect 3943 1250 3960 1263
rect 3912 1248 3960 1250
rect 3554 1244 3587 1248
rect 3550 1242 3587 1244
rect 3550 1241 3617 1242
rect 3550 1236 3581 1241
rect 3587 1236 3617 1241
rect 3550 1232 3617 1236
rect 3523 1229 3617 1232
rect 3523 1222 3572 1229
rect 3523 1216 3553 1222
rect 3572 1217 3577 1222
rect 3489 1200 3569 1216
rect 3581 1208 3617 1229
rect 3678 1224 3867 1248
rect 3912 1247 3959 1248
rect 3925 1242 3959 1247
rect 3693 1221 3867 1224
rect 3686 1218 3867 1221
rect 3895 1241 3959 1242
rect 3489 1198 3508 1200
rect 3523 1198 3557 1200
rect 3489 1182 3569 1198
rect 3489 1176 3508 1182
rect 3205 1150 3308 1160
rect 3159 1148 3308 1150
rect 3329 1148 3364 1160
rect 2998 1146 3160 1148
rect 3010 1126 3029 1146
rect 3044 1144 3074 1146
rect 2893 1118 2934 1126
rect 3016 1122 3029 1126
rect 3081 1130 3160 1146
rect 3192 1146 3364 1148
rect 3192 1130 3271 1146
rect 3278 1144 3308 1146
rect 2856 1108 2885 1118
rect 2899 1108 2928 1118
rect 2943 1108 2973 1122
rect 3016 1108 3059 1122
rect 3081 1118 3271 1130
rect 3336 1126 3342 1146
rect 3066 1108 3096 1118
rect 3097 1108 3255 1118
rect 3259 1108 3289 1118
rect 3293 1108 3323 1122
rect 3351 1108 3364 1146
rect 3436 1160 3465 1176
rect 3479 1160 3508 1176
rect 3523 1166 3553 1182
rect 3581 1160 3587 1208
rect 3590 1202 3609 1208
rect 3624 1202 3654 1210
rect 3590 1194 3654 1202
rect 3590 1178 3670 1194
rect 3686 1187 3748 1218
rect 3764 1187 3826 1218
rect 3895 1216 3944 1241
rect 3959 1216 3989 1232
rect 3858 1202 3888 1210
rect 3895 1208 4005 1216
rect 3858 1194 3903 1202
rect 3590 1176 3609 1178
rect 3624 1176 3670 1178
rect 3590 1160 3670 1176
rect 3697 1174 3732 1187
rect 3773 1184 3810 1187
rect 3773 1182 3815 1184
rect 3702 1171 3732 1174
rect 3711 1167 3718 1171
rect 3718 1166 3719 1167
rect 3677 1160 3687 1166
rect 3436 1152 3471 1160
rect 3436 1126 3437 1152
rect 3444 1126 3471 1152
rect 3379 1108 3409 1122
rect 3436 1118 3471 1126
rect 3473 1152 3514 1160
rect 3473 1126 3488 1152
rect 3495 1126 3514 1152
rect 3578 1148 3609 1160
rect 3624 1148 3727 1160
rect 3739 1150 3765 1176
rect 3780 1171 3810 1182
rect 3842 1178 3904 1194
rect 3842 1176 3888 1178
rect 3842 1160 3904 1176
rect 3916 1160 3922 1208
rect 3925 1200 4005 1208
rect 3925 1198 3944 1200
rect 3959 1198 3993 1200
rect 3925 1182 4005 1198
rect 3925 1160 3944 1182
rect 3959 1166 3989 1182
rect 4017 1176 4023 1250
rect 4026 1176 4045 1320
rect 4060 1176 4066 1320
rect 4075 1250 4088 1320
rect 4140 1316 4162 1320
rect 4133 1294 4162 1308
rect 4215 1294 4231 1308
rect 4269 1304 4275 1306
rect 4282 1304 4390 1320
rect 4397 1304 4403 1306
rect 4411 1304 4426 1320
rect 4492 1314 4511 1317
rect 4133 1292 4231 1294
rect 4258 1292 4426 1304
rect 4441 1294 4457 1308
rect 4492 1295 4514 1314
rect 4524 1308 4540 1309
rect 4523 1306 4540 1308
rect 4524 1301 4540 1306
rect 4514 1294 4520 1295
rect 4523 1294 4552 1301
rect 4441 1293 4552 1294
rect 4441 1292 4558 1293
rect 4117 1284 4168 1292
rect 4215 1284 4249 1292
rect 4117 1272 4142 1284
rect 4149 1272 4168 1284
rect 4222 1282 4249 1284
rect 4258 1282 4479 1292
rect 4514 1289 4520 1292
rect 4222 1278 4479 1282
rect 4117 1264 4168 1272
rect 4215 1264 4479 1278
rect 4523 1284 4558 1292
rect 4069 1216 4088 1250
rect 4133 1256 4162 1264
rect 4133 1250 4150 1256
rect 4133 1248 4167 1250
rect 4215 1248 4231 1264
rect 4232 1254 4440 1264
rect 4441 1254 4457 1264
rect 4505 1260 4520 1275
rect 4523 1272 4524 1284
rect 4531 1272 4558 1284
rect 4523 1264 4558 1272
rect 4523 1263 4552 1264
rect 4243 1250 4457 1254
rect 4258 1248 4457 1250
rect 4492 1250 4505 1260
rect 4523 1250 4540 1263
rect 4492 1248 4540 1250
rect 4134 1244 4167 1248
rect 4130 1242 4167 1244
rect 4130 1241 4197 1242
rect 4130 1236 4161 1241
rect 4167 1236 4197 1241
rect 4130 1232 4197 1236
rect 4103 1229 4197 1232
rect 4103 1222 4152 1229
rect 4103 1216 4133 1222
rect 4152 1217 4157 1222
rect 4069 1200 4149 1216
rect 4161 1208 4197 1229
rect 4258 1224 4447 1248
rect 4492 1247 4539 1248
rect 4505 1242 4539 1247
rect 4273 1221 4447 1224
rect 4266 1218 4447 1221
rect 4475 1241 4539 1242
rect 4069 1198 4088 1200
rect 4103 1198 4137 1200
rect 4069 1182 4149 1198
rect 4069 1176 4088 1182
rect 3785 1150 3888 1160
rect 3739 1148 3888 1150
rect 3909 1148 3944 1160
rect 3578 1146 3740 1148
rect 3590 1126 3609 1146
rect 3624 1144 3654 1146
rect 3473 1118 3514 1126
rect 3596 1122 3609 1126
rect 3661 1130 3740 1146
rect 3772 1146 3944 1148
rect 3772 1130 3851 1146
rect 3858 1144 3888 1146
rect 3436 1108 3465 1118
rect 3479 1108 3508 1118
rect 3523 1108 3553 1122
rect 3596 1108 3639 1122
rect 3661 1118 3851 1130
rect 3916 1126 3922 1146
rect 3646 1108 3676 1118
rect 3677 1108 3835 1118
rect 3839 1108 3869 1118
rect 3873 1108 3903 1122
rect 3931 1108 3944 1146
rect 4016 1160 4045 1176
rect 4059 1160 4088 1176
rect 4103 1166 4133 1182
rect 4161 1160 4167 1208
rect 4170 1202 4189 1208
rect 4204 1202 4234 1210
rect 4170 1194 4234 1202
rect 4170 1178 4250 1194
rect 4266 1187 4328 1218
rect 4344 1187 4406 1218
rect 4475 1216 4524 1241
rect 4539 1216 4569 1232
rect 4438 1202 4468 1210
rect 4475 1208 4585 1216
rect 4438 1194 4483 1202
rect 4170 1176 4189 1178
rect 4204 1176 4250 1178
rect 4170 1160 4250 1176
rect 4277 1174 4312 1187
rect 4353 1184 4390 1187
rect 4353 1182 4395 1184
rect 4282 1171 4312 1174
rect 4291 1167 4298 1171
rect 4298 1166 4299 1167
rect 4257 1160 4267 1166
rect 4016 1152 4051 1160
rect 4016 1126 4017 1152
rect 4024 1126 4051 1152
rect 3959 1108 3989 1122
rect 4016 1118 4051 1126
rect 4053 1152 4094 1160
rect 4053 1126 4068 1152
rect 4075 1126 4094 1152
rect 4158 1148 4189 1160
rect 4204 1148 4307 1160
rect 4319 1150 4345 1176
rect 4360 1171 4390 1182
rect 4422 1178 4484 1194
rect 4422 1176 4468 1178
rect 4422 1160 4484 1176
rect 4496 1160 4502 1208
rect 4505 1200 4585 1208
rect 4505 1198 4524 1200
rect 4539 1198 4573 1200
rect 4505 1182 4585 1198
rect 4505 1160 4524 1182
rect 4539 1166 4569 1182
rect 4597 1176 4603 1250
rect 4606 1176 4625 1320
rect 4640 1176 4646 1320
rect 4655 1250 4668 1320
rect 4720 1316 4742 1320
rect 4713 1294 4742 1308
rect 4795 1294 4811 1308
rect 4849 1304 4855 1306
rect 4862 1304 4970 1320
rect 4977 1304 4983 1306
rect 4991 1304 5006 1320
rect 5072 1314 5091 1317
rect 4713 1292 4811 1294
rect 4838 1292 5006 1304
rect 5021 1294 5037 1308
rect 5072 1295 5094 1314
rect 5104 1308 5120 1309
rect 5103 1306 5120 1308
rect 5104 1301 5120 1306
rect 5094 1294 5100 1295
rect 5103 1294 5132 1301
rect 5021 1293 5132 1294
rect 5021 1292 5138 1293
rect 4697 1284 4748 1292
rect 4795 1284 4829 1292
rect 4697 1272 4722 1284
rect 4729 1272 4748 1284
rect 4802 1282 4829 1284
rect 4838 1282 5059 1292
rect 5094 1289 5100 1292
rect 4802 1278 5059 1282
rect 4697 1264 4748 1272
rect 4795 1264 5059 1278
rect 5103 1284 5138 1292
rect 4649 1216 4668 1250
rect 4713 1256 4742 1264
rect 4713 1250 4730 1256
rect 4713 1248 4747 1250
rect 4795 1248 4811 1264
rect 4812 1254 5020 1264
rect 5021 1254 5037 1264
rect 5085 1260 5100 1275
rect 5103 1272 5104 1284
rect 5111 1272 5138 1284
rect 5103 1264 5138 1272
rect 5103 1263 5132 1264
rect 4823 1250 5037 1254
rect 4838 1248 5037 1250
rect 5072 1250 5085 1260
rect 5103 1250 5120 1263
rect 5072 1248 5120 1250
rect 4714 1244 4747 1248
rect 4710 1242 4747 1244
rect 4710 1241 4777 1242
rect 4710 1236 4741 1241
rect 4747 1236 4777 1241
rect 4710 1232 4777 1236
rect 4683 1229 4777 1232
rect 4683 1222 4732 1229
rect 4683 1216 4713 1222
rect 4732 1217 4737 1222
rect 4649 1200 4729 1216
rect 4741 1208 4777 1229
rect 4838 1224 5027 1248
rect 5072 1247 5119 1248
rect 5085 1242 5119 1247
rect 4853 1221 5027 1224
rect 4846 1218 5027 1221
rect 5055 1241 5119 1242
rect 4649 1198 4668 1200
rect 4683 1198 4717 1200
rect 4649 1182 4729 1198
rect 4649 1176 4668 1182
rect 4365 1150 4468 1160
rect 4319 1148 4468 1150
rect 4489 1148 4524 1160
rect 4158 1146 4320 1148
rect 4170 1126 4189 1146
rect 4204 1144 4234 1146
rect 4053 1118 4094 1126
rect 4176 1122 4189 1126
rect 4241 1130 4320 1146
rect 4352 1146 4524 1148
rect 4352 1130 4431 1146
rect 4438 1144 4468 1146
rect 4016 1108 4045 1118
rect 4059 1108 4088 1118
rect 4103 1108 4133 1122
rect 4176 1108 4219 1122
rect 4241 1118 4431 1130
rect 4496 1126 4502 1146
rect 4226 1108 4256 1118
rect 4257 1108 4415 1118
rect 4419 1108 4449 1118
rect 4453 1108 4483 1122
rect 4511 1108 4524 1146
rect 4596 1160 4625 1176
rect 4639 1160 4668 1176
rect 4683 1166 4713 1182
rect 4741 1160 4747 1208
rect 4750 1202 4769 1208
rect 4784 1202 4814 1210
rect 4750 1194 4814 1202
rect 4750 1178 4830 1194
rect 4846 1187 4908 1218
rect 4924 1187 4986 1218
rect 5055 1216 5104 1241
rect 5119 1216 5149 1232
rect 5018 1202 5048 1210
rect 5055 1208 5165 1216
rect 5018 1194 5063 1202
rect 4750 1176 4769 1178
rect 4784 1176 4830 1178
rect 4750 1160 4830 1176
rect 4857 1174 4892 1187
rect 4933 1184 4970 1187
rect 4933 1182 4975 1184
rect 4862 1171 4892 1174
rect 4871 1167 4878 1171
rect 4878 1166 4879 1167
rect 4837 1160 4847 1166
rect 4596 1152 4631 1160
rect 4596 1126 4597 1152
rect 4604 1126 4631 1152
rect 4539 1108 4569 1122
rect 4596 1118 4631 1126
rect 4633 1152 4674 1160
rect 4633 1126 4648 1152
rect 4655 1126 4674 1152
rect 4738 1148 4769 1160
rect 4784 1148 4887 1160
rect 4899 1150 4925 1176
rect 4940 1171 4970 1182
rect 5002 1178 5064 1194
rect 5002 1176 5048 1178
rect 5002 1160 5064 1176
rect 5076 1160 5082 1208
rect 5085 1200 5165 1208
rect 5085 1198 5104 1200
rect 5119 1198 5153 1200
rect 5085 1182 5165 1198
rect 5085 1160 5104 1182
rect 5119 1166 5149 1182
rect 5177 1176 5183 1250
rect 5186 1176 5205 1320
rect 5220 1176 5226 1320
rect 5235 1250 5248 1320
rect 5300 1316 5322 1320
rect 5293 1294 5322 1308
rect 5375 1294 5391 1308
rect 5429 1304 5435 1306
rect 5442 1304 5550 1320
rect 5557 1304 5563 1306
rect 5571 1304 5586 1320
rect 5652 1314 5671 1317
rect 5293 1292 5391 1294
rect 5418 1292 5586 1304
rect 5601 1294 5617 1308
rect 5652 1295 5674 1314
rect 5684 1308 5700 1309
rect 5683 1306 5700 1308
rect 5684 1301 5700 1306
rect 5674 1294 5680 1295
rect 5683 1294 5712 1301
rect 5601 1293 5712 1294
rect 5601 1292 5718 1293
rect 5277 1284 5328 1292
rect 5375 1284 5409 1292
rect 5277 1272 5302 1284
rect 5309 1272 5328 1284
rect 5382 1282 5409 1284
rect 5418 1282 5639 1292
rect 5674 1289 5680 1292
rect 5382 1278 5639 1282
rect 5277 1264 5328 1272
rect 5375 1264 5639 1278
rect 5683 1284 5718 1292
rect 5229 1216 5248 1250
rect 5293 1256 5322 1264
rect 5293 1250 5310 1256
rect 5293 1248 5327 1250
rect 5375 1248 5391 1264
rect 5392 1254 5600 1264
rect 5601 1254 5617 1264
rect 5665 1260 5680 1275
rect 5683 1272 5684 1284
rect 5691 1272 5718 1284
rect 5683 1264 5718 1272
rect 5683 1263 5712 1264
rect 5403 1250 5617 1254
rect 5418 1248 5617 1250
rect 5652 1250 5665 1260
rect 5683 1250 5700 1263
rect 5652 1248 5700 1250
rect 5294 1244 5327 1248
rect 5290 1242 5327 1244
rect 5290 1241 5357 1242
rect 5290 1236 5321 1241
rect 5327 1236 5357 1241
rect 5290 1232 5357 1236
rect 5263 1229 5357 1232
rect 5263 1222 5312 1229
rect 5263 1216 5293 1222
rect 5312 1217 5317 1222
rect 5229 1200 5309 1216
rect 5321 1208 5357 1229
rect 5418 1224 5607 1248
rect 5652 1247 5699 1248
rect 5665 1242 5699 1247
rect 5433 1221 5607 1224
rect 5426 1218 5607 1221
rect 5635 1241 5699 1242
rect 5229 1198 5248 1200
rect 5263 1198 5297 1200
rect 5229 1182 5309 1198
rect 5229 1176 5248 1182
rect 4945 1150 5048 1160
rect 4899 1148 5048 1150
rect 5069 1148 5104 1160
rect 4738 1146 4900 1148
rect 4750 1126 4769 1146
rect 4784 1144 4814 1146
rect 4633 1118 4674 1126
rect 4756 1122 4769 1126
rect 4821 1130 4900 1146
rect 4932 1146 5104 1148
rect 4932 1130 5011 1146
rect 5018 1144 5048 1146
rect 4596 1108 4625 1118
rect 4639 1108 4668 1118
rect 4683 1108 4713 1122
rect 4756 1108 4799 1122
rect 4821 1118 5011 1130
rect 5076 1126 5082 1146
rect 4806 1108 4836 1118
rect 4837 1108 4995 1118
rect 4999 1108 5029 1118
rect 5033 1108 5063 1122
rect 5091 1108 5104 1146
rect 5176 1160 5205 1176
rect 5219 1160 5248 1176
rect 5263 1166 5293 1182
rect 5321 1160 5327 1208
rect 5330 1202 5349 1208
rect 5364 1202 5394 1210
rect 5330 1194 5394 1202
rect 5330 1178 5410 1194
rect 5426 1187 5488 1218
rect 5504 1187 5566 1218
rect 5635 1216 5684 1241
rect 5699 1216 5729 1232
rect 5598 1202 5628 1210
rect 5635 1208 5745 1216
rect 5598 1194 5643 1202
rect 5330 1176 5349 1178
rect 5364 1176 5410 1178
rect 5330 1160 5410 1176
rect 5437 1174 5472 1187
rect 5513 1184 5550 1187
rect 5513 1182 5555 1184
rect 5442 1171 5472 1174
rect 5451 1167 5458 1171
rect 5458 1166 5459 1167
rect 5417 1160 5427 1166
rect 5176 1152 5211 1160
rect 5176 1126 5177 1152
rect 5184 1126 5211 1152
rect 5119 1108 5149 1122
rect 5176 1118 5211 1126
rect 5213 1152 5254 1160
rect 5213 1126 5228 1152
rect 5235 1126 5254 1152
rect 5318 1148 5349 1160
rect 5364 1148 5467 1160
rect 5479 1150 5505 1176
rect 5520 1171 5550 1182
rect 5582 1178 5644 1194
rect 5582 1176 5628 1178
rect 5582 1160 5644 1176
rect 5656 1160 5662 1208
rect 5665 1200 5745 1208
rect 5665 1198 5684 1200
rect 5699 1198 5733 1200
rect 5665 1182 5745 1198
rect 5665 1160 5684 1182
rect 5699 1166 5729 1182
rect 5757 1176 5763 1250
rect 5766 1176 5785 1320
rect 5800 1176 5806 1320
rect 5815 1250 5828 1320
rect 5880 1316 5902 1320
rect 5873 1294 5902 1308
rect 5955 1294 5971 1308
rect 6009 1304 6015 1306
rect 6022 1304 6130 1320
rect 6137 1304 6143 1306
rect 6151 1304 6166 1320
rect 6232 1314 6251 1317
rect 5873 1292 5971 1294
rect 5998 1292 6166 1304
rect 6181 1294 6197 1308
rect 6232 1295 6254 1314
rect 6264 1308 6280 1309
rect 6263 1306 6280 1308
rect 6264 1301 6280 1306
rect 6254 1294 6260 1295
rect 6263 1294 6292 1301
rect 6181 1293 6292 1294
rect 6181 1292 6298 1293
rect 5857 1284 5908 1292
rect 5955 1284 5989 1292
rect 5857 1272 5882 1284
rect 5889 1272 5908 1284
rect 5962 1282 5989 1284
rect 5998 1282 6219 1292
rect 6254 1289 6260 1292
rect 5962 1278 6219 1282
rect 5857 1264 5908 1272
rect 5955 1264 6219 1278
rect 6263 1284 6298 1292
rect 5809 1216 5828 1250
rect 5873 1256 5902 1264
rect 5873 1250 5890 1256
rect 5873 1248 5907 1250
rect 5955 1248 5971 1264
rect 5972 1254 6180 1264
rect 6181 1254 6197 1264
rect 6245 1260 6260 1275
rect 6263 1272 6264 1284
rect 6271 1272 6298 1284
rect 6263 1264 6298 1272
rect 6263 1263 6292 1264
rect 5983 1250 6197 1254
rect 5998 1248 6197 1250
rect 6232 1250 6245 1260
rect 6263 1250 6280 1263
rect 6232 1248 6280 1250
rect 5874 1244 5907 1248
rect 5870 1242 5907 1244
rect 5870 1241 5937 1242
rect 5870 1236 5901 1241
rect 5907 1236 5937 1241
rect 5870 1232 5937 1236
rect 5843 1229 5937 1232
rect 5843 1222 5892 1229
rect 5843 1216 5873 1222
rect 5892 1217 5897 1222
rect 5809 1200 5889 1216
rect 5901 1208 5937 1229
rect 5998 1224 6187 1248
rect 6232 1247 6279 1248
rect 6245 1242 6279 1247
rect 6013 1221 6187 1224
rect 6006 1218 6187 1221
rect 6215 1241 6279 1242
rect 5809 1198 5828 1200
rect 5843 1198 5877 1200
rect 5809 1182 5889 1198
rect 5809 1176 5828 1182
rect 5525 1150 5628 1160
rect 5479 1148 5628 1150
rect 5649 1148 5684 1160
rect 5318 1146 5480 1148
rect 5330 1126 5349 1146
rect 5364 1144 5394 1146
rect 5213 1118 5254 1126
rect 5336 1122 5349 1126
rect 5401 1130 5480 1146
rect 5512 1146 5684 1148
rect 5512 1130 5591 1146
rect 5598 1144 5628 1146
rect 5176 1108 5205 1118
rect 5219 1108 5248 1118
rect 5263 1108 5293 1122
rect 5336 1108 5379 1122
rect 5401 1118 5591 1130
rect 5656 1126 5662 1146
rect 5386 1108 5416 1118
rect 5417 1108 5575 1118
rect 5579 1108 5609 1118
rect 5613 1108 5643 1122
rect 5671 1108 5684 1146
rect 5756 1160 5785 1176
rect 5799 1160 5828 1176
rect 5843 1166 5873 1182
rect 5901 1160 5907 1208
rect 5910 1202 5929 1208
rect 5944 1202 5974 1210
rect 5910 1194 5974 1202
rect 5910 1178 5990 1194
rect 6006 1187 6068 1218
rect 6084 1187 6146 1218
rect 6215 1216 6264 1241
rect 6279 1216 6309 1232
rect 6178 1202 6208 1210
rect 6215 1208 6325 1216
rect 6178 1194 6223 1202
rect 5910 1176 5929 1178
rect 5944 1176 5990 1178
rect 5910 1160 5990 1176
rect 6017 1174 6052 1187
rect 6093 1184 6130 1187
rect 6093 1182 6135 1184
rect 6022 1171 6052 1174
rect 6031 1167 6038 1171
rect 6038 1166 6039 1167
rect 5997 1160 6007 1166
rect 5756 1152 5791 1160
rect 5756 1126 5757 1152
rect 5764 1126 5791 1152
rect 5699 1108 5729 1122
rect 5756 1118 5791 1126
rect 5793 1152 5834 1160
rect 5793 1126 5808 1152
rect 5815 1126 5834 1152
rect 5898 1148 5929 1160
rect 5944 1148 6047 1160
rect 6059 1150 6085 1176
rect 6100 1171 6130 1182
rect 6162 1178 6224 1194
rect 6162 1176 6208 1178
rect 6162 1160 6224 1176
rect 6236 1160 6242 1208
rect 6245 1200 6325 1208
rect 6245 1198 6264 1200
rect 6279 1198 6313 1200
rect 6245 1182 6325 1198
rect 6245 1160 6264 1182
rect 6279 1166 6309 1182
rect 6337 1176 6343 1250
rect 6346 1176 6365 1320
rect 6380 1176 6386 1320
rect 6395 1250 6408 1320
rect 6460 1316 6482 1320
rect 6453 1294 6482 1308
rect 6535 1294 6551 1308
rect 6589 1304 6595 1306
rect 6602 1304 6710 1320
rect 6717 1304 6723 1306
rect 6731 1304 6746 1320
rect 6812 1314 6831 1317
rect 6453 1292 6551 1294
rect 6578 1292 6746 1304
rect 6761 1294 6777 1308
rect 6812 1295 6834 1314
rect 6844 1308 6860 1309
rect 6843 1306 6860 1308
rect 6844 1301 6860 1306
rect 6834 1294 6840 1295
rect 6843 1294 6872 1301
rect 6761 1293 6872 1294
rect 6761 1292 6878 1293
rect 6437 1284 6488 1292
rect 6535 1284 6569 1292
rect 6437 1272 6462 1284
rect 6469 1272 6488 1284
rect 6542 1282 6569 1284
rect 6578 1282 6799 1292
rect 6834 1289 6840 1292
rect 6542 1278 6799 1282
rect 6437 1264 6488 1272
rect 6535 1264 6799 1278
rect 6843 1284 6878 1292
rect 6389 1216 6408 1250
rect 6453 1256 6482 1264
rect 6453 1250 6470 1256
rect 6453 1248 6487 1250
rect 6535 1248 6551 1264
rect 6552 1254 6760 1264
rect 6761 1254 6777 1264
rect 6825 1260 6840 1275
rect 6843 1272 6844 1284
rect 6851 1272 6878 1284
rect 6843 1264 6878 1272
rect 6843 1263 6872 1264
rect 6563 1250 6777 1254
rect 6578 1248 6777 1250
rect 6812 1250 6825 1260
rect 6843 1250 6860 1263
rect 6812 1248 6860 1250
rect 6454 1244 6487 1248
rect 6450 1242 6487 1244
rect 6450 1241 6517 1242
rect 6450 1236 6481 1241
rect 6487 1236 6517 1241
rect 6450 1232 6517 1236
rect 6423 1229 6517 1232
rect 6423 1222 6472 1229
rect 6423 1216 6453 1222
rect 6472 1217 6477 1222
rect 6389 1200 6469 1216
rect 6481 1208 6517 1229
rect 6578 1224 6767 1248
rect 6812 1247 6859 1248
rect 6825 1242 6859 1247
rect 6593 1221 6767 1224
rect 6586 1218 6767 1221
rect 6795 1241 6859 1242
rect 6389 1198 6408 1200
rect 6423 1198 6457 1200
rect 6389 1182 6469 1198
rect 6389 1176 6408 1182
rect 6105 1150 6208 1160
rect 6059 1148 6208 1150
rect 6229 1148 6264 1160
rect 5898 1146 6060 1148
rect 5910 1126 5929 1146
rect 5944 1144 5974 1146
rect 5793 1118 5834 1126
rect 5916 1122 5929 1126
rect 5981 1130 6060 1146
rect 6092 1146 6264 1148
rect 6092 1130 6171 1146
rect 6178 1144 6208 1146
rect 5756 1108 5785 1118
rect 5799 1108 5828 1118
rect 5843 1108 5873 1122
rect 5916 1108 5959 1122
rect 5981 1118 6171 1130
rect 6236 1126 6242 1146
rect 5966 1108 5996 1118
rect 5997 1108 6155 1118
rect 6159 1108 6189 1118
rect 6193 1108 6223 1122
rect 6251 1108 6264 1146
rect 6336 1160 6365 1176
rect 6379 1160 6408 1176
rect 6423 1166 6453 1182
rect 6481 1160 6487 1208
rect 6490 1202 6509 1208
rect 6524 1202 6554 1210
rect 6490 1194 6554 1202
rect 6490 1178 6570 1194
rect 6586 1187 6648 1218
rect 6664 1187 6726 1218
rect 6795 1216 6844 1241
rect 6859 1216 6889 1232
rect 6758 1202 6788 1210
rect 6795 1208 6905 1216
rect 6758 1194 6803 1202
rect 6490 1176 6509 1178
rect 6524 1176 6570 1178
rect 6490 1160 6570 1176
rect 6597 1174 6632 1187
rect 6673 1184 6710 1187
rect 6673 1182 6715 1184
rect 6602 1171 6632 1174
rect 6611 1167 6618 1171
rect 6618 1166 6619 1167
rect 6577 1160 6587 1166
rect 6336 1152 6371 1160
rect 6336 1126 6337 1152
rect 6344 1126 6371 1152
rect 6279 1108 6309 1122
rect 6336 1118 6371 1126
rect 6373 1152 6414 1160
rect 6373 1126 6388 1152
rect 6395 1126 6414 1152
rect 6478 1148 6509 1160
rect 6524 1148 6627 1160
rect 6639 1150 6665 1176
rect 6680 1171 6710 1182
rect 6742 1178 6804 1194
rect 6742 1176 6788 1178
rect 6742 1160 6804 1176
rect 6816 1160 6822 1208
rect 6825 1200 6905 1208
rect 6825 1198 6844 1200
rect 6859 1198 6893 1200
rect 6825 1182 6905 1198
rect 6825 1160 6844 1182
rect 6859 1166 6889 1182
rect 6917 1176 6923 1250
rect 6926 1176 6945 1320
rect 6960 1176 6966 1320
rect 6975 1250 6988 1320
rect 7040 1316 7062 1320
rect 7033 1294 7062 1308
rect 7115 1294 7131 1308
rect 7169 1304 7175 1306
rect 7182 1304 7290 1320
rect 7297 1304 7303 1306
rect 7311 1304 7326 1320
rect 7392 1314 7411 1317
rect 7033 1292 7131 1294
rect 7158 1292 7326 1304
rect 7341 1294 7357 1308
rect 7392 1295 7414 1314
rect 7424 1308 7440 1309
rect 7423 1306 7440 1308
rect 7424 1301 7440 1306
rect 7414 1294 7420 1295
rect 7423 1294 7452 1301
rect 7341 1293 7452 1294
rect 7341 1292 7458 1293
rect 7017 1284 7068 1292
rect 7115 1284 7149 1292
rect 7017 1272 7042 1284
rect 7049 1272 7068 1284
rect 7122 1282 7149 1284
rect 7158 1282 7379 1292
rect 7414 1289 7420 1292
rect 7122 1278 7379 1282
rect 7017 1264 7068 1272
rect 7115 1264 7379 1278
rect 7423 1284 7458 1292
rect 6969 1216 6988 1250
rect 7033 1256 7062 1264
rect 7033 1250 7050 1256
rect 7033 1248 7067 1250
rect 7115 1248 7131 1264
rect 7132 1254 7340 1264
rect 7341 1254 7357 1264
rect 7405 1260 7420 1275
rect 7423 1272 7424 1284
rect 7431 1272 7458 1284
rect 7423 1264 7458 1272
rect 7423 1263 7452 1264
rect 7151 1250 7357 1254
rect 7158 1248 7357 1250
rect 7392 1250 7405 1260
rect 7423 1250 7440 1263
rect 7392 1248 7440 1250
rect 7034 1244 7067 1248
rect 7030 1242 7067 1244
rect 7030 1241 7097 1242
rect 7030 1236 7061 1241
rect 7067 1236 7097 1241
rect 7030 1232 7097 1236
rect 7003 1229 7097 1232
rect 7003 1222 7052 1229
rect 7003 1216 7033 1222
rect 7052 1217 7057 1222
rect 6969 1200 7049 1216
rect 7061 1208 7097 1229
rect 7158 1224 7347 1248
rect 7392 1247 7439 1248
rect 7405 1242 7439 1247
rect 7173 1221 7347 1224
rect 7166 1218 7347 1221
rect 7375 1241 7439 1242
rect 6969 1198 6988 1200
rect 7003 1198 7037 1200
rect 6969 1182 7049 1198
rect 6969 1176 6988 1182
rect 6685 1150 6788 1160
rect 6639 1148 6788 1150
rect 6809 1148 6844 1160
rect 6478 1146 6640 1148
rect 6490 1126 6509 1146
rect 6524 1144 6554 1146
rect 6373 1118 6414 1126
rect 6496 1122 6509 1126
rect 6561 1130 6640 1146
rect 6672 1146 6844 1148
rect 6672 1130 6751 1146
rect 6758 1144 6788 1146
rect 6336 1108 6365 1118
rect 6379 1108 6408 1118
rect 6423 1108 6453 1122
rect 6496 1108 6539 1122
rect 6561 1118 6751 1130
rect 6816 1126 6822 1146
rect 6546 1108 6576 1118
rect 6577 1108 6735 1118
rect 6739 1108 6769 1118
rect 6773 1108 6803 1122
rect 6831 1108 6844 1146
rect 6916 1160 6945 1176
rect 6959 1160 6988 1176
rect 7003 1166 7033 1182
rect 7061 1160 7067 1208
rect 7070 1202 7089 1208
rect 7104 1202 7134 1210
rect 7070 1194 7134 1202
rect 7070 1178 7150 1194
rect 7166 1187 7228 1218
rect 7244 1187 7306 1218
rect 7375 1216 7424 1241
rect 7439 1216 7469 1232
rect 7338 1202 7368 1210
rect 7375 1208 7485 1216
rect 7338 1194 7383 1202
rect 7070 1176 7089 1178
rect 7104 1176 7150 1178
rect 7070 1160 7150 1176
rect 7177 1174 7212 1187
rect 7253 1184 7290 1187
rect 7253 1182 7295 1184
rect 7182 1171 7212 1174
rect 7191 1167 7198 1171
rect 7198 1166 7199 1167
rect 7157 1160 7167 1166
rect 6916 1152 6951 1160
rect 6916 1126 6917 1152
rect 6924 1126 6951 1152
rect 6859 1108 6889 1122
rect 6916 1118 6951 1126
rect 6953 1152 6994 1160
rect 6953 1126 6968 1152
rect 6975 1126 6994 1152
rect 7058 1148 7089 1160
rect 7104 1148 7207 1160
rect 7219 1150 7245 1176
rect 7260 1171 7290 1182
rect 7322 1178 7384 1194
rect 7322 1176 7368 1178
rect 7322 1160 7384 1176
rect 7396 1160 7402 1208
rect 7405 1200 7485 1208
rect 7405 1198 7424 1200
rect 7439 1198 7473 1200
rect 7405 1182 7485 1198
rect 7405 1160 7424 1182
rect 7439 1166 7469 1182
rect 7497 1176 7503 1250
rect 7506 1176 7525 1320
rect 7540 1176 7546 1320
rect 7555 1250 7568 1320
rect 7620 1316 7642 1320
rect 7613 1294 7642 1308
rect 7695 1294 7711 1308
rect 7749 1304 7755 1306
rect 7762 1304 7870 1320
rect 7877 1304 7883 1306
rect 7891 1304 7906 1320
rect 7972 1314 7991 1317
rect 7613 1292 7711 1294
rect 7738 1292 7906 1304
rect 7921 1294 7937 1308
rect 7972 1295 7994 1314
rect 8004 1308 8020 1309
rect 8003 1306 8020 1308
rect 8004 1301 8020 1306
rect 7994 1294 8000 1295
rect 8003 1294 8032 1301
rect 7921 1293 8032 1294
rect 7921 1292 8038 1293
rect 7597 1284 7648 1292
rect 7695 1284 7729 1292
rect 7597 1272 7622 1284
rect 7629 1272 7648 1284
rect 7702 1282 7729 1284
rect 7738 1282 7959 1292
rect 7994 1289 8000 1292
rect 7702 1278 7959 1282
rect 7597 1264 7648 1272
rect 7695 1264 7959 1278
rect 8003 1284 8038 1292
rect 7549 1216 7568 1250
rect 7613 1256 7642 1264
rect 7613 1250 7630 1256
rect 7613 1248 7647 1250
rect 7695 1248 7711 1264
rect 7712 1254 7920 1264
rect 7921 1254 7937 1264
rect 7985 1260 8000 1275
rect 8003 1272 8004 1284
rect 8011 1272 8038 1284
rect 8003 1264 8038 1272
rect 8003 1263 8032 1264
rect 7723 1250 7937 1254
rect 7738 1248 7937 1250
rect 7972 1250 7985 1260
rect 8003 1250 8020 1263
rect 7972 1248 8020 1250
rect 7614 1244 7647 1248
rect 7610 1242 7647 1244
rect 7610 1241 7677 1242
rect 7610 1236 7641 1241
rect 7647 1236 7677 1241
rect 7610 1232 7677 1236
rect 7583 1229 7677 1232
rect 7583 1222 7632 1229
rect 7583 1216 7613 1222
rect 7632 1217 7637 1222
rect 7549 1200 7629 1216
rect 7641 1208 7677 1229
rect 7738 1224 7927 1248
rect 7972 1247 8019 1248
rect 7985 1242 8019 1247
rect 7753 1221 7927 1224
rect 7746 1218 7927 1221
rect 7955 1241 8019 1242
rect 7549 1198 7568 1200
rect 7583 1198 7617 1200
rect 7549 1182 7629 1198
rect 7549 1176 7568 1182
rect 7265 1150 7368 1160
rect 7219 1148 7368 1150
rect 7389 1148 7424 1160
rect 7058 1146 7220 1148
rect 7070 1126 7089 1146
rect 7104 1144 7134 1146
rect 6953 1118 6994 1126
rect 7076 1122 7089 1126
rect 7141 1130 7220 1146
rect 7252 1146 7424 1148
rect 7252 1130 7331 1146
rect 7338 1144 7368 1146
rect 6916 1108 6945 1118
rect 6959 1108 6988 1118
rect 7003 1108 7033 1122
rect 7076 1108 7119 1122
rect 7141 1118 7331 1130
rect 7396 1126 7402 1146
rect 7126 1108 7156 1118
rect 7157 1108 7315 1118
rect 7319 1108 7349 1118
rect 7353 1108 7383 1122
rect 7411 1108 7424 1146
rect 7496 1160 7525 1176
rect 7539 1160 7568 1176
rect 7583 1166 7613 1182
rect 7641 1160 7647 1208
rect 7650 1202 7669 1208
rect 7684 1202 7714 1210
rect 7650 1194 7714 1202
rect 7650 1178 7730 1194
rect 7746 1187 7808 1218
rect 7824 1187 7886 1218
rect 7955 1216 8004 1241
rect 8019 1216 8049 1232
rect 7918 1202 7948 1210
rect 7955 1208 8065 1216
rect 7918 1194 7963 1202
rect 7650 1176 7669 1178
rect 7684 1176 7730 1178
rect 7650 1160 7730 1176
rect 7757 1174 7792 1187
rect 7833 1184 7870 1187
rect 7833 1182 7875 1184
rect 7762 1171 7792 1174
rect 7771 1167 7778 1171
rect 7778 1166 7779 1167
rect 7737 1160 7747 1166
rect 7496 1152 7531 1160
rect 7496 1126 7497 1152
rect 7504 1126 7531 1152
rect 7439 1108 7469 1122
rect 7496 1118 7531 1126
rect 7533 1152 7574 1160
rect 7533 1126 7548 1152
rect 7555 1126 7574 1152
rect 7638 1148 7669 1160
rect 7684 1148 7787 1160
rect 7799 1150 7825 1176
rect 7840 1171 7870 1182
rect 7902 1178 7964 1194
rect 7902 1176 7948 1178
rect 7902 1160 7964 1176
rect 7976 1160 7982 1208
rect 7985 1200 8065 1208
rect 7985 1198 8004 1200
rect 8019 1198 8053 1200
rect 7985 1182 8065 1198
rect 7985 1160 8004 1182
rect 8019 1166 8049 1182
rect 8077 1176 8083 1250
rect 8086 1176 8105 1320
rect 8120 1176 8126 1320
rect 8135 1250 8148 1320
rect 8200 1316 8222 1320
rect 8193 1294 8222 1308
rect 8275 1294 8291 1308
rect 8329 1304 8335 1306
rect 8342 1304 8450 1320
rect 8457 1304 8463 1306
rect 8471 1304 8486 1320
rect 8552 1314 8571 1317
rect 8193 1292 8291 1294
rect 8318 1292 8486 1304
rect 8501 1294 8517 1308
rect 8552 1295 8574 1314
rect 8584 1308 8600 1309
rect 8583 1306 8600 1308
rect 8584 1301 8600 1306
rect 8574 1294 8580 1295
rect 8583 1294 8612 1301
rect 8501 1293 8612 1294
rect 8501 1292 8618 1293
rect 8177 1284 8228 1292
rect 8275 1284 8309 1292
rect 8177 1272 8202 1284
rect 8209 1272 8228 1284
rect 8282 1282 8309 1284
rect 8318 1282 8539 1292
rect 8574 1289 8580 1292
rect 8282 1278 8539 1282
rect 8177 1264 8228 1272
rect 8275 1264 8539 1278
rect 8583 1284 8618 1292
rect 8129 1216 8148 1250
rect 8193 1256 8222 1264
rect 8193 1250 8210 1256
rect 8193 1248 8227 1250
rect 8275 1248 8291 1264
rect 8292 1254 8500 1264
rect 8501 1254 8517 1264
rect 8565 1260 8580 1275
rect 8583 1272 8584 1284
rect 8591 1272 8618 1284
rect 8583 1264 8618 1272
rect 8583 1263 8612 1264
rect 8303 1250 8517 1254
rect 8318 1248 8517 1250
rect 8552 1250 8565 1260
rect 8583 1250 8600 1263
rect 8552 1248 8600 1250
rect 8194 1244 8227 1248
rect 8190 1242 8227 1244
rect 8190 1241 8257 1242
rect 8190 1236 8221 1241
rect 8227 1236 8257 1241
rect 8190 1232 8257 1236
rect 8163 1229 8257 1232
rect 8163 1222 8212 1229
rect 8163 1216 8193 1222
rect 8212 1217 8217 1222
rect 8129 1200 8209 1216
rect 8221 1208 8257 1229
rect 8318 1224 8507 1248
rect 8552 1247 8599 1248
rect 8565 1242 8599 1247
rect 8333 1221 8507 1224
rect 8326 1218 8507 1221
rect 8535 1241 8599 1242
rect 8129 1198 8148 1200
rect 8163 1198 8197 1200
rect 8129 1182 8209 1198
rect 8129 1176 8148 1182
rect 7845 1150 7948 1160
rect 7799 1148 7948 1150
rect 7969 1148 8004 1160
rect 7638 1146 7800 1148
rect 7650 1126 7669 1146
rect 7684 1144 7714 1146
rect 7533 1118 7574 1126
rect 7656 1122 7669 1126
rect 7721 1130 7800 1146
rect 7832 1146 8004 1148
rect 7832 1130 7911 1146
rect 7918 1144 7948 1146
rect 7496 1108 7525 1118
rect 7539 1108 7568 1118
rect 7583 1108 7613 1122
rect 7656 1108 7699 1122
rect 7721 1118 7911 1130
rect 7976 1126 7982 1146
rect 7706 1108 7736 1118
rect 7737 1108 7895 1118
rect 7899 1108 7929 1118
rect 7933 1108 7963 1122
rect 7991 1108 8004 1146
rect 8076 1160 8105 1176
rect 8119 1160 8148 1176
rect 8163 1166 8193 1182
rect 8221 1160 8227 1208
rect 8230 1202 8249 1208
rect 8264 1202 8294 1210
rect 8230 1194 8294 1202
rect 8230 1178 8310 1194
rect 8326 1187 8388 1218
rect 8404 1187 8466 1218
rect 8535 1216 8584 1241
rect 8599 1216 8629 1232
rect 8498 1202 8528 1210
rect 8535 1208 8645 1216
rect 8498 1194 8543 1202
rect 8230 1176 8249 1178
rect 8264 1176 8310 1178
rect 8230 1160 8310 1176
rect 8337 1174 8372 1187
rect 8413 1184 8450 1187
rect 8413 1182 8455 1184
rect 8342 1171 8372 1174
rect 8351 1167 8358 1171
rect 8358 1166 8359 1167
rect 8317 1160 8327 1166
rect 8076 1152 8111 1160
rect 8076 1126 8077 1152
rect 8084 1126 8111 1152
rect 8019 1108 8049 1122
rect 8076 1118 8111 1126
rect 8113 1152 8154 1160
rect 8113 1126 8128 1152
rect 8135 1126 8154 1152
rect 8218 1148 8249 1160
rect 8264 1148 8367 1160
rect 8379 1150 8405 1176
rect 8420 1171 8450 1182
rect 8482 1178 8544 1194
rect 8482 1176 8528 1178
rect 8482 1160 8544 1176
rect 8556 1160 8562 1208
rect 8565 1200 8645 1208
rect 8565 1198 8584 1200
rect 8599 1198 8633 1200
rect 8565 1182 8645 1198
rect 8565 1160 8584 1182
rect 8599 1166 8629 1182
rect 8657 1176 8663 1250
rect 8666 1176 8685 1320
rect 8700 1176 8706 1320
rect 8715 1250 8728 1320
rect 8780 1316 8802 1320
rect 8773 1294 8802 1308
rect 8855 1294 8871 1308
rect 8909 1304 8915 1306
rect 8922 1304 9030 1320
rect 9037 1304 9043 1306
rect 9051 1304 9066 1320
rect 9132 1314 9151 1317
rect 8773 1292 8871 1294
rect 8898 1292 9066 1304
rect 9081 1294 9097 1308
rect 9132 1295 9154 1314
rect 9164 1308 9180 1309
rect 9163 1306 9180 1308
rect 9164 1301 9180 1306
rect 9154 1294 9160 1295
rect 9163 1294 9192 1301
rect 9081 1293 9192 1294
rect 9081 1292 9198 1293
rect 8757 1284 8808 1292
rect 8855 1284 8889 1292
rect 8757 1272 8782 1284
rect 8789 1272 8808 1284
rect 8862 1282 8889 1284
rect 8898 1282 9119 1292
rect 9154 1289 9160 1292
rect 8862 1278 9119 1282
rect 8757 1264 8808 1272
rect 8855 1264 9119 1278
rect 9163 1284 9198 1292
rect 8709 1216 8728 1250
rect 8773 1256 8802 1264
rect 8773 1250 8790 1256
rect 8773 1248 8807 1250
rect 8855 1248 8871 1264
rect 8872 1254 9080 1264
rect 9081 1254 9097 1264
rect 9145 1260 9160 1275
rect 9163 1272 9164 1284
rect 9171 1272 9198 1284
rect 9163 1264 9198 1272
rect 9163 1263 9192 1264
rect 8883 1250 9097 1254
rect 8898 1248 9097 1250
rect 9132 1250 9145 1260
rect 9163 1250 9180 1263
rect 9132 1248 9180 1250
rect 8774 1244 8807 1248
rect 8770 1242 8807 1244
rect 8770 1241 8837 1242
rect 8770 1236 8801 1241
rect 8807 1236 8837 1241
rect 8770 1232 8837 1236
rect 8743 1229 8837 1232
rect 8743 1222 8792 1229
rect 8743 1216 8773 1222
rect 8792 1217 8797 1222
rect 8709 1200 8789 1216
rect 8801 1208 8837 1229
rect 8898 1224 9087 1248
rect 9132 1247 9179 1248
rect 9145 1242 9179 1247
rect 8913 1221 9087 1224
rect 8906 1218 9087 1221
rect 9115 1241 9179 1242
rect 8709 1198 8728 1200
rect 8743 1198 8777 1200
rect 8709 1182 8789 1198
rect 8709 1176 8728 1182
rect 8425 1150 8528 1160
rect 8379 1148 8528 1150
rect 8549 1148 8584 1160
rect 8218 1146 8380 1148
rect 8230 1126 8249 1146
rect 8264 1144 8294 1146
rect 8113 1118 8154 1126
rect 8236 1122 8249 1126
rect 8301 1130 8380 1146
rect 8412 1146 8584 1148
rect 8412 1130 8491 1146
rect 8498 1144 8528 1146
rect 8076 1108 8105 1118
rect 8119 1108 8148 1118
rect 8163 1108 8193 1122
rect 8236 1108 8279 1122
rect 8301 1118 8491 1130
rect 8556 1126 8562 1146
rect 8286 1108 8316 1118
rect 8317 1108 8475 1118
rect 8479 1108 8509 1118
rect 8513 1108 8543 1122
rect 8571 1108 8584 1146
rect 8656 1160 8685 1176
rect 8699 1160 8728 1176
rect 8743 1166 8773 1182
rect 8801 1160 8807 1208
rect 8810 1202 8829 1208
rect 8844 1202 8874 1210
rect 8810 1194 8874 1202
rect 8810 1178 8890 1194
rect 8906 1187 8968 1218
rect 8984 1187 9046 1218
rect 9115 1216 9164 1241
rect 9179 1216 9209 1232
rect 9078 1202 9108 1210
rect 9115 1208 9225 1216
rect 9078 1194 9123 1202
rect 8810 1176 8829 1178
rect 8844 1176 8890 1178
rect 8810 1160 8890 1176
rect 8917 1174 8952 1187
rect 8993 1184 9030 1187
rect 8993 1182 9035 1184
rect 8922 1171 8952 1174
rect 8931 1167 8938 1171
rect 8938 1166 8939 1167
rect 8897 1160 8907 1166
rect 8656 1152 8691 1160
rect 8656 1126 8657 1152
rect 8664 1126 8691 1152
rect 8599 1108 8629 1122
rect 8656 1118 8691 1126
rect 8693 1152 8734 1160
rect 8693 1126 8708 1152
rect 8715 1126 8734 1152
rect 8798 1148 8829 1160
rect 8844 1148 8947 1160
rect 8959 1150 8985 1176
rect 9000 1171 9030 1182
rect 9062 1178 9124 1194
rect 9062 1176 9108 1178
rect 9062 1160 9124 1176
rect 9136 1160 9142 1208
rect 9145 1200 9225 1208
rect 9145 1198 9164 1200
rect 9179 1198 9213 1200
rect 9145 1182 9225 1198
rect 9145 1160 9164 1182
rect 9179 1166 9209 1182
rect 9237 1176 9243 1250
rect 9246 1176 9265 1320
rect 9280 1176 9286 1320
rect 9295 1250 9308 1320
rect 9360 1316 9382 1320
rect 9353 1294 9382 1308
rect 9435 1294 9451 1308
rect 9489 1304 9495 1306
rect 9502 1304 9610 1320
rect 9617 1304 9623 1306
rect 9631 1304 9646 1320
rect 9712 1314 9731 1317
rect 9353 1292 9451 1294
rect 9478 1292 9646 1304
rect 9661 1294 9677 1308
rect 9712 1295 9734 1314
rect 9744 1308 9760 1309
rect 9743 1306 9760 1308
rect 9744 1301 9760 1306
rect 9734 1294 9740 1295
rect 9743 1294 9772 1301
rect 9661 1293 9772 1294
rect 9661 1292 9778 1293
rect 9337 1284 9388 1292
rect 9435 1284 9469 1292
rect 9337 1272 9362 1284
rect 9369 1272 9388 1284
rect 9442 1282 9469 1284
rect 9478 1282 9699 1292
rect 9734 1289 9740 1292
rect 9442 1278 9699 1282
rect 9337 1264 9388 1272
rect 9435 1264 9699 1278
rect 9743 1284 9778 1292
rect 9289 1216 9308 1250
rect 9353 1256 9382 1264
rect 9353 1250 9370 1256
rect 9353 1248 9387 1250
rect 9435 1248 9451 1264
rect 9452 1254 9660 1264
rect 9661 1254 9677 1264
rect 9725 1260 9740 1275
rect 9743 1272 9744 1284
rect 9751 1272 9778 1284
rect 9743 1264 9778 1272
rect 9743 1263 9772 1264
rect 9463 1250 9677 1254
rect 9478 1248 9677 1250
rect 9712 1250 9725 1260
rect 9743 1250 9760 1263
rect 9712 1248 9760 1250
rect 9354 1244 9387 1248
rect 9350 1242 9387 1244
rect 9350 1241 9417 1242
rect 9350 1236 9381 1241
rect 9387 1236 9417 1241
rect 9350 1232 9417 1236
rect 9323 1229 9417 1232
rect 9323 1222 9372 1229
rect 9323 1216 9353 1222
rect 9372 1217 9377 1222
rect 9289 1200 9369 1216
rect 9381 1208 9417 1229
rect 9478 1224 9667 1248
rect 9712 1247 9759 1248
rect 9725 1242 9759 1247
rect 9493 1221 9667 1224
rect 9486 1218 9667 1221
rect 9695 1241 9759 1242
rect 9289 1198 9308 1200
rect 9323 1198 9357 1200
rect 9289 1182 9369 1198
rect 9289 1176 9308 1182
rect 9005 1150 9108 1160
rect 8959 1148 9108 1150
rect 9129 1148 9164 1160
rect 8798 1146 8960 1148
rect 8810 1126 8829 1146
rect 8844 1144 8874 1146
rect 8693 1118 8734 1126
rect 8816 1122 8829 1126
rect 8881 1130 8960 1146
rect 8992 1146 9164 1148
rect 8992 1130 9071 1146
rect 9078 1144 9108 1146
rect 8656 1108 8685 1118
rect 8699 1108 8728 1118
rect 8743 1108 8773 1122
rect 8816 1108 8859 1122
rect 8881 1118 9071 1130
rect 9136 1126 9142 1146
rect 8866 1108 8896 1118
rect 8897 1108 9055 1118
rect 9059 1108 9089 1118
rect 9093 1108 9123 1122
rect 9151 1108 9164 1146
rect 9236 1160 9265 1176
rect 9279 1160 9308 1176
rect 9323 1166 9353 1182
rect 9381 1160 9387 1208
rect 9390 1202 9409 1208
rect 9424 1202 9454 1210
rect 9390 1194 9454 1202
rect 9390 1178 9470 1194
rect 9486 1187 9548 1218
rect 9564 1187 9626 1218
rect 9695 1216 9744 1241
rect 9759 1216 9789 1232
rect 9658 1202 9688 1210
rect 9695 1208 9805 1216
rect 9658 1194 9703 1202
rect 9390 1176 9409 1178
rect 9424 1176 9470 1178
rect 9390 1160 9470 1176
rect 9497 1174 9532 1187
rect 9573 1184 9610 1187
rect 9573 1182 9615 1184
rect 9502 1171 9532 1174
rect 9511 1167 9518 1171
rect 9518 1166 9519 1167
rect 9477 1160 9487 1166
rect 9236 1152 9271 1160
rect 9236 1126 9237 1152
rect 9244 1126 9271 1152
rect 9179 1108 9209 1122
rect 9236 1118 9271 1126
rect 9273 1152 9314 1160
rect 9273 1126 9288 1152
rect 9295 1126 9314 1152
rect 9378 1148 9409 1160
rect 9424 1148 9527 1160
rect 9539 1150 9565 1176
rect 9580 1171 9610 1182
rect 9642 1178 9704 1194
rect 9642 1176 9688 1178
rect 9642 1160 9704 1176
rect 9716 1160 9722 1208
rect 9725 1200 9805 1208
rect 9725 1198 9744 1200
rect 9759 1198 9793 1200
rect 9725 1182 9805 1198
rect 9725 1160 9744 1182
rect 9759 1166 9789 1182
rect 9817 1176 9823 1250
rect 9826 1176 9845 1320
rect 9860 1176 9866 1320
rect 9875 1250 9888 1320
rect 9940 1316 9962 1320
rect 9933 1294 9962 1308
rect 10015 1294 10031 1308
rect 10069 1304 10075 1306
rect 10082 1304 10190 1320
rect 10197 1304 10203 1306
rect 10211 1304 10226 1320
rect 10292 1314 10311 1317
rect 9933 1292 10031 1294
rect 10058 1292 10226 1304
rect 10241 1294 10257 1308
rect 10292 1295 10314 1314
rect 10324 1308 10340 1309
rect 10323 1306 10340 1308
rect 10324 1301 10340 1306
rect 10314 1294 10320 1295
rect 10323 1294 10352 1301
rect 10241 1293 10352 1294
rect 10241 1292 10358 1293
rect 9917 1284 9968 1292
rect 10015 1284 10049 1292
rect 9917 1272 9942 1284
rect 9949 1272 9968 1284
rect 10022 1282 10049 1284
rect 10058 1282 10279 1292
rect 10314 1289 10320 1292
rect 10022 1278 10279 1282
rect 9917 1264 9968 1272
rect 10015 1264 10279 1278
rect 10323 1284 10358 1292
rect 9869 1216 9888 1250
rect 9933 1256 9962 1264
rect 9933 1250 9950 1256
rect 9933 1248 9967 1250
rect 10015 1248 10031 1264
rect 10032 1254 10240 1264
rect 10241 1254 10257 1264
rect 10305 1260 10320 1275
rect 10323 1272 10324 1284
rect 10331 1272 10358 1284
rect 10323 1264 10358 1272
rect 10323 1263 10352 1264
rect 10043 1250 10257 1254
rect 10058 1248 10257 1250
rect 10292 1250 10305 1260
rect 10323 1250 10340 1263
rect 10292 1248 10340 1250
rect 9934 1244 9967 1248
rect 9930 1242 9967 1244
rect 9930 1241 9997 1242
rect 9930 1236 9961 1241
rect 9967 1236 9997 1241
rect 9930 1232 9997 1236
rect 9903 1229 9997 1232
rect 9903 1222 9952 1229
rect 9903 1216 9933 1222
rect 9952 1217 9957 1222
rect 9869 1200 9949 1216
rect 9961 1208 9997 1229
rect 10058 1224 10247 1248
rect 10292 1247 10339 1248
rect 10305 1242 10339 1247
rect 10073 1221 10247 1224
rect 10066 1218 10247 1221
rect 10275 1241 10339 1242
rect 9869 1198 9888 1200
rect 9903 1198 9937 1200
rect 9869 1182 9949 1198
rect 9869 1176 9888 1182
rect 9585 1150 9688 1160
rect 9539 1148 9688 1150
rect 9709 1148 9744 1160
rect 9378 1146 9540 1148
rect 9390 1126 9409 1146
rect 9424 1144 9454 1146
rect 9273 1118 9314 1126
rect 9396 1122 9409 1126
rect 9461 1130 9540 1146
rect 9572 1146 9744 1148
rect 9572 1130 9651 1146
rect 9658 1144 9688 1146
rect 9236 1108 9265 1118
rect 9279 1108 9308 1118
rect 9323 1108 9353 1122
rect 9396 1108 9439 1122
rect 9461 1118 9651 1130
rect 9716 1126 9722 1146
rect 9446 1108 9476 1118
rect 9477 1108 9635 1118
rect 9639 1108 9669 1118
rect 9673 1108 9703 1122
rect 9731 1108 9744 1146
rect 9816 1160 9845 1176
rect 9859 1160 9888 1176
rect 9903 1166 9933 1182
rect 9961 1160 9967 1208
rect 9970 1202 9989 1208
rect 10004 1202 10034 1210
rect 9970 1194 10034 1202
rect 9970 1178 10050 1194
rect 10066 1187 10128 1218
rect 10144 1187 10206 1218
rect 10275 1216 10324 1241
rect 10339 1216 10369 1232
rect 10238 1202 10268 1210
rect 10275 1208 10385 1216
rect 10238 1194 10283 1202
rect 9970 1176 9989 1178
rect 10004 1176 10050 1178
rect 9970 1160 10050 1176
rect 10077 1174 10112 1187
rect 10153 1184 10190 1187
rect 10153 1182 10195 1184
rect 10082 1171 10112 1174
rect 10091 1167 10098 1171
rect 10098 1166 10099 1167
rect 10057 1160 10067 1166
rect 9816 1152 9851 1160
rect 9816 1126 9817 1152
rect 9824 1126 9851 1152
rect 9759 1108 9789 1122
rect 9816 1118 9851 1126
rect 9853 1152 9894 1160
rect 9853 1126 9868 1152
rect 9875 1126 9894 1152
rect 9958 1148 9989 1160
rect 10004 1148 10107 1160
rect 10119 1150 10145 1176
rect 10160 1171 10190 1182
rect 10222 1178 10284 1194
rect 10222 1176 10268 1178
rect 10222 1160 10284 1176
rect 10296 1160 10302 1208
rect 10305 1200 10385 1208
rect 10305 1198 10324 1200
rect 10339 1198 10373 1200
rect 10305 1182 10385 1198
rect 10305 1160 10324 1182
rect 10339 1166 10369 1182
rect 10397 1176 10403 1250
rect 10406 1176 10425 1320
rect 10440 1176 10446 1320
rect 10455 1250 10468 1320
rect 10520 1316 10542 1320
rect 10513 1294 10542 1308
rect 10595 1294 10611 1308
rect 10649 1304 10655 1306
rect 10662 1304 10770 1320
rect 10777 1304 10783 1306
rect 10791 1304 10806 1320
rect 10872 1314 10891 1317
rect 10513 1292 10611 1294
rect 10638 1292 10806 1304
rect 10821 1294 10837 1308
rect 10872 1295 10894 1314
rect 10904 1308 10920 1309
rect 10903 1306 10920 1308
rect 10904 1301 10920 1306
rect 10894 1294 10900 1295
rect 10903 1294 10932 1301
rect 10821 1293 10932 1294
rect 10821 1292 10938 1293
rect 10497 1284 10548 1292
rect 10595 1284 10629 1292
rect 10497 1272 10522 1284
rect 10529 1272 10548 1284
rect 10602 1282 10629 1284
rect 10638 1282 10859 1292
rect 10894 1289 10900 1292
rect 10602 1278 10859 1282
rect 10497 1264 10548 1272
rect 10595 1264 10859 1278
rect 10903 1284 10938 1292
rect 10449 1216 10468 1250
rect 10513 1256 10542 1264
rect 10513 1250 10530 1256
rect 10513 1248 10547 1250
rect 10595 1248 10611 1264
rect 10612 1254 10820 1264
rect 10821 1254 10837 1264
rect 10885 1260 10900 1275
rect 10903 1272 10904 1284
rect 10911 1272 10938 1284
rect 10903 1264 10938 1272
rect 10903 1263 10932 1264
rect 10623 1250 10837 1254
rect 10638 1248 10837 1250
rect 10872 1250 10885 1260
rect 10903 1250 10920 1263
rect 10872 1248 10920 1250
rect 10514 1244 10547 1248
rect 10510 1242 10547 1244
rect 10510 1241 10577 1242
rect 10510 1236 10541 1241
rect 10547 1236 10577 1241
rect 10510 1232 10577 1236
rect 10483 1229 10577 1232
rect 10483 1222 10532 1229
rect 10483 1216 10513 1222
rect 10532 1217 10537 1222
rect 10449 1200 10529 1216
rect 10541 1208 10577 1229
rect 10638 1224 10827 1248
rect 10872 1247 10919 1248
rect 10885 1242 10919 1247
rect 10653 1221 10827 1224
rect 10646 1218 10827 1221
rect 10855 1241 10919 1242
rect 10449 1198 10468 1200
rect 10483 1198 10517 1200
rect 10449 1182 10529 1198
rect 10449 1176 10468 1182
rect 10165 1150 10268 1160
rect 10119 1148 10268 1150
rect 10289 1148 10324 1160
rect 9958 1146 10120 1148
rect 9970 1126 9989 1146
rect 10004 1144 10034 1146
rect 9853 1118 9894 1126
rect 9976 1122 9989 1126
rect 10041 1130 10120 1146
rect 10152 1146 10324 1148
rect 10152 1130 10231 1146
rect 10238 1144 10268 1146
rect 9816 1108 9845 1118
rect 9859 1108 9888 1118
rect 9903 1108 9933 1122
rect 9976 1108 10019 1122
rect 10041 1118 10231 1130
rect 10296 1126 10302 1146
rect 10026 1108 10056 1118
rect 10057 1108 10215 1118
rect 10219 1108 10249 1118
rect 10253 1108 10283 1122
rect 10311 1108 10324 1146
rect 10396 1160 10425 1176
rect 10439 1160 10468 1176
rect 10483 1166 10513 1182
rect 10541 1160 10547 1208
rect 10550 1202 10569 1208
rect 10584 1202 10614 1210
rect 10550 1194 10614 1202
rect 10550 1178 10630 1194
rect 10646 1187 10708 1218
rect 10724 1187 10786 1218
rect 10855 1216 10904 1241
rect 10919 1216 10949 1232
rect 10818 1202 10848 1210
rect 10855 1208 10965 1216
rect 10818 1194 10863 1202
rect 10550 1176 10569 1178
rect 10584 1176 10630 1178
rect 10550 1160 10630 1176
rect 10657 1174 10692 1187
rect 10733 1184 10770 1187
rect 10733 1182 10775 1184
rect 10662 1171 10692 1174
rect 10671 1167 10678 1171
rect 10678 1166 10679 1167
rect 10637 1160 10647 1166
rect 10396 1152 10431 1160
rect 10396 1126 10397 1152
rect 10404 1126 10431 1152
rect 10339 1108 10369 1122
rect 10396 1118 10431 1126
rect 10433 1152 10474 1160
rect 10433 1126 10448 1152
rect 10455 1126 10474 1152
rect 10538 1148 10569 1160
rect 10584 1148 10687 1160
rect 10699 1150 10725 1176
rect 10740 1171 10770 1182
rect 10802 1178 10864 1194
rect 10802 1176 10848 1178
rect 10802 1160 10864 1176
rect 10876 1160 10882 1208
rect 10885 1200 10965 1208
rect 10885 1198 10904 1200
rect 10919 1198 10953 1200
rect 10885 1182 10965 1198
rect 10885 1160 10904 1182
rect 10919 1166 10949 1182
rect 10977 1176 10983 1250
rect 10986 1176 11005 1320
rect 11020 1176 11026 1320
rect 11035 1250 11048 1320
rect 11100 1316 11122 1320
rect 11093 1294 11122 1308
rect 11175 1294 11191 1308
rect 11229 1304 11235 1306
rect 11242 1304 11350 1320
rect 11357 1304 11363 1306
rect 11371 1304 11386 1320
rect 11452 1314 11471 1317
rect 11093 1292 11191 1294
rect 11218 1292 11386 1304
rect 11401 1294 11417 1308
rect 11452 1295 11474 1314
rect 11484 1308 11500 1309
rect 11483 1306 11500 1308
rect 11484 1301 11500 1306
rect 11474 1294 11480 1295
rect 11483 1294 11512 1301
rect 11401 1293 11512 1294
rect 11401 1292 11518 1293
rect 11077 1284 11128 1292
rect 11175 1284 11209 1292
rect 11077 1272 11102 1284
rect 11109 1272 11128 1284
rect 11182 1282 11209 1284
rect 11218 1282 11439 1292
rect 11474 1289 11480 1292
rect 11182 1278 11439 1282
rect 11077 1264 11128 1272
rect 11175 1264 11439 1278
rect 11483 1284 11518 1292
rect 11029 1216 11048 1250
rect 11093 1256 11122 1264
rect 11093 1250 11110 1256
rect 11093 1248 11127 1250
rect 11175 1248 11191 1264
rect 11192 1254 11400 1264
rect 11401 1254 11417 1264
rect 11465 1260 11480 1275
rect 11483 1272 11484 1284
rect 11491 1272 11518 1284
rect 11483 1264 11518 1272
rect 11483 1263 11512 1264
rect 11203 1250 11417 1254
rect 11218 1248 11417 1250
rect 11452 1250 11465 1260
rect 11483 1250 11500 1263
rect 11452 1248 11500 1250
rect 11094 1244 11127 1248
rect 11090 1242 11127 1244
rect 11090 1241 11157 1242
rect 11090 1236 11121 1241
rect 11127 1236 11157 1241
rect 11090 1232 11157 1236
rect 11063 1229 11157 1232
rect 11063 1222 11112 1229
rect 11063 1216 11093 1222
rect 11112 1217 11117 1222
rect 11029 1200 11109 1216
rect 11121 1208 11157 1229
rect 11218 1224 11407 1248
rect 11452 1247 11499 1248
rect 11465 1242 11499 1247
rect 11233 1221 11407 1224
rect 11226 1218 11407 1221
rect 11435 1241 11499 1242
rect 11029 1198 11048 1200
rect 11063 1198 11097 1200
rect 11029 1182 11109 1198
rect 11029 1176 11048 1182
rect 10745 1150 10848 1160
rect 10699 1148 10848 1150
rect 10869 1148 10904 1160
rect 10538 1146 10700 1148
rect 10550 1126 10569 1146
rect 10584 1144 10614 1146
rect 10433 1118 10474 1126
rect 10556 1122 10569 1126
rect 10621 1130 10700 1146
rect 10732 1146 10904 1148
rect 10732 1130 10811 1146
rect 10818 1144 10848 1146
rect 10396 1108 10425 1118
rect 10439 1108 10468 1118
rect 10483 1108 10513 1122
rect 10556 1108 10599 1122
rect 10621 1118 10811 1130
rect 10876 1126 10882 1146
rect 10606 1108 10636 1118
rect 10637 1108 10795 1118
rect 10799 1108 10829 1118
rect 10833 1108 10863 1122
rect 10891 1108 10904 1146
rect 10976 1160 11005 1176
rect 11019 1160 11048 1176
rect 11063 1166 11093 1182
rect 11121 1160 11127 1208
rect 11130 1202 11149 1208
rect 11164 1202 11194 1210
rect 11130 1194 11194 1202
rect 11130 1178 11210 1194
rect 11226 1187 11288 1218
rect 11304 1187 11366 1218
rect 11435 1216 11484 1241
rect 11499 1216 11529 1232
rect 11398 1202 11428 1210
rect 11435 1208 11545 1216
rect 11398 1194 11443 1202
rect 11130 1176 11149 1178
rect 11164 1176 11210 1178
rect 11130 1160 11210 1176
rect 11237 1174 11272 1187
rect 11313 1184 11350 1187
rect 11313 1182 11355 1184
rect 11242 1171 11272 1174
rect 11251 1167 11258 1171
rect 11258 1166 11259 1167
rect 11217 1160 11227 1166
rect 10976 1152 11011 1160
rect 10976 1126 10977 1152
rect 10984 1126 11011 1152
rect 10919 1108 10949 1122
rect 10976 1118 11011 1126
rect 11013 1152 11054 1160
rect 11013 1126 11028 1152
rect 11035 1126 11054 1152
rect 11118 1148 11149 1160
rect 11164 1148 11267 1160
rect 11279 1150 11305 1176
rect 11320 1171 11350 1182
rect 11382 1178 11444 1194
rect 11382 1176 11428 1178
rect 11382 1160 11444 1176
rect 11456 1160 11462 1208
rect 11465 1200 11545 1208
rect 11465 1198 11484 1200
rect 11499 1198 11533 1200
rect 11465 1182 11545 1198
rect 11465 1160 11484 1182
rect 11499 1166 11529 1182
rect 11557 1176 11563 1250
rect 11566 1176 11585 1320
rect 11600 1176 11606 1320
rect 11615 1250 11628 1320
rect 11680 1316 11702 1320
rect 11673 1294 11702 1308
rect 11755 1294 11771 1308
rect 11809 1304 11815 1306
rect 11822 1304 11930 1320
rect 11937 1304 11943 1306
rect 11951 1304 11966 1320
rect 12032 1314 12051 1317
rect 11673 1292 11771 1294
rect 11798 1292 11966 1304
rect 11981 1294 11997 1308
rect 12032 1295 12054 1314
rect 12064 1308 12080 1309
rect 12063 1306 12080 1308
rect 12064 1301 12080 1306
rect 12054 1294 12060 1295
rect 12063 1294 12092 1301
rect 11981 1293 12092 1294
rect 11981 1292 12098 1293
rect 11657 1284 11708 1292
rect 11755 1284 11789 1292
rect 11657 1272 11682 1284
rect 11689 1272 11708 1284
rect 11762 1282 11789 1284
rect 11798 1282 12019 1292
rect 12054 1289 12060 1292
rect 11762 1278 12019 1282
rect 11657 1264 11708 1272
rect 11755 1264 12019 1278
rect 12063 1284 12098 1292
rect 11609 1216 11628 1250
rect 11673 1256 11702 1264
rect 11673 1250 11690 1256
rect 11673 1248 11707 1250
rect 11755 1248 11771 1264
rect 11772 1254 11980 1264
rect 11981 1254 11997 1264
rect 12045 1260 12060 1275
rect 12063 1272 12064 1284
rect 12071 1272 12098 1284
rect 12063 1264 12098 1272
rect 12063 1263 12092 1264
rect 11783 1250 11997 1254
rect 11798 1248 11997 1250
rect 12032 1250 12045 1260
rect 12063 1250 12080 1263
rect 12032 1248 12080 1250
rect 11674 1244 11707 1248
rect 11670 1242 11707 1244
rect 11670 1241 11737 1242
rect 11670 1236 11701 1241
rect 11707 1236 11737 1241
rect 11670 1232 11737 1236
rect 11643 1229 11737 1232
rect 11643 1222 11692 1229
rect 11643 1216 11673 1222
rect 11692 1217 11697 1222
rect 11609 1200 11689 1216
rect 11701 1208 11737 1229
rect 11798 1224 11987 1248
rect 12032 1247 12079 1248
rect 12045 1242 12079 1247
rect 11813 1221 11987 1224
rect 11806 1218 11987 1221
rect 12015 1241 12079 1242
rect 11609 1198 11628 1200
rect 11643 1198 11677 1200
rect 11609 1182 11689 1198
rect 11609 1176 11628 1182
rect 11325 1150 11428 1160
rect 11279 1148 11428 1150
rect 11449 1148 11484 1160
rect 11118 1146 11280 1148
rect 11130 1126 11149 1146
rect 11164 1144 11194 1146
rect 11013 1118 11054 1126
rect 11136 1122 11149 1126
rect 11201 1130 11280 1146
rect 11312 1146 11484 1148
rect 11312 1130 11391 1146
rect 11398 1144 11428 1146
rect 10976 1108 11005 1118
rect 11019 1108 11048 1118
rect 11063 1108 11093 1122
rect 11136 1108 11179 1122
rect 11201 1118 11391 1130
rect 11456 1126 11462 1146
rect 11186 1108 11216 1118
rect 11217 1108 11375 1118
rect 11379 1108 11409 1118
rect 11413 1108 11443 1122
rect 11471 1108 11484 1146
rect 11556 1160 11585 1176
rect 11599 1160 11628 1176
rect 11643 1166 11673 1182
rect 11701 1160 11707 1208
rect 11710 1202 11729 1208
rect 11744 1202 11774 1210
rect 11710 1194 11774 1202
rect 11710 1178 11790 1194
rect 11806 1187 11868 1218
rect 11884 1187 11946 1218
rect 12015 1216 12064 1241
rect 12079 1216 12109 1232
rect 11978 1202 12008 1210
rect 12015 1208 12125 1216
rect 11978 1194 12023 1202
rect 11710 1176 11729 1178
rect 11744 1176 11790 1178
rect 11710 1160 11790 1176
rect 11817 1174 11852 1187
rect 11893 1184 11930 1187
rect 11893 1182 11935 1184
rect 11822 1171 11852 1174
rect 11831 1167 11838 1171
rect 11838 1166 11839 1167
rect 11797 1160 11807 1166
rect 11556 1152 11591 1160
rect 11556 1126 11557 1152
rect 11564 1126 11591 1152
rect 11499 1108 11529 1122
rect 11556 1118 11591 1126
rect 11593 1152 11634 1160
rect 11593 1126 11608 1152
rect 11615 1126 11634 1152
rect 11698 1148 11729 1160
rect 11744 1148 11847 1160
rect 11859 1150 11885 1176
rect 11900 1171 11930 1182
rect 11962 1178 12024 1194
rect 11962 1176 12008 1178
rect 11962 1160 12024 1176
rect 12036 1160 12042 1208
rect 12045 1200 12125 1208
rect 12045 1198 12064 1200
rect 12079 1198 12113 1200
rect 12045 1182 12125 1198
rect 12045 1160 12064 1182
rect 12079 1166 12109 1182
rect 12137 1176 12143 1250
rect 12146 1176 12165 1320
rect 12180 1176 12186 1320
rect 12195 1250 12208 1320
rect 12260 1316 12282 1320
rect 12253 1294 12282 1308
rect 12335 1294 12351 1308
rect 12389 1304 12395 1306
rect 12402 1304 12510 1320
rect 12517 1304 12523 1306
rect 12531 1304 12546 1320
rect 12612 1314 12631 1317
rect 12253 1292 12351 1294
rect 12378 1292 12546 1304
rect 12561 1294 12577 1308
rect 12612 1295 12634 1314
rect 12644 1308 12660 1309
rect 12643 1306 12660 1308
rect 12644 1301 12660 1306
rect 12634 1294 12640 1295
rect 12643 1294 12672 1301
rect 12561 1293 12672 1294
rect 12561 1292 12678 1293
rect 12237 1284 12288 1292
rect 12335 1284 12369 1292
rect 12237 1272 12262 1284
rect 12269 1272 12288 1284
rect 12342 1282 12369 1284
rect 12378 1282 12599 1292
rect 12634 1289 12640 1292
rect 12342 1278 12599 1282
rect 12237 1264 12288 1272
rect 12335 1264 12599 1278
rect 12643 1284 12678 1292
rect 12189 1216 12208 1250
rect 12253 1256 12282 1264
rect 12253 1250 12270 1256
rect 12253 1248 12287 1250
rect 12335 1248 12351 1264
rect 12352 1254 12560 1264
rect 12561 1254 12577 1264
rect 12625 1260 12640 1275
rect 12643 1272 12644 1284
rect 12651 1272 12678 1284
rect 12643 1264 12678 1272
rect 12643 1263 12672 1264
rect 12363 1250 12577 1254
rect 12378 1248 12577 1250
rect 12612 1250 12625 1260
rect 12643 1250 12660 1263
rect 12612 1248 12660 1250
rect 12254 1244 12287 1248
rect 12250 1242 12287 1244
rect 12250 1241 12317 1242
rect 12250 1236 12281 1241
rect 12287 1236 12317 1241
rect 12250 1232 12317 1236
rect 12223 1229 12317 1232
rect 12223 1222 12272 1229
rect 12223 1216 12253 1222
rect 12272 1217 12277 1222
rect 12189 1200 12269 1216
rect 12281 1208 12317 1229
rect 12378 1224 12567 1248
rect 12612 1247 12659 1248
rect 12625 1242 12659 1247
rect 12393 1221 12567 1224
rect 12386 1218 12567 1221
rect 12595 1241 12659 1242
rect 12189 1198 12208 1200
rect 12223 1198 12257 1200
rect 12189 1182 12269 1198
rect 12189 1176 12208 1182
rect 11905 1150 12008 1160
rect 11859 1148 12008 1150
rect 12029 1148 12064 1160
rect 11698 1146 11860 1148
rect 11710 1126 11729 1146
rect 11744 1144 11774 1146
rect 11593 1118 11634 1126
rect 11716 1122 11729 1126
rect 11781 1130 11860 1146
rect 11892 1146 12064 1148
rect 11892 1130 11971 1146
rect 11978 1144 12008 1146
rect 11556 1108 11585 1118
rect 11599 1108 11628 1118
rect 11643 1108 11673 1122
rect 11716 1108 11759 1122
rect 11781 1118 11971 1130
rect 12036 1126 12042 1146
rect 11766 1108 11796 1118
rect 11797 1108 11955 1118
rect 11959 1108 11989 1118
rect 11993 1108 12023 1122
rect 12051 1108 12064 1146
rect 12136 1160 12165 1176
rect 12179 1160 12208 1176
rect 12223 1166 12253 1182
rect 12281 1160 12287 1208
rect 12290 1202 12309 1208
rect 12324 1202 12354 1210
rect 12290 1194 12354 1202
rect 12290 1178 12370 1194
rect 12386 1187 12448 1218
rect 12464 1187 12526 1218
rect 12595 1216 12644 1241
rect 12659 1216 12689 1232
rect 12558 1202 12588 1210
rect 12595 1208 12705 1216
rect 12558 1194 12603 1202
rect 12290 1176 12309 1178
rect 12324 1176 12370 1178
rect 12290 1160 12370 1176
rect 12397 1174 12432 1187
rect 12473 1184 12510 1187
rect 12473 1182 12515 1184
rect 12402 1171 12432 1174
rect 12411 1167 12418 1171
rect 12418 1166 12419 1167
rect 12377 1160 12387 1166
rect 12136 1152 12171 1160
rect 12136 1126 12137 1152
rect 12144 1126 12171 1152
rect 12079 1108 12109 1122
rect 12136 1118 12171 1126
rect 12173 1152 12214 1160
rect 12173 1126 12188 1152
rect 12195 1126 12214 1152
rect 12278 1148 12309 1160
rect 12324 1148 12427 1160
rect 12439 1150 12465 1176
rect 12480 1171 12510 1182
rect 12542 1178 12604 1194
rect 12542 1176 12588 1178
rect 12542 1160 12604 1176
rect 12616 1160 12622 1208
rect 12625 1200 12705 1208
rect 12625 1198 12644 1200
rect 12659 1198 12693 1200
rect 12625 1182 12705 1198
rect 12625 1160 12644 1182
rect 12659 1166 12689 1182
rect 12717 1176 12723 1250
rect 12726 1176 12745 1320
rect 12760 1176 12766 1320
rect 12775 1250 12788 1320
rect 12840 1316 12862 1320
rect 12833 1294 12862 1308
rect 12915 1294 12931 1308
rect 12969 1304 12975 1306
rect 12982 1304 13090 1320
rect 13097 1304 13103 1306
rect 13111 1304 13126 1320
rect 13192 1314 13211 1317
rect 12833 1292 12931 1294
rect 12958 1292 13126 1304
rect 13141 1294 13157 1308
rect 13192 1295 13214 1314
rect 13224 1308 13240 1309
rect 13223 1306 13240 1308
rect 13224 1301 13240 1306
rect 13214 1294 13220 1295
rect 13223 1294 13252 1301
rect 13141 1293 13252 1294
rect 13141 1292 13258 1293
rect 12817 1284 12868 1292
rect 12915 1284 12949 1292
rect 12817 1272 12842 1284
rect 12849 1272 12868 1284
rect 12922 1282 12949 1284
rect 12958 1282 13179 1292
rect 13214 1289 13220 1292
rect 12922 1278 13179 1282
rect 12817 1264 12868 1272
rect 12915 1264 13179 1278
rect 13223 1284 13258 1292
rect 12769 1216 12788 1250
rect 12833 1256 12862 1264
rect 12833 1250 12850 1256
rect 12833 1248 12867 1250
rect 12915 1248 12931 1264
rect 12932 1254 13140 1264
rect 13141 1254 13157 1264
rect 13205 1260 13220 1275
rect 13223 1272 13224 1284
rect 13231 1272 13258 1284
rect 13223 1264 13258 1272
rect 13223 1263 13252 1264
rect 12943 1250 13157 1254
rect 12958 1248 13157 1250
rect 13192 1250 13205 1260
rect 13223 1250 13240 1263
rect 13192 1248 13240 1250
rect 12834 1244 12867 1248
rect 12830 1242 12867 1244
rect 12830 1241 12897 1242
rect 12830 1236 12861 1241
rect 12867 1236 12897 1241
rect 12830 1232 12897 1236
rect 12803 1229 12897 1232
rect 12803 1222 12852 1229
rect 12803 1216 12833 1222
rect 12852 1217 12857 1222
rect 12769 1200 12849 1216
rect 12861 1208 12897 1229
rect 12958 1224 13147 1248
rect 13192 1247 13239 1248
rect 13205 1242 13239 1247
rect 12973 1221 13147 1224
rect 12966 1218 13147 1221
rect 13175 1241 13239 1242
rect 12769 1198 12788 1200
rect 12803 1198 12837 1200
rect 12769 1182 12849 1198
rect 12769 1176 12788 1182
rect 12485 1150 12588 1160
rect 12439 1148 12588 1150
rect 12609 1148 12644 1160
rect 12278 1146 12440 1148
rect 12290 1126 12309 1146
rect 12324 1144 12354 1146
rect 12173 1118 12214 1126
rect 12296 1122 12309 1126
rect 12361 1130 12440 1146
rect 12472 1146 12644 1148
rect 12472 1130 12551 1146
rect 12558 1144 12588 1146
rect 12136 1108 12165 1118
rect 12179 1108 12208 1118
rect 12223 1108 12253 1122
rect 12296 1108 12339 1122
rect 12361 1118 12551 1130
rect 12616 1126 12622 1146
rect 12346 1108 12376 1118
rect 12377 1108 12535 1118
rect 12539 1108 12569 1118
rect 12573 1108 12603 1122
rect 12631 1108 12644 1146
rect 12716 1160 12745 1176
rect 12759 1160 12788 1176
rect 12803 1166 12833 1182
rect 12861 1160 12867 1208
rect 12870 1202 12889 1208
rect 12904 1202 12934 1210
rect 12870 1194 12934 1202
rect 12870 1178 12950 1194
rect 12966 1187 13028 1218
rect 13044 1187 13106 1218
rect 13175 1216 13224 1241
rect 13239 1216 13269 1232
rect 13138 1202 13168 1210
rect 13175 1208 13285 1216
rect 13138 1194 13183 1202
rect 12870 1176 12889 1178
rect 12904 1176 12950 1178
rect 12870 1160 12950 1176
rect 12977 1174 13012 1187
rect 13053 1184 13090 1187
rect 13053 1182 13095 1184
rect 12982 1171 13012 1174
rect 12991 1167 12998 1171
rect 12998 1166 12999 1167
rect 12957 1160 12967 1166
rect 12716 1152 12751 1160
rect 12716 1126 12717 1152
rect 12724 1126 12751 1152
rect 12659 1108 12689 1122
rect 12716 1118 12751 1126
rect 12753 1152 12794 1160
rect 12753 1126 12768 1152
rect 12775 1126 12794 1152
rect 12858 1148 12889 1160
rect 12904 1148 13007 1160
rect 13019 1150 13045 1176
rect 13060 1171 13090 1182
rect 13122 1178 13184 1194
rect 13122 1176 13168 1178
rect 13122 1160 13184 1176
rect 13196 1160 13202 1208
rect 13205 1200 13285 1208
rect 13205 1198 13224 1200
rect 13239 1198 13273 1200
rect 13205 1182 13285 1198
rect 13205 1160 13224 1182
rect 13239 1166 13269 1182
rect 13297 1176 13303 1250
rect 13306 1176 13325 1320
rect 13340 1176 13346 1320
rect 13355 1250 13368 1320
rect 13420 1316 13442 1320
rect 13413 1294 13442 1308
rect 13495 1294 13511 1308
rect 13549 1304 13555 1306
rect 13562 1304 13670 1320
rect 13677 1304 13683 1306
rect 13691 1304 13706 1320
rect 13772 1314 13791 1317
rect 13413 1292 13511 1294
rect 13538 1292 13706 1304
rect 13721 1294 13737 1308
rect 13772 1295 13794 1314
rect 13804 1308 13820 1309
rect 13803 1306 13820 1308
rect 13804 1301 13820 1306
rect 13794 1294 13800 1295
rect 13803 1294 13832 1301
rect 13721 1293 13832 1294
rect 13721 1292 13838 1293
rect 13397 1284 13448 1292
rect 13495 1284 13529 1292
rect 13397 1272 13422 1284
rect 13429 1272 13448 1284
rect 13502 1282 13529 1284
rect 13538 1282 13759 1292
rect 13794 1289 13800 1292
rect 13502 1278 13759 1282
rect 13397 1264 13448 1272
rect 13495 1264 13759 1278
rect 13803 1284 13838 1292
rect 13349 1216 13368 1250
rect 13413 1256 13442 1264
rect 13413 1250 13430 1256
rect 13413 1248 13447 1250
rect 13495 1248 13511 1264
rect 13512 1254 13720 1264
rect 13721 1254 13737 1264
rect 13785 1260 13800 1275
rect 13803 1272 13804 1284
rect 13811 1272 13838 1284
rect 13803 1264 13838 1272
rect 13803 1263 13832 1264
rect 13523 1250 13737 1254
rect 13538 1248 13737 1250
rect 13772 1250 13785 1260
rect 13803 1250 13820 1263
rect 13772 1248 13820 1250
rect 13414 1244 13447 1248
rect 13410 1242 13447 1244
rect 13410 1241 13477 1242
rect 13410 1236 13441 1241
rect 13447 1236 13477 1241
rect 13410 1232 13477 1236
rect 13383 1229 13477 1232
rect 13383 1222 13432 1229
rect 13383 1216 13413 1222
rect 13432 1217 13437 1222
rect 13349 1200 13429 1216
rect 13441 1208 13477 1229
rect 13538 1224 13727 1248
rect 13772 1247 13819 1248
rect 13785 1242 13819 1247
rect 13553 1221 13727 1224
rect 13546 1218 13727 1221
rect 13755 1241 13819 1242
rect 13349 1198 13368 1200
rect 13383 1198 13417 1200
rect 13349 1182 13429 1198
rect 13349 1176 13368 1182
rect 13065 1150 13168 1160
rect 13019 1148 13168 1150
rect 13189 1148 13224 1160
rect 12858 1146 13020 1148
rect 12870 1126 12889 1146
rect 12904 1144 12934 1146
rect 12753 1118 12794 1126
rect 12876 1122 12889 1126
rect 12941 1130 13020 1146
rect 13052 1146 13224 1148
rect 13052 1130 13131 1146
rect 13138 1144 13168 1146
rect 12716 1108 12745 1118
rect 12759 1108 12788 1118
rect 12803 1108 12833 1122
rect 12876 1108 12919 1122
rect 12941 1118 13131 1130
rect 13196 1126 13202 1146
rect 12926 1108 12956 1118
rect 12957 1108 13115 1118
rect 13119 1108 13149 1118
rect 13153 1108 13183 1122
rect 13211 1108 13224 1146
rect 13296 1160 13325 1176
rect 13339 1160 13368 1176
rect 13383 1166 13413 1182
rect 13441 1160 13447 1208
rect 13450 1202 13469 1208
rect 13484 1202 13514 1210
rect 13450 1194 13514 1202
rect 13450 1178 13530 1194
rect 13546 1187 13608 1218
rect 13624 1187 13686 1218
rect 13755 1216 13804 1241
rect 13819 1216 13849 1232
rect 13718 1202 13748 1210
rect 13755 1208 13865 1216
rect 13718 1194 13763 1202
rect 13450 1176 13469 1178
rect 13484 1176 13530 1178
rect 13450 1160 13530 1176
rect 13557 1174 13592 1187
rect 13633 1184 13670 1187
rect 13633 1182 13675 1184
rect 13562 1171 13592 1174
rect 13571 1167 13578 1171
rect 13578 1166 13579 1167
rect 13537 1160 13547 1166
rect 13296 1152 13331 1160
rect 13296 1126 13297 1152
rect 13304 1126 13331 1152
rect 13239 1108 13269 1122
rect 13296 1118 13331 1126
rect 13333 1152 13374 1160
rect 13333 1126 13348 1152
rect 13355 1126 13374 1152
rect 13438 1148 13469 1160
rect 13484 1148 13587 1160
rect 13599 1150 13625 1176
rect 13640 1171 13670 1182
rect 13702 1178 13764 1194
rect 13702 1176 13748 1178
rect 13702 1160 13764 1176
rect 13776 1160 13782 1208
rect 13785 1200 13865 1208
rect 13785 1198 13804 1200
rect 13819 1198 13853 1200
rect 13785 1182 13865 1198
rect 13785 1160 13804 1182
rect 13819 1166 13849 1182
rect 13877 1176 13883 1250
rect 13886 1176 13905 1320
rect 13920 1176 13926 1320
rect 13935 1250 13948 1320
rect 14000 1316 14022 1320
rect 13993 1294 14022 1308
rect 14075 1294 14091 1308
rect 14129 1304 14135 1306
rect 14142 1304 14250 1320
rect 14257 1304 14263 1306
rect 14271 1304 14286 1320
rect 14352 1314 14371 1317
rect 13993 1292 14091 1294
rect 14118 1292 14286 1304
rect 14301 1294 14317 1308
rect 14352 1295 14374 1314
rect 14384 1308 14400 1309
rect 14383 1306 14400 1308
rect 14384 1301 14400 1306
rect 14374 1294 14380 1295
rect 14383 1294 14412 1301
rect 14301 1293 14412 1294
rect 14301 1292 14418 1293
rect 13977 1284 14028 1292
rect 14075 1284 14109 1292
rect 13977 1272 14002 1284
rect 14009 1272 14028 1284
rect 14082 1282 14109 1284
rect 14118 1282 14339 1292
rect 14374 1289 14380 1292
rect 14082 1278 14339 1282
rect 13977 1264 14028 1272
rect 14075 1264 14339 1278
rect 14383 1284 14418 1292
rect 13929 1216 13948 1250
rect 13993 1256 14022 1264
rect 13993 1250 14010 1256
rect 13993 1248 14027 1250
rect 14075 1248 14091 1264
rect 14092 1254 14300 1264
rect 14301 1254 14317 1264
rect 14365 1260 14380 1275
rect 14383 1272 14384 1284
rect 14391 1272 14418 1284
rect 14383 1264 14418 1272
rect 14383 1263 14412 1264
rect 14103 1250 14317 1254
rect 14118 1248 14317 1250
rect 14352 1250 14365 1260
rect 14383 1250 14400 1263
rect 14352 1248 14400 1250
rect 13994 1244 14027 1248
rect 13990 1242 14027 1244
rect 13990 1241 14057 1242
rect 13990 1236 14021 1241
rect 14027 1236 14057 1241
rect 13990 1232 14057 1236
rect 13963 1229 14057 1232
rect 13963 1222 14012 1229
rect 13963 1216 13993 1222
rect 14012 1217 14017 1222
rect 13929 1200 14009 1216
rect 14021 1208 14057 1229
rect 14118 1224 14307 1248
rect 14352 1247 14399 1248
rect 14365 1242 14399 1247
rect 14133 1221 14307 1224
rect 14126 1218 14307 1221
rect 14335 1241 14399 1242
rect 13929 1198 13948 1200
rect 13963 1198 13997 1200
rect 13929 1182 14009 1198
rect 13929 1176 13948 1182
rect 13645 1150 13748 1160
rect 13599 1148 13748 1150
rect 13769 1148 13804 1160
rect 13438 1146 13600 1148
rect 13450 1126 13469 1146
rect 13484 1144 13514 1146
rect 13333 1118 13374 1126
rect 13456 1122 13469 1126
rect 13521 1130 13600 1146
rect 13632 1146 13804 1148
rect 13632 1130 13711 1146
rect 13718 1144 13748 1146
rect 13296 1108 13325 1118
rect 13339 1108 13368 1118
rect 13383 1108 13413 1122
rect 13456 1108 13499 1122
rect 13521 1118 13711 1130
rect 13776 1126 13782 1146
rect 13506 1108 13536 1118
rect 13537 1108 13695 1118
rect 13699 1108 13729 1118
rect 13733 1108 13763 1122
rect 13791 1108 13804 1146
rect 13876 1160 13905 1176
rect 13919 1160 13948 1176
rect 13963 1166 13993 1182
rect 14021 1160 14027 1208
rect 14030 1202 14049 1208
rect 14064 1202 14094 1210
rect 14030 1194 14094 1202
rect 14030 1178 14110 1194
rect 14126 1187 14188 1218
rect 14204 1187 14266 1218
rect 14335 1216 14384 1241
rect 14399 1216 14429 1232
rect 14298 1202 14328 1210
rect 14335 1208 14445 1216
rect 14298 1194 14343 1202
rect 14030 1176 14049 1178
rect 14064 1176 14110 1178
rect 14030 1160 14110 1176
rect 14137 1174 14172 1187
rect 14213 1184 14250 1187
rect 14213 1182 14255 1184
rect 14142 1171 14172 1174
rect 14151 1167 14158 1171
rect 14158 1166 14159 1167
rect 14117 1160 14127 1166
rect 13876 1152 13911 1160
rect 13876 1126 13877 1152
rect 13884 1126 13911 1152
rect 13819 1108 13849 1122
rect 13876 1118 13911 1126
rect 13913 1152 13954 1160
rect 13913 1126 13928 1152
rect 13935 1126 13954 1152
rect 14018 1148 14049 1160
rect 14064 1148 14167 1160
rect 14179 1150 14205 1176
rect 14220 1171 14250 1182
rect 14282 1178 14344 1194
rect 14282 1176 14328 1178
rect 14282 1160 14344 1176
rect 14356 1160 14362 1208
rect 14365 1200 14445 1208
rect 14365 1198 14384 1200
rect 14399 1198 14433 1200
rect 14365 1182 14445 1198
rect 14365 1160 14384 1182
rect 14399 1166 14429 1182
rect 14457 1176 14463 1250
rect 14466 1176 14485 1320
rect 14500 1176 14506 1320
rect 14515 1250 14528 1320
rect 14580 1316 14602 1320
rect 14573 1294 14602 1308
rect 14655 1294 14671 1308
rect 14709 1304 14715 1306
rect 14722 1304 14830 1320
rect 14837 1304 14843 1306
rect 14851 1304 14866 1320
rect 14932 1314 14951 1317
rect 14573 1292 14671 1294
rect 14698 1292 14866 1304
rect 14881 1294 14897 1308
rect 14932 1295 14954 1314
rect 14964 1308 14980 1309
rect 14963 1306 14980 1308
rect 14964 1301 14980 1306
rect 14954 1294 14960 1295
rect 14963 1294 14992 1301
rect 14881 1293 14992 1294
rect 14881 1292 14998 1293
rect 14557 1284 14608 1292
rect 14655 1284 14689 1292
rect 14557 1272 14582 1284
rect 14589 1272 14608 1284
rect 14662 1282 14689 1284
rect 14698 1282 14919 1292
rect 14954 1289 14960 1292
rect 14662 1278 14919 1282
rect 14557 1264 14608 1272
rect 14655 1264 14919 1278
rect 14963 1284 14998 1292
rect 14509 1216 14528 1250
rect 14573 1256 14602 1264
rect 14573 1250 14590 1256
rect 14573 1248 14607 1250
rect 14655 1248 14671 1264
rect 14672 1254 14880 1264
rect 14881 1254 14897 1264
rect 14945 1260 14960 1275
rect 14963 1272 14964 1284
rect 14971 1272 14998 1284
rect 14963 1264 14998 1272
rect 14963 1263 14992 1264
rect 14683 1250 14897 1254
rect 14698 1248 14897 1250
rect 14932 1250 14945 1260
rect 14963 1250 14980 1263
rect 14932 1248 14980 1250
rect 14574 1244 14607 1248
rect 14570 1242 14607 1244
rect 14570 1241 14637 1242
rect 14570 1236 14601 1241
rect 14607 1236 14637 1241
rect 14570 1232 14637 1236
rect 14543 1229 14637 1232
rect 14543 1222 14592 1229
rect 14543 1216 14573 1222
rect 14592 1217 14597 1222
rect 14509 1200 14589 1216
rect 14601 1208 14637 1229
rect 14698 1224 14887 1248
rect 14932 1247 14979 1248
rect 14945 1242 14979 1247
rect 14713 1221 14887 1224
rect 14706 1218 14887 1221
rect 14915 1241 14979 1242
rect 14509 1198 14528 1200
rect 14543 1198 14577 1200
rect 14509 1182 14589 1198
rect 14509 1176 14528 1182
rect 14225 1150 14328 1160
rect 14179 1148 14328 1150
rect 14349 1148 14384 1160
rect 14018 1146 14180 1148
rect 14030 1126 14049 1146
rect 14064 1144 14094 1146
rect 13913 1118 13954 1126
rect 14036 1122 14049 1126
rect 14101 1130 14180 1146
rect 14212 1146 14384 1148
rect 14212 1130 14291 1146
rect 14298 1144 14328 1146
rect 13876 1108 13905 1118
rect 13919 1108 13948 1118
rect 13963 1108 13993 1122
rect 14036 1108 14079 1122
rect 14101 1118 14291 1130
rect 14356 1126 14362 1146
rect 14086 1108 14116 1118
rect 14117 1108 14275 1118
rect 14279 1108 14309 1118
rect 14313 1108 14343 1122
rect 14371 1108 14384 1146
rect 14456 1160 14485 1176
rect 14499 1160 14528 1176
rect 14543 1166 14573 1182
rect 14601 1160 14607 1208
rect 14610 1202 14629 1208
rect 14644 1202 14674 1210
rect 14610 1194 14674 1202
rect 14610 1178 14690 1194
rect 14706 1187 14768 1218
rect 14784 1187 14846 1218
rect 14915 1216 14964 1241
rect 14979 1216 15009 1232
rect 14878 1202 14908 1210
rect 14915 1208 15025 1216
rect 14878 1194 14923 1202
rect 14610 1176 14629 1178
rect 14644 1176 14690 1178
rect 14610 1160 14690 1176
rect 14717 1174 14752 1187
rect 14793 1184 14830 1187
rect 14793 1182 14835 1184
rect 14722 1171 14752 1174
rect 14731 1167 14738 1171
rect 14738 1166 14739 1167
rect 14697 1160 14707 1166
rect 14456 1152 14491 1160
rect 14456 1126 14457 1152
rect 14464 1126 14491 1152
rect 14399 1108 14429 1122
rect 14456 1118 14491 1126
rect 14493 1152 14534 1160
rect 14493 1126 14508 1152
rect 14515 1126 14534 1152
rect 14598 1148 14629 1160
rect 14644 1148 14747 1160
rect 14759 1150 14785 1176
rect 14800 1171 14830 1182
rect 14862 1178 14924 1194
rect 14862 1176 14908 1178
rect 14862 1160 14924 1176
rect 14936 1160 14942 1208
rect 14945 1200 15025 1208
rect 14945 1198 14964 1200
rect 14979 1198 15013 1200
rect 14945 1182 15025 1198
rect 14945 1160 14964 1182
rect 14979 1166 15009 1182
rect 15037 1176 15043 1250
rect 15046 1176 15065 1320
rect 15080 1176 15086 1320
rect 15095 1250 15108 1320
rect 15160 1316 15182 1320
rect 15153 1294 15182 1308
rect 15235 1294 15251 1308
rect 15289 1304 15295 1306
rect 15302 1304 15410 1320
rect 15417 1304 15423 1306
rect 15431 1304 15446 1320
rect 15512 1314 15531 1317
rect 15153 1292 15251 1294
rect 15278 1292 15446 1304
rect 15461 1294 15477 1308
rect 15512 1295 15534 1314
rect 15544 1308 15560 1309
rect 15543 1306 15560 1308
rect 15544 1301 15560 1306
rect 15534 1294 15540 1295
rect 15543 1294 15572 1301
rect 15461 1293 15572 1294
rect 15461 1292 15578 1293
rect 15137 1284 15188 1292
rect 15235 1284 15269 1292
rect 15137 1272 15162 1284
rect 15169 1272 15188 1284
rect 15242 1282 15269 1284
rect 15278 1282 15499 1292
rect 15534 1289 15540 1292
rect 15242 1278 15499 1282
rect 15137 1264 15188 1272
rect 15235 1264 15499 1278
rect 15543 1284 15578 1292
rect 15089 1216 15108 1250
rect 15153 1256 15182 1264
rect 15153 1250 15170 1256
rect 15153 1248 15187 1250
rect 15235 1248 15251 1264
rect 15252 1254 15460 1264
rect 15461 1254 15477 1264
rect 15525 1260 15540 1275
rect 15543 1272 15544 1284
rect 15551 1272 15578 1284
rect 15543 1264 15578 1272
rect 15543 1263 15572 1264
rect 15263 1250 15477 1254
rect 15278 1248 15477 1250
rect 15512 1250 15525 1260
rect 15543 1250 15560 1263
rect 15512 1248 15560 1250
rect 15154 1244 15187 1248
rect 15150 1242 15187 1244
rect 15150 1241 15217 1242
rect 15150 1236 15181 1241
rect 15187 1236 15217 1241
rect 15150 1232 15217 1236
rect 15123 1229 15217 1232
rect 15123 1222 15172 1229
rect 15123 1216 15153 1222
rect 15172 1217 15177 1222
rect 15089 1200 15169 1216
rect 15181 1208 15217 1229
rect 15278 1224 15467 1248
rect 15512 1247 15559 1248
rect 15525 1242 15559 1247
rect 15293 1221 15467 1224
rect 15286 1218 15467 1221
rect 15495 1241 15559 1242
rect 15089 1198 15108 1200
rect 15123 1198 15157 1200
rect 15089 1182 15169 1198
rect 15089 1176 15108 1182
rect 14805 1150 14908 1160
rect 14759 1148 14908 1150
rect 14929 1148 14964 1160
rect 14598 1146 14760 1148
rect 14610 1126 14629 1146
rect 14644 1144 14674 1146
rect 14493 1118 14534 1126
rect 14616 1122 14629 1126
rect 14681 1130 14760 1146
rect 14792 1146 14964 1148
rect 14792 1130 14871 1146
rect 14878 1144 14908 1146
rect 14456 1108 14485 1118
rect 14499 1108 14528 1118
rect 14543 1108 14573 1122
rect 14616 1108 14659 1122
rect 14681 1118 14871 1130
rect 14936 1126 14942 1146
rect 14666 1108 14696 1118
rect 14697 1108 14855 1118
rect 14859 1108 14889 1118
rect 14893 1108 14923 1122
rect 14951 1108 14964 1146
rect 15036 1160 15065 1176
rect 15079 1160 15108 1176
rect 15123 1166 15153 1182
rect 15181 1160 15187 1208
rect 15190 1202 15209 1208
rect 15224 1202 15254 1210
rect 15190 1194 15254 1202
rect 15190 1178 15270 1194
rect 15286 1187 15348 1218
rect 15364 1187 15426 1218
rect 15495 1216 15544 1241
rect 15559 1216 15589 1232
rect 15458 1202 15488 1210
rect 15495 1208 15605 1216
rect 15458 1194 15503 1202
rect 15190 1176 15209 1178
rect 15224 1176 15270 1178
rect 15190 1160 15270 1176
rect 15297 1174 15332 1187
rect 15373 1184 15410 1187
rect 15373 1182 15415 1184
rect 15302 1171 15332 1174
rect 15311 1167 15318 1171
rect 15318 1166 15319 1167
rect 15277 1160 15287 1166
rect 15036 1152 15071 1160
rect 15036 1126 15037 1152
rect 15044 1126 15071 1152
rect 14979 1108 15009 1122
rect 15036 1118 15071 1126
rect 15073 1152 15114 1160
rect 15073 1126 15088 1152
rect 15095 1126 15114 1152
rect 15178 1148 15209 1160
rect 15224 1148 15327 1160
rect 15339 1150 15365 1176
rect 15380 1171 15410 1182
rect 15442 1178 15504 1194
rect 15442 1176 15488 1178
rect 15442 1160 15504 1176
rect 15516 1160 15522 1208
rect 15525 1200 15605 1208
rect 15525 1198 15544 1200
rect 15559 1198 15593 1200
rect 15525 1182 15605 1198
rect 15525 1160 15544 1182
rect 15559 1166 15589 1182
rect 15617 1176 15623 1250
rect 15626 1176 15645 1320
rect 15660 1176 15666 1320
rect 15675 1250 15688 1320
rect 15740 1316 15762 1320
rect 15733 1294 15762 1308
rect 15815 1294 15831 1308
rect 15869 1304 15875 1306
rect 15882 1304 15990 1320
rect 15997 1304 16003 1306
rect 16011 1304 16026 1320
rect 16092 1314 16111 1317
rect 15733 1292 15831 1294
rect 15858 1292 16026 1304
rect 16041 1294 16057 1308
rect 16092 1295 16114 1314
rect 16124 1308 16140 1309
rect 16123 1306 16140 1308
rect 16124 1301 16140 1306
rect 16114 1294 16120 1295
rect 16123 1294 16152 1301
rect 16041 1293 16152 1294
rect 16041 1292 16158 1293
rect 15717 1284 15768 1292
rect 15815 1284 15849 1292
rect 15717 1272 15742 1284
rect 15749 1272 15768 1284
rect 15822 1282 15849 1284
rect 15858 1282 16079 1292
rect 16114 1289 16120 1292
rect 15822 1278 16079 1282
rect 15717 1264 15768 1272
rect 15815 1264 16079 1278
rect 16123 1284 16158 1292
rect 15669 1216 15688 1250
rect 15733 1256 15762 1264
rect 15733 1250 15750 1256
rect 15733 1248 15767 1250
rect 15815 1248 15831 1264
rect 15832 1254 16040 1264
rect 16041 1254 16057 1264
rect 16105 1260 16120 1275
rect 16123 1272 16124 1284
rect 16131 1272 16158 1284
rect 16123 1264 16158 1272
rect 16123 1263 16152 1264
rect 15843 1250 16057 1254
rect 15858 1248 16057 1250
rect 16092 1250 16105 1260
rect 16123 1250 16140 1263
rect 16092 1248 16140 1250
rect 15734 1244 15767 1248
rect 15730 1242 15767 1244
rect 15730 1241 15797 1242
rect 15730 1236 15761 1241
rect 15767 1236 15797 1241
rect 15730 1232 15797 1236
rect 15703 1229 15797 1232
rect 15703 1222 15752 1229
rect 15703 1216 15733 1222
rect 15752 1217 15757 1222
rect 15669 1200 15749 1216
rect 15761 1208 15797 1229
rect 15858 1224 16047 1248
rect 16092 1247 16139 1248
rect 16105 1242 16139 1247
rect 15873 1221 16047 1224
rect 15866 1218 16047 1221
rect 16075 1241 16139 1242
rect 15669 1198 15688 1200
rect 15703 1198 15737 1200
rect 15669 1182 15749 1198
rect 15669 1176 15688 1182
rect 15385 1150 15488 1160
rect 15339 1148 15488 1150
rect 15509 1148 15544 1160
rect 15178 1146 15340 1148
rect 15190 1126 15209 1146
rect 15224 1144 15254 1146
rect 15073 1118 15114 1126
rect 15196 1122 15209 1126
rect 15261 1130 15340 1146
rect 15372 1146 15544 1148
rect 15372 1130 15451 1146
rect 15458 1144 15488 1146
rect 15036 1108 15065 1118
rect 15079 1108 15108 1118
rect 15123 1108 15153 1122
rect 15196 1108 15239 1122
rect 15261 1118 15451 1130
rect 15516 1126 15522 1146
rect 15246 1108 15276 1118
rect 15277 1108 15435 1118
rect 15439 1108 15469 1118
rect 15473 1108 15503 1122
rect 15531 1108 15544 1146
rect 15616 1160 15645 1176
rect 15659 1160 15688 1176
rect 15703 1166 15733 1182
rect 15761 1160 15767 1208
rect 15770 1202 15789 1208
rect 15804 1202 15834 1210
rect 15770 1194 15834 1202
rect 15770 1178 15850 1194
rect 15866 1187 15928 1218
rect 15944 1187 16006 1218
rect 16075 1216 16124 1241
rect 16139 1216 16169 1232
rect 16038 1202 16068 1210
rect 16075 1208 16185 1216
rect 16038 1194 16083 1202
rect 15770 1176 15789 1178
rect 15804 1176 15850 1178
rect 15770 1160 15850 1176
rect 15877 1174 15912 1187
rect 15953 1184 15990 1187
rect 15953 1182 15995 1184
rect 15882 1171 15912 1174
rect 15891 1167 15898 1171
rect 15898 1166 15899 1167
rect 15857 1160 15867 1166
rect 15616 1152 15651 1160
rect 15616 1126 15617 1152
rect 15624 1126 15651 1152
rect 15559 1108 15589 1122
rect 15616 1118 15651 1126
rect 15653 1152 15694 1160
rect 15653 1126 15668 1152
rect 15675 1126 15694 1152
rect 15758 1148 15789 1160
rect 15804 1148 15907 1160
rect 15919 1150 15945 1176
rect 15960 1171 15990 1182
rect 16022 1178 16084 1194
rect 16022 1176 16068 1178
rect 16022 1160 16084 1176
rect 16096 1160 16102 1208
rect 16105 1200 16185 1208
rect 16105 1198 16124 1200
rect 16139 1198 16173 1200
rect 16105 1182 16185 1198
rect 16105 1160 16124 1182
rect 16139 1166 16169 1182
rect 16197 1176 16203 1250
rect 16206 1176 16225 1320
rect 16240 1176 16246 1320
rect 16255 1250 16268 1320
rect 16320 1316 16342 1320
rect 16313 1294 16342 1308
rect 16395 1294 16411 1308
rect 16449 1304 16455 1306
rect 16462 1304 16570 1320
rect 16577 1304 16583 1306
rect 16591 1304 16606 1320
rect 16672 1314 16691 1317
rect 16313 1292 16411 1294
rect 16438 1292 16606 1304
rect 16621 1294 16637 1308
rect 16672 1295 16694 1314
rect 16704 1308 16720 1309
rect 16703 1306 16720 1308
rect 16704 1301 16720 1306
rect 16694 1294 16700 1295
rect 16703 1294 16732 1301
rect 16621 1293 16732 1294
rect 16621 1292 16738 1293
rect 16297 1284 16348 1292
rect 16395 1284 16429 1292
rect 16297 1272 16322 1284
rect 16329 1272 16348 1284
rect 16402 1282 16429 1284
rect 16438 1282 16659 1292
rect 16694 1289 16700 1292
rect 16402 1278 16659 1282
rect 16297 1264 16348 1272
rect 16395 1264 16659 1278
rect 16703 1284 16738 1292
rect 16249 1216 16268 1250
rect 16313 1256 16342 1264
rect 16313 1250 16330 1256
rect 16313 1248 16347 1250
rect 16395 1248 16411 1264
rect 16412 1254 16620 1264
rect 16621 1254 16637 1264
rect 16685 1260 16700 1275
rect 16703 1272 16704 1284
rect 16711 1272 16738 1284
rect 16703 1264 16738 1272
rect 16703 1263 16732 1264
rect 16423 1250 16637 1254
rect 16438 1248 16637 1250
rect 16672 1250 16685 1260
rect 16703 1250 16720 1263
rect 16672 1248 16720 1250
rect 16314 1244 16347 1248
rect 16310 1242 16347 1244
rect 16310 1241 16377 1242
rect 16310 1236 16341 1241
rect 16347 1236 16377 1241
rect 16310 1232 16377 1236
rect 16283 1229 16377 1232
rect 16283 1222 16332 1229
rect 16283 1216 16313 1222
rect 16332 1217 16337 1222
rect 16249 1200 16329 1216
rect 16341 1208 16377 1229
rect 16438 1224 16627 1248
rect 16672 1247 16719 1248
rect 16685 1242 16719 1247
rect 16453 1221 16627 1224
rect 16446 1218 16627 1221
rect 16655 1241 16719 1242
rect 16249 1198 16268 1200
rect 16283 1198 16317 1200
rect 16249 1182 16329 1198
rect 16249 1176 16268 1182
rect 15965 1150 16068 1160
rect 15919 1148 16068 1150
rect 16089 1148 16124 1160
rect 15758 1146 15920 1148
rect 15770 1126 15789 1146
rect 15804 1144 15834 1146
rect 15653 1118 15694 1126
rect 15776 1122 15789 1126
rect 15841 1130 15920 1146
rect 15952 1146 16124 1148
rect 15952 1130 16031 1146
rect 16038 1144 16068 1146
rect 15616 1108 15645 1118
rect 15659 1108 15688 1118
rect 15703 1108 15733 1122
rect 15776 1108 15819 1122
rect 15841 1118 16031 1130
rect 16096 1126 16102 1146
rect 15826 1108 15856 1118
rect 15857 1108 16015 1118
rect 16019 1108 16049 1118
rect 16053 1108 16083 1122
rect 16111 1108 16124 1146
rect 16196 1160 16225 1176
rect 16239 1160 16268 1176
rect 16283 1166 16313 1182
rect 16341 1160 16347 1208
rect 16350 1202 16369 1208
rect 16384 1202 16414 1210
rect 16350 1194 16414 1202
rect 16350 1178 16430 1194
rect 16446 1187 16508 1218
rect 16524 1187 16586 1218
rect 16655 1216 16704 1241
rect 16719 1216 16749 1232
rect 16618 1202 16648 1210
rect 16655 1208 16765 1216
rect 16618 1194 16663 1202
rect 16350 1176 16369 1178
rect 16384 1176 16430 1178
rect 16350 1160 16430 1176
rect 16457 1174 16492 1187
rect 16533 1184 16570 1187
rect 16533 1182 16575 1184
rect 16462 1171 16492 1174
rect 16471 1167 16478 1171
rect 16478 1166 16479 1167
rect 16437 1160 16447 1166
rect 16196 1152 16231 1160
rect 16196 1126 16197 1152
rect 16204 1126 16231 1152
rect 16139 1108 16169 1122
rect 16196 1118 16231 1126
rect 16233 1152 16274 1160
rect 16233 1126 16248 1152
rect 16255 1126 16274 1152
rect 16338 1148 16369 1160
rect 16384 1148 16487 1160
rect 16499 1150 16525 1176
rect 16540 1171 16570 1182
rect 16602 1178 16664 1194
rect 16602 1176 16648 1178
rect 16602 1160 16664 1176
rect 16676 1160 16682 1208
rect 16685 1200 16765 1208
rect 16685 1198 16704 1200
rect 16719 1198 16753 1200
rect 16685 1182 16765 1198
rect 16685 1160 16704 1182
rect 16719 1166 16749 1182
rect 16777 1176 16783 1250
rect 16786 1176 16805 1320
rect 16820 1176 16826 1320
rect 16835 1250 16848 1320
rect 16900 1316 16922 1320
rect 16893 1294 16922 1308
rect 16975 1294 16991 1308
rect 17029 1304 17035 1306
rect 17042 1304 17150 1320
rect 17157 1304 17163 1306
rect 17171 1304 17186 1320
rect 17252 1314 17271 1317
rect 16893 1292 16991 1294
rect 17018 1292 17186 1304
rect 17201 1294 17217 1308
rect 17252 1295 17274 1314
rect 17284 1308 17300 1309
rect 17283 1306 17300 1308
rect 17284 1301 17300 1306
rect 17274 1294 17280 1295
rect 17283 1294 17312 1301
rect 17201 1293 17312 1294
rect 17201 1292 17318 1293
rect 16877 1284 16928 1292
rect 16975 1284 17009 1292
rect 16877 1272 16902 1284
rect 16909 1272 16928 1284
rect 16982 1282 17009 1284
rect 17018 1282 17239 1292
rect 17274 1289 17280 1292
rect 16982 1278 17239 1282
rect 16877 1264 16928 1272
rect 16975 1264 17239 1278
rect 17283 1284 17318 1292
rect 16829 1216 16848 1250
rect 16893 1256 16922 1264
rect 16893 1250 16910 1256
rect 16893 1248 16927 1250
rect 16975 1248 16991 1264
rect 16992 1254 17200 1264
rect 17201 1254 17217 1264
rect 17265 1260 17280 1275
rect 17283 1272 17284 1284
rect 17291 1272 17318 1284
rect 17283 1264 17318 1272
rect 17283 1263 17312 1264
rect 17003 1250 17217 1254
rect 17018 1248 17217 1250
rect 17252 1250 17265 1260
rect 17283 1250 17300 1263
rect 17252 1248 17300 1250
rect 16894 1244 16927 1248
rect 16890 1242 16927 1244
rect 16890 1241 16957 1242
rect 16890 1236 16921 1241
rect 16927 1236 16957 1241
rect 16890 1232 16957 1236
rect 16863 1229 16957 1232
rect 16863 1222 16912 1229
rect 16863 1216 16893 1222
rect 16912 1217 16917 1222
rect 16829 1200 16909 1216
rect 16921 1208 16957 1229
rect 17018 1224 17207 1248
rect 17252 1247 17299 1248
rect 17265 1242 17299 1247
rect 17033 1221 17207 1224
rect 17026 1218 17207 1221
rect 17235 1241 17299 1242
rect 16829 1198 16848 1200
rect 16863 1198 16897 1200
rect 16829 1182 16909 1198
rect 16829 1176 16848 1182
rect 16545 1150 16648 1160
rect 16499 1148 16648 1150
rect 16669 1148 16704 1160
rect 16338 1146 16500 1148
rect 16350 1126 16369 1146
rect 16384 1144 16414 1146
rect 16233 1118 16274 1126
rect 16356 1122 16369 1126
rect 16421 1130 16500 1146
rect 16532 1146 16704 1148
rect 16532 1130 16611 1146
rect 16618 1144 16648 1146
rect 16196 1108 16225 1118
rect 16239 1108 16268 1118
rect 16283 1108 16313 1122
rect 16356 1108 16399 1122
rect 16421 1118 16611 1130
rect 16676 1126 16682 1146
rect 16406 1108 16436 1118
rect 16437 1108 16595 1118
rect 16599 1108 16629 1118
rect 16633 1108 16663 1122
rect 16691 1108 16704 1146
rect 16776 1160 16805 1176
rect 16819 1160 16848 1176
rect 16863 1166 16893 1182
rect 16921 1160 16927 1208
rect 16930 1202 16949 1208
rect 16964 1202 16994 1210
rect 16930 1194 16994 1202
rect 16930 1178 17010 1194
rect 17026 1187 17088 1218
rect 17104 1187 17166 1218
rect 17235 1216 17284 1241
rect 17299 1216 17329 1232
rect 17198 1202 17228 1210
rect 17235 1208 17345 1216
rect 17198 1194 17243 1202
rect 16930 1176 16949 1178
rect 16964 1176 17010 1178
rect 16930 1160 17010 1176
rect 17037 1174 17072 1187
rect 17113 1184 17150 1187
rect 17113 1182 17155 1184
rect 17042 1171 17072 1174
rect 17051 1167 17058 1171
rect 17058 1166 17059 1167
rect 17017 1160 17027 1166
rect 16776 1152 16811 1160
rect 16776 1126 16777 1152
rect 16784 1126 16811 1152
rect 16719 1108 16749 1122
rect 16776 1118 16811 1126
rect 16813 1152 16854 1160
rect 16813 1126 16828 1152
rect 16835 1126 16854 1152
rect 16918 1148 16949 1160
rect 16964 1148 17067 1160
rect 17079 1150 17105 1176
rect 17120 1171 17150 1182
rect 17182 1178 17244 1194
rect 17182 1176 17228 1178
rect 17182 1160 17244 1176
rect 17256 1160 17262 1208
rect 17265 1200 17345 1208
rect 17265 1198 17284 1200
rect 17299 1198 17333 1200
rect 17265 1182 17345 1198
rect 17265 1160 17284 1182
rect 17299 1166 17329 1182
rect 17357 1176 17363 1250
rect 17366 1176 17385 1320
rect 17400 1176 17406 1320
rect 17415 1250 17428 1320
rect 17480 1316 17502 1320
rect 17473 1294 17502 1308
rect 17555 1294 17571 1308
rect 17609 1304 17615 1306
rect 17622 1304 17730 1320
rect 17737 1304 17743 1306
rect 17751 1304 17766 1320
rect 17832 1314 17851 1317
rect 17473 1292 17571 1294
rect 17598 1292 17766 1304
rect 17781 1294 17797 1308
rect 17832 1295 17854 1314
rect 17864 1308 17880 1309
rect 17863 1306 17880 1308
rect 17864 1301 17880 1306
rect 17854 1294 17860 1295
rect 17863 1294 17892 1301
rect 17781 1293 17892 1294
rect 17781 1292 17898 1293
rect 17457 1284 17508 1292
rect 17555 1284 17589 1292
rect 17457 1272 17482 1284
rect 17489 1272 17508 1284
rect 17562 1282 17589 1284
rect 17598 1282 17819 1292
rect 17854 1289 17860 1292
rect 17562 1278 17819 1282
rect 17457 1264 17508 1272
rect 17555 1264 17819 1278
rect 17863 1284 17898 1292
rect 17409 1216 17428 1250
rect 17473 1256 17502 1264
rect 17473 1250 17490 1256
rect 17473 1248 17507 1250
rect 17555 1248 17571 1264
rect 17572 1254 17780 1264
rect 17781 1254 17797 1264
rect 17845 1260 17860 1275
rect 17863 1272 17864 1284
rect 17871 1272 17898 1284
rect 17863 1264 17898 1272
rect 17863 1263 17892 1264
rect 17583 1250 17797 1254
rect 17598 1248 17797 1250
rect 17832 1250 17845 1260
rect 17863 1250 17880 1263
rect 17832 1248 17880 1250
rect 17474 1244 17507 1248
rect 17470 1242 17507 1244
rect 17470 1241 17537 1242
rect 17470 1236 17501 1241
rect 17507 1236 17537 1241
rect 17470 1232 17537 1236
rect 17443 1229 17537 1232
rect 17443 1222 17492 1229
rect 17443 1216 17473 1222
rect 17492 1217 17497 1222
rect 17409 1200 17489 1216
rect 17501 1208 17537 1229
rect 17598 1224 17787 1248
rect 17832 1247 17879 1248
rect 17845 1242 17879 1247
rect 17613 1221 17787 1224
rect 17606 1218 17787 1221
rect 17815 1241 17879 1242
rect 17409 1198 17428 1200
rect 17443 1198 17477 1200
rect 17409 1182 17489 1198
rect 17409 1176 17428 1182
rect 17125 1150 17228 1160
rect 17079 1148 17228 1150
rect 17249 1148 17284 1160
rect 16918 1146 17080 1148
rect 16930 1126 16949 1146
rect 16964 1144 16994 1146
rect 16813 1118 16854 1126
rect 16936 1122 16949 1126
rect 17001 1130 17080 1146
rect 17112 1146 17284 1148
rect 17112 1130 17191 1146
rect 17198 1144 17228 1146
rect 16776 1108 16805 1118
rect 16819 1108 16848 1118
rect 16863 1108 16893 1122
rect 16936 1108 16979 1122
rect 17001 1118 17191 1130
rect 17256 1126 17262 1146
rect 16986 1108 17016 1118
rect 17017 1108 17175 1118
rect 17179 1108 17209 1118
rect 17213 1108 17243 1122
rect 17271 1108 17284 1146
rect 17356 1160 17385 1176
rect 17399 1160 17428 1176
rect 17443 1166 17473 1182
rect 17501 1160 17507 1208
rect 17510 1202 17529 1208
rect 17544 1202 17574 1210
rect 17510 1194 17574 1202
rect 17510 1178 17590 1194
rect 17606 1187 17668 1218
rect 17684 1187 17746 1218
rect 17815 1216 17864 1241
rect 17879 1216 17909 1232
rect 17778 1202 17808 1210
rect 17815 1208 17925 1216
rect 17778 1194 17823 1202
rect 17510 1176 17529 1178
rect 17544 1176 17590 1178
rect 17510 1160 17590 1176
rect 17617 1174 17652 1187
rect 17693 1184 17730 1187
rect 17693 1182 17735 1184
rect 17622 1171 17652 1174
rect 17631 1167 17638 1171
rect 17638 1166 17639 1167
rect 17597 1160 17607 1166
rect 17356 1152 17391 1160
rect 17356 1126 17357 1152
rect 17364 1126 17391 1152
rect 17299 1108 17329 1122
rect 17356 1118 17391 1126
rect 17393 1152 17434 1160
rect 17393 1126 17408 1152
rect 17415 1126 17434 1152
rect 17498 1148 17529 1160
rect 17544 1148 17647 1160
rect 17659 1150 17685 1176
rect 17700 1171 17730 1182
rect 17762 1178 17824 1194
rect 17762 1176 17808 1178
rect 17762 1160 17824 1176
rect 17836 1160 17842 1208
rect 17845 1200 17925 1208
rect 17845 1198 17864 1200
rect 17879 1198 17913 1200
rect 17845 1182 17925 1198
rect 17845 1160 17864 1182
rect 17879 1166 17909 1182
rect 17937 1176 17943 1250
rect 17946 1176 17965 1320
rect 17980 1176 17986 1320
rect 17995 1250 18008 1320
rect 18060 1316 18082 1320
rect 18053 1294 18082 1308
rect 18135 1294 18151 1308
rect 18189 1304 18195 1306
rect 18202 1304 18310 1320
rect 18317 1304 18323 1306
rect 18331 1304 18346 1320
rect 18412 1314 18431 1317
rect 18053 1292 18151 1294
rect 18178 1292 18346 1304
rect 18361 1294 18377 1308
rect 18412 1295 18434 1314
rect 18444 1308 18460 1309
rect 18443 1306 18460 1308
rect 18444 1301 18460 1306
rect 18434 1294 18440 1295
rect 18443 1294 18472 1301
rect 18361 1293 18472 1294
rect 18361 1292 18478 1293
rect 18037 1284 18088 1292
rect 18135 1284 18169 1292
rect 18037 1272 18062 1284
rect 18069 1272 18088 1284
rect 18142 1282 18169 1284
rect 18178 1282 18399 1292
rect 18434 1289 18440 1292
rect 18142 1278 18399 1282
rect 18037 1264 18088 1272
rect 18135 1264 18399 1278
rect 18443 1284 18478 1292
rect 17989 1216 18008 1250
rect 18053 1256 18082 1264
rect 18053 1250 18070 1256
rect 18053 1248 18087 1250
rect 18135 1248 18151 1264
rect 18152 1254 18360 1264
rect 18361 1254 18377 1264
rect 18425 1260 18440 1275
rect 18443 1272 18444 1284
rect 18451 1272 18478 1284
rect 18443 1264 18478 1272
rect 18443 1263 18472 1264
rect 18163 1250 18377 1254
rect 18178 1248 18377 1250
rect 18412 1250 18425 1260
rect 18443 1250 18460 1263
rect 18412 1248 18460 1250
rect 18054 1244 18087 1248
rect 18050 1242 18087 1244
rect 18050 1241 18117 1242
rect 18050 1236 18081 1241
rect 18087 1236 18117 1241
rect 18050 1232 18117 1236
rect 18023 1229 18117 1232
rect 18023 1222 18072 1229
rect 18023 1216 18053 1222
rect 18072 1217 18077 1222
rect 17989 1200 18069 1216
rect 18081 1208 18117 1229
rect 18178 1224 18367 1248
rect 18412 1247 18459 1248
rect 18425 1242 18459 1247
rect 18193 1221 18367 1224
rect 18186 1218 18367 1221
rect 18395 1241 18459 1242
rect 17989 1198 18008 1200
rect 18023 1198 18057 1200
rect 17989 1182 18069 1198
rect 17989 1176 18008 1182
rect 17705 1150 17808 1160
rect 17659 1148 17808 1150
rect 17829 1148 17864 1160
rect 17498 1146 17660 1148
rect 17510 1126 17529 1146
rect 17544 1144 17574 1146
rect 17393 1118 17434 1126
rect 17516 1122 17529 1126
rect 17581 1130 17660 1146
rect 17692 1146 17864 1148
rect 17692 1130 17771 1146
rect 17778 1144 17808 1146
rect 17356 1108 17385 1118
rect 17399 1108 17428 1118
rect 17443 1108 17473 1122
rect 17516 1108 17559 1122
rect 17581 1118 17771 1130
rect 17836 1126 17842 1146
rect 17566 1108 17596 1118
rect 17597 1108 17755 1118
rect 17759 1108 17789 1118
rect 17793 1108 17823 1122
rect 17851 1108 17864 1146
rect 17936 1160 17965 1176
rect 17979 1160 18008 1176
rect 18023 1166 18053 1182
rect 18081 1160 18087 1208
rect 18090 1202 18109 1208
rect 18124 1202 18154 1210
rect 18090 1194 18154 1202
rect 18090 1178 18170 1194
rect 18186 1187 18248 1218
rect 18264 1187 18326 1218
rect 18395 1216 18444 1241
rect 18459 1216 18489 1232
rect 18358 1202 18388 1210
rect 18395 1208 18505 1216
rect 18358 1194 18403 1202
rect 18090 1176 18109 1178
rect 18124 1176 18170 1178
rect 18090 1160 18170 1176
rect 18197 1174 18232 1187
rect 18273 1184 18310 1187
rect 18273 1182 18315 1184
rect 18202 1171 18232 1174
rect 18211 1167 18218 1171
rect 18218 1166 18219 1167
rect 18177 1160 18187 1166
rect 17936 1152 17971 1160
rect 17936 1126 17937 1152
rect 17944 1126 17971 1152
rect 17879 1108 17909 1122
rect 17936 1118 17971 1126
rect 17973 1152 18014 1160
rect 17973 1126 17988 1152
rect 17995 1126 18014 1152
rect 18078 1148 18109 1160
rect 18124 1148 18227 1160
rect 18239 1150 18265 1176
rect 18280 1171 18310 1182
rect 18342 1178 18404 1194
rect 18342 1176 18388 1178
rect 18342 1160 18404 1176
rect 18416 1160 18422 1208
rect 18425 1200 18505 1208
rect 18425 1198 18444 1200
rect 18459 1198 18493 1200
rect 18425 1182 18505 1198
rect 18425 1160 18444 1182
rect 18459 1166 18489 1182
rect 18517 1176 18523 1250
rect 18532 1176 18545 1320
rect 18285 1150 18388 1160
rect 18239 1148 18388 1150
rect 18409 1148 18444 1160
rect 18078 1146 18240 1148
rect 18090 1126 18109 1146
rect 18124 1144 18154 1146
rect 17973 1118 18014 1126
rect 18096 1122 18109 1126
rect 18161 1130 18240 1146
rect 18272 1146 18444 1148
rect 18272 1130 18351 1146
rect 18358 1144 18388 1146
rect 17936 1108 17965 1118
rect 17979 1108 18008 1118
rect 18023 1108 18053 1122
rect 18096 1108 18139 1122
rect 18161 1118 18351 1130
rect 18416 1126 18422 1146
rect 18146 1108 18176 1118
rect 18177 1108 18335 1118
rect 18339 1108 18369 1118
rect 18373 1108 18403 1122
rect 18431 1108 18444 1146
rect 18516 1160 18545 1176
rect 18516 1152 18551 1160
rect 18516 1126 18517 1152
rect 18524 1126 18551 1152
rect 18459 1108 18489 1122
rect 18516 1118 18551 1126
rect 18516 1108 18545 1118
rect -1 1102 18545 1108
rect 0 1094 18545 1102
rect 15 1064 28 1094
rect 43 1080 73 1094
rect 116 1080 159 1094
rect 166 1080 386 1094
rect 393 1080 423 1094
rect 83 1066 98 1078
rect 117 1066 130 1080
rect 198 1076 351 1080
rect 80 1064 102 1066
rect 180 1064 372 1076
rect 451 1064 464 1094
rect 479 1080 509 1094
rect 546 1064 565 1094
rect 580 1064 586 1094
rect 595 1064 608 1094
rect 623 1080 653 1094
rect 696 1080 739 1094
rect 746 1080 966 1094
rect 973 1080 1003 1094
rect 663 1066 678 1078
rect 697 1066 710 1080
rect 778 1076 931 1080
rect 660 1064 682 1066
rect 760 1064 952 1076
rect 1031 1064 1044 1094
rect 1059 1080 1089 1094
rect 1126 1064 1145 1094
rect 1160 1064 1166 1094
rect 1175 1064 1188 1094
rect 1203 1080 1233 1094
rect 1276 1080 1319 1094
rect 1326 1080 1546 1094
rect 1553 1080 1583 1094
rect 1243 1066 1258 1078
rect 1277 1066 1290 1080
rect 1358 1076 1511 1080
rect 1240 1064 1262 1066
rect 1340 1064 1532 1076
rect 1611 1064 1624 1094
rect 1639 1080 1669 1094
rect 1706 1064 1725 1094
rect 1740 1064 1746 1094
rect 1755 1064 1768 1094
rect 1783 1080 1813 1094
rect 1856 1080 1899 1094
rect 1906 1080 2126 1094
rect 2133 1080 2163 1094
rect 1823 1066 1838 1078
rect 1857 1066 1870 1080
rect 1938 1076 2091 1080
rect 1820 1064 1842 1066
rect 1920 1064 2112 1076
rect 2191 1064 2204 1094
rect 2219 1080 2249 1094
rect 2286 1064 2305 1094
rect 2320 1064 2326 1094
rect 2335 1064 2348 1094
rect 2363 1080 2393 1094
rect 2436 1080 2479 1094
rect 2486 1080 2706 1094
rect 2713 1080 2743 1094
rect 2403 1066 2418 1078
rect 2437 1066 2450 1080
rect 2518 1076 2671 1080
rect 2400 1064 2422 1066
rect 2500 1064 2692 1076
rect 2771 1064 2784 1094
rect 2799 1080 2829 1094
rect 2866 1064 2885 1094
rect 2900 1064 2906 1094
rect 2915 1064 2928 1094
rect 2943 1080 2973 1094
rect 3016 1080 3059 1094
rect 3066 1080 3286 1094
rect 3293 1080 3323 1094
rect 2983 1066 2998 1078
rect 3017 1066 3030 1080
rect 3098 1076 3251 1080
rect 2980 1064 3002 1066
rect 3080 1064 3272 1076
rect 3351 1064 3364 1094
rect 3379 1080 3409 1094
rect 3446 1064 3465 1094
rect 3480 1064 3486 1094
rect 3495 1064 3508 1094
rect 3523 1080 3553 1094
rect 3596 1080 3639 1094
rect 3646 1080 3866 1094
rect 3873 1080 3903 1094
rect 3563 1066 3578 1078
rect 3597 1066 3610 1080
rect 3678 1076 3831 1080
rect 3560 1064 3582 1066
rect 3660 1064 3852 1076
rect 3931 1064 3944 1094
rect 3959 1080 3989 1094
rect 4026 1064 4045 1094
rect 4060 1064 4066 1094
rect 4075 1064 4088 1094
rect 4103 1080 4133 1094
rect 4176 1080 4219 1094
rect 4226 1080 4446 1094
rect 4453 1080 4483 1094
rect 4143 1066 4158 1078
rect 4177 1066 4190 1080
rect 4258 1076 4411 1080
rect 4140 1064 4162 1066
rect 4240 1064 4432 1076
rect 4511 1064 4524 1094
rect 4539 1080 4569 1094
rect 4606 1064 4625 1094
rect 4640 1064 4646 1094
rect 4655 1064 4668 1094
rect 4683 1080 4713 1094
rect 4756 1080 4799 1094
rect 4806 1080 5026 1094
rect 5033 1080 5063 1094
rect 4723 1066 4738 1078
rect 4757 1066 4770 1080
rect 4838 1076 4991 1080
rect 4720 1064 4742 1066
rect 4820 1064 5012 1076
rect 5091 1064 5104 1094
rect 5119 1080 5149 1094
rect 5186 1064 5205 1094
rect 5220 1064 5226 1094
rect 5235 1064 5248 1094
rect 5263 1080 5293 1094
rect 5336 1080 5379 1094
rect 5386 1080 5606 1094
rect 5613 1080 5643 1094
rect 5303 1066 5318 1078
rect 5337 1066 5350 1080
rect 5418 1076 5571 1080
rect 5300 1064 5322 1066
rect 5400 1064 5592 1076
rect 5671 1064 5684 1094
rect 5699 1080 5729 1094
rect 5766 1064 5785 1094
rect 5800 1064 5806 1094
rect 5815 1064 5828 1094
rect 5843 1080 5873 1094
rect 5916 1080 5959 1094
rect 5966 1080 6186 1094
rect 6193 1080 6223 1094
rect 5883 1066 5898 1078
rect 5917 1066 5930 1080
rect 5998 1076 6151 1080
rect 5880 1064 5902 1066
rect 5980 1064 6172 1076
rect 6251 1064 6264 1094
rect 6279 1080 6309 1094
rect 6346 1064 6365 1094
rect 6380 1064 6386 1094
rect 6395 1064 6408 1094
rect 6423 1080 6453 1094
rect 6496 1080 6539 1094
rect 6546 1080 6766 1094
rect 6773 1080 6803 1094
rect 6463 1066 6478 1078
rect 6497 1066 6510 1080
rect 6578 1076 6731 1080
rect 6460 1064 6482 1066
rect 6560 1064 6752 1076
rect 6831 1064 6844 1094
rect 6859 1080 6889 1094
rect 6926 1064 6945 1094
rect 6960 1064 6966 1094
rect 6975 1064 6988 1094
rect 7003 1080 7033 1094
rect 7076 1080 7119 1094
rect 7126 1080 7346 1094
rect 7353 1080 7383 1094
rect 7043 1066 7058 1078
rect 7077 1066 7090 1080
rect 7158 1076 7311 1080
rect 7040 1064 7062 1066
rect 7140 1064 7332 1076
rect 7411 1064 7424 1094
rect 7439 1080 7469 1094
rect 7506 1064 7525 1094
rect 7540 1064 7546 1094
rect 7555 1064 7568 1094
rect 7583 1080 7613 1094
rect 7656 1080 7699 1094
rect 7706 1080 7926 1094
rect 7933 1080 7963 1094
rect 7623 1066 7638 1078
rect 7657 1066 7670 1080
rect 7738 1076 7891 1080
rect 7620 1064 7642 1066
rect 7720 1064 7912 1076
rect 7991 1064 8004 1094
rect 8019 1080 8049 1094
rect 8086 1064 8105 1094
rect 8120 1064 8126 1094
rect 8135 1064 8148 1094
rect 8163 1080 8193 1094
rect 8236 1080 8279 1094
rect 8286 1080 8506 1094
rect 8513 1080 8543 1094
rect 8203 1066 8218 1078
rect 8237 1066 8250 1080
rect 8318 1076 8471 1080
rect 8200 1064 8222 1066
rect 8300 1064 8492 1076
rect 8571 1064 8584 1094
rect 8599 1080 8629 1094
rect 8666 1064 8685 1094
rect 8700 1064 8706 1094
rect 8715 1064 8728 1094
rect 8743 1080 8773 1094
rect 8816 1080 8859 1094
rect 8866 1080 9086 1094
rect 9093 1080 9123 1094
rect 8783 1066 8798 1078
rect 8817 1066 8830 1080
rect 8898 1076 9051 1080
rect 8780 1064 8802 1066
rect 8880 1064 9072 1076
rect 9151 1064 9164 1094
rect 9179 1080 9209 1094
rect 9246 1064 9265 1094
rect 9280 1064 9286 1094
rect 9295 1064 9308 1094
rect 9323 1080 9353 1094
rect 9396 1080 9439 1094
rect 9446 1080 9666 1094
rect 9673 1080 9703 1094
rect 9363 1066 9378 1078
rect 9397 1066 9410 1080
rect 9478 1076 9631 1080
rect 9360 1064 9382 1066
rect 9460 1064 9652 1076
rect 9731 1064 9744 1094
rect 9759 1080 9789 1094
rect 9826 1064 9845 1094
rect 9860 1064 9866 1094
rect 9875 1064 9888 1094
rect 9903 1080 9933 1094
rect 9976 1080 10019 1094
rect 10026 1080 10246 1094
rect 10253 1080 10283 1094
rect 9943 1066 9958 1078
rect 9977 1066 9990 1080
rect 10058 1076 10211 1080
rect 9940 1064 9962 1066
rect 10040 1064 10232 1076
rect 10311 1064 10324 1094
rect 10339 1080 10369 1094
rect 10406 1064 10425 1094
rect 10440 1064 10446 1094
rect 10455 1064 10468 1094
rect 10483 1080 10513 1094
rect 10556 1080 10599 1094
rect 10606 1080 10826 1094
rect 10833 1080 10863 1094
rect 10523 1066 10538 1078
rect 10557 1066 10570 1080
rect 10638 1076 10791 1080
rect 10520 1064 10542 1066
rect 10620 1064 10812 1076
rect 10891 1064 10904 1094
rect 10919 1080 10949 1094
rect 10986 1064 11005 1094
rect 11020 1064 11026 1094
rect 11035 1064 11048 1094
rect 11063 1080 11093 1094
rect 11136 1080 11179 1094
rect 11186 1080 11406 1094
rect 11413 1080 11443 1094
rect 11103 1066 11118 1078
rect 11137 1066 11150 1080
rect 11218 1076 11371 1080
rect 11100 1064 11122 1066
rect 11200 1064 11392 1076
rect 11471 1064 11484 1094
rect 11499 1080 11529 1094
rect 11566 1064 11585 1094
rect 11600 1064 11606 1094
rect 11615 1064 11628 1094
rect 11643 1080 11673 1094
rect 11716 1080 11759 1094
rect 11766 1080 11986 1094
rect 11993 1080 12023 1094
rect 11683 1066 11698 1078
rect 11717 1066 11730 1080
rect 11798 1076 11951 1080
rect 11680 1064 11702 1066
rect 11780 1064 11972 1076
rect 12051 1064 12064 1094
rect 12079 1080 12109 1094
rect 12146 1064 12165 1094
rect 12180 1064 12186 1094
rect 12195 1064 12208 1094
rect 12223 1080 12253 1094
rect 12296 1080 12339 1094
rect 12346 1080 12566 1094
rect 12573 1080 12603 1094
rect 12263 1066 12278 1078
rect 12297 1066 12310 1080
rect 12378 1076 12531 1080
rect 12260 1064 12282 1066
rect 12360 1064 12552 1076
rect 12631 1064 12644 1094
rect 12659 1080 12689 1094
rect 12726 1064 12745 1094
rect 12760 1064 12766 1094
rect 12775 1064 12788 1094
rect 12803 1080 12833 1094
rect 12876 1080 12919 1094
rect 12926 1080 13146 1094
rect 13153 1080 13183 1094
rect 12843 1066 12858 1078
rect 12877 1066 12890 1080
rect 12958 1076 13111 1080
rect 12840 1064 12862 1066
rect 12940 1064 13132 1076
rect 13211 1064 13224 1094
rect 13239 1080 13269 1094
rect 13306 1064 13325 1094
rect 13340 1064 13346 1094
rect 13355 1064 13368 1094
rect 13383 1080 13413 1094
rect 13456 1080 13499 1094
rect 13506 1080 13726 1094
rect 13733 1080 13763 1094
rect 13423 1066 13438 1078
rect 13457 1066 13470 1080
rect 13538 1076 13691 1080
rect 13420 1064 13442 1066
rect 13520 1064 13712 1076
rect 13791 1064 13804 1094
rect 13819 1080 13849 1094
rect 13886 1064 13905 1094
rect 13920 1064 13926 1094
rect 13935 1064 13948 1094
rect 13963 1080 13993 1094
rect 14036 1080 14079 1094
rect 14086 1080 14306 1094
rect 14313 1080 14343 1094
rect 14003 1066 14018 1078
rect 14037 1066 14050 1080
rect 14118 1076 14271 1080
rect 14000 1064 14022 1066
rect 14100 1064 14292 1076
rect 14371 1064 14384 1094
rect 14399 1080 14429 1094
rect 14466 1064 14485 1094
rect 14500 1064 14506 1094
rect 14515 1064 14528 1094
rect 14543 1080 14573 1094
rect 14616 1080 14659 1094
rect 14666 1080 14886 1094
rect 14893 1080 14923 1094
rect 14583 1066 14598 1078
rect 14617 1066 14630 1080
rect 14698 1076 14851 1080
rect 14580 1064 14602 1066
rect 14680 1064 14872 1076
rect 14951 1064 14964 1094
rect 14979 1080 15009 1094
rect 15046 1064 15065 1094
rect 15080 1064 15086 1094
rect 15095 1064 15108 1094
rect 15123 1080 15153 1094
rect 15196 1080 15239 1094
rect 15246 1080 15466 1094
rect 15473 1080 15503 1094
rect 15163 1066 15178 1078
rect 15197 1066 15210 1080
rect 15278 1076 15431 1080
rect 15160 1064 15182 1066
rect 15260 1064 15452 1076
rect 15531 1064 15544 1094
rect 15559 1080 15589 1094
rect 15626 1064 15645 1094
rect 15660 1064 15666 1094
rect 15675 1064 15688 1094
rect 15703 1080 15733 1094
rect 15776 1080 15819 1094
rect 15826 1080 16046 1094
rect 16053 1080 16083 1094
rect 15743 1066 15758 1078
rect 15777 1066 15790 1080
rect 15858 1076 16011 1080
rect 15740 1064 15762 1066
rect 15840 1064 16032 1076
rect 16111 1064 16124 1094
rect 16139 1080 16169 1094
rect 16206 1064 16225 1094
rect 16240 1064 16246 1094
rect 16255 1064 16268 1094
rect 16283 1080 16313 1094
rect 16356 1080 16399 1094
rect 16406 1080 16626 1094
rect 16633 1080 16663 1094
rect 16323 1066 16338 1078
rect 16357 1066 16370 1080
rect 16438 1076 16591 1080
rect 16320 1064 16342 1066
rect 16420 1064 16612 1076
rect 16691 1064 16704 1094
rect 16719 1080 16749 1094
rect 16786 1064 16805 1094
rect 16820 1064 16826 1094
rect 16835 1064 16848 1094
rect 16863 1080 16893 1094
rect 16936 1080 16979 1094
rect 16986 1080 17206 1094
rect 17213 1080 17243 1094
rect 16903 1066 16918 1078
rect 16937 1066 16950 1080
rect 17018 1076 17171 1080
rect 16900 1064 16922 1066
rect 17000 1064 17192 1076
rect 17271 1064 17284 1094
rect 17299 1080 17329 1094
rect 17366 1064 17385 1094
rect 17400 1064 17406 1094
rect 17415 1064 17428 1094
rect 17443 1080 17473 1094
rect 17516 1080 17559 1094
rect 17566 1080 17786 1094
rect 17793 1080 17823 1094
rect 17483 1066 17498 1078
rect 17517 1066 17530 1080
rect 17598 1076 17751 1080
rect 17480 1064 17502 1066
rect 17580 1064 17772 1076
rect 17851 1064 17864 1094
rect 17879 1080 17909 1094
rect 17946 1064 17965 1094
rect 17980 1064 17986 1094
rect 17995 1064 18008 1094
rect 18023 1080 18053 1094
rect 18096 1080 18139 1094
rect 18146 1080 18366 1094
rect 18373 1080 18403 1094
rect 18063 1066 18078 1078
rect 18097 1066 18110 1080
rect 18178 1076 18331 1080
rect 18060 1064 18082 1066
rect 18160 1064 18352 1076
rect 18431 1064 18444 1094
rect 18459 1080 18489 1094
rect 18532 1064 18545 1094
rect 0 1050 18545 1064
rect 15 980 28 1050
rect 80 1046 102 1050
rect 73 1024 102 1038
rect 155 1024 171 1038
rect 209 1034 215 1036
rect 222 1034 330 1050
rect 337 1034 343 1036
rect 351 1034 366 1050
rect 432 1044 451 1047
rect 73 1022 171 1024
rect 198 1022 366 1034
rect 381 1024 397 1038
rect 432 1025 454 1044
rect 464 1038 480 1039
rect 463 1036 480 1038
rect 464 1031 480 1036
rect 454 1024 460 1025
rect 463 1024 492 1031
rect 381 1023 492 1024
rect 381 1022 498 1023
rect 57 1014 108 1022
rect 155 1014 189 1022
rect 57 1002 82 1014
rect 89 1002 108 1014
rect 162 1012 189 1014
rect 198 1012 419 1022
rect 454 1019 460 1022
rect 162 1008 419 1012
rect 57 994 108 1002
rect 155 994 419 1008
rect 463 1014 498 1022
rect 9 946 28 980
rect 73 986 102 994
rect 73 980 90 986
rect 73 978 107 980
rect 155 978 171 994
rect 172 984 380 994
rect 381 984 397 994
rect 445 990 460 1005
rect 463 1002 464 1014
rect 471 1002 498 1014
rect 463 994 498 1002
rect 463 993 492 994
rect 183 980 397 984
rect 198 978 397 980
rect 432 980 445 990
rect 463 980 480 993
rect 432 978 480 980
rect 74 974 107 978
rect 70 972 107 974
rect 70 971 137 972
rect 70 966 101 971
rect 107 966 137 971
rect 70 962 137 966
rect 43 959 137 962
rect 43 952 92 959
rect 43 946 73 952
rect 92 947 97 952
rect 9 930 89 946
rect 101 938 137 959
rect 198 954 387 978
rect 432 977 479 978
rect 445 972 479 977
rect 213 951 387 954
rect 206 948 387 951
rect 415 971 479 972
rect 9 928 28 930
rect 43 928 77 930
rect 9 912 89 928
rect 9 906 28 912
rect -1 890 28 906
rect 43 896 73 912
rect 101 890 107 938
rect 110 932 129 938
rect 144 932 174 940
rect 110 924 174 932
rect 110 908 190 924
rect 206 917 268 948
rect 284 917 346 948
rect 415 946 464 971
rect 479 946 509 962
rect 378 932 408 940
rect 415 938 525 946
rect 378 924 423 932
rect 110 906 129 908
rect 144 906 190 908
rect 110 890 190 906
rect 217 904 252 917
rect 293 914 330 917
rect 293 912 335 914
rect 222 901 252 904
rect 231 897 238 901
rect 238 896 239 897
rect 197 890 207 896
rect -7 882 34 890
rect -7 856 8 882
rect 15 856 34 882
rect 98 878 129 890
rect 144 878 247 890
rect 259 880 285 906
rect 300 901 330 912
rect 362 908 424 924
rect 362 906 408 908
rect 362 890 424 906
rect 436 890 442 938
rect 445 930 525 938
rect 445 928 464 930
rect 479 928 513 930
rect 445 912 525 928
rect 445 890 464 912
rect 479 896 509 912
rect 537 906 543 980
rect 546 906 565 1050
rect 580 906 586 1050
rect 595 980 608 1050
rect 660 1046 682 1050
rect 653 1024 682 1038
rect 735 1024 751 1038
rect 789 1034 795 1036
rect 802 1034 910 1050
rect 917 1034 923 1036
rect 931 1034 946 1050
rect 1012 1044 1031 1047
rect 653 1022 751 1024
rect 778 1022 946 1034
rect 961 1024 977 1038
rect 1012 1025 1034 1044
rect 1044 1038 1060 1039
rect 1043 1036 1060 1038
rect 1044 1031 1060 1036
rect 1034 1024 1040 1025
rect 1043 1024 1072 1031
rect 961 1023 1072 1024
rect 961 1022 1078 1023
rect 637 1014 688 1022
rect 735 1014 769 1022
rect 637 1002 662 1014
rect 669 1002 688 1014
rect 742 1012 769 1014
rect 778 1012 999 1022
rect 1034 1019 1040 1022
rect 742 1008 999 1012
rect 637 994 688 1002
rect 735 994 999 1008
rect 1043 1014 1078 1022
rect 589 946 608 980
rect 653 986 682 994
rect 653 980 670 986
rect 653 978 687 980
rect 735 978 751 994
rect 752 984 960 994
rect 961 984 977 994
rect 1025 990 1040 1005
rect 1043 1002 1044 1014
rect 1051 1002 1078 1014
rect 1043 994 1078 1002
rect 1043 993 1072 994
rect 763 980 977 984
rect 778 978 977 980
rect 1012 980 1025 990
rect 1043 980 1060 993
rect 1012 978 1060 980
rect 654 974 687 978
rect 650 972 687 974
rect 650 971 717 972
rect 650 966 681 971
rect 687 966 717 971
rect 650 962 717 966
rect 623 959 717 962
rect 623 952 672 959
rect 623 946 653 952
rect 672 947 677 952
rect 589 930 669 946
rect 681 938 717 959
rect 778 954 967 978
rect 1012 977 1059 978
rect 1025 972 1059 977
rect 793 951 967 954
rect 786 948 967 951
rect 995 971 1059 972
rect 589 928 608 930
rect 623 928 657 930
rect 589 912 669 928
rect 589 906 608 912
rect 305 880 408 890
rect 259 878 408 880
rect 429 878 464 890
rect 98 876 260 878
rect 110 856 129 876
rect 144 874 174 876
rect -7 848 34 856
rect 116 852 129 856
rect 181 860 260 876
rect 292 876 464 878
rect 292 860 371 876
rect 378 874 408 876
rect -1 838 28 848
rect 43 838 73 852
rect 116 838 159 852
rect 181 848 371 860
rect 436 856 442 876
rect 166 838 196 848
rect 197 838 355 848
rect 359 838 389 848
rect 393 838 423 852
rect 451 838 464 876
rect 536 890 565 906
rect 579 890 608 906
rect 623 896 653 912
rect 681 890 687 938
rect 690 932 709 938
rect 724 932 754 940
rect 690 924 754 932
rect 690 908 770 924
rect 786 917 848 948
rect 864 917 926 948
rect 995 946 1044 971
rect 1059 946 1089 962
rect 958 932 988 940
rect 995 938 1105 946
rect 958 924 1003 932
rect 690 906 709 908
rect 724 906 770 908
rect 690 890 770 906
rect 797 904 832 917
rect 873 914 910 917
rect 873 912 915 914
rect 802 901 832 904
rect 811 897 818 901
rect 818 896 819 897
rect 777 890 787 896
rect 536 882 571 890
rect 536 856 537 882
rect 544 856 571 882
rect 479 838 509 852
rect 536 848 571 856
rect 573 882 614 890
rect 573 856 588 882
rect 595 856 614 882
rect 678 878 709 890
rect 724 878 827 890
rect 839 880 865 906
rect 880 901 910 912
rect 942 908 1004 924
rect 942 906 988 908
rect 942 890 1004 906
rect 1016 890 1022 938
rect 1025 930 1105 938
rect 1025 928 1044 930
rect 1059 928 1093 930
rect 1025 912 1105 928
rect 1025 890 1044 912
rect 1059 896 1089 912
rect 1117 906 1123 980
rect 1126 906 1145 1050
rect 1160 906 1166 1050
rect 1175 980 1188 1050
rect 1240 1046 1262 1050
rect 1233 1024 1262 1038
rect 1315 1024 1331 1038
rect 1369 1034 1375 1036
rect 1382 1034 1490 1050
rect 1497 1034 1503 1036
rect 1511 1034 1526 1050
rect 1592 1044 1611 1047
rect 1233 1022 1331 1024
rect 1358 1022 1526 1034
rect 1541 1024 1557 1038
rect 1592 1025 1614 1044
rect 1624 1038 1640 1039
rect 1623 1036 1640 1038
rect 1624 1031 1640 1036
rect 1614 1024 1620 1025
rect 1623 1024 1652 1031
rect 1541 1023 1652 1024
rect 1541 1022 1658 1023
rect 1217 1014 1268 1022
rect 1315 1014 1349 1022
rect 1217 1002 1242 1014
rect 1249 1002 1268 1014
rect 1322 1012 1349 1014
rect 1358 1012 1579 1022
rect 1614 1019 1620 1022
rect 1322 1008 1579 1012
rect 1217 994 1268 1002
rect 1315 994 1579 1008
rect 1623 1014 1658 1022
rect 1169 946 1188 980
rect 1233 986 1262 994
rect 1233 980 1250 986
rect 1233 978 1267 980
rect 1315 978 1331 994
rect 1332 984 1540 994
rect 1541 984 1557 994
rect 1605 990 1620 1005
rect 1623 1002 1624 1014
rect 1631 1002 1658 1014
rect 1623 994 1658 1002
rect 1623 993 1652 994
rect 1343 980 1557 984
rect 1358 978 1557 980
rect 1592 980 1605 990
rect 1623 980 1640 993
rect 1592 978 1640 980
rect 1234 974 1267 978
rect 1230 972 1267 974
rect 1230 971 1297 972
rect 1230 966 1261 971
rect 1267 966 1297 971
rect 1230 962 1297 966
rect 1203 959 1297 962
rect 1203 952 1252 959
rect 1203 946 1233 952
rect 1252 947 1257 952
rect 1169 930 1249 946
rect 1261 938 1297 959
rect 1358 954 1547 978
rect 1592 977 1639 978
rect 1605 972 1639 977
rect 1373 951 1547 954
rect 1366 948 1547 951
rect 1575 971 1639 972
rect 1169 928 1188 930
rect 1203 928 1237 930
rect 1169 912 1249 928
rect 1169 906 1188 912
rect 885 880 988 890
rect 839 878 988 880
rect 1009 878 1044 890
rect 678 876 840 878
rect 690 856 709 876
rect 724 874 754 876
rect 573 848 614 856
rect 696 852 709 856
rect 761 860 840 876
rect 872 876 1044 878
rect 872 860 951 876
rect 958 874 988 876
rect 536 838 565 848
rect 579 838 608 848
rect 623 838 653 852
rect 696 838 739 852
rect 761 848 951 860
rect 1016 856 1022 876
rect 746 838 776 848
rect 777 838 935 848
rect 939 838 969 848
rect 973 838 1003 852
rect 1031 838 1044 876
rect 1116 890 1145 906
rect 1159 890 1188 906
rect 1203 896 1233 912
rect 1261 890 1267 938
rect 1270 932 1289 938
rect 1304 932 1334 940
rect 1270 924 1334 932
rect 1270 908 1350 924
rect 1366 917 1428 948
rect 1444 917 1506 948
rect 1575 946 1624 971
rect 1639 946 1669 962
rect 1538 932 1568 940
rect 1575 938 1685 946
rect 1538 924 1583 932
rect 1270 906 1289 908
rect 1304 906 1350 908
rect 1270 890 1350 906
rect 1377 904 1412 917
rect 1453 914 1490 917
rect 1453 912 1495 914
rect 1382 901 1412 904
rect 1391 897 1398 901
rect 1398 896 1399 897
rect 1357 890 1367 896
rect 1116 882 1151 890
rect 1116 856 1117 882
rect 1124 856 1151 882
rect 1059 838 1089 852
rect 1116 848 1151 856
rect 1153 882 1194 890
rect 1153 856 1168 882
rect 1175 856 1194 882
rect 1258 878 1289 890
rect 1304 878 1407 890
rect 1419 880 1445 906
rect 1460 901 1490 912
rect 1522 908 1584 924
rect 1522 906 1568 908
rect 1522 890 1584 906
rect 1596 890 1602 938
rect 1605 930 1685 938
rect 1605 928 1624 930
rect 1639 928 1673 930
rect 1605 912 1685 928
rect 1605 890 1624 912
rect 1639 896 1669 912
rect 1697 906 1703 980
rect 1706 906 1725 1050
rect 1740 906 1746 1050
rect 1755 980 1768 1050
rect 1820 1046 1842 1050
rect 1813 1024 1842 1038
rect 1895 1024 1911 1038
rect 1949 1034 1955 1036
rect 1962 1034 2070 1050
rect 2077 1034 2083 1036
rect 2091 1034 2106 1050
rect 2172 1044 2191 1047
rect 1813 1022 1911 1024
rect 1938 1022 2106 1034
rect 2121 1024 2137 1038
rect 2172 1025 2194 1044
rect 2204 1038 2220 1039
rect 2203 1036 2220 1038
rect 2204 1031 2220 1036
rect 2194 1024 2200 1025
rect 2203 1024 2232 1031
rect 2121 1023 2232 1024
rect 2121 1022 2238 1023
rect 1797 1014 1848 1022
rect 1895 1014 1929 1022
rect 1797 1002 1822 1014
rect 1829 1002 1848 1014
rect 1902 1012 1929 1014
rect 1938 1012 2159 1022
rect 2194 1019 2200 1022
rect 1902 1008 2159 1012
rect 1797 994 1848 1002
rect 1895 994 2159 1008
rect 2203 1014 2238 1022
rect 1749 946 1768 980
rect 1813 986 1842 994
rect 1813 980 1830 986
rect 1813 978 1847 980
rect 1895 978 1911 994
rect 1912 984 2120 994
rect 2121 984 2137 994
rect 2185 990 2200 1005
rect 2203 1002 2204 1014
rect 2211 1002 2238 1014
rect 2203 994 2238 1002
rect 2203 993 2232 994
rect 1923 980 2137 984
rect 1938 978 2137 980
rect 2172 980 2185 990
rect 2203 980 2220 993
rect 2172 978 2220 980
rect 1814 974 1847 978
rect 1810 972 1847 974
rect 1810 971 1877 972
rect 1810 966 1841 971
rect 1847 966 1877 971
rect 1810 962 1877 966
rect 1783 959 1877 962
rect 1783 952 1832 959
rect 1783 946 1813 952
rect 1832 947 1837 952
rect 1749 930 1829 946
rect 1841 938 1877 959
rect 1938 954 2127 978
rect 2172 977 2219 978
rect 2185 972 2219 977
rect 1953 951 2127 954
rect 1946 948 2127 951
rect 2155 971 2219 972
rect 1749 928 1768 930
rect 1783 928 1817 930
rect 1749 912 1829 928
rect 1749 906 1768 912
rect 1465 880 1568 890
rect 1419 878 1568 880
rect 1589 878 1624 890
rect 1258 876 1420 878
rect 1270 856 1289 876
rect 1304 874 1334 876
rect 1153 848 1194 856
rect 1276 852 1289 856
rect 1341 860 1420 876
rect 1452 876 1624 878
rect 1452 860 1531 876
rect 1538 874 1568 876
rect 1116 838 1145 848
rect 1159 838 1188 848
rect 1203 838 1233 852
rect 1276 838 1319 852
rect 1341 848 1531 860
rect 1596 856 1602 876
rect 1326 838 1356 848
rect 1357 838 1515 848
rect 1519 838 1549 848
rect 1553 838 1583 852
rect 1611 838 1624 876
rect 1696 890 1725 906
rect 1739 890 1768 906
rect 1783 896 1813 912
rect 1841 890 1847 938
rect 1850 932 1869 938
rect 1884 932 1914 940
rect 1850 924 1914 932
rect 1850 908 1930 924
rect 1946 917 2008 948
rect 2024 917 2086 948
rect 2155 946 2204 971
rect 2219 946 2249 962
rect 2118 932 2148 940
rect 2155 938 2265 946
rect 2118 924 2163 932
rect 1850 906 1869 908
rect 1884 906 1930 908
rect 1850 890 1930 906
rect 1957 904 1992 917
rect 2033 914 2070 917
rect 2033 912 2075 914
rect 1962 901 1992 904
rect 1971 897 1978 901
rect 1978 896 1979 897
rect 1937 890 1947 896
rect 1696 882 1731 890
rect 1696 856 1697 882
rect 1704 856 1731 882
rect 1639 838 1669 852
rect 1696 848 1731 856
rect 1733 882 1774 890
rect 1733 856 1748 882
rect 1755 856 1774 882
rect 1838 878 1869 890
rect 1884 878 1987 890
rect 1999 880 2025 906
rect 2040 901 2070 912
rect 2102 908 2164 924
rect 2102 906 2148 908
rect 2102 890 2164 906
rect 2176 890 2182 938
rect 2185 930 2265 938
rect 2185 928 2204 930
rect 2219 928 2253 930
rect 2185 912 2265 928
rect 2185 890 2204 912
rect 2219 896 2249 912
rect 2277 906 2283 980
rect 2286 906 2305 1050
rect 2320 906 2326 1050
rect 2335 980 2348 1050
rect 2400 1046 2422 1050
rect 2393 1024 2422 1038
rect 2475 1024 2491 1038
rect 2529 1034 2535 1036
rect 2542 1034 2650 1050
rect 2657 1034 2663 1036
rect 2671 1034 2686 1050
rect 2752 1044 2771 1047
rect 2393 1022 2491 1024
rect 2518 1022 2686 1034
rect 2701 1024 2717 1038
rect 2752 1025 2774 1044
rect 2784 1038 2800 1039
rect 2783 1036 2800 1038
rect 2784 1031 2800 1036
rect 2774 1024 2780 1025
rect 2783 1024 2812 1031
rect 2701 1023 2812 1024
rect 2701 1022 2818 1023
rect 2377 1014 2428 1022
rect 2475 1014 2509 1022
rect 2377 1002 2402 1014
rect 2409 1002 2428 1014
rect 2482 1012 2509 1014
rect 2518 1012 2739 1022
rect 2774 1019 2780 1022
rect 2482 1008 2739 1012
rect 2377 994 2428 1002
rect 2475 994 2739 1008
rect 2783 1014 2818 1022
rect 2329 946 2348 980
rect 2393 986 2422 994
rect 2393 980 2410 986
rect 2393 978 2427 980
rect 2475 978 2491 994
rect 2492 984 2700 994
rect 2701 984 2717 994
rect 2765 990 2780 1005
rect 2783 1002 2784 1014
rect 2791 1002 2818 1014
rect 2783 994 2818 1002
rect 2783 993 2812 994
rect 2503 980 2717 984
rect 2518 978 2717 980
rect 2752 980 2765 990
rect 2783 980 2800 993
rect 2752 978 2800 980
rect 2394 974 2427 978
rect 2390 972 2427 974
rect 2390 971 2457 972
rect 2390 966 2421 971
rect 2427 966 2457 971
rect 2390 962 2457 966
rect 2363 959 2457 962
rect 2363 952 2412 959
rect 2363 946 2393 952
rect 2412 947 2417 952
rect 2329 930 2409 946
rect 2421 938 2457 959
rect 2518 954 2707 978
rect 2752 977 2799 978
rect 2765 972 2799 977
rect 2533 951 2707 954
rect 2526 948 2707 951
rect 2735 971 2799 972
rect 2329 928 2348 930
rect 2363 928 2397 930
rect 2329 912 2409 928
rect 2329 906 2348 912
rect 2045 880 2148 890
rect 1999 878 2148 880
rect 2169 878 2204 890
rect 1838 876 2000 878
rect 1850 856 1869 876
rect 1884 874 1914 876
rect 1733 848 1774 856
rect 1856 852 1869 856
rect 1921 860 2000 876
rect 2032 876 2204 878
rect 2032 860 2111 876
rect 2118 874 2148 876
rect 1696 838 1725 848
rect 1739 838 1768 848
rect 1783 838 1813 852
rect 1856 838 1899 852
rect 1921 848 2111 860
rect 2176 856 2182 876
rect 1906 838 1936 848
rect 1937 838 2095 848
rect 2099 838 2129 848
rect 2133 838 2163 852
rect 2191 838 2204 876
rect 2276 890 2305 906
rect 2319 890 2348 906
rect 2363 896 2393 912
rect 2421 890 2427 938
rect 2430 932 2449 938
rect 2464 932 2494 940
rect 2430 924 2494 932
rect 2430 908 2510 924
rect 2526 917 2588 948
rect 2604 917 2666 948
rect 2735 946 2784 971
rect 2799 946 2829 962
rect 2698 932 2728 940
rect 2735 938 2845 946
rect 2698 924 2743 932
rect 2430 906 2449 908
rect 2464 906 2510 908
rect 2430 890 2510 906
rect 2537 904 2572 917
rect 2613 914 2650 917
rect 2613 912 2655 914
rect 2542 901 2572 904
rect 2551 897 2558 901
rect 2558 896 2559 897
rect 2517 890 2527 896
rect 2276 882 2311 890
rect 2276 856 2277 882
rect 2284 856 2311 882
rect 2219 838 2249 852
rect 2276 848 2311 856
rect 2313 882 2354 890
rect 2313 856 2328 882
rect 2335 856 2354 882
rect 2418 878 2449 890
rect 2464 878 2567 890
rect 2579 880 2605 906
rect 2620 901 2650 912
rect 2682 908 2744 924
rect 2682 906 2728 908
rect 2682 890 2744 906
rect 2756 890 2762 938
rect 2765 930 2845 938
rect 2765 928 2784 930
rect 2799 928 2833 930
rect 2765 912 2845 928
rect 2765 890 2784 912
rect 2799 896 2829 912
rect 2857 906 2863 980
rect 2866 906 2885 1050
rect 2900 906 2906 1050
rect 2915 980 2928 1050
rect 2980 1046 3002 1050
rect 2973 1024 3002 1038
rect 3055 1024 3071 1038
rect 3109 1034 3115 1036
rect 3122 1034 3230 1050
rect 3237 1034 3243 1036
rect 3251 1034 3266 1050
rect 3332 1044 3351 1047
rect 2973 1022 3071 1024
rect 3098 1022 3266 1034
rect 3281 1024 3297 1038
rect 3332 1025 3354 1044
rect 3364 1038 3380 1039
rect 3363 1036 3380 1038
rect 3364 1031 3380 1036
rect 3354 1024 3360 1025
rect 3363 1024 3392 1031
rect 3281 1023 3392 1024
rect 3281 1022 3398 1023
rect 2957 1014 3008 1022
rect 3055 1014 3089 1022
rect 2957 1002 2982 1014
rect 2989 1002 3008 1014
rect 3062 1012 3089 1014
rect 3098 1012 3319 1022
rect 3354 1019 3360 1022
rect 3062 1008 3319 1012
rect 2957 994 3008 1002
rect 3055 994 3319 1008
rect 3363 1014 3398 1022
rect 2909 946 2928 980
rect 2973 986 3002 994
rect 2973 980 2990 986
rect 2973 978 3007 980
rect 3055 978 3071 994
rect 3072 984 3280 994
rect 3281 984 3297 994
rect 3345 990 3360 1005
rect 3363 1002 3364 1014
rect 3371 1002 3398 1014
rect 3363 994 3398 1002
rect 3363 993 3392 994
rect 3083 980 3297 984
rect 3098 978 3297 980
rect 3332 980 3345 990
rect 3363 980 3380 993
rect 3332 978 3380 980
rect 2974 974 3007 978
rect 2970 972 3007 974
rect 2970 971 3037 972
rect 2970 966 3001 971
rect 3007 966 3037 971
rect 2970 962 3037 966
rect 2943 959 3037 962
rect 2943 952 2992 959
rect 2943 946 2973 952
rect 2992 947 2997 952
rect 2909 930 2989 946
rect 3001 938 3037 959
rect 3098 954 3287 978
rect 3332 977 3379 978
rect 3345 972 3379 977
rect 3113 951 3287 954
rect 3106 948 3287 951
rect 3315 971 3379 972
rect 2909 928 2928 930
rect 2943 928 2977 930
rect 2909 912 2989 928
rect 2909 906 2928 912
rect 2625 880 2728 890
rect 2579 878 2728 880
rect 2749 878 2784 890
rect 2418 876 2580 878
rect 2430 856 2449 876
rect 2464 874 2494 876
rect 2313 848 2354 856
rect 2436 852 2449 856
rect 2501 860 2580 876
rect 2612 876 2784 878
rect 2612 860 2691 876
rect 2698 874 2728 876
rect 2276 838 2305 848
rect 2319 838 2348 848
rect 2363 838 2393 852
rect 2436 838 2479 852
rect 2501 848 2691 860
rect 2756 856 2762 876
rect 2486 838 2516 848
rect 2517 838 2675 848
rect 2679 838 2709 848
rect 2713 838 2743 852
rect 2771 838 2784 876
rect 2856 890 2885 906
rect 2899 890 2928 906
rect 2943 896 2973 912
rect 3001 890 3007 938
rect 3010 932 3029 938
rect 3044 932 3074 940
rect 3010 924 3074 932
rect 3010 908 3090 924
rect 3106 917 3168 948
rect 3184 917 3246 948
rect 3315 946 3364 971
rect 3379 946 3409 962
rect 3278 932 3308 940
rect 3315 938 3425 946
rect 3278 924 3323 932
rect 3010 906 3029 908
rect 3044 906 3090 908
rect 3010 890 3090 906
rect 3117 904 3152 917
rect 3193 914 3230 917
rect 3193 912 3235 914
rect 3122 901 3152 904
rect 3131 897 3138 901
rect 3138 896 3139 897
rect 3097 890 3107 896
rect 2856 882 2891 890
rect 2856 856 2857 882
rect 2864 856 2891 882
rect 2799 838 2829 852
rect 2856 848 2891 856
rect 2893 882 2934 890
rect 2893 856 2908 882
rect 2915 856 2934 882
rect 2998 878 3029 890
rect 3044 878 3147 890
rect 3159 880 3185 906
rect 3200 901 3230 912
rect 3262 908 3324 924
rect 3262 906 3308 908
rect 3262 890 3324 906
rect 3336 890 3342 938
rect 3345 930 3425 938
rect 3345 928 3364 930
rect 3379 928 3413 930
rect 3345 912 3425 928
rect 3345 890 3364 912
rect 3379 896 3409 912
rect 3437 906 3443 980
rect 3446 906 3465 1050
rect 3480 906 3486 1050
rect 3495 980 3508 1050
rect 3560 1046 3582 1050
rect 3553 1024 3582 1038
rect 3635 1024 3651 1038
rect 3689 1034 3695 1036
rect 3702 1034 3810 1050
rect 3817 1034 3823 1036
rect 3831 1034 3846 1050
rect 3912 1044 3931 1047
rect 3553 1022 3651 1024
rect 3678 1022 3846 1034
rect 3861 1024 3877 1038
rect 3912 1025 3934 1044
rect 3944 1038 3960 1039
rect 3943 1036 3960 1038
rect 3944 1031 3960 1036
rect 3934 1024 3940 1025
rect 3943 1024 3972 1031
rect 3861 1023 3972 1024
rect 3861 1022 3978 1023
rect 3537 1014 3588 1022
rect 3635 1014 3669 1022
rect 3537 1002 3562 1014
rect 3569 1002 3588 1014
rect 3642 1012 3669 1014
rect 3678 1012 3899 1022
rect 3934 1019 3940 1022
rect 3642 1008 3899 1012
rect 3537 994 3588 1002
rect 3635 994 3899 1008
rect 3943 1014 3978 1022
rect 3489 946 3508 980
rect 3553 986 3582 994
rect 3553 980 3570 986
rect 3553 978 3587 980
rect 3635 978 3651 994
rect 3652 984 3860 994
rect 3861 984 3877 994
rect 3925 990 3940 1005
rect 3943 1002 3944 1014
rect 3951 1002 3978 1014
rect 3943 994 3978 1002
rect 3943 993 3972 994
rect 3663 980 3877 984
rect 3678 978 3877 980
rect 3912 980 3925 990
rect 3943 980 3960 993
rect 3912 978 3960 980
rect 3554 974 3587 978
rect 3550 972 3587 974
rect 3550 971 3617 972
rect 3550 966 3581 971
rect 3587 966 3617 971
rect 3550 962 3617 966
rect 3523 959 3617 962
rect 3523 952 3572 959
rect 3523 946 3553 952
rect 3572 947 3577 952
rect 3489 930 3569 946
rect 3581 938 3617 959
rect 3678 954 3867 978
rect 3912 977 3959 978
rect 3925 972 3959 977
rect 3693 951 3867 954
rect 3686 948 3867 951
rect 3895 971 3959 972
rect 3489 928 3508 930
rect 3523 928 3557 930
rect 3489 912 3569 928
rect 3489 906 3508 912
rect 3205 880 3308 890
rect 3159 878 3308 880
rect 3329 878 3364 890
rect 2998 876 3160 878
rect 3010 856 3029 876
rect 3044 874 3074 876
rect 2893 848 2934 856
rect 3016 852 3029 856
rect 3081 860 3160 876
rect 3192 876 3364 878
rect 3192 860 3271 876
rect 3278 874 3308 876
rect 2856 838 2885 848
rect 2899 838 2928 848
rect 2943 838 2973 852
rect 3016 838 3059 852
rect 3081 848 3271 860
rect 3336 856 3342 876
rect 3066 838 3096 848
rect 3097 838 3255 848
rect 3259 838 3289 848
rect 3293 838 3323 852
rect 3351 838 3364 876
rect 3436 890 3465 906
rect 3479 890 3508 906
rect 3523 896 3553 912
rect 3581 890 3587 938
rect 3590 932 3609 938
rect 3624 932 3654 940
rect 3590 924 3654 932
rect 3590 908 3670 924
rect 3686 917 3748 948
rect 3764 917 3826 948
rect 3895 946 3944 971
rect 3959 946 3989 962
rect 3858 932 3888 940
rect 3895 938 4005 946
rect 3858 924 3903 932
rect 3590 906 3609 908
rect 3624 906 3670 908
rect 3590 890 3670 906
rect 3697 904 3732 917
rect 3773 914 3810 917
rect 3773 912 3815 914
rect 3702 901 3732 904
rect 3711 897 3718 901
rect 3718 896 3719 897
rect 3677 890 3687 896
rect 3436 882 3471 890
rect 3436 856 3437 882
rect 3444 856 3471 882
rect 3379 838 3409 852
rect 3436 848 3471 856
rect 3473 882 3514 890
rect 3473 856 3488 882
rect 3495 856 3514 882
rect 3578 878 3609 890
rect 3624 878 3727 890
rect 3739 880 3765 906
rect 3780 901 3810 912
rect 3842 908 3904 924
rect 3842 906 3888 908
rect 3842 890 3904 906
rect 3916 890 3922 938
rect 3925 930 4005 938
rect 3925 928 3944 930
rect 3959 928 3993 930
rect 3925 912 4005 928
rect 3925 890 3944 912
rect 3959 896 3989 912
rect 4017 906 4023 980
rect 4026 906 4045 1050
rect 4060 906 4066 1050
rect 4075 980 4088 1050
rect 4140 1046 4162 1050
rect 4133 1024 4162 1038
rect 4215 1024 4231 1038
rect 4269 1034 4275 1036
rect 4282 1034 4390 1050
rect 4397 1034 4403 1036
rect 4411 1034 4426 1050
rect 4492 1044 4511 1047
rect 4133 1022 4231 1024
rect 4258 1022 4426 1034
rect 4441 1024 4457 1038
rect 4492 1025 4514 1044
rect 4524 1038 4540 1039
rect 4523 1036 4540 1038
rect 4524 1031 4540 1036
rect 4514 1024 4520 1025
rect 4523 1024 4552 1031
rect 4441 1023 4552 1024
rect 4441 1022 4558 1023
rect 4117 1014 4168 1022
rect 4215 1014 4249 1022
rect 4117 1002 4142 1014
rect 4149 1002 4168 1014
rect 4222 1012 4249 1014
rect 4258 1012 4479 1022
rect 4514 1019 4520 1022
rect 4222 1008 4479 1012
rect 4117 994 4168 1002
rect 4215 994 4479 1008
rect 4523 1014 4558 1022
rect 4069 946 4088 980
rect 4133 986 4162 994
rect 4133 980 4150 986
rect 4133 978 4167 980
rect 4215 978 4231 994
rect 4232 984 4440 994
rect 4441 984 4457 994
rect 4505 990 4520 1005
rect 4523 1002 4524 1014
rect 4531 1002 4558 1014
rect 4523 994 4558 1002
rect 4523 993 4552 994
rect 4243 980 4457 984
rect 4258 978 4457 980
rect 4492 980 4505 990
rect 4523 980 4540 993
rect 4492 978 4540 980
rect 4134 974 4167 978
rect 4130 972 4167 974
rect 4130 971 4197 972
rect 4130 966 4161 971
rect 4167 966 4197 971
rect 4130 962 4197 966
rect 4103 959 4197 962
rect 4103 952 4152 959
rect 4103 946 4133 952
rect 4152 947 4157 952
rect 4069 930 4149 946
rect 4161 938 4197 959
rect 4258 954 4447 978
rect 4492 977 4539 978
rect 4505 972 4539 977
rect 4273 951 4447 954
rect 4266 948 4447 951
rect 4475 971 4539 972
rect 4069 928 4088 930
rect 4103 928 4137 930
rect 4069 912 4149 928
rect 4069 906 4088 912
rect 3785 880 3888 890
rect 3739 878 3888 880
rect 3909 878 3944 890
rect 3578 876 3740 878
rect 3590 856 3609 876
rect 3624 874 3654 876
rect 3473 848 3514 856
rect 3596 852 3609 856
rect 3661 860 3740 876
rect 3772 876 3944 878
rect 3772 860 3851 876
rect 3858 874 3888 876
rect 3436 838 3465 848
rect 3479 838 3508 848
rect 3523 838 3553 852
rect 3596 838 3639 852
rect 3661 848 3851 860
rect 3916 856 3922 876
rect 3646 838 3676 848
rect 3677 838 3835 848
rect 3839 838 3869 848
rect 3873 838 3903 852
rect 3931 838 3944 876
rect 4016 890 4045 906
rect 4059 890 4088 906
rect 4103 896 4133 912
rect 4161 890 4167 938
rect 4170 932 4189 938
rect 4204 932 4234 940
rect 4170 924 4234 932
rect 4170 908 4250 924
rect 4266 917 4328 948
rect 4344 917 4406 948
rect 4475 946 4524 971
rect 4539 946 4569 962
rect 4438 932 4468 940
rect 4475 938 4585 946
rect 4438 924 4483 932
rect 4170 906 4189 908
rect 4204 906 4250 908
rect 4170 890 4250 906
rect 4277 904 4312 917
rect 4353 914 4390 917
rect 4353 912 4395 914
rect 4282 901 4312 904
rect 4291 897 4298 901
rect 4298 896 4299 897
rect 4257 890 4267 896
rect 4016 882 4051 890
rect 4016 856 4017 882
rect 4024 856 4051 882
rect 3959 838 3989 852
rect 4016 848 4051 856
rect 4053 882 4094 890
rect 4053 856 4068 882
rect 4075 856 4094 882
rect 4158 878 4189 890
rect 4204 878 4307 890
rect 4319 880 4345 906
rect 4360 901 4390 912
rect 4422 908 4484 924
rect 4422 906 4468 908
rect 4422 890 4484 906
rect 4496 890 4502 938
rect 4505 930 4585 938
rect 4505 928 4524 930
rect 4539 928 4573 930
rect 4505 912 4585 928
rect 4505 890 4524 912
rect 4539 896 4569 912
rect 4597 906 4603 980
rect 4606 906 4625 1050
rect 4640 906 4646 1050
rect 4655 980 4668 1050
rect 4720 1046 4742 1050
rect 4713 1024 4742 1038
rect 4795 1024 4811 1038
rect 4849 1034 4855 1036
rect 4862 1034 4970 1050
rect 4977 1034 4983 1036
rect 4991 1034 5006 1050
rect 5072 1044 5091 1047
rect 4713 1022 4811 1024
rect 4838 1022 5006 1034
rect 5021 1024 5037 1038
rect 5072 1025 5094 1044
rect 5104 1038 5120 1039
rect 5103 1036 5120 1038
rect 5104 1031 5120 1036
rect 5094 1024 5100 1025
rect 5103 1024 5132 1031
rect 5021 1023 5132 1024
rect 5021 1022 5138 1023
rect 4697 1014 4748 1022
rect 4795 1014 4829 1022
rect 4697 1002 4722 1014
rect 4729 1002 4748 1014
rect 4802 1012 4829 1014
rect 4838 1012 5059 1022
rect 5094 1019 5100 1022
rect 4802 1008 5059 1012
rect 4697 994 4748 1002
rect 4795 994 5059 1008
rect 5103 1014 5138 1022
rect 4649 946 4668 980
rect 4713 986 4742 994
rect 4713 980 4730 986
rect 4713 978 4747 980
rect 4795 978 4811 994
rect 4812 984 5020 994
rect 5021 984 5037 994
rect 5085 990 5100 1005
rect 5103 1002 5104 1014
rect 5111 1002 5138 1014
rect 5103 994 5138 1002
rect 5103 993 5132 994
rect 4823 980 5037 984
rect 4838 978 5037 980
rect 5072 980 5085 990
rect 5103 980 5120 993
rect 5072 978 5120 980
rect 4714 974 4747 978
rect 4710 972 4747 974
rect 4710 971 4777 972
rect 4710 966 4741 971
rect 4747 966 4777 971
rect 4710 962 4777 966
rect 4683 959 4777 962
rect 4683 952 4732 959
rect 4683 946 4713 952
rect 4732 947 4737 952
rect 4649 930 4729 946
rect 4741 938 4777 959
rect 4838 954 5027 978
rect 5072 977 5119 978
rect 5085 972 5119 977
rect 4853 951 5027 954
rect 4846 948 5027 951
rect 5055 971 5119 972
rect 4649 928 4668 930
rect 4683 928 4717 930
rect 4649 912 4729 928
rect 4649 906 4668 912
rect 4365 880 4468 890
rect 4319 878 4468 880
rect 4489 878 4524 890
rect 4158 876 4320 878
rect 4170 856 4189 876
rect 4204 874 4234 876
rect 4053 848 4094 856
rect 4176 852 4189 856
rect 4241 860 4320 876
rect 4352 876 4524 878
rect 4352 860 4431 876
rect 4438 874 4468 876
rect 4016 838 4045 848
rect 4059 838 4088 848
rect 4103 838 4133 852
rect 4176 838 4219 852
rect 4241 848 4431 860
rect 4496 856 4502 876
rect 4226 838 4256 848
rect 4257 838 4415 848
rect 4419 838 4449 848
rect 4453 838 4483 852
rect 4511 838 4524 876
rect 4596 890 4625 906
rect 4639 890 4668 906
rect 4683 896 4713 912
rect 4741 890 4747 938
rect 4750 932 4769 938
rect 4784 932 4814 940
rect 4750 924 4814 932
rect 4750 908 4830 924
rect 4846 917 4908 948
rect 4924 917 4986 948
rect 5055 946 5104 971
rect 5119 946 5149 962
rect 5018 932 5048 940
rect 5055 938 5165 946
rect 5018 924 5063 932
rect 4750 906 4769 908
rect 4784 906 4830 908
rect 4750 890 4830 906
rect 4857 904 4892 917
rect 4933 914 4970 917
rect 4933 912 4975 914
rect 4862 901 4892 904
rect 4871 897 4878 901
rect 4878 896 4879 897
rect 4837 890 4847 896
rect 4596 882 4631 890
rect 4596 856 4597 882
rect 4604 856 4631 882
rect 4539 838 4569 852
rect 4596 848 4631 856
rect 4633 882 4674 890
rect 4633 856 4648 882
rect 4655 856 4674 882
rect 4738 878 4769 890
rect 4784 878 4887 890
rect 4899 880 4925 906
rect 4940 901 4970 912
rect 5002 908 5064 924
rect 5002 906 5048 908
rect 5002 890 5064 906
rect 5076 890 5082 938
rect 5085 930 5165 938
rect 5085 928 5104 930
rect 5119 928 5153 930
rect 5085 912 5165 928
rect 5085 890 5104 912
rect 5119 896 5149 912
rect 5177 906 5183 980
rect 5186 906 5205 1050
rect 5220 906 5226 1050
rect 5235 980 5248 1050
rect 5300 1046 5322 1050
rect 5293 1024 5322 1038
rect 5375 1024 5391 1038
rect 5429 1034 5435 1036
rect 5442 1034 5550 1050
rect 5557 1034 5563 1036
rect 5571 1034 5586 1050
rect 5652 1044 5671 1047
rect 5293 1022 5391 1024
rect 5418 1022 5586 1034
rect 5601 1024 5617 1038
rect 5652 1025 5674 1044
rect 5684 1038 5700 1039
rect 5683 1036 5700 1038
rect 5684 1031 5700 1036
rect 5674 1024 5680 1025
rect 5683 1024 5712 1031
rect 5601 1023 5712 1024
rect 5601 1022 5718 1023
rect 5277 1014 5328 1022
rect 5375 1014 5409 1022
rect 5277 1002 5302 1014
rect 5309 1002 5328 1014
rect 5382 1012 5409 1014
rect 5418 1012 5639 1022
rect 5674 1019 5680 1022
rect 5382 1008 5639 1012
rect 5277 994 5328 1002
rect 5375 994 5639 1008
rect 5683 1014 5718 1022
rect 5229 946 5248 980
rect 5293 986 5322 994
rect 5293 980 5310 986
rect 5293 978 5327 980
rect 5375 978 5391 994
rect 5392 984 5600 994
rect 5601 984 5617 994
rect 5665 990 5680 1005
rect 5683 1002 5684 1014
rect 5691 1002 5718 1014
rect 5683 994 5718 1002
rect 5683 993 5712 994
rect 5403 980 5617 984
rect 5418 978 5617 980
rect 5652 980 5665 990
rect 5683 980 5700 993
rect 5652 978 5700 980
rect 5294 974 5327 978
rect 5290 972 5327 974
rect 5290 971 5357 972
rect 5290 966 5321 971
rect 5327 966 5357 971
rect 5290 962 5357 966
rect 5263 959 5357 962
rect 5263 952 5312 959
rect 5263 946 5293 952
rect 5312 947 5317 952
rect 5229 930 5309 946
rect 5321 938 5357 959
rect 5418 954 5607 978
rect 5652 977 5699 978
rect 5665 972 5699 977
rect 5433 951 5607 954
rect 5426 948 5607 951
rect 5635 971 5699 972
rect 5229 928 5248 930
rect 5263 928 5297 930
rect 5229 912 5309 928
rect 5229 906 5248 912
rect 4945 880 5048 890
rect 4899 878 5048 880
rect 5069 878 5104 890
rect 4738 876 4900 878
rect 4750 856 4769 876
rect 4784 874 4814 876
rect 4633 848 4674 856
rect 4756 852 4769 856
rect 4821 860 4900 876
rect 4932 876 5104 878
rect 4932 860 5011 876
rect 5018 874 5048 876
rect 4596 838 4625 848
rect 4639 838 4668 848
rect 4683 838 4713 852
rect 4756 838 4799 852
rect 4821 848 5011 860
rect 5076 856 5082 876
rect 4806 838 4836 848
rect 4837 838 4995 848
rect 4999 838 5029 848
rect 5033 838 5063 852
rect 5091 838 5104 876
rect 5176 890 5205 906
rect 5219 890 5248 906
rect 5263 896 5293 912
rect 5321 890 5327 938
rect 5330 932 5349 938
rect 5364 932 5394 940
rect 5330 924 5394 932
rect 5330 908 5410 924
rect 5426 917 5488 948
rect 5504 917 5566 948
rect 5635 946 5684 971
rect 5699 946 5729 962
rect 5598 932 5628 940
rect 5635 938 5745 946
rect 5598 924 5643 932
rect 5330 906 5349 908
rect 5364 906 5410 908
rect 5330 890 5410 906
rect 5437 904 5472 917
rect 5513 914 5550 917
rect 5513 912 5555 914
rect 5442 901 5472 904
rect 5451 897 5458 901
rect 5458 896 5459 897
rect 5417 890 5427 896
rect 5176 882 5211 890
rect 5176 856 5177 882
rect 5184 856 5211 882
rect 5119 838 5149 852
rect 5176 848 5211 856
rect 5213 882 5254 890
rect 5213 856 5228 882
rect 5235 856 5254 882
rect 5318 878 5349 890
rect 5364 878 5467 890
rect 5479 880 5505 906
rect 5520 901 5550 912
rect 5582 908 5644 924
rect 5582 906 5628 908
rect 5582 890 5644 906
rect 5656 890 5662 938
rect 5665 930 5745 938
rect 5665 928 5684 930
rect 5699 928 5733 930
rect 5665 912 5745 928
rect 5665 890 5684 912
rect 5699 896 5729 912
rect 5757 906 5763 980
rect 5766 906 5785 1050
rect 5800 906 5806 1050
rect 5815 980 5828 1050
rect 5880 1046 5902 1050
rect 5873 1024 5902 1038
rect 5955 1024 5971 1038
rect 6009 1034 6015 1036
rect 6022 1034 6130 1050
rect 6137 1034 6143 1036
rect 6151 1034 6166 1050
rect 6232 1044 6251 1047
rect 5873 1022 5971 1024
rect 5998 1022 6166 1034
rect 6181 1024 6197 1038
rect 6232 1025 6254 1044
rect 6264 1038 6280 1039
rect 6263 1036 6280 1038
rect 6264 1031 6280 1036
rect 6254 1024 6260 1025
rect 6263 1024 6292 1031
rect 6181 1023 6292 1024
rect 6181 1022 6298 1023
rect 5857 1014 5908 1022
rect 5955 1014 5989 1022
rect 5857 1002 5882 1014
rect 5889 1002 5908 1014
rect 5962 1012 5989 1014
rect 5998 1012 6219 1022
rect 6254 1019 6260 1022
rect 5962 1008 6219 1012
rect 5857 994 5908 1002
rect 5955 994 6219 1008
rect 6263 1014 6298 1022
rect 5809 946 5828 980
rect 5873 986 5902 994
rect 5873 980 5890 986
rect 5873 978 5907 980
rect 5955 978 5971 994
rect 5972 984 6180 994
rect 6181 984 6197 994
rect 6245 990 6260 1005
rect 6263 1002 6264 1014
rect 6271 1002 6298 1014
rect 6263 994 6298 1002
rect 6263 993 6292 994
rect 5983 980 6197 984
rect 5998 978 6197 980
rect 6232 980 6245 990
rect 6263 980 6280 993
rect 6232 978 6280 980
rect 5874 974 5907 978
rect 5870 972 5907 974
rect 5870 971 5937 972
rect 5870 966 5901 971
rect 5907 966 5937 971
rect 5870 962 5937 966
rect 5843 959 5937 962
rect 5843 952 5892 959
rect 5843 946 5873 952
rect 5892 947 5897 952
rect 5809 930 5889 946
rect 5901 938 5937 959
rect 5998 954 6187 978
rect 6232 977 6279 978
rect 6245 972 6279 977
rect 6013 951 6187 954
rect 6006 948 6187 951
rect 6215 971 6279 972
rect 5809 928 5828 930
rect 5843 928 5877 930
rect 5809 912 5889 928
rect 5809 906 5828 912
rect 5525 880 5628 890
rect 5479 878 5628 880
rect 5649 878 5684 890
rect 5318 876 5480 878
rect 5330 856 5349 876
rect 5364 874 5394 876
rect 5213 848 5254 856
rect 5336 852 5349 856
rect 5401 860 5480 876
rect 5512 876 5684 878
rect 5512 860 5591 876
rect 5598 874 5628 876
rect 5176 838 5205 848
rect 5219 838 5248 848
rect 5263 838 5293 852
rect 5336 838 5379 852
rect 5401 848 5591 860
rect 5656 856 5662 876
rect 5386 838 5416 848
rect 5417 838 5575 848
rect 5579 838 5609 848
rect 5613 838 5643 852
rect 5671 838 5684 876
rect 5756 890 5785 906
rect 5799 890 5828 906
rect 5843 896 5873 912
rect 5901 890 5907 938
rect 5910 932 5929 938
rect 5944 932 5974 940
rect 5910 924 5974 932
rect 5910 908 5990 924
rect 6006 917 6068 948
rect 6084 917 6146 948
rect 6215 946 6264 971
rect 6279 946 6309 962
rect 6178 932 6208 940
rect 6215 938 6325 946
rect 6178 924 6223 932
rect 5910 906 5929 908
rect 5944 906 5990 908
rect 5910 890 5990 906
rect 6017 904 6052 917
rect 6093 914 6130 917
rect 6093 912 6135 914
rect 6022 901 6052 904
rect 6031 897 6038 901
rect 6038 896 6039 897
rect 5997 890 6007 896
rect 5756 882 5791 890
rect 5756 856 5757 882
rect 5764 856 5791 882
rect 5699 838 5729 852
rect 5756 848 5791 856
rect 5793 882 5834 890
rect 5793 856 5808 882
rect 5815 856 5834 882
rect 5898 878 5929 890
rect 5944 878 6047 890
rect 6059 880 6085 906
rect 6100 901 6130 912
rect 6162 908 6224 924
rect 6162 906 6208 908
rect 6162 890 6224 906
rect 6236 890 6242 938
rect 6245 930 6325 938
rect 6245 928 6264 930
rect 6279 928 6313 930
rect 6245 912 6325 928
rect 6245 890 6264 912
rect 6279 896 6309 912
rect 6337 906 6343 980
rect 6346 906 6365 1050
rect 6380 906 6386 1050
rect 6395 980 6408 1050
rect 6460 1046 6482 1050
rect 6453 1024 6482 1038
rect 6535 1024 6551 1038
rect 6589 1034 6595 1036
rect 6602 1034 6710 1050
rect 6717 1034 6723 1036
rect 6731 1034 6746 1050
rect 6812 1044 6831 1047
rect 6453 1022 6551 1024
rect 6578 1022 6746 1034
rect 6761 1024 6777 1038
rect 6812 1025 6834 1044
rect 6844 1038 6860 1039
rect 6843 1036 6860 1038
rect 6844 1031 6860 1036
rect 6834 1024 6840 1025
rect 6843 1024 6872 1031
rect 6761 1023 6872 1024
rect 6761 1022 6878 1023
rect 6437 1014 6488 1022
rect 6535 1014 6569 1022
rect 6437 1002 6462 1014
rect 6469 1002 6488 1014
rect 6542 1012 6569 1014
rect 6578 1012 6799 1022
rect 6834 1019 6840 1022
rect 6542 1008 6799 1012
rect 6437 994 6488 1002
rect 6535 994 6799 1008
rect 6843 1014 6878 1022
rect 6389 946 6408 980
rect 6453 986 6482 994
rect 6453 980 6470 986
rect 6453 978 6487 980
rect 6535 978 6551 994
rect 6552 984 6760 994
rect 6761 984 6777 994
rect 6825 990 6840 1005
rect 6843 1002 6844 1014
rect 6851 1002 6878 1014
rect 6843 994 6878 1002
rect 6843 993 6872 994
rect 6563 980 6777 984
rect 6578 978 6777 980
rect 6812 980 6825 990
rect 6843 980 6860 993
rect 6812 978 6860 980
rect 6454 974 6487 978
rect 6450 972 6487 974
rect 6450 971 6517 972
rect 6450 966 6481 971
rect 6487 966 6517 971
rect 6450 962 6517 966
rect 6423 959 6517 962
rect 6423 952 6472 959
rect 6423 946 6453 952
rect 6472 947 6477 952
rect 6389 930 6469 946
rect 6481 938 6517 959
rect 6578 954 6767 978
rect 6812 977 6859 978
rect 6825 972 6859 977
rect 6593 951 6767 954
rect 6586 948 6767 951
rect 6795 971 6859 972
rect 6389 928 6408 930
rect 6423 928 6457 930
rect 6389 912 6469 928
rect 6389 906 6408 912
rect 6105 880 6208 890
rect 6059 878 6208 880
rect 6229 878 6264 890
rect 5898 876 6060 878
rect 5910 856 5929 876
rect 5944 874 5974 876
rect 5793 848 5834 856
rect 5916 852 5929 856
rect 5981 860 6060 876
rect 6092 876 6264 878
rect 6092 860 6171 876
rect 6178 874 6208 876
rect 5756 838 5785 848
rect 5799 838 5828 848
rect 5843 838 5873 852
rect 5916 838 5959 852
rect 5981 848 6171 860
rect 6236 856 6242 876
rect 5966 838 5996 848
rect 5997 838 6155 848
rect 6159 838 6189 848
rect 6193 838 6223 852
rect 6251 838 6264 876
rect 6336 890 6365 906
rect 6379 890 6408 906
rect 6423 896 6453 912
rect 6481 890 6487 938
rect 6490 932 6509 938
rect 6524 932 6554 940
rect 6490 924 6554 932
rect 6490 908 6570 924
rect 6586 917 6648 948
rect 6664 917 6726 948
rect 6795 946 6844 971
rect 6859 946 6889 962
rect 6758 932 6788 940
rect 6795 938 6905 946
rect 6758 924 6803 932
rect 6490 906 6509 908
rect 6524 906 6570 908
rect 6490 890 6570 906
rect 6597 904 6632 917
rect 6673 914 6710 917
rect 6673 912 6715 914
rect 6602 901 6632 904
rect 6611 897 6618 901
rect 6618 896 6619 897
rect 6577 890 6587 896
rect 6336 882 6371 890
rect 6336 856 6337 882
rect 6344 856 6371 882
rect 6279 838 6309 852
rect 6336 848 6371 856
rect 6373 882 6414 890
rect 6373 856 6388 882
rect 6395 856 6414 882
rect 6478 878 6509 890
rect 6524 878 6627 890
rect 6639 880 6665 906
rect 6680 901 6710 912
rect 6742 908 6804 924
rect 6742 906 6788 908
rect 6742 890 6804 906
rect 6816 890 6822 938
rect 6825 930 6905 938
rect 6825 928 6844 930
rect 6859 928 6893 930
rect 6825 912 6905 928
rect 6825 890 6844 912
rect 6859 896 6889 912
rect 6917 906 6923 980
rect 6926 906 6945 1050
rect 6960 906 6966 1050
rect 6975 980 6988 1050
rect 7040 1046 7062 1050
rect 7033 1024 7062 1038
rect 7115 1024 7131 1038
rect 7169 1034 7175 1036
rect 7182 1034 7290 1050
rect 7297 1034 7303 1036
rect 7311 1034 7326 1050
rect 7392 1044 7411 1047
rect 7033 1022 7131 1024
rect 7158 1022 7326 1034
rect 7341 1024 7357 1038
rect 7392 1025 7414 1044
rect 7424 1038 7440 1039
rect 7423 1036 7440 1038
rect 7424 1031 7440 1036
rect 7414 1024 7420 1025
rect 7423 1024 7452 1031
rect 7341 1023 7452 1024
rect 7341 1022 7458 1023
rect 7017 1014 7068 1022
rect 7115 1014 7149 1022
rect 7017 1002 7042 1014
rect 7049 1002 7068 1014
rect 7122 1012 7149 1014
rect 7158 1012 7379 1022
rect 7414 1019 7420 1022
rect 7122 1008 7379 1012
rect 7017 994 7068 1002
rect 7115 994 7379 1008
rect 7423 1014 7458 1022
rect 6969 946 6988 980
rect 7033 986 7062 994
rect 7033 980 7050 986
rect 7033 978 7067 980
rect 7115 978 7131 994
rect 7132 984 7340 994
rect 7341 984 7357 994
rect 7405 990 7420 1005
rect 7423 1002 7424 1014
rect 7431 1002 7458 1014
rect 7423 994 7458 1002
rect 7423 993 7452 994
rect 7151 980 7357 984
rect 7158 978 7357 980
rect 7392 980 7405 990
rect 7423 980 7440 993
rect 7392 978 7440 980
rect 7034 974 7067 978
rect 7030 972 7067 974
rect 7030 971 7097 972
rect 7030 966 7061 971
rect 7067 966 7097 971
rect 7030 962 7097 966
rect 7003 959 7097 962
rect 7003 952 7052 959
rect 7003 946 7033 952
rect 7052 947 7057 952
rect 6969 930 7049 946
rect 7061 938 7097 959
rect 7158 954 7347 978
rect 7392 977 7439 978
rect 7405 972 7439 977
rect 7173 951 7347 954
rect 7166 948 7347 951
rect 7375 971 7439 972
rect 6969 928 6988 930
rect 7003 928 7037 930
rect 6969 912 7049 928
rect 6969 906 6988 912
rect 6685 880 6788 890
rect 6639 878 6788 880
rect 6809 878 6844 890
rect 6478 876 6640 878
rect 6490 856 6509 876
rect 6524 874 6554 876
rect 6373 848 6414 856
rect 6496 852 6509 856
rect 6561 860 6640 876
rect 6672 876 6844 878
rect 6672 860 6751 876
rect 6758 874 6788 876
rect 6336 838 6365 848
rect 6379 838 6408 848
rect 6423 838 6453 852
rect 6496 838 6539 852
rect 6561 848 6751 860
rect 6816 856 6822 876
rect 6546 838 6576 848
rect 6577 838 6735 848
rect 6739 838 6769 848
rect 6773 838 6803 852
rect 6831 838 6844 876
rect 6916 890 6945 906
rect 6959 890 6988 906
rect 7003 896 7033 912
rect 7061 890 7067 938
rect 7070 932 7089 938
rect 7104 932 7134 940
rect 7070 924 7134 932
rect 7070 908 7150 924
rect 7166 917 7228 948
rect 7244 917 7306 948
rect 7375 946 7424 971
rect 7439 946 7469 962
rect 7338 932 7368 940
rect 7375 938 7485 946
rect 7338 924 7383 932
rect 7070 906 7089 908
rect 7104 906 7150 908
rect 7070 890 7150 906
rect 7177 904 7212 917
rect 7253 914 7290 917
rect 7253 912 7295 914
rect 7182 901 7212 904
rect 7191 897 7198 901
rect 7198 896 7199 897
rect 7157 890 7167 896
rect 6916 882 6951 890
rect 6916 856 6917 882
rect 6924 856 6951 882
rect 6859 838 6889 852
rect 6916 848 6951 856
rect 6953 882 6994 890
rect 6953 856 6968 882
rect 6975 856 6994 882
rect 7058 878 7089 890
rect 7104 878 7207 890
rect 7219 880 7245 906
rect 7260 901 7290 912
rect 7322 908 7384 924
rect 7322 906 7368 908
rect 7322 890 7384 906
rect 7396 890 7402 938
rect 7405 930 7485 938
rect 7405 928 7424 930
rect 7439 928 7473 930
rect 7405 912 7485 928
rect 7405 890 7424 912
rect 7439 896 7469 912
rect 7497 906 7503 980
rect 7506 906 7525 1050
rect 7540 906 7546 1050
rect 7555 980 7568 1050
rect 7620 1046 7642 1050
rect 7613 1024 7642 1038
rect 7695 1024 7711 1038
rect 7749 1034 7755 1036
rect 7762 1034 7870 1050
rect 7877 1034 7883 1036
rect 7891 1034 7906 1050
rect 7972 1044 7991 1047
rect 7613 1022 7711 1024
rect 7738 1022 7906 1034
rect 7921 1024 7937 1038
rect 7972 1025 7994 1044
rect 8004 1038 8020 1039
rect 8003 1036 8020 1038
rect 8004 1031 8020 1036
rect 7994 1024 8000 1025
rect 8003 1024 8032 1031
rect 7921 1023 8032 1024
rect 7921 1022 8038 1023
rect 7597 1014 7648 1022
rect 7695 1014 7729 1022
rect 7597 1002 7622 1014
rect 7629 1002 7648 1014
rect 7702 1012 7729 1014
rect 7738 1012 7959 1022
rect 7994 1019 8000 1022
rect 7702 1008 7959 1012
rect 7597 994 7648 1002
rect 7695 994 7959 1008
rect 8003 1014 8038 1022
rect 7549 946 7568 980
rect 7613 986 7642 994
rect 7613 980 7630 986
rect 7613 978 7647 980
rect 7695 978 7711 994
rect 7712 984 7920 994
rect 7921 984 7937 994
rect 7985 990 8000 1005
rect 8003 1002 8004 1014
rect 8011 1002 8038 1014
rect 8003 994 8038 1002
rect 8003 993 8032 994
rect 7723 980 7937 984
rect 7738 978 7937 980
rect 7972 980 7985 990
rect 8003 980 8020 993
rect 7972 978 8020 980
rect 7614 974 7647 978
rect 7610 972 7647 974
rect 7610 971 7677 972
rect 7610 966 7641 971
rect 7647 966 7677 971
rect 7610 962 7677 966
rect 7583 959 7677 962
rect 7583 952 7632 959
rect 7583 946 7613 952
rect 7632 947 7637 952
rect 7549 930 7629 946
rect 7641 938 7677 959
rect 7738 954 7927 978
rect 7972 977 8019 978
rect 7985 972 8019 977
rect 7753 951 7927 954
rect 7746 948 7927 951
rect 7955 971 8019 972
rect 7549 928 7568 930
rect 7583 928 7617 930
rect 7549 912 7629 928
rect 7549 906 7568 912
rect 7265 880 7368 890
rect 7219 878 7368 880
rect 7389 878 7424 890
rect 7058 876 7220 878
rect 7070 856 7089 876
rect 7104 874 7134 876
rect 6953 848 6994 856
rect 7076 852 7089 856
rect 7141 860 7220 876
rect 7252 876 7424 878
rect 7252 860 7331 876
rect 7338 874 7368 876
rect 6916 838 6945 848
rect 6959 838 6988 848
rect 7003 838 7033 852
rect 7076 838 7119 852
rect 7141 848 7331 860
rect 7396 856 7402 876
rect 7126 838 7156 848
rect 7157 838 7315 848
rect 7319 838 7349 848
rect 7353 838 7383 852
rect 7411 838 7424 876
rect 7496 890 7525 906
rect 7539 890 7568 906
rect 7583 896 7613 912
rect 7641 890 7647 938
rect 7650 932 7669 938
rect 7684 932 7714 940
rect 7650 924 7714 932
rect 7650 908 7730 924
rect 7746 917 7808 948
rect 7824 917 7886 948
rect 7955 946 8004 971
rect 8019 946 8049 962
rect 7918 932 7948 940
rect 7955 938 8065 946
rect 7918 924 7963 932
rect 7650 906 7669 908
rect 7684 906 7730 908
rect 7650 890 7730 906
rect 7757 904 7792 917
rect 7833 914 7870 917
rect 7833 912 7875 914
rect 7762 901 7792 904
rect 7771 897 7778 901
rect 7778 896 7779 897
rect 7737 890 7747 896
rect 7496 882 7531 890
rect 7496 856 7497 882
rect 7504 856 7531 882
rect 7439 838 7469 852
rect 7496 848 7531 856
rect 7533 882 7574 890
rect 7533 856 7548 882
rect 7555 856 7574 882
rect 7638 878 7669 890
rect 7684 878 7787 890
rect 7799 880 7825 906
rect 7840 901 7870 912
rect 7902 908 7964 924
rect 7902 906 7948 908
rect 7902 890 7964 906
rect 7976 890 7982 938
rect 7985 930 8065 938
rect 7985 928 8004 930
rect 8019 928 8053 930
rect 7985 912 8065 928
rect 7985 890 8004 912
rect 8019 896 8049 912
rect 8077 906 8083 980
rect 8086 906 8105 1050
rect 8120 906 8126 1050
rect 8135 980 8148 1050
rect 8200 1046 8222 1050
rect 8193 1024 8222 1038
rect 8275 1024 8291 1038
rect 8329 1034 8335 1036
rect 8342 1034 8450 1050
rect 8457 1034 8463 1036
rect 8471 1034 8486 1050
rect 8552 1044 8571 1047
rect 8193 1022 8291 1024
rect 8318 1022 8486 1034
rect 8501 1024 8517 1038
rect 8552 1025 8574 1044
rect 8584 1038 8600 1039
rect 8583 1036 8600 1038
rect 8584 1031 8600 1036
rect 8574 1024 8580 1025
rect 8583 1024 8612 1031
rect 8501 1023 8612 1024
rect 8501 1022 8618 1023
rect 8177 1014 8228 1022
rect 8275 1014 8309 1022
rect 8177 1002 8202 1014
rect 8209 1002 8228 1014
rect 8282 1012 8309 1014
rect 8318 1012 8539 1022
rect 8574 1019 8580 1022
rect 8282 1008 8539 1012
rect 8177 994 8228 1002
rect 8275 994 8539 1008
rect 8583 1014 8618 1022
rect 8129 946 8148 980
rect 8193 986 8222 994
rect 8193 980 8210 986
rect 8193 978 8227 980
rect 8275 978 8291 994
rect 8292 984 8500 994
rect 8501 984 8517 994
rect 8565 990 8580 1005
rect 8583 1002 8584 1014
rect 8591 1002 8618 1014
rect 8583 994 8618 1002
rect 8583 993 8612 994
rect 8303 980 8517 984
rect 8318 978 8517 980
rect 8552 980 8565 990
rect 8583 980 8600 993
rect 8552 978 8600 980
rect 8194 974 8227 978
rect 8190 972 8227 974
rect 8190 971 8257 972
rect 8190 966 8221 971
rect 8227 966 8257 971
rect 8190 962 8257 966
rect 8163 959 8257 962
rect 8163 952 8212 959
rect 8163 946 8193 952
rect 8212 947 8217 952
rect 8129 930 8209 946
rect 8221 938 8257 959
rect 8318 954 8507 978
rect 8552 977 8599 978
rect 8565 972 8599 977
rect 8333 951 8507 954
rect 8326 948 8507 951
rect 8535 971 8599 972
rect 8129 928 8148 930
rect 8163 928 8197 930
rect 8129 912 8209 928
rect 8129 906 8148 912
rect 7845 880 7948 890
rect 7799 878 7948 880
rect 7969 878 8004 890
rect 7638 876 7800 878
rect 7650 856 7669 876
rect 7684 874 7714 876
rect 7533 848 7574 856
rect 7656 852 7669 856
rect 7721 860 7800 876
rect 7832 876 8004 878
rect 7832 860 7911 876
rect 7918 874 7948 876
rect 7496 838 7525 848
rect 7539 838 7568 848
rect 7583 838 7613 852
rect 7656 838 7699 852
rect 7721 848 7911 860
rect 7976 856 7982 876
rect 7706 838 7736 848
rect 7737 838 7895 848
rect 7899 838 7929 848
rect 7933 838 7963 852
rect 7991 838 8004 876
rect 8076 890 8105 906
rect 8119 890 8148 906
rect 8163 896 8193 912
rect 8221 890 8227 938
rect 8230 932 8249 938
rect 8264 932 8294 940
rect 8230 924 8294 932
rect 8230 908 8310 924
rect 8326 917 8388 948
rect 8404 917 8466 948
rect 8535 946 8584 971
rect 8599 946 8629 962
rect 8498 932 8528 940
rect 8535 938 8645 946
rect 8498 924 8543 932
rect 8230 906 8249 908
rect 8264 906 8310 908
rect 8230 890 8310 906
rect 8337 904 8372 917
rect 8413 914 8450 917
rect 8413 912 8455 914
rect 8342 901 8372 904
rect 8351 897 8358 901
rect 8358 896 8359 897
rect 8317 890 8327 896
rect 8076 882 8111 890
rect 8076 856 8077 882
rect 8084 856 8111 882
rect 8019 838 8049 852
rect 8076 848 8111 856
rect 8113 882 8154 890
rect 8113 856 8128 882
rect 8135 856 8154 882
rect 8218 878 8249 890
rect 8264 878 8367 890
rect 8379 880 8405 906
rect 8420 901 8450 912
rect 8482 908 8544 924
rect 8482 906 8528 908
rect 8482 890 8544 906
rect 8556 890 8562 938
rect 8565 930 8645 938
rect 8565 928 8584 930
rect 8599 928 8633 930
rect 8565 912 8645 928
rect 8565 890 8584 912
rect 8599 896 8629 912
rect 8657 906 8663 980
rect 8666 906 8685 1050
rect 8700 906 8706 1050
rect 8715 980 8728 1050
rect 8780 1046 8802 1050
rect 8773 1024 8802 1038
rect 8855 1024 8871 1038
rect 8909 1034 8915 1036
rect 8922 1034 9030 1050
rect 9037 1034 9043 1036
rect 9051 1034 9066 1050
rect 9132 1044 9151 1047
rect 8773 1022 8871 1024
rect 8898 1022 9066 1034
rect 9081 1024 9097 1038
rect 9132 1025 9154 1044
rect 9164 1038 9180 1039
rect 9163 1036 9180 1038
rect 9164 1031 9180 1036
rect 9154 1024 9160 1025
rect 9163 1024 9192 1031
rect 9081 1023 9192 1024
rect 9081 1022 9198 1023
rect 8757 1014 8808 1022
rect 8855 1014 8889 1022
rect 8757 1002 8782 1014
rect 8789 1002 8808 1014
rect 8862 1012 8889 1014
rect 8898 1012 9119 1022
rect 9154 1019 9160 1022
rect 8862 1008 9119 1012
rect 8757 994 8808 1002
rect 8855 994 9119 1008
rect 9163 1014 9198 1022
rect 8709 946 8728 980
rect 8773 986 8802 994
rect 8773 980 8790 986
rect 8773 978 8807 980
rect 8855 978 8871 994
rect 8872 984 9080 994
rect 9081 984 9097 994
rect 9145 990 9160 1005
rect 9163 1002 9164 1014
rect 9171 1002 9198 1014
rect 9163 994 9198 1002
rect 9163 993 9192 994
rect 8883 980 9097 984
rect 8898 978 9097 980
rect 9132 980 9145 990
rect 9163 980 9180 993
rect 9132 978 9180 980
rect 8774 974 8807 978
rect 8770 972 8807 974
rect 8770 971 8837 972
rect 8770 966 8801 971
rect 8807 966 8837 971
rect 8770 962 8837 966
rect 8743 959 8837 962
rect 8743 952 8792 959
rect 8743 946 8773 952
rect 8792 947 8797 952
rect 8709 930 8789 946
rect 8801 938 8837 959
rect 8898 954 9087 978
rect 9132 977 9179 978
rect 9145 972 9179 977
rect 8913 951 9087 954
rect 8906 948 9087 951
rect 9115 971 9179 972
rect 8709 928 8728 930
rect 8743 928 8777 930
rect 8709 912 8789 928
rect 8709 906 8728 912
rect 8425 880 8528 890
rect 8379 878 8528 880
rect 8549 878 8584 890
rect 8218 876 8380 878
rect 8230 856 8249 876
rect 8264 874 8294 876
rect 8113 848 8154 856
rect 8236 852 8249 856
rect 8301 860 8380 876
rect 8412 876 8584 878
rect 8412 860 8491 876
rect 8498 874 8528 876
rect 8076 838 8105 848
rect 8119 838 8148 848
rect 8163 838 8193 852
rect 8236 838 8279 852
rect 8301 848 8491 860
rect 8556 856 8562 876
rect 8286 838 8316 848
rect 8317 838 8475 848
rect 8479 838 8509 848
rect 8513 838 8543 852
rect 8571 838 8584 876
rect 8656 890 8685 906
rect 8699 890 8728 906
rect 8743 896 8773 912
rect 8801 890 8807 938
rect 8810 932 8829 938
rect 8844 932 8874 940
rect 8810 924 8874 932
rect 8810 908 8890 924
rect 8906 917 8968 948
rect 8984 917 9046 948
rect 9115 946 9164 971
rect 9179 946 9209 962
rect 9078 932 9108 940
rect 9115 938 9225 946
rect 9078 924 9123 932
rect 8810 906 8829 908
rect 8844 906 8890 908
rect 8810 890 8890 906
rect 8917 904 8952 917
rect 8993 914 9030 917
rect 8993 912 9035 914
rect 8922 901 8952 904
rect 8931 897 8938 901
rect 8938 896 8939 897
rect 8897 890 8907 896
rect 8656 882 8691 890
rect 8656 856 8657 882
rect 8664 856 8691 882
rect 8599 838 8629 852
rect 8656 848 8691 856
rect 8693 882 8734 890
rect 8693 856 8708 882
rect 8715 856 8734 882
rect 8798 878 8829 890
rect 8844 878 8947 890
rect 8959 880 8985 906
rect 9000 901 9030 912
rect 9062 908 9124 924
rect 9062 906 9108 908
rect 9062 890 9124 906
rect 9136 890 9142 938
rect 9145 930 9225 938
rect 9145 928 9164 930
rect 9179 928 9213 930
rect 9145 912 9225 928
rect 9145 890 9164 912
rect 9179 896 9209 912
rect 9237 906 9243 980
rect 9246 906 9265 1050
rect 9280 906 9286 1050
rect 9295 980 9308 1050
rect 9360 1046 9382 1050
rect 9353 1024 9382 1038
rect 9435 1024 9451 1038
rect 9489 1034 9495 1036
rect 9502 1034 9610 1050
rect 9617 1034 9623 1036
rect 9631 1034 9646 1050
rect 9712 1044 9731 1047
rect 9353 1022 9451 1024
rect 9478 1022 9646 1034
rect 9661 1024 9677 1038
rect 9712 1025 9734 1044
rect 9744 1038 9760 1039
rect 9743 1036 9760 1038
rect 9744 1031 9760 1036
rect 9734 1024 9740 1025
rect 9743 1024 9772 1031
rect 9661 1023 9772 1024
rect 9661 1022 9778 1023
rect 9337 1014 9388 1022
rect 9435 1014 9469 1022
rect 9337 1002 9362 1014
rect 9369 1002 9388 1014
rect 9442 1012 9469 1014
rect 9478 1012 9699 1022
rect 9734 1019 9740 1022
rect 9442 1008 9699 1012
rect 9337 994 9388 1002
rect 9435 994 9699 1008
rect 9743 1014 9778 1022
rect 9289 946 9308 980
rect 9353 986 9382 994
rect 9353 980 9370 986
rect 9353 978 9387 980
rect 9435 978 9451 994
rect 9452 984 9660 994
rect 9661 984 9677 994
rect 9725 990 9740 1005
rect 9743 1002 9744 1014
rect 9751 1002 9778 1014
rect 9743 994 9778 1002
rect 9743 993 9772 994
rect 9463 980 9677 984
rect 9478 978 9677 980
rect 9712 980 9725 990
rect 9743 980 9760 993
rect 9712 978 9760 980
rect 9354 974 9387 978
rect 9350 972 9387 974
rect 9350 971 9417 972
rect 9350 966 9381 971
rect 9387 966 9417 971
rect 9350 962 9417 966
rect 9323 959 9417 962
rect 9323 952 9372 959
rect 9323 946 9353 952
rect 9372 947 9377 952
rect 9289 930 9369 946
rect 9381 938 9417 959
rect 9478 954 9667 978
rect 9712 977 9759 978
rect 9725 972 9759 977
rect 9493 951 9667 954
rect 9486 948 9667 951
rect 9695 971 9759 972
rect 9289 928 9308 930
rect 9323 928 9357 930
rect 9289 912 9369 928
rect 9289 906 9308 912
rect 9005 880 9108 890
rect 8959 878 9108 880
rect 9129 878 9164 890
rect 8798 876 8960 878
rect 8810 856 8829 876
rect 8844 874 8874 876
rect 8693 848 8734 856
rect 8816 852 8829 856
rect 8881 860 8960 876
rect 8992 876 9164 878
rect 8992 860 9071 876
rect 9078 874 9108 876
rect 8656 838 8685 848
rect 8699 838 8728 848
rect 8743 838 8773 852
rect 8816 838 8859 852
rect 8881 848 9071 860
rect 9136 856 9142 876
rect 8866 838 8896 848
rect 8897 838 9055 848
rect 9059 838 9089 848
rect 9093 838 9123 852
rect 9151 838 9164 876
rect 9236 890 9265 906
rect 9279 890 9308 906
rect 9323 896 9353 912
rect 9381 890 9387 938
rect 9390 932 9409 938
rect 9424 932 9454 940
rect 9390 924 9454 932
rect 9390 908 9470 924
rect 9486 917 9548 948
rect 9564 917 9626 948
rect 9695 946 9744 971
rect 9759 946 9789 962
rect 9658 932 9688 940
rect 9695 938 9805 946
rect 9658 924 9703 932
rect 9390 906 9409 908
rect 9424 906 9470 908
rect 9390 890 9470 906
rect 9497 904 9532 917
rect 9573 914 9610 917
rect 9573 912 9615 914
rect 9502 901 9532 904
rect 9511 897 9518 901
rect 9518 896 9519 897
rect 9477 890 9487 896
rect 9236 882 9271 890
rect 9236 856 9237 882
rect 9244 856 9271 882
rect 9179 838 9209 852
rect 9236 848 9271 856
rect 9273 882 9314 890
rect 9273 856 9288 882
rect 9295 856 9314 882
rect 9378 878 9409 890
rect 9424 878 9527 890
rect 9539 880 9565 906
rect 9580 901 9610 912
rect 9642 908 9704 924
rect 9642 906 9688 908
rect 9642 890 9704 906
rect 9716 890 9722 938
rect 9725 930 9805 938
rect 9725 928 9744 930
rect 9759 928 9793 930
rect 9725 912 9805 928
rect 9725 890 9744 912
rect 9759 896 9789 912
rect 9817 906 9823 980
rect 9826 906 9845 1050
rect 9860 906 9866 1050
rect 9875 980 9888 1050
rect 9940 1046 9962 1050
rect 9933 1024 9962 1038
rect 10015 1024 10031 1038
rect 10069 1034 10075 1036
rect 10082 1034 10190 1050
rect 10197 1034 10203 1036
rect 10211 1034 10226 1050
rect 10292 1044 10311 1047
rect 9933 1022 10031 1024
rect 10058 1022 10226 1034
rect 10241 1024 10257 1038
rect 10292 1025 10314 1044
rect 10324 1038 10340 1039
rect 10323 1036 10340 1038
rect 10324 1031 10340 1036
rect 10314 1024 10320 1025
rect 10323 1024 10352 1031
rect 10241 1023 10352 1024
rect 10241 1022 10358 1023
rect 9917 1014 9968 1022
rect 10015 1014 10049 1022
rect 9917 1002 9942 1014
rect 9949 1002 9968 1014
rect 10022 1012 10049 1014
rect 10058 1012 10279 1022
rect 10314 1019 10320 1022
rect 10022 1008 10279 1012
rect 9917 994 9968 1002
rect 10015 994 10279 1008
rect 10323 1014 10358 1022
rect 9869 946 9888 980
rect 9933 986 9962 994
rect 9933 980 9950 986
rect 9933 978 9967 980
rect 10015 978 10031 994
rect 10032 984 10240 994
rect 10241 984 10257 994
rect 10305 990 10320 1005
rect 10323 1002 10324 1014
rect 10331 1002 10358 1014
rect 10323 994 10358 1002
rect 10323 993 10352 994
rect 10043 980 10257 984
rect 10058 978 10257 980
rect 10292 980 10305 990
rect 10323 980 10340 993
rect 10292 978 10340 980
rect 9934 974 9967 978
rect 9930 972 9967 974
rect 9930 971 9997 972
rect 9930 966 9961 971
rect 9967 966 9997 971
rect 9930 962 9997 966
rect 9903 959 9997 962
rect 9903 952 9952 959
rect 9903 946 9933 952
rect 9952 947 9957 952
rect 9869 930 9949 946
rect 9961 938 9997 959
rect 10058 954 10247 978
rect 10292 977 10339 978
rect 10305 972 10339 977
rect 10073 951 10247 954
rect 10066 948 10247 951
rect 10275 971 10339 972
rect 9869 928 9888 930
rect 9903 928 9937 930
rect 9869 912 9949 928
rect 9869 906 9888 912
rect 9585 880 9688 890
rect 9539 878 9688 880
rect 9709 878 9744 890
rect 9378 876 9540 878
rect 9390 856 9409 876
rect 9424 874 9454 876
rect 9273 848 9314 856
rect 9396 852 9409 856
rect 9461 860 9540 876
rect 9572 876 9744 878
rect 9572 860 9651 876
rect 9658 874 9688 876
rect 9236 838 9265 848
rect 9279 838 9308 848
rect 9323 838 9353 852
rect 9396 838 9439 852
rect 9461 848 9651 860
rect 9716 856 9722 876
rect 9446 838 9476 848
rect 9477 838 9635 848
rect 9639 838 9669 848
rect 9673 838 9703 852
rect 9731 838 9744 876
rect 9816 890 9845 906
rect 9859 890 9888 906
rect 9903 896 9933 912
rect 9961 890 9967 938
rect 9970 932 9989 938
rect 10004 932 10034 940
rect 9970 924 10034 932
rect 9970 908 10050 924
rect 10066 917 10128 948
rect 10144 917 10206 948
rect 10275 946 10324 971
rect 10339 946 10369 962
rect 10238 932 10268 940
rect 10275 938 10385 946
rect 10238 924 10283 932
rect 9970 906 9989 908
rect 10004 906 10050 908
rect 9970 890 10050 906
rect 10077 904 10112 917
rect 10153 914 10190 917
rect 10153 912 10195 914
rect 10082 901 10112 904
rect 10091 897 10098 901
rect 10098 896 10099 897
rect 10057 890 10067 896
rect 9816 882 9851 890
rect 9816 856 9817 882
rect 9824 856 9851 882
rect 9759 838 9789 852
rect 9816 848 9851 856
rect 9853 882 9894 890
rect 9853 856 9868 882
rect 9875 856 9894 882
rect 9958 878 9989 890
rect 10004 878 10107 890
rect 10119 880 10145 906
rect 10160 901 10190 912
rect 10222 908 10284 924
rect 10222 906 10268 908
rect 10222 890 10284 906
rect 10296 890 10302 938
rect 10305 930 10385 938
rect 10305 928 10324 930
rect 10339 928 10373 930
rect 10305 912 10385 928
rect 10305 890 10324 912
rect 10339 896 10369 912
rect 10397 906 10403 980
rect 10406 906 10425 1050
rect 10440 906 10446 1050
rect 10455 980 10468 1050
rect 10520 1046 10542 1050
rect 10513 1024 10542 1038
rect 10595 1024 10611 1038
rect 10649 1034 10655 1036
rect 10662 1034 10770 1050
rect 10777 1034 10783 1036
rect 10791 1034 10806 1050
rect 10872 1044 10891 1047
rect 10513 1022 10611 1024
rect 10638 1022 10806 1034
rect 10821 1024 10837 1038
rect 10872 1025 10894 1044
rect 10904 1038 10920 1039
rect 10903 1036 10920 1038
rect 10904 1031 10920 1036
rect 10894 1024 10900 1025
rect 10903 1024 10932 1031
rect 10821 1023 10932 1024
rect 10821 1022 10938 1023
rect 10497 1014 10548 1022
rect 10595 1014 10629 1022
rect 10497 1002 10522 1014
rect 10529 1002 10548 1014
rect 10602 1012 10629 1014
rect 10638 1012 10859 1022
rect 10894 1019 10900 1022
rect 10602 1008 10859 1012
rect 10497 994 10548 1002
rect 10595 994 10859 1008
rect 10903 1014 10938 1022
rect 10449 946 10468 980
rect 10513 986 10542 994
rect 10513 980 10530 986
rect 10513 978 10547 980
rect 10595 978 10611 994
rect 10612 984 10820 994
rect 10821 984 10837 994
rect 10885 990 10900 1005
rect 10903 1002 10904 1014
rect 10911 1002 10938 1014
rect 10903 994 10938 1002
rect 10903 993 10932 994
rect 10623 980 10837 984
rect 10638 978 10837 980
rect 10872 980 10885 990
rect 10903 980 10920 993
rect 10872 978 10920 980
rect 10514 974 10547 978
rect 10510 972 10547 974
rect 10510 971 10577 972
rect 10510 966 10541 971
rect 10547 966 10577 971
rect 10510 962 10577 966
rect 10483 959 10577 962
rect 10483 952 10532 959
rect 10483 946 10513 952
rect 10532 947 10537 952
rect 10449 930 10529 946
rect 10541 938 10577 959
rect 10638 954 10827 978
rect 10872 977 10919 978
rect 10885 972 10919 977
rect 10653 951 10827 954
rect 10646 948 10827 951
rect 10855 971 10919 972
rect 10449 928 10468 930
rect 10483 928 10517 930
rect 10449 912 10529 928
rect 10449 906 10468 912
rect 10165 880 10268 890
rect 10119 878 10268 880
rect 10289 878 10324 890
rect 9958 876 10120 878
rect 9970 856 9989 876
rect 10004 874 10034 876
rect 9853 848 9894 856
rect 9976 852 9989 856
rect 10041 860 10120 876
rect 10152 876 10324 878
rect 10152 860 10231 876
rect 10238 874 10268 876
rect 9816 838 9845 848
rect 9859 838 9888 848
rect 9903 838 9933 852
rect 9976 838 10019 852
rect 10041 848 10231 860
rect 10296 856 10302 876
rect 10026 838 10056 848
rect 10057 838 10215 848
rect 10219 838 10249 848
rect 10253 838 10283 852
rect 10311 838 10324 876
rect 10396 890 10425 906
rect 10439 890 10468 906
rect 10483 896 10513 912
rect 10541 890 10547 938
rect 10550 932 10569 938
rect 10584 932 10614 940
rect 10550 924 10614 932
rect 10550 908 10630 924
rect 10646 917 10708 948
rect 10724 917 10786 948
rect 10855 946 10904 971
rect 10919 946 10949 962
rect 10818 932 10848 940
rect 10855 938 10965 946
rect 10818 924 10863 932
rect 10550 906 10569 908
rect 10584 906 10630 908
rect 10550 890 10630 906
rect 10657 904 10692 917
rect 10733 914 10770 917
rect 10733 912 10775 914
rect 10662 901 10692 904
rect 10671 897 10678 901
rect 10678 896 10679 897
rect 10637 890 10647 896
rect 10396 882 10431 890
rect 10396 856 10397 882
rect 10404 856 10431 882
rect 10339 838 10369 852
rect 10396 848 10431 856
rect 10433 882 10474 890
rect 10433 856 10448 882
rect 10455 856 10474 882
rect 10538 878 10569 890
rect 10584 878 10687 890
rect 10699 880 10725 906
rect 10740 901 10770 912
rect 10802 908 10864 924
rect 10802 906 10848 908
rect 10802 890 10864 906
rect 10876 890 10882 938
rect 10885 930 10965 938
rect 10885 928 10904 930
rect 10919 928 10953 930
rect 10885 912 10965 928
rect 10885 890 10904 912
rect 10919 896 10949 912
rect 10977 906 10983 980
rect 10986 906 11005 1050
rect 11020 906 11026 1050
rect 11035 980 11048 1050
rect 11100 1046 11122 1050
rect 11093 1024 11122 1038
rect 11175 1024 11191 1038
rect 11229 1034 11235 1036
rect 11242 1034 11350 1050
rect 11357 1034 11363 1036
rect 11371 1034 11386 1050
rect 11452 1044 11471 1047
rect 11093 1022 11191 1024
rect 11218 1022 11386 1034
rect 11401 1024 11417 1038
rect 11452 1025 11474 1044
rect 11484 1038 11500 1039
rect 11483 1036 11500 1038
rect 11484 1031 11500 1036
rect 11474 1024 11480 1025
rect 11483 1024 11512 1031
rect 11401 1023 11512 1024
rect 11401 1022 11518 1023
rect 11077 1014 11128 1022
rect 11175 1014 11209 1022
rect 11077 1002 11102 1014
rect 11109 1002 11128 1014
rect 11182 1012 11209 1014
rect 11218 1012 11439 1022
rect 11474 1019 11480 1022
rect 11182 1008 11439 1012
rect 11077 994 11128 1002
rect 11175 994 11439 1008
rect 11483 1014 11518 1022
rect 11029 946 11048 980
rect 11093 986 11122 994
rect 11093 980 11110 986
rect 11093 978 11127 980
rect 11175 978 11191 994
rect 11192 984 11400 994
rect 11401 984 11417 994
rect 11465 990 11480 1005
rect 11483 1002 11484 1014
rect 11491 1002 11518 1014
rect 11483 994 11518 1002
rect 11483 993 11512 994
rect 11203 980 11417 984
rect 11218 978 11417 980
rect 11452 980 11465 990
rect 11483 980 11500 993
rect 11452 978 11500 980
rect 11094 974 11127 978
rect 11090 972 11127 974
rect 11090 971 11157 972
rect 11090 966 11121 971
rect 11127 966 11157 971
rect 11090 962 11157 966
rect 11063 959 11157 962
rect 11063 952 11112 959
rect 11063 946 11093 952
rect 11112 947 11117 952
rect 11029 930 11109 946
rect 11121 938 11157 959
rect 11218 954 11407 978
rect 11452 977 11499 978
rect 11465 972 11499 977
rect 11233 951 11407 954
rect 11226 948 11407 951
rect 11435 971 11499 972
rect 11029 928 11048 930
rect 11063 928 11097 930
rect 11029 912 11109 928
rect 11029 906 11048 912
rect 10745 880 10848 890
rect 10699 878 10848 880
rect 10869 878 10904 890
rect 10538 876 10700 878
rect 10550 856 10569 876
rect 10584 874 10614 876
rect 10433 848 10474 856
rect 10556 852 10569 856
rect 10621 860 10700 876
rect 10732 876 10904 878
rect 10732 860 10811 876
rect 10818 874 10848 876
rect 10396 838 10425 848
rect 10439 838 10468 848
rect 10483 838 10513 852
rect 10556 838 10599 852
rect 10621 848 10811 860
rect 10876 856 10882 876
rect 10606 838 10636 848
rect 10637 838 10795 848
rect 10799 838 10829 848
rect 10833 838 10863 852
rect 10891 838 10904 876
rect 10976 890 11005 906
rect 11019 890 11048 906
rect 11063 896 11093 912
rect 11121 890 11127 938
rect 11130 932 11149 938
rect 11164 932 11194 940
rect 11130 924 11194 932
rect 11130 908 11210 924
rect 11226 917 11288 948
rect 11304 917 11366 948
rect 11435 946 11484 971
rect 11499 946 11529 962
rect 11398 932 11428 940
rect 11435 938 11545 946
rect 11398 924 11443 932
rect 11130 906 11149 908
rect 11164 906 11210 908
rect 11130 890 11210 906
rect 11237 904 11272 917
rect 11313 914 11350 917
rect 11313 912 11355 914
rect 11242 901 11272 904
rect 11251 897 11258 901
rect 11258 896 11259 897
rect 11217 890 11227 896
rect 10976 882 11011 890
rect 10976 856 10977 882
rect 10984 856 11011 882
rect 10919 838 10949 852
rect 10976 848 11011 856
rect 11013 882 11054 890
rect 11013 856 11028 882
rect 11035 856 11054 882
rect 11118 878 11149 890
rect 11164 878 11267 890
rect 11279 880 11305 906
rect 11320 901 11350 912
rect 11382 908 11444 924
rect 11382 906 11428 908
rect 11382 890 11444 906
rect 11456 890 11462 938
rect 11465 930 11545 938
rect 11465 928 11484 930
rect 11499 928 11533 930
rect 11465 912 11545 928
rect 11465 890 11484 912
rect 11499 896 11529 912
rect 11557 906 11563 980
rect 11566 906 11585 1050
rect 11600 906 11606 1050
rect 11615 980 11628 1050
rect 11680 1046 11702 1050
rect 11673 1024 11702 1038
rect 11755 1024 11771 1038
rect 11809 1034 11815 1036
rect 11822 1034 11930 1050
rect 11937 1034 11943 1036
rect 11951 1034 11966 1050
rect 12032 1044 12051 1047
rect 11673 1022 11771 1024
rect 11798 1022 11966 1034
rect 11981 1024 11997 1038
rect 12032 1025 12054 1044
rect 12064 1038 12080 1039
rect 12063 1036 12080 1038
rect 12064 1031 12080 1036
rect 12054 1024 12060 1025
rect 12063 1024 12092 1031
rect 11981 1023 12092 1024
rect 11981 1022 12098 1023
rect 11657 1014 11708 1022
rect 11755 1014 11789 1022
rect 11657 1002 11682 1014
rect 11689 1002 11708 1014
rect 11762 1012 11789 1014
rect 11798 1012 12019 1022
rect 12054 1019 12060 1022
rect 11762 1008 12019 1012
rect 11657 994 11708 1002
rect 11755 994 12019 1008
rect 12063 1014 12098 1022
rect 11609 946 11628 980
rect 11673 986 11702 994
rect 11673 980 11690 986
rect 11673 978 11707 980
rect 11755 978 11771 994
rect 11772 984 11980 994
rect 11981 984 11997 994
rect 12045 990 12060 1005
rect 12063 1002 12064 1014
rect 12071 1002 12098 1014
rect 12063 994 12098 1002
rect 12063 993 12092 994
rect 11783 980 11997 984
rect 11798 978 11997 980
rect 12032 980 12045 990
rect 12063 980 12080 993
rect 12032 978 12080 980
rect 11674 974 11707 978
rect 11670 972 11707 974
rect 11670 971 11737 972
rect 11670 966 11701 971
rect 11707 966 11737 971
rect 11670 962 11737 966
rect 11643 959 11737 962
rect 11643 952 11692 959
rect 11643 946 11673 952
rect 11692 947 11697 952
rect 11609 930 11689 946
rect 11701 938 11737 959
rect 11798 954 11987 978
rect 12032 977 12079 978
rect 12045 972 12079 977
rect 11813 951 11987 954
rect 11806 948 11987 951
rect 12015 971 12079 972
rect 11609 928 11628 930
rect 11643 928 11677 930
rect 11609 912 11689 928
rect 11609 906 11628 912
rect 11325 880 11428 890
rect 11279 878 11428 880
rect 11449 878 11484 890
rect 11118 876 11280 878
rect 11130 856 11149 876
rect 11164 874 11194 876
rect 11013 848 11054 856
rect 11136 852 11149 856
rect 11201 860 11280 876
rect 11312 876 11484 878
rect 11312 860 11391 876
rect 11398 874 11428 876
rect 10976 838 11005 848
rect 11019 838 11048 848
rect 11063 838 11093 852
rect 11136 838 11179 852
rect 11201 848 11391 860
rect 11456 856 11462 876
rect 11186 838 11216 848
rect 11217 838 11375 848
rect 11379 838 11409 848
rect 11413 838 11443 852
rect 11471 838 11484 876
rect 11556 890 11585 906
rect 11599 890 11628 906
rect 11643 896 11673 912
rect 11701 890 11707 938
rect 11710 932 11729 938
rect 11744 932 11774 940
rect 11710 924 11774 932
rect 11710 908 11790 924
rect 11806 917 11868 948
rect 11884 917 11946 948
rect 12015 946 12064 971
rect 12079 946 12109 962
rect 11978 932 12008 940
rect 12015 938 12125 946
rect 11978 924 12023 932
rect 11710 906 11729 908
rect 11744 906 11790 908
rect 11710 890 11790 906
rect 11817 904 11852 917
rect 11893 914 11930 917
rect 11893 912 11935 914
rect 11822 901 11852 904
rect 11831 897 11838 901
rect 11838 896 11839 897
rect 11797 890 11807 896
rect 11556 882 11591 890
rect 11556 856 11557 882
rect 11564 856 11591 882
rect 11499 838 11529 852
rect 11556 848 11591 856
rect 11593 882 11634 890
rect 11593 856 11608 882
rect 11615 856 11634 882
rect 11698 878 11729 890
rect 11744 878 11847 890
rect 11859 880 11885 906
rect 11900 901 11930 912
rect 11962 908 12024 924
rect 11962 906 12008 908
rect 11962 890 12024 906
rect 12036 890 12042 938
rect 12045 930 12125 938
rect 12045 928 12064 930
rect 12079 928 12113 930
rect 12045 912 12125 928
rect 12045 890 12064 912
rect 12079 896 12109 912
rect 12137 906 12143 980
rect 12146 906 12165 1050
rect 12180 906 12186 1050
rect 12195 980 12208 1050
rect 12260 1046 12282 1050
rect 12253 1024 12282 1038
rect 12335 1024 12351 1038
rect 12389 1034 12395 1036
rect 12402 1034 12510 1050
rect 12517 1034 12523 1036
rect 12531 1034 12546 1050
rect 12612 1044 12631 1047
rect 12253 1022 12351 1024
rect 12378 1022 12546 1034
rect 12561 1024 12577 1038
rect 12612 1025 12634 1044
rect 12644 1038 12660 1039
rect 12643 1036 12660 1038
rect 12644 1031 12660 1036
rect 12634 1024 12640 1025
rect 12643 1024 12672 1031
rect 12561 1023 12672 1024
rect 12561 1022 12678 1023
rect 12237 1014 12288 1022
rect 12335 1014 12369 1022
rect 12237 1002 12262 1014
rect 12269 1002 12288 1014
rect 12342 1012 12369 1014
rect 12378 1012 12599 1022
rect 12634 1019 12640 1022
rect 12342 1008 12599 1012
rect 12237 994 12288 1002
rect 12335 994 12599 1008
rect 12643 1014 12678 1022
rect 12189 946 12208 980
rect 12253 986 12282 994
rect 12253 980 12270 986
rect 12253 978 12287 980
rect 12335 978 12351 994
rect 12352 984 12560 994
rect 12561 984 12577 994
rect 12625 990 12640 1005
rect 12643 1002 12644 1014
rect 12651 1002 12678 1014
rect 12643 994 12678 1002
rect 12643 993 12672 994
rect 12363 980 12577 984
rect 12378 978 12577 980
rect 12612 980 12625 990
rect 12643 980 12660 993
rect 12612 978 12660 980
rect 12254 974 12287 978
rect 12250 972 12287 974
rect 12250 971 12317 972
rect 12250 966 12281 971
rect 12287 966 12317 971
rect 12250 962 12317 966
rect 12223 959 12317 962
rect 12223 952 12272 959
rect 12223 946 12253 952
rect 12272 947 12277 952
rect 12189 930 12269 946
rect 12281 938 12317 959
rect 12378 954 12567 978
rect 12612 977 12659 978
rect 12625 972 12659 977
rect 12393 951 12567 954
rect 12386 948 12567 951
rect 12595 971 12659 972
rect 12189 928 12208 930
rect 12223 928 12257 930
rect 12189 912 12269 928
rect 12189 906 12208 912
rect 11905 880 12008 890
rect 11859 878 12008 880
rect 12029 878 12064 890
rect 11698 876 11860 878
rect 11710 856 11729 876
rect 11744 874 11774 876
rect 11593 848 11634 856
rect 11716 852 11729 856
rect 11781 860 11860 876
rect 11892 876 12064 878
rect 11892 860 11971 876
rect 11978 874 12008 876
rect 11556 838 11585 848
rect 11599 838 11628 848
rect 11643 838 11673 852
rect 11716 838 11759 852
rect 11781 848 11971 860
rect 12036 856 12042 876
rect 11766 838 11796 848
rect 11797 838 11955 848
rect 11959 838 11989 848
rect 11993 838 12023 852
rect 12051 838 12064 876
rect 12136 890 12165 906
rect 12179 890 12208 906
rect 12223 896 12253 912
rect 12281 890 12287 938
rect 12290 932 12309 938
rect 12324 932 12354 940
rect 12290 924 12354 932
rect 12290 908 12370 924
rect 12386 917 12448 948
rect 12464 917 12526 948
rect 12595 946 12644 971
rect 12659 946 12689 962
rect 12558 932 12588 940
rect 12595 938 12705 946
rect 12558 924 12603 932
rect 12290 906 12309 908
rect 12324 906 12370 908
rect 12290 890 12370 906
rect 12397 904 12432 917
rect 12473 914 12510 917
rect 12473 912 12515 914
rect 12402 901 12432 904
rect 12411 897 12418 901
rect 12418 896 12419 897
rect 12377 890 12387 896
rect 12136 882 12171 890
rect 12136 856 12137 882
rect 12144 856 12171 882
rect 12079 838 12109 852
rect 12136 848 12171 856
rect 12173 882 12214 890
rect 12173 856 12188 882
rect 12195 856 12214 882
rect 12278 878 12309 890
rect 12324 878 12427 890
rect 12439 880 12465 906
rect 12480 901 12510 912
rect 12542 908 12604 924
rect 12542 906 12588 908
rect 12542 890 12604 906
rect 12616 890 12622 938
rect 12625 930 12705 938
rect 12625 928 12644 930
rect 12659 928 12693 930
rect 12625 912 12705 928
rect 12625 890 12644 912
rect 12659 896 12689 912
rect 12717 906 12723 980
rect 12726 906 12745 1050
rect 12760 906 12766 1050
rect 12775 980 12788 1050
rect 12840 1046 12862 1050
rect 12833 1024 12862 1038
rect 12915 1024 12931 1038
rect 12969 1034 12975 1036
rect 12982 1034 13090 1050
rect 13097 1034 13103 1036
rect 13111 1034 13126 1050
rect 13192 1044 13211 1047
rect 12833 1022 12931 1024
rect 12958 1022 13126 1034
rect 13141 1024 13157 1038
rect 13192 1025 13214 1044
rect 13224 1038 13240 1039
rect 13223 1036 13240 1038
rect 13224 1031 13240 1036
rect 13214 1024 13220 1025
rect 13223 1024 13252 1031
rect 13141 1023 13252 1024
rect 13141 1022 13258 1023
rect 12817 1014 12868 1022
rect 12915 1014 12949 1022
rect 12817 1002 12842 1014
rect 12849 1002 12868 1014
rect 12922 1012 12949 1014
rect 12958 1012 13179 1022
rect 13214 1019 13220 1022
rect 12922 1008 13179 1012
rect 12817 994 12868 1002
rect 12915 994 13179 1008
rect 13223 1014 13258 1022
rect 12769 946 12788 980
rect 12833 986 12862 994
rect 12833 980 12850 986
rect 12833 978 12867 980
rect 12915 978 12931 994
rect 12932 984 13140 994
rect 13141 984 13157 994
rect 13205 990 13220 1005
rect 13223 1002 13224 1014
rect 13231 1002 13258 1014
rect 13223 994 13258 1002
rect 13223 993 13252 994
rect 12943 980 13157 984
rect 12958 978 13157 980
rect 13192 980 13205 990
rect 13223 980 13240 993
rect 13192 978 13240 980
rect 12834 974 12867 978
rect 12830 972 12867 974
rect 12830 971 12897 972
rect 12830 966 12861 971
rect 12867 966 12897 971
rect 12830 962 12897 966
rect 12803 959 12897 962
rect 12803 952 12852 959
rect 12803 946 12833 952
rect 12852 947 12857 952
rect 12769 930 12849 946
rect 12861 938 12897 959
rect 12958 954 13147 978
rect 13192 977 13239 978
rect 13205 972 13239 977
rect 12973 951 13147 954
rect 12966 948 13147 951
rect 13175 971 13239 972
rect 12769 928 12788 930
rect 12803 928 12837 930
rect 12769 912 12849 928
rect 12769 906 12788 912
rect 12485 880 12588 890
rect 12439 878 12588 880
rect 12609 878 12644 890
rect 12278 876 12440 878
rect 12290 856 12309 876
rect 12324 874 12354 876
rect 12173 848 12214 856
rect 12296 852 12309 856
rect 12361 860 12440 876
rect 12472 876 12644 878
rect 12472 860 12551 876
rect 12558 874 12588 876
rect 12136 838 12165 848
rect 12179 838 12208 848
rect 12223 838 12253 852
rect 12296 838 12339 852
rect 12361 848 12551 860
rect 12616 856 12622 876
rect 12346 838 12376 848
rect 12377 838 12535 848
rect 12539 838 12569 848
rect 12573 838 12603 852
rect 12631 838 12644 876
rect 12716 890 12745 906
rect 12759 890 12788 906
rect 12803 896 12833 912
rect 12861 890 12867 938
rect 12870 932 12889 938
rect 12904 932 12934 940
rect 12870 924 12934 932
rect 12870 908 12950 924
rect 12966 917 13028 948
rect 13044 917 13106 948
rect 13175 946 13224 971
rect 13239 946 13269 962
rect 13138 932 13168 940
rect 13175 938 13285 946
rect 13138 924 13183 932
rect 12870 906 12889 908
rect 12904 906 12950 908
rect 12870 890 12950 906
rect 12977 904 13012 917
rect 13053 914 13090 917
rect 13053 912 13095 914
rect 12982 901 13012 904
rect 12991 897 12998 901
rect 12998 896 12999 897
rect 12957 890 12967 896
rect 12716 882 12751 890
rect 12716 856 12717 882
rect 12724 856 12751 882
rect 12659 838 12689 852
rect 12716 848 12751 856
rect 12753 882 12794 890
rect 12753 856 12768 882
rect 12775 856 12794 882
rect 12858 878 12889 890
rect 12904 878 13007 890
rect 13019 880 13045 906
rect 13060 901 13090 912
rect 13122 908 13184 924
rect 13122 906 13168 908
rect 13122 890 13184 906
rect 13196 890 13202 938
rect 13205 930 13285 938
rect 13205 928 13224 930
rect 13239 928 13273 930
rect 13205 912 13285 928
rect 13205 890 13224 912
rect 13239 896 13269 912
rect 13297 906 13303 980
rect 13306 906 13325 1050
rect 13340 906 13346 1050
rect 13355 980 13368 1050
rect 13420 1046 13442 1050
rect 13413 1024 13442 1038
rect 13495 1024 13511 1038
rect 13549 1034 13555 1036
rect 13562 1034 13670 1050
rect 13677 1034 13683 1036
rect 13691 1034 13706 1050
rect 13772 1044 13791 1047
rect 13413 1022 13511 1024
rect 13538 1022 13706 1034
rect 13721 1024 13737 1038
rect 13772 1025 13794 1044
rect 13804 1038 13820 1039
rect 13803 1036 13820 1038
rect 13804 1031 13820 1036
rect 13794 1024 13800 1025
rect 13803 1024 13832 1031
rect 13721 1023 13832 1024
rect 13721 1022 13838 1023
rect 13397 1014 13448 1022
rect 13495 1014 13529 1022
rect 13397 1002 13422 1014
rect 13429 1002 13448 1014
rect 13502 1012 13529 1014
rect 13538 1012 13759 1022
rect 13794 1019 13800 1022
rect 13502 1008 13759 1012
rect 13397 994 13448 1002
rect 13495 994 13759 1008
rect 13803 1014 13838 1022
rect 13349 946 13368 980
rect 13413 986 13442 994
rect 13413 980 13430 986
rect 13413 978 13447 980
rect 13495 978 13511 994
rect 13512 984 13720 994
rect 13721 984 13737 994
rect 13785 990 13800 1005
rect 13803 1002 13804 1014
rect 13811 1002 13838 1014
rect 13803 994 13838 1002
rect 13803 993 13832 994
rect 13523 980 13737 984
rect 13538 978 13737 980
rect 13772 980 13785 990
rect 13803 980 13820 993
rect 13772 978 13820 980
rect 13414 974 13447 978
rect 13410 972 13447 974
rect 13410 971 13477 972
rect 13410 966 13441 971
rect 13447 966 13477 971
rect 13410 962 13477 966
rect 13383 959 13477 962
rect 13383 952 13432 959
rect 13383 946 13413 952
rect 13432 947 13437 952
rect 13349 930 13429 946
rect 13441 938 13477 959
rect 13538 954 13727 978
rect 13772 977 13819 978
rect 13785 972 13819 977
rect 13553 951 13727 954
rect 13546 948 13727 951
rect 13755 971 13819 972
rect 13349 928 13368 930
rect 13383 928 13417 930
rect 13349 912 13429 928
rect 13349 906 13368 912
rect 13065 880 13168 890
rect 13019 878 13168 880
rect 13189 878 13224 890
rect 12858 876 13020 878
rect 12870 856 12889 876
rect 12904 874 12934 876
rect 12753 848 12794 856
rect 12876 852 12889 856
rect 12941 860 13020 876
rect 13052 876 13224 878
rect 13052 860 13131 876
rect 13138 874 13168 876
rect 12716 838 12745 848
rect 12759 838 12788 848
rect 12803 838 12833 852
rect 12876 838 12919 852
rect 12941 848 13131 860
rect 13196 856 13202 876
rect 12926 838 12956 848
rect 12957 838 13115 848
rect 13119 838 13149 848
rect 13153 838 13183 852
rect 13211 838 13224 876
rect 13296 890 13325 906
rect 13339 890 13368 906
rect 13383 896 13413 912
rect 13441 890 13447 938
rect 13450 932 13469 938
rect 13484 932 13514 940
rect 13450 924 13514 932
rect 13450 908 13530 924
rect 13546 917 13608 948
rect 13624 917 13686 948
rect 13755 946 13804 971
rect 13819 946 13849 962
rect 13718 932 13748 940
rect 13755 938 13865 946
rect 13718 924 13763 932
rect 13450 906 13469 908
rect 13484 906 13530 908
rect 13450 890 13530 906
rect 13557 904 13592 917
rect 13633 914 13670 917
rect 13633 912 13675 914
rect 13562 901 13592 904
rect 13571 897 13578 901
rect 13578 896 13579 897
rect 13537 890 13547 896
rect 13296 882 13331 890
rect 13296 856 13297 882
rect 13304 856 13331 882
rect 13239 838 13269 852
rect 13296 848 13331 856
rect 13333 882 13374 890
rect 13333 856 13348 882
rect 13355 856 13374 882
rect 13438 878 13469 890
rect 13484 878 13587 890
rect 13599 880 13625 906
rect 13640 901 13670 912
rect 13702 908 13764 924
rect 13702 906 13748 908
rect 13702 890 13764 906
rect 13776 890 13782 938
rect 13785 930 13865 938
rect 13785 928 13804 930
rect 13819 928 13853 930
rect 13785 912 13865 928
rect 13785 890 13804 912
rect 13819 896 13849 912
rect 13877 906 13883 980
rect 13886 906 13905 1050
rect 13920 906 13926 1050
rect 13935 980 13948 1050
rect 14000 1046 14022 1050
rect 13993 1024 14022 1038
rect 14075 1024 14091 1038
rect 14129 1034 14135 1036
rect 14142 1034 14250 1050
rect 14257 1034 14263 1036
rect 14271 1034 14286 1050
rect 14352 1044 14371 1047
rect 13993 1022 14091 1024
rect 14118 1022 14286 1034
rect 14301 1024 14317 1038
rect 14352 1025 14374 1044
rect 14384 1038 14400 1039
rect 14383 1036 14400 1038
rect 14384 1031 14400 1036
rect 14374 1024 14380 1025
rect 14383 1024 14412 1031
rect 14301 1023 14412 1024
rect 14301 1022 14418 1023
rect 13977 1014 14028 1022
rect 14075 1014 14109 1022
rect 13977 1002 14002 1014
rect 14009 1002 14028 1014
rect 14082 1012 14109 1014
rect 14118 1012 14339 1022
rect 14374 1019 14380 1022
rect 14082 1008 14339 1012
rect 13977 994 14028 1002
rect 14075 994 14339 1008
rect 14383 1014 14418 1022
rect 13929 946 13948 980
rect 13993 986 14022 994
rect 13993 980 14010 986
rect 13993 978 14027 980
rect 14075 978 14091 994
rect 14092 984 14300 994
rect 14301 984 14317 994
rect 14365 990 14380 1005
rect 14383 1002 14384 1014
rect 14391 1002 14418 1014
rect 14383 994 14418 1002
rect 14383 993 14412 994
rect 14103 980 14317 984
rect 14118 978 14317 980
rect 14352 980 14365 990
rect 14383 980 14400 993
rect 14352 978 14400 980
rect 13994 974 14027 978
rect 13990 972 14027 974
rect 13990 971 14057 972
rect 13990 966 14021 971
rect 14027 966 14057 971
rect 13990 962 14057 966
rect 13963 959 14057 962
rect 13963 952 14012 959
rect 13963 946 13993 952
rect 14012 947 14017 952
rect 13929 930 14009 946
rect 14021 938 14057 959
rect 14118 954 14307 978
rect 14352 977 14399 978
rect 14365 972 14399 977
rect 14133 951 14307 954
rect 14126 948 14307 951
rect 14335 971 14399 972
rect 13929 928 13948 930
rect 13963 928 13997 930
rect 13929 912 14009 928
rect 13929 906 13948 912
rect 13645 880 13748 890
rect 13599 878 13748 880
rect 13769 878 13804 890
rect 13438 876 13600 878
rect 13450 856 13469 876
rect 13484 874 13514 876
rect 13333 848 13374 856
rect 13456 852 13469 856
rect 13521 860 13600 876
rect 13632 876 13804 878
rect 13632 860 13711 876
rect 13718 874 13748 876
rect 13296 838 13325 848
rect 13339 838 13368 848
rect 13383 838 13413 852
rect 13456 838 13499 852
rect 13521 848 13711 860
rect 13776 856 13782 876
rect 13506 838 13536 848
rect 13537 838 13695 848
rect 13699 838 13729 848
rect 13733 838 13763 852
rect 13791 838 13804 876
rect 13876 890 13905 906
rect 13919 890 13948 906
rect 13963 896 13993 912
rect 14021 890 14027 938
rect 14030 932 14049 938
rect 14064 932 14094 940
rect 14030 924 14094 932
rect 14030 908 14110 924
rect 14126 917 14188 948
rect 14204 917 14266 948
rect 14335 946 14384 971
rect 14399 946 14429 962
rect 14298 932 14328 940
rect 14335 938 14445 946
rect 14298 924 14343 932
rect 14030 906 14049 908
rect 14064 906 14110 908
rect 14030 890 14110 906
rect 14137 904 14172 917
rect 14213 914 14250 917
rect 14213 912 14255 914
rect 14142 901 14172 904
rect 14151 897 14158 901
rect 14158 896 14159 897
rect 14117 890 14127 896
rect 13876 882 13911 890
rect 13876 856 13877 882
rect 13884 856 13911 882
rect 13819 838 13849 852
rect 13876 848 13911 856
rect 13913 882 13954 890
rect 13913 856 13928 882
rect 13935 856 13954 882
rect 14018 878 14049 890
rect 14064 878 14167 890
rect 14179 880 14205 906
rect 14220 901 14250 912
rect 14282 908 14344 924
rect 14282 906 14328 908
rect 14282 890 14344 906
rect 14356 890 14362 938
rect 14365 930 14445 938
rect 14365 928 14384 930
rect 14399 928 14433 930
rect 14365 912 14445 928
rect 14365 890 14384 912
rect 14399 896 14429 912
rect 14457 906 14463 980
rect 14466 906 14485 1050
rect 14500 906 14506 1050
rect 14515 980 14528 1050
rect 14580 1046 14602 1050
rect 14573 1024 14602 1038
rect 14655 1024 14671 1038
rect 14709 1034 14715 1036
rect 14722 1034 14830 1050
rect 14837 1034 14843 1036
rect 14851 1034 14866 1050
rect 14932 1044 14951 1047
rect 14573 1022 14671 1024
rect 14698 1022 14866 1034
rect 14881 1024 14897 1038
rect 14932 1025 14954 1044
rect 14964 1038 14980 1039
rect 14963 1036 14980 1038
rect 14964 1031 14980 1036
rect 14954 1024 14960 1025
rect 14963 1024 14992 1031
rect 14881 1023 14992 1024
rect 14881 1022 14998 1023
rect 14557 1014 14608 1022
rect 14655 1014 14689 1022
rect 14557 1002 14582 1014
rect 14589 1002 14608 1014
rect 14662 1012 14689 1014
rect 14698 1012 14919 1022
rect 14954 1019 14960 1022
rect 14662 1008 14919 1012
rect 14557 994 14608 1002
rect 14655 994 14919 1008
rect 14963 1014 14998 1022
rect 14509 946 14528 980
rect 14573 986 14602 994
rect 14573 980 14590 986
rect 14573 978 14607 980
rect 14655 978 14671 994
rect 14672 984 14880 994
rect 14881 984 14897 994
rect 14945 990 14960 1005
rect 14963 1002 14964 1014
rect 14971 1002 14998 1014
rect 14963 994 14998 1002
rect 14963 993 14992 994
rect 14683 980 14897 984
rect 14698 978 14897 980
rect 14932 980 14945 990
rect 14963 980 14980 993
rect 14932 978 14980 980
rect 14574 974 14607 978
rect 14570 972 14607 974
rect 14570 971 14637 972
rect 14570 966 14601 971
rect 14607 966 14637 971
rect 14570 962 14637 966
rect 14543 959 14637 962
rect 14543 952 14592 959
rect 14543 946 14573 952
rect 14592 947 14597 952
rect 14509 930 14589 946
rect 14601 938 14637 959
rect 14698 954 14887 978
rect 14932 977 14979 978
rect 14945 972 14979 977
rect 14713 951 14887 954
rect 14706 948 14887 951
rect 14915 971 14979 972
rect 14509 928 14528 930
rect 14543 928 14577 930
rect 14509 912 14589 928
rect 14509 906 14528 912
rect 14225 880 14328 890
rect 14179 878 14328 880
rect 14349 878 14384 890
rect 14018 876 14180 878
rect 14030 856 14049 876
rect 14064 874 14094 876
rect 13913 848 13954 856
rect 14036 852 14049 856
rect 14101 860 14180 876
rect 14212 876 14384 878
rect 14212 860 14291 876
rect 14298 874 14328 876
rect 13876 838 13905 848
rect 13919 838 13948 848
rect 13963 838 13993 852
rect 14036 838 14079 852
rect 14101 848 14291 860
rect 14356 856 14362 876
rect 14086 838 14116 848
rect 14117 838 14275 848
rect 14279 838 14309 848
rect 14313 838 14343 852
rect 14371 838 14384 876
rect 14456 890 14485 906
rect 14499 890 14528 906
rect 14543 896 14573 912
rect 14601 890 14607 938
rect 14610 932 14629 938
rect 14644 932 14674 940
rect 14610 924 14674 932
rect 14610 908 14690 924
rect 14706 917 14768 948
rect 14784 917 14846 948
rect 14915 946 14964 971
rect 14979 946 15009 962
rect 14878 932 14908 940
rect 14915 938 15025 946
rect 14878 924 14923 932
rect 14610 906 14629 908
rect 14644 906 14690 908
rect 14610 890 14690 906
rect 14717 904 14752 917
rect 14793 914 14830 917
rect 14793 912 14835 914
rect 14722 901 14752 904
rect 14731 897 14738 901
rect 14738 896 14739 897
rect 14697 890 14707 896
rect 14456 882 14491 890
rect 14456 856 14457 882
rect 14464 856 14491 882
rect 14399 838 14429 852
rect 14456 848 14491 856
rect 14493 882 14534 890
rect 14493 856 14508 882
rect 14515 856 14534 882
rect 14598 878 14629 890
rect 14644 878 14747 890
rect 14759 880 14785 906
rect 14800 901 14830 912
rect 14862 908 14924 924
rect 14862 906 14908 908
rect 14862 890 14924 906
rect 14936 890 14942 938
rect 14945 930 15025 938
rect 14945 928 14964 930
rect 14979 928 15013 930
rect 14945 912 15025 928
rect 14945 890 14964 912
rect 14979 896 15009 912
rect 15037 906 15043 980
rect 15046 906 15065 1050
rect 15080 906 15086 1050
rect 15095 980 15108 1050
rect 15160 1046 15182 1050
rect 15153 1024 15182 1038
rect 15235 1024 15251 1038
rect 15289 1034 15295 1036
rect 15302 1034 15410 1050
rect 15417 1034 15423 1036
rect 15431 1034 15446 1050
rect 15512 1044 15531 1047
rect 15153 1022 15251 1024
rect 15278 1022 15446 1034
rect 15461 1024 15477 1038
rect 15512 1025 15534 1044
rect 15544 1038 15560 1039
rect 15543 1036 15560 1038
rect 15544 1031 15560 1036
rect 15534 1024 15540 1025
rect 15543 1024 15572 1031
rect 15461 1023 15572 1024
rect 15461 1022 15578 1023
rect 15137 1014 15188 1022
rect 15235 1014 15269 1022
rect 15137 1002 15162 1014
rect 15169 1002 15188 1014
rect 15242 1012 15269 1014
rect 15278 1012 15499 1022
rect 15534 1019 15540 1022
rect 15242 1008 15499 1012
rect 15137 994 15188 1002
rect 15235 994 15499 1008
rect 15543 1014 15578 1022
rect 15089 946 15108 980
rect 15153 986 15182 994
rect 15153 980 15170 986
rect 15153 978 15187 980
rect 15235 978 15251 994
rect 15252 984 15460 994
rect 15461 984 15477 994
rect 15525 990 15540 1005
rect 15543 1002 15544 1014
rect 15551 1002 15578 1014
rect 15543 994 15578 1002
rect 15543 993 15572 994
rect 15263 980 15477 984
rect 15278 978 15477 980
rect 15512 980 15525 990
rect 15543 980 15560 993
rect 15512 978 15560 980
rect 15154 974 15187 978
rect 15150 972 15187 974
rect 15150 971 15217 972
rect 15150 966 15181 971
rect 15187 966 15217 971
rect 15150 962 15217 966
rect 15123 959 15217 962
rect 15123 952 15172 959
rect 15123 946 15153 952
rect 15172 947 15177 952
rect 15089 930 15169 946
rect 15181 938 15217 959
rect 15278 954 15467 978
rect 15512 977 15559 978
rect 15525 972 15559 977
rect 15293 951 15467 954
rect 15286 948 15467 951
rect 15495 971 15559 972
rect 15089 928 15108 930
rect 15123 928 15157 930
rect 15089 912 15169 928
rect 15089 906 15108 912
rect 14805 880 14908 890
rect 14759 878 14908 880
rect 14929 878 14964 890
rect 14598 876 14760 878
rect 14610 856 14629 876
rect 14644 874 14674 876
rect 14493 848 14534 856
rect 14616 852 14629 856
rect 14681 860 14760 876
rect 14792 876 14964 878
rect 14792 860 14871 876
rect 14878 874 14908 876
rect 14456 838 14485 848
rect 14499 838 14528 848
rect 14543 838 14573 852
rect 14616 838 14659 852
rect 14681 848 14871 860
rect 14936 856 14942 876
rect 14666 838 14696 848
rect 14697 838 14855 848
rect 14859 838 14889 848
rect 14893 838 14923 852
rect 14951 838 14964 876
rect 15036 890 15065 906
rect 15079 890 15108 906
rect 15123 896 15153 912
rect 15181 890 15187 938
rect 15190 932 15209 938
rect 15224 932 15254 940
rect 15190 924 15254 932
rect 15190 908 15270 924
rect 15286 917 15348 948
rect 15364 917 15426 948
rect 15495 946 15544 971
rect 15559 946 15589 962
rect 15458 932 15488 940
rect 15495 938 15605 946
rect 15458 924 15503 932
rect 15190 906 15209 908
rect 15224 906 15270 908
rect 15190 890 15270 906
rect 15297 904 15332 917
rect 15373 914 15410 917
rect 15373 912 15415 914
rect 15302 901 15332 904
rect 15311 897 15318 901
rect 15318 896 15319 897
rect 15277 890 15287 896
rect 15036 882 15071 890
rect 15036 856 15037 882
rect 15044 856 15071 882
rect 14979 838 15009 852
rect 15036 848 15071 856
rect 15073 882 15114 890
rect 15073 856 15088 882
rect 15095 856 15114 882
rect 15178 878 15209 890
rect 15224 878 15327 890
rect 15339 880 15365 906
rect 15380 901 15410 912
rect 15442 908 15504 924
rect 15442 906 15488 908
rect 15442 890 15504 906
rect 15516 890 15522 938
rect 15525 930 15605 938
rect 15525 928 15544 930
rect 15559 928 15593 930
rect 15525 912 15605 928
rect 15525 890 15544 912
rect 15559 896 15589 912
rect 15617 906 15623 980
rect 15626 906 15645 1050
rect 15660 906 15666 1050
rect 15675 980 15688 1050
rect 15740 1046 15762 1050
rect 15733 1024 15762 1038
rect 15815 1024 15831 1038
rect 15869 1034 15875 1036
rect 15882 1034 15990 1050
rect 15997 1034 16003 1036
rect 16011 1034 16026 1050
rect 16092 1044 16111 1047
rect 15733 1022 15831 1024
rect 15858 1022 16026 1034
rect 16041 1024 16057 1038
rect 16092 1025 16114 1044
rect 16124 1038 16140 1039
rect 16123 1036 16140 1038
rect 16124 1031 16140 1036
rect 16114 1024 16120 1025
rect 16123 1024 16152 1031
rect 16041 1023 16152 1024
rect 16041 1022 16158 1023
rect 15717 1014 15768 1022
rect 15815 1014 15849 1022
rect 15717 1002 15742 1014
rect 15749 1002 15768 1014
rect 15822 1012 15849 1014
rect 15858 1012 16079 1022
rect 16114 1019 16120 1022
rect 15822 1008 16079 1012
rect 15717 994 15768 1002
rect 15815 994 16079 1008
rect 16123 1014 16158 1022
rect 15669 946 15688 980
rect 15733 986 15762 994
rect 15733 980 15750 986
rect 15733 978 15767 980
rect 15815 978 15831 994
rect 15832 984 16040 994
rect 16041 984 16057 994
rect 16105 990 16120 1005
rect 16123 1002 16124 1014
rect 16131 1002 16158 1014
rect 16123 994 16158 1002
rect 16123 993 16152 994
rect 15843 980 16057 984
rect 15858 978 16057 980
rect 16092 980 16105 990
rect 16123 980 16140 993
rect 16092 978 16140 980
rect 15734 974 15767 978
rect 15730 972 15767 974
rect 15730 971 15797 972
rect 15730 966 15761 971
rect 15767 966 15797 971
rect 15730 962 15797 966
rect 15703 959 15797 962
rect 15703 952 15752 959
rect 15703 946 15733 952
rect 15752 947 15757 952
rect 15669 930 15749 946
rect 15761 938 15797 959
rect 15858 954 16047 978
rect 16092 977 16139 978
rect 16105 972 16139 977
rect 15873 951 16047 954
rect 15866 948 16047 951
rect 16075 971 16139 972
rect 15669 928 15688 930
rect 15703 928 15737 930
rect 15669 912 15749 928
rect 15669 906 15688 912
rect 15385 880 15488 890
rect 15339 878 15488 880
rect 15509 878 15544 890
rect 15178 876 15340 878
rect 15190 856 15209 876
rect 15224 874 15254 876
rect 15073 848 15114 856
rect 15196 852 15209 856
rect 15261 860 15340 876
rect 15372 876 15544 878
rect 15372 860 15451 876
rect 15458 874 15488 876
rect 15036 838 15065 848
rect 15079 838 15108 848
rect 15123 838 15153 852
rect 15196 838 15239 852
rect 15261 848 15451 860
rect 15516 856 15522 876
rect 15246 838 15276 848
rect 15277 838 15435 848
rect 15439 838 15469 848
rect 15473 838 15503 852
rect 15531 838 15544 876
rect 15616 890 15645 906
rect 15659 890 15688 906
rect 15703 896 15733 912
rect 15761 890 15767 938
rect 15770 932 15789 938
rect 15804 932 15834 940
rect 15770 924 15834 932
rect 15770 908 15850 924
rect 15866 917 15928 948
rect 15944 917 16006 948
rect 16075 946 16124 971
rect 16139 946 16169 962
rect 16038 932 16068 940
rect 16075 938 16185 946
rect 16038 924 16083 932
rect 15770 906 15789 908
rect 15804 906 15850 908
rect 15770 890 15850 906
rect 15877 904 15912 917
rect 15953 914 15990 917
rect 15953 912 15995 914
rect 15882 901 15912 904
rect 15891 897 15898 901
rect 15898 896 15899 897
rect 15857 890 15867 896
rect 15616 882 15651 890
rect 15616 856 15617 882
rect 15624 856 15651 882
rect 15559 838 15589 852
rect 15616 848 15651 856
rect 15653 882 15694 890
rect 15653 856 15668 882
rect 15675 856 15694 882
rect 15758 878 15789 890
rect 15804 878 15907 890
rect 15919 880 15945 906
rect 15960 901 15990 912
rect 16022 908 16084 924
rect 16022 906 16068 908
rect 16022 890 16084 906
rect 16096 890 16102 938
rect 16105 930 16185 938
rect 16105 928 16124 930
rect 16139 928 16173 930
rect 16105 912 16185 928
rect 16105 890 16124 912
rect 16139 896 16169 912
rect 16197 906 16203 980
rect 16206 906 16225 1050
rect 16240 906 16246 1050
rect 16255 980 16268 1050
rect 16320 1046 16342 1050
rect 16313 1024 16342 1038
rect 16395 1024 16411 1038
rect 16449 1034 16455 1036
rect 16462 1034 16570 1050
rect 16577 1034 16583 1036
rect 16591 1034 16606 1050
rect 16672 1044 16691 1047
rect 16313 1022 16411 1024
rect 16438 1022 16606 1034
rect 16621 1024 16637 1038
rect 16672 1025 16694 1044
rect 16704 1038 16720 1039
rect 16703 1036 16720 1038
rect 16704 1031 16720 1036
rect 16694 1024 16700 1025
rect 16703 1024 16732 1031
rect 16621 1023 16732 1024
rect 16621 1022 16738 1023
rect 16297 1014 16348 1022
rect 16395 1014 16429 1022
rect 16297 1002 16322 1014
rect 16329 1002 16348 1014
rect 16402 1012 16429 1014
rect 16438 1012 16659 1022
rect 16694 1019 16700 1022
rect 16402 1008 16659 1012
rect 16297 994 16348 1002
rect 16395 994 16659 1008
rect 16703 1014 16738 1022
rect 16249 946 16268 980
rect 16313 986 16342 994
rect 16313 980 16330 986
rect 16313 978 16347 980
rect 16395 978 16411 994
rect 16412 984 16620 994
rect 16621 984 16637 994
rect 16685 990 16700 1005
rect 16703 1002 16704 1014
rect 16711 1002 16738 1014
rect 16703 994 16738 1002
rect 16703 993 16732 994
rect 16423 980 16637 984
rect 16438 978 16637 980
rect 16672 980 16685 990
rect 16703 980 16720 993
rect 16672 978 16720 980
rect 16314 974 16347 978
rect 16310 972 16347 974
rect 16310 971 16377 972
rect 16310 966 16341 971
rect 16347 966 16377 971
rect 16310 962 16377 966
rect 16283 959 16377 962
rect 16283 952 16332 959
rect 16283 946 16313 952
rect 16332 947 16337 952
rect 16249 930 16329 946
rect 16341 938 16377 959
rect 16438 954 16627 978
rect 16672 977 16719 978
rect 16685 972 16719 977
rect 16453 951 16627 954
rect 16446 948 16627 951
rect 16655 971 16719 972
rect 16249 928 16268 930
rect 16283 928 16317 930
rect 16249 912 16329 928
rect 16249 906 16268 912
rect 15965 880 16068 890
rect 15919 878 16068 880
rect 16089 878 16124 890
rect 15758 876 15920 878
rect 15770 856 15789 876
rect 15804 874 15834 876
rect 15653 848 15694 856
rect 15776 852 15789 856
rect 15841 860 15920 876
rect 15952 876 16124 878
rect 15952 860 16031 876
rect 16038 874 16068 876
rect 15616 838 15645 848
rect 15659 838 15688 848
rect 15703 838 15733 852
rect 15776 838 15819 852
rect 15841 848 16031 860
rect 16096 856 16102 876
rect 15826 838 15856 848
rect 15857 838 16015 848
rect 16019 838 16049 848
rect 16053 838 16083 852
rect 16111 838 16124 876
rect 16196 890 16225 906
rect 16239 890 16268 906
rect 16283 896 16313 912
rect 16341 890 16347 938
rect 16350 932 16369 938
rect 16384 932 16414 940
rect 16350 924 16414 932
rect 16350 908 16430 924
rect 16446 917 16508 948
rect 16524 917 16586 948
rect 16655 946 16704 971
rect 16719 946 16749 962
rect 16618 932 16648 940
rect 16655 938 16765 946
rect 16618 924 16663 932
rect 16350 906 16369 908
rect 16384 906 16430 908
rect 16350 890 16430 906
rect 16457 904 16492 917
rect 16533 914 16570 917
rect 16533 912 16575 914
rect 16462 901 16492 904
rect 16471 897 16478 901
rect 16478 896 16479 897
rect 16437 890 16447 896
rect 16196 882 16231 890
rect 16196 856 16197 882
rect 16204 856 16231 882
rect 16139 838 16169 852
rect 16196 848 16231 856
rect 16233 882 16274 890
rect 16233 856 16248 882
rect 16255 856 16274 882
rect 16338 878 16369 890
rect 16384 878 16487 890
rect 16499 880 16525 906
rect 16540 901 16570 912
rect 16602 908 16664 924
rect 16602 906 16648 908
rect 16602 890 16664 906
rect 16676 890 16682 938
rect 16685 930 16765 938
rect 16685 928 16704 930
rect 16719 928 16753 930
rect 16685 912 16765 928
rect 16685 890 16704 912
rect 16719 896 16749 912
rect 16777 906 16783 980
rect 16786 906 16805 1050
rect 16820 906 16826 1050
rect 16835 980 16848 1050
rect 16900 1046 16922 1050
rect 16893 1024 16922 1038
rect 16975 1024 16991 1038
rect 17029 1034 17035 1036
rect 17042 1034 17150 1050
rect 17157 1034 17163 1036
rect 17171 1034 17186 1050
rect 17252 1044 17271 1047
rect 16893 1022 16991 1024
rect 17018 1022 17186 1034
rect 17201 1024 17217 1038
rect 17252 1025 17274 1044
rect 17284 1038 17300 1039
rect 17283 1036 17300 1038
rect 17284 1031 17300 1036
rect 17274 1024 17280 1025
rect 17283 1024 17312 1031
rect 17201 1023 17312 1024
rect 17201 1022 17318 1023
rect 16877 1014 16928 1022
rect 16975 1014 17009 1022
rect 16877 1002 16902 1014
rect 16909 1002 16928 1014
rect 16982 1012 17009 1014
rect 17018 1012 17239 1022
rect 17274 1019 17280 1022
rect 16982 1008 17239 1012
rect 16877 994 16928 1002
rect 16975 994 17239 1008
rect 17283 1014 17318 1022
rect 16829 946 16848 980
rect 16893 986 16922 994
rect 16893 980 16910 986
rect 16893 978 16927 980
rect 16975 978 16991 994
rect 16992 984 17200 994
rect 17201 984 17217 994
rect 17265 990 17280 1005
rect 17283 1002 17284 1014
rect 17291 1002 17318 1014
rect 17283 994 17318 1002
rect 17283 993 17312 994
rect 17003 980 17217 984
rect 17018 978 17217 980
rect 17252 980 17265 990
rect 17283 980 17300 993
rect 17252 978 17300 980
rect 16894 974 16927 978
rect 16890 972 16927 974
rect 16890 971 16957 972
rect 16890 966 16921 971
rect 16927 966 16957 971
rect 16890 962 16957 966
rect 16863 959 16957 962
rect 16863 952 16912 959
rect 16863 946 16893 952
rect 16912 947 16917 952
rect 16829 930 16909 946
rect 16921 938 16957 959
rect 17018 954 17207 978
rect 17252 977 17299 978
rect 17265 972 17299 977
rect 17033 951 17207 954
rect 17026 948 17207 951
rect 17235 971 17299 972
rect 16829 928 16848 930
rect 16863 928 16897 930
rect 16829 912 16909 928
rect 16829 906 16848 912
rect 16545 880 16648 890
rect 16499 878 16648 880
rect 16669 878 16704 890
rect 16338 876 16500 878
rect 16350 856 16369 876
rect 16384 874 16414 876
rect 16233 848 16274 856
rect 16356 852 16369 856
rect 16421 860 16500 876
rect 16532 876 16704 878
rect 16532 860 16611 876
rect 16618 874 16648 876
rect 16196 838 16225 848
rect 16239 838 16268 848
rect 16283 838 16313 852
rect 16356 838 16399 852
rect 16421 848 16611 860
rect 16676 856 16682 876
rect 16406 838 16436 848
rect 16437 838 16595 848
rect 16599 838 16629 848
rect 16633 838 16663 852
rect 16691 838 16704 876
rect 16776 890 16805 906
rect 16819 890 16848 906
rect 16863 896 16893 912
rect 16921 890 16927 938
rect 16930 932 16949 938
rect 16964 932 16994 940
rect 16930 924 16994 932
rect 16930 908 17010 924
rect 17026 917 17088 948
rect 17104 917 17166 948
rect 17235 946 17284 971
rect 17299 946 17329 962
rect 17198 932 17228 940
rect 17235 938 17345 946
rect 17198 924 17243 932
rect 16930 906 16949 908
rect 16964 906 17010 908
rect 16930 890 17010 906
rect 17037 904 17072 917
rect 17113 914 17150 917
rect 17113 912 17155 914
rect 17042 901 17072 904
rect 17051 897 17058 901
rect 17058 896 17059 897
rect 17017 890 17027 896
rect 16776 882 16811 890
rect 16776 856 16777 882
rect 16784 856 16811 882
rect 16719 838 16749 852
rect 16776 848 16811 856
rect 16813 882 16854 890
rect 16813 856 16828 882
rect 16835 856 16854 882
rect 16918 878 16949 890
rect 16964 878 17067 890
rect 17079 880 17105 906
rect 17120 901 17150 912
rect 17182 908 17244 924
rect 17182 906 17228 908
rect 17182 890 17244 906
rect 17256 890 17262 938
rect 17265 930 17345 938
rect 17265 928 17284 930
rect 17299 928 17333 930
rect 17265 912 17345 928
rect 17265 890 17284 912
rect 17299 896 17329 912
rect 17357 906 17363 980
rect 17366 906 17385 1050
rect 17400 906 17406 1050
rect 17415 980 17428 1050
rect 17480 1046 17502 1050
rect 17473 1024 17502 1038
rect 17555 1024 17571 1038
rect 17609 1034 17615 1036
rect 17622 1034 17730 1050
rect 17737 1034 17743 1036
rect 17751 1034 17766 1050
rect 17832 1044 17851 1047
rect 17473 1022 17571 1024
rect 17598 1022 17766 1034
rect 17781 1024 17797 1038
rect 17832 1025 17854 1044
rect 17864 1038 17880 1039
rect 17863 1036 17880 1038
rect 17864 1031 17880 1036
rect 17854 1024 17860 1025
rect 17863 1024 17892 1031
rect 17781 1023 17892 1024
rect 17781 1022 17898 1023
rect 17457 1014 17508 1022
rect 17555 1014 17589 1022
rect 17457 1002 17482 1014
rect 17489 1002 17508 1014
rect 17562 1012 17589 1014
rect 17598 1012 17819 1022
rect 17854 1019 17860 1022
rect 17562 1008 17819 1012
rect 17457 994 17508 1002
rect 17555 994 17819 1008
rect 17863 1014 17898 1022
rect 17409 946 17428 980
rect 17473 986 17502 994
rect 17473 980 17490 986
rect 17473 978 17507 980
rect 17555 978 17571 994
rect 17572 984 17780 994
rect 17781 984 17797 994
rect 17845 990 17860 1005
rect 17863 1002 17864 1014
rect 17871 1002 17898 1014
rect 17863 994 17898 1002
rect 17863 993 17892 994
rect 17583 980 17797 984
rect 17598 978 17797 980
rect 17832 980 17845 990
rect 17863 980 17880 993
rect 17832 978 17880 980
rect 17474 974 17507 978
rect 17470 972 17507 974
rect 17470 971 17537 972
rect 17470 966 17501 971
rect 17507 966 17537 971
rect 17470 962 17537 966
rect 17443 959 17537 962
rect 17443 952 17492 959
rect 17443 946 17473 952
rect 17492 947 17497 952
rect 17409 930 17489 946
rect 17501 938 17537 959
rect 17598 954 17787 978
rect 17832 977 17879 978
rect 17845 972 17879 977
rect 17613 951 17787 954
rect 17606 948 17787 951
rect 17815 971 17879 972
rect 17409 928 17428 930
rect 17443 928 17477 930
rect 17409 912 17489 928
rect 17409 906 17428 912
rect 17125 880 17228 890
rect 17079 878 17228 880
rect 17249 878 17284 890
rect 16918 876 17080 878
rect 16930 856 16949 876
rect 16964 874 16994 876
rect 16813 848 16854 856
rect 16936 852 16949 856
rect 17001 860 17080 876
rect 17112 876 17284 878
rect 17112 860 17191 876
rect 17198 874 17228 876
rect 16776 838 16805 848
rect 16819 838 16848 848
rect 16863 838 16893 852
rect 16936 838 16979 852
rect 17001 848 17191 860
rect 17256 856 17262 876
rect 16986 838 17016 848
rect 17017 838 17175 848
rect 17179 838 17209 848
rect 17213 838 17243 852
rect 17271 838 17284 876
rect 17356 890 17385 906
rect 17399 890 17428 906
rect 17443 896 17473 912
rect 17501 890 17507 938
rect 17510 932 17529 938
rect 17544 932 17574 940
rect 17510 924 17574 932
rect 17510 908 17590 924
rect 17606 917 17668 948
rect 17684 917 17746 948
rect 17815 946 17864 971
rect 17879 946 17909 962
rect 17778 932 17808 940
rect 17815 938 17925 946
rect 17778 924 17823 932
rect 17510 906 17529 908
rect 17544 906 17590 908
rect 17510 890 17590 906
rect 17617 904 17652 917
rect 17693 914 17730 917
rect 17693 912 17735 914
rect 17622 901 17652 904
rect 17631 897 17638 901
rect 17638 896 17639 897
rect 17597 890 17607 896
rect 17356 882 17391 890
rect 17356 856 17357 882
rect 17364 856 17391 882
rect 17299 838 17329 852
rect 17356 848 17391 856
rect 17393 882 17434 890
rect 17393 856 17408 882
rect 17415 856 17434 882
rect 17498 878 17529 890
rect 17544 878 17647 890
rect 17659 880 17685 906
rect 17700 901 17730 912
rect 17762 908 17824 924
rect 17762 906 17808 908
rect 17762 890 17824 906
rect 17836 890 17842 938
rect 17845 930 17925 938
rect 17845 928 17864 930
rect 17879 928 17913 930
rect 17845 912 17925 928
rect 17845 890 17864 912
rect 17879 896 17909 912
rect 17937 906 17943 980
rect 17946 906 17965 1050
rect 17980 906 17986 1050
rect 17995 980 18008 1050
rect 18060 1046 18082 1050
rect 18053 1024 18082 1038
rect 18135 1024 18151 1038
rect 18189 1034 18195 1036
rect 18202 1034 18310 1050
rect 18317 1034 18323 1036
rect 18331 1034 18346 1050
rect 18412 1044 18431 1047
rect 18053 1022 18151 1024
rect 18178 1022 18346 1034
rect 18361 1024 18377 1038
rect 18412 1025 18434 1044
rect 18444 1038 18460 1039
rect 18443 1036 18460 1038
rect 18444 1031 18460 1036
rect 18434 1024 18440 1025
rect 18443 1024 18472 1031
rect 18361 1023 18472 1024
rect 18361 1022 18478 1023
rect 18037 1014 18088 1022
rect 18135 1014 18169 1022
rect 18037 1002 18062 1014
rect 18069 1002 18088 1014
rect 18142 1012 18169 1014
rect 18178 1012 18399 1022
rect 18434 1019 18440 1022
rect 18142 1008 18399 1012
rect 18037 994 18088 1002
rect 18135 994 18399 1008
rect 18443 1014 18478 1022
rect 17989 946 18008 980
rect 18053 986 18082 994
rect 18053 980 18070 986
rect 18053 978 18087 980
rect 18135 978 18151 994
rect 18152 984 18360 994
rect 18361 984 18377 994
rect 18425 990 18440 1005
rect 18443 1002 18444 1014
rect 18451 1002 18478 1014
rect 18443 994 18478 1002
rect 18443 993 18472 994
rect 18163 980 18377 984
rect 18178 978 18377 980
rect 18412 980 18425 990
rect 18443 980 18460 993
rect 18412 978 18460 980
rect 18054 974 18087 978
rect 18050 972 18087 974
rect 18050 971 18117 972
rect 18050 966 18081 971
rect 18087 966 18117 971
rect 18050 962 18117 966
rect 18023 959 18117 962
rect 18023 952 18072 959
rect 18023 946 18053 952
rect 18072 947 18077 952
rect 17989 930 18069 946
rect 18081 938 18117 959
rect 18178 954 18367 978
rect 18412 977 18459 978
rect 18425 972 18459 977
rect 18193 951 18367 954
rect 18186 948 18367 951
rect 18395 971 18459 972
rect 17989 928 18008 930
rect 18023 928 18057 930
rect 17989 912 18069 928
rect 17989 906 18008 912
rect 17705 880 17808 890
rect 17659 878 17808 880
rect 17829 878 17864 890
rect 17498 876 17660 878
rect 17510 856 17529 876
rect 17544 874 17574 876
rect 17393 848 17434 856
rect 17516 852 17529 856
rect 17581 860 17660 876
rect 17692 876 17864 878
rect 17692 860 17771 876
rect 17778 874 17808 876
rect 17356 838 17385 848
rect 17399 838 17428 848
rect 17443 838 17473 852
rect 17516 838 17559 852
rect 17581 848 17771 860
rect 17836 856 17842 876
rect 17566 838 17596 848
rect 17597 838 17755 848
rect 17759 838 17789 848
rect 17793 838 17823 852
rect 17851 838 17864 876
rect 17936 890 17965 906
rect 17979 890 18008 906
rect 18023 896 18053 912
rect 18081 890 18087 938
rect 18090 932 18109 938
rect 18124 932 18154 940
rect 18090 924 18154 932
rect 18090 908 18170 924
rect 18186 917 18248 948
rect 18264 917 18326 948
rect 18395 946 18444 971
rect 18459 946 18489 962
rect 18358 932 18388 940
rect 18395 938 18505 946
rect 18358 924 18403 932
rect 18090 906 18109 908
rect 18124 906 18170 908
rect 18090 890 18170 906
rect 18197 904 18232 917
rect 18273 914 18310 917
rect 18273 912 18315 914
rect 18202 901 18232 904
rect 18211 897 18218 901
rect 18218 896 18219 897
rect 18177 890 18187 896
rect 17936 882 17971 890
rect 17936 856 17937 882
rect 17944 856 17971 882
rect 17879 838 17909 852
rect 17936 848 17971 856
rect 17973 882 18014 890
rect 17973 856 17988 882
rect 17995 856 18014 882
rect 18078 878 18109 890
rect 18124 878 18227 890
rect 18239 880 18265 906
rect 18280 901 18310 912
rect 18342 908 18404 924
rect 18342 906 18388 908
rect 18342 890 18404 906
rect 18416 890 18422 938
rect 18425 930 18505 938
rect 18425 928 18444 930
rect 18459 928 18493 930
rect 18425 912 18505 928
rect 18425 890 18444 912
rect 18459 896 18489 912
rect 18517 906 18523 980
rect 18532 906 18545 1050
rect 18285 880 18388 890
rect 18239 878 18388 880
rect 18409 878 18444 890
rect 18078 876 18240 878
rect 18090 856 18109 876
rect 18124 874 18154 876
rect 17973 848 18014 856
rect 18096 852 18109 856
rect 18161 860 18240 876
rect 18272 876 18444 878
rect 18272 860 18351 876
rect 18358 874 18388 876
rect 17936 838 17965 848
rect 17979 838 18008 848
rect 18023 838 18053 852
rect 18096 838 18139 852
rect 18161 848 18351 860
rect 18416 856 18422 876
rect 18146 838 18176 848
rect 18177 838 18335 848
rect 18339 838 18369 848
rect 18373 838 18403 852
rect 18431 838 18444 876
rect 18516 890 18545 906
rect 18516 882 18551 890
rect 18516 856 18517 882
rect 18524 856 18551 882
rect 18459 838 18489 852
rect 18516 848 18551 856
rect 18516 838 18545 848
rect -1 832 18545 838
rect 0 824 18545 832
rect 15 794 28 824
rect 43 810 73 824
rect 116 810 159 824
rect 166 810 386 824
rect 393 810 423 824
rect 83 796 98 808
rect 117 796 130 810
rect 198 806 351 810
rect 80 794 102 796
rect 180 794 372 806
rect 451 794 464 824
rect 479 810 509 824
rect 546 794 565 824
rect 580 794 586 824
rect 595 794 608 824
rect 623 810 653 824
rect 696 810 739 824
rect 746 810 966 824
rect 973 810 1003 824
rect 663 796 678 808
rect 697 796 710 810
rect 778 806 931 810
rect 660 794 682 796
rect 760 794 952 806
rect 1031 794 1044 824
rect 1059 810 1089 824
rect 1126 794 1145 824
rect 1160 794 1166 824
rect 1175 794 1188 824
rect 1203 810 1233 824
rect 1276 810 1319 824
rect 1326 810 1546 824
rect 1553 810 1583 824
rect 1243 796 1258 808
rect 1277 796 1290 810
rect 1358 806 1511 810
rect 1240 794 1262 796
rect 1340 794 1532 806
rect 1611 794 1624 824
rect 1639 810 1669 824
rect 1706 794 1725 824
rect 1740 794 1746 824
rect 1755 794 1768 824
rect 1783 810 1813 824
rect 1856 810 1899 824
rect 1906 810 2126 824
rect 2133 810 2163 824
rect 1823 796 1838 808
rect 1857 796 1870 810
rect 1938 806 2091 810
rect 1820 794 1842 796
rect 1920 794 2112 806
rect 2191 794 2204 824
rect 2219 810 2249 824
rect 2286 794 2305 824
rect 2320 794 2326 824
rect 2335 794 2348 824
rect 2363 810 2393 824
rect 2436 810 2479 824
rect 2486 810 2706 824
rect 2713 810 2743 824
rect 2403 796 2418 808
rect 2437 796 2450 810
rect 2518 806 2671 810
rect 2400 794 2422 796
rect 2500 794 2692 806
rect 2771 794 2784 824
rect 2799 810 2829 824
rect 2866 794 2885 824
rect 2900 794 2906 824
rect 2915 794 2928 824
rect 2943 810 2973 824
rect 3016 810 3059 824
rect 3066 810 3286 824
rect 3293 810 3323 824
rect 2983 796 2998 808
rect 3017 796 3030 810
rect 3098 806 3251 810
rect 2980 794 3002 796
rect 3080 794 3272 806
rect 3351 794 3364 824
rect 3379 810 3409 824
rect 3446 794 3465 824
rect 3480 794 3486 824
rect 3495 794 3508 824
rect 3523 810 3553 824
rect 3596 810 3639 824
rect 3646 810 3866 824
rect 3873 810 3903 824
rect 3563 796 3578 808
rect 3597 796 3610 810
rect 3678 806 3831 810
rect 3560 794 3582 796
rect 3660 794 3852 806
rect 3931 794 3944 824
rect 3959 810 3989 824
rect 4026 794 4045 824
rect 4060 794 4066 824
rect 4075 794 4088 824
rect 4103 810 4133 824
rect 4176 810 4219 824
rect 4226 810 4446 824
rect 4453 810 4483 824
rect 4143 796 4158 808
rect 4177 796 4190 810
rect 4258 806 4411 810
rect 4140 794 4162 796
rect 4240 794 4432 806
rect 4511 794 4524 824
rect 4539 810 4569 824
rect 4606 794 4625 824
rect 4640 794 4646 824
rect 4655 794 4668 824
rect 4683 810 4713 824
rect 4756 810 4799 824
rect 4806 810 5026 824
rect 5033 810 5063 824
rect 4723 796 4738 808
rect 4757 796 4770 810
rect 4838 806 4991 810
rect 4720 794 4742 796
rect 4820 794 5012 806
rect 5091 794 5104 824
rect 5119 810 5149 824
rect 5186 794 5205 824
rect 5220 794 5226 824
rect 5235 794 5248 824
rect 5263 810 5293 824
rect 5336 810 5379 824
rect 5386 810 5606 824
rect 5613 810 5643 824
rect 5303 796 5318 808
rect 5337 796 5350 810
rect 5418 806 5571 810
rect 5300 794 5322 796
rect 5400 794 5592 806
rect 5671 794 5684 824
rect 5699 810 5729 824
rect 5766 794 5785 824
rect 5800 794 5806 824
rect 5815 794 5828 824
rect 5843 810 5873 824
rect 5916 810 5959 824
rect 5966 810 6186 824
rect 6193 810 6223 824
rect 5883 796 5898 808
rect 5917 796 5930 810
rect 5998 806 6151 810
rect 5880 794 5902 796
rect 5980 794 6172 806
rect 6251 794 6264 824
rect 6279 810 6309 824
rect 6346 794 6365 824
rect 6380 794 6386 824
rect 6395 794 6408 824
rect 6423 810 6453 824
rect 6496 810 6539 824
rect 6546 810 6766 824
rect 6773 810 6803 824
rect 6463 796 6478 808
rect 6497 796 6510 810
rect 6578 806 6731 810
rect 6460 794 6482 796
rect 6560 794 6752 806
rect 6831 794 6844 824
rect 6859 810 6889 824
rect 6926 794 6945 824
rect 6960 794 6966 824
rect 6975 794 6988 824
rect 7003 810 7033 824
rect 7076 810 7119 824
rect 7126 810 7346 824
rect 7353 810 7383 824
rect 7043 796 7058 808
rect 7077 796 7090 810
rect 7158 806 7311 810
rect 7040 794 7062 796
rect 7140 794 7332 806
rect 7411 794 7424 824
rect 7439 810 7469 824
rect 7506 794 7525 824
rect 7540 794 7546 824
rect 7555 794 7568 824
rect 7583 810 7613 824
rect 7656 810 7699 824
rect 7706 810 7926 824
rect 7933 810 7963 824
rect 7623 796 7638 808
rect 7657 796 7670 810
rect 7738 806 7891 810
rect 7620 794 7642 796
rect 7720 794 7912 806
rect 7991 794 8004 824
rect 8019 810 8049 824
rect 8086 794 8105 824
rect 8120 794 8126 824
rect 8135 794 8148 824
rect 8163 810 8193 824
rect 8236 810 8279 824
rect 8286 810 8506 824
rect 8513 810 8543 824
rect 8203 796 8218 808
rect 8237 796 8250 810
rect 8318 806 8471 810
rect 8200 794 8222 796
rect 8300 794 8492 806
rect 8571 794 8584 824
rect 8599 810 8629 824
rect 8666 794 8685 824
rect 8700 794 8706 824
rect 8715 794 8728 824
rect 8743 810 8773 824
rect 8816 810 8859 824
rect 8866 810 9086 824
rect 9093 810 9123 824
rect 8783 796 8798 808
rect 8817 796 8830 810
rect 8898 806 9051 810
rect 8780 794 8802 796
rect 8880 794 9072 806
rect 9151 794 9164 824
rect 9179 810 9209 824
rect 9246 794 9265 824
rect 9280 794 9286 824
rect 9295 794 9308 824
rect 9323 810 9353 824
rect 9396 810 9439 824
rect 9446 810 9666 824
rect 9673 810 9703 824
rect 9363 796 9378 808
rect 9397 796 9410 810
rect 9478 806 9631 810
rect 9360 794 9382 796
rect 9460 794 9652 806
rect 9731 794 9744 824
rect 9759 810 9789 824
rect 9826 794 9845 824
rect 9860 794 9866 824
rect 9875 794 9888 824
rect 9903 810 9933 824
rect 9976 810 10019 824
rect 10026 810 10246 824
rect 10253 810 10283 824
rect 9943 796 9958 808
rect 9977 796 9990 810
rect 10058 806 10211 810
rect 9940 794 9962 796
rect 10040 794 10232 806
rect 10311 794 10324 824
rect 10339 810 10369 824
rect 10406 794 10425 824
rect 10440 794 10446 824
rect 10455 794 10468 824
rect 10483 810 10513 824
rect 10556 810 10599 824
rect 10606 810 10826 824
rect 10833 810 10863 824
rect 10523 796 10538 808
rect 10557 796 10570 810
rect 10638 806 10791 810
rect 10520 794 10542 796
rect 10620 794 10812 806
rect 10891 794 10904 824
rect 10919 810 10949 824
rect 10986 794 11005 824
rect 11020 794 11026 824
rect 11035 794 11048 824
rect 11063 810 11093 824
rect 11136 810 11179 824
rect 11186 810 11406 824
rect 11413 810 11443 824
rect 11103 796 11118 808
rect 11137 796 11150 810
rect 11218 806 11371 810
rect 11100 794 11122 796
rect 11200 794 11392 806
rect 11471 794 11484 824
rect 11499 810 11529 824
rect 11566 794 11585 824
rect 11600 794 11606 824
rect 11615 794 11628 824
rect 11643 810 11673 824
rect 11716 810 11759 824
rect 11766 810 11986 824
rect 11993 810 12023 824
rect 11683 796 11698 808
rect 11717 796 11730 810
rect 11798 806 11951 810
rect 11680 794 11702 796
rect 11780 794 11972 806
rect 12051 794 12064 824
rect 12079 810 12109 824
rect 12146 794 12165 824
rect 12180 794 12186 824
rect 12195 794 12208 824
rect 12223 810 12253 824
rect 12296 810 12339 824
rect 12346 810 12566 824
rect 12573 810 12603 824
rect 12263 796 12278 808
rect 12297 796 12310 810
rect 12378 806 12531 810
rect 12260 794 12282 796
rect 12360 794 12552 806
rect 12631 794 12644 824
rect 12659 810 12689 824
rect 12726 794 12745 824
rect 12760 794 12766 824
rect 12775 794 12788 824
rect 12803 810 12833 824
rect 12876 810 12919 824
rect 12926 810 13146 824
rect 13153 810 13183 824
rect 12843 796 12858 808
rect 12877 796 12890 810
rect 12958 806 13111 810
rect 12840 794 12862 796
rect 12940 794 13132 806
rect 13211 794 13224 824
rect 13239 810 13269 824
rect 13306 794 13325 824
rect 13340 794 13346 824
rect 13355 794 13368 824
rect 13383 810 13413 824
rect 13456 810 13499 824
rect 13506 810 13726 824
rect 13733 810 13763 824
rect 13423 796 13438 808
rect 13457 796 13470 810
rect 13538 806 13691 810
rect 13420 794 13442 796
rect 13520 794 13712 806
rect 13791 794 13804 824
rect 13819 810 13849 824
rect 13886 794 13905 824
rect 13920 794 13926 824
rect 13935 794 13948 824
rect 13963 810 13993 824
rect 14036 810 14079 824
rect 14086 810 14306 824
rect 14313 810 14343 824
rect 14003 796 14018 808
rect 14037 796 14050 810
rect 14118 806 14271 810
rect 14000 794 14022 796
rect 14100 794 14292 806
rect 14371 794 14384 824
rect 14399 810 14429 824
rect 14466 794 14485 824
rect 14500 794 14506 824
rect 14515 794 14528 824
rect 14543 810 14573 824
rect 14616 810 14659 824
rect 14666 810 14886 824
rect 14893 810 14923 824
rect 14583 796 14598 808
rect 14617 796 14630 810
rect 14698 806 14851 810
rect 14580 794 14602 796
rect 14680 794 14872 806
rect 14951 794 14964 824
rect 14979 810 15009 824
rect 15046 794 15065 824
rect 15080 794 15086 824
rect 15095 794 15108 824
rect 15123 810 15153 824
rect 15196 810 15239 824
rect 15246 810 15466 824
rect 15473 810 15503 824
rect 15163 796 15178 808
rect 15197 796 15210 810
rect 15278 806 15431 810
rect 15160 794 15182 796
rect 15260 794 15452 806
rect 15531 794 15544 824
rect 15559 810 15589 824
rect 15626 794 15645 824
rect 15660 794 15666 824
rect 15675 794 15688 824
rect 15703 810 15733 824
rect 15776 810 15819 824
rect 15826 810 16046 824
rect 16053 810 16083 824
rect 15743 796 15758 808
rect 15777 796 15790 810
rect 15858 806 16011 810
rect 15740 794 15762 796
rect 15840 794 16032 806
rect 16111 794 16124 824
rect 16139 810 16169 824
rect 16206 794 16225 824
rect 16240 794 16246 824
rect 16255 794 16268 824
rect 16283 810 16313 824
rect 16356 810 16399 824
rect 16406 810 16626 824
rect 16633 810 16663 824
rect 16323 796 16338 808
rect 16357 796 16370 810
rect 16438 806 16591 810
rect 16320 794 16342 796
rect 16420 794 16612 806
rect 16691 794 16704 824
rect 16719 810 16749 824
rect 16786 794 16805 824
rect 16820 794 16826 824
rect 16835 794 16848 824
rect 16863 810 16893 824
rect 16936 810 16979 824
rect 16986 810 17206 824
rect 17213 810 17243 824
rect 16903 796 16918 808
rect 16937 796 16950 810
rect 17018 806 17171 810
rect 16900 794 16922 796
rect 17000 794 17192 806
rect 17271 794 17284 824
rect 17299 810 17329 824
rect 17366 794 17385 824
rect 17400 794 17406 824
rect 17415 794 17428 824
rect 17443 810 17473 824
rect 17516 810 17559 824
rect 17566 810 17786 824
rect 17793 810 17823 824
rect 17483 796 17498 808
rect 17517 796 17530 810
rect 17598 806 17751 810
rect 17480 794 17502 796
rect 17580 794 17772 806
rect 17851 794 17864 824
rect 17879 810 17909 824
rect 17946 794 17965 824
rect 17980 794 17986 824
rect 17995 794 18008 824
rect 18023 810 18053 824
rect 18096 810 18139 824
rect 18146 810 18366 824
rect 18373 810 18403 824
rect 18063 796 18078 808
rect 18097 796 18110 810
rect 18178 806 18331 810
rect 18060 794 18082 796
rect 18160 794 18352 806
rect 18431 794 18444 824
rect 18459 810 18489 824
rect 18532 794 18545 824
rect 0 780 18545 794
rect 15 710 28 780
rect 80 776 102 780
rect 73 754 102 768
rect 155 754 171 768
rect 209 764 215 766
rect 222 764 330 780
rect 337 764 343 766
rect 351 764 366 780
rect 432 774 451 777
rect 73 752 171 754
rect 198 752 366 764
rect 381 754 397 768
rect 432 755 454 774
rect 464 768 480 769
rect 463 766 480 768
rect 464 761 480 766
rect 454 754 460 755
rect 463 754 492 761
rect 381 753 492 754
rect 381 752 498 753
rect 57 744 108 752
rect 155 744 189 752
rect 57 732 82 744
rect 89 732 108 744
rect 162 742 189 744
rect 198 742 419 752
rect 454 749 460 752
rect 162 738 419 742
rect 57 724 108 732
rect 155 724 419 738
rect 463 744 498 752
rect 9 676 28 710
rect 73 716 102 724
rect 73 710 90 716
rect 73 708 107 710
rect 155 708 171 724
rect 172 714 380 724
rect 381 714 397 724
rect 445 720 460 735
rect 463 732 464 744
rect 471 732 498 744
rect 463 724 498 732
rect 463 723 492 724
rect 183 710 397 714
rect 198 708 397 710
rect 432 710 445 720
rect 463 710 480 723
rect 432 708 480 710
rect 74 704 107 708
rect 70 702 107 704
rect 70 701 137 702
rect 70 696 101 701
rect 107 696 137 701
rect 70 692 137 696
rect 43 689 137 692
rect 43 682 92 689
rect 43 676 73 682
rect 92 677 97 682
rect 9 660 89 676
rect 101 668 137 689
rect 198 684 387 708
rect 432 707 479 708
rect 445 702 479 707
rect 213 681 387 684
rect 206 678 387 681
rect 415 701 479 702
rect 9 658 28 660
rect 43 658 77 660
rect 9 642 89 658
rect 9 636 28 642
rect -1 620 28 636
rect 43 626 73 642
rect 101 620 107 668
rect 110 662 129 668
rect 144 662 174 670
rect 110 654 174 662
rect 110 638 190 654
rect 206 647 268 678
rect 284 647 346 678
rect 415 676 464 701
rect 479 676 509 692
rect 378 662 408 670
rect 415 668 525 676
rect 378 654 423 662
rect 110 636 129 638
rect 144 636 190 638
rect 110 620 190 636
rect 217 634 252 647
rect 293 644 330 647
rect 293 642 335 644
rect 222 631 252 634
rect 231 627 238 631
rect 238 626 239 627
rect 197 620 207 626
rect -7 612 34 620
rect -7 586 8 612
rect 15 586 34 612
rect 98 608 129 620
rect 144 608 247 620
rect 259 610 285 636
rect 300 631 330 642
rect 362 638 424 654
rect 362 636 408 638
rect 362 620 424 636
rect 436 620 442 668
rect 445 660 525 668
rect 445 658 464 660
rect 479 658 513 660
rect 445 642 525 658
rect 445 620 464 642
rect 479 626 509 642
rect 537 636 543 710
rect 546 636 565 780
rect 580 636 586 780
rect 595 710 608 780
rect 660 776 682 780
rect 653 754 682 768
rect 735 754 751 768
rect 789 764 795 766
rect 802 764 910 780
rect 917 764 923 766
rect 931 764 946 780
rect 1012 774 1031 777
rect 653 752 751 754
rect 778 752 946 764
rect 961 754 977 768
rect 1012 755 1034 774
rect 1044 768 1060 769
rect 1043 766 1060 768
rect 1044 761 1060 766
rect 1034 754 1040 755
rect 1043 754 1072 761
rect 961 753 1072 754
rect 961 752 1078 753
rect 637 744 688 752
rect 735 744 769 752
rect 637 732 662 744
rect 669 732 688 744
rect 742 742 769 744
rect 778 742 999 752
rect 1034 749 1040 752
rect 742 738 999 742
rect 637 724 688 732
rect 735 724 999 738
rect 1043 744 1078 752
rect 589 676 608 710
rect 653 716 682 724
rect 653 710 670 716
rect 653 708 687 710
rect 735 708 751 724
rect 752 714 960 724
rect 961 714 977 724
rect 1025 720 1040 735
rect 1043 732 1044 744
rect 1051 732 1078 744
rect 1043 724 1078 732
rect 1043 723 1072 724
rect 763 710 977 714
rect 778 708 977 710
rect 1012 710 1025 720
rect 1043 710 1060 723
rect 1012 708 1060 710
rect 654 704 687 708
rect 650 702 687 704
rect 650 701 717 702
rect 650 696 681 701
rect 687 696 717 701
rect 650 692 717 696
rect 623 689 717 692
rect 623 682 672 689
rect 623 676 653 682
rect 672 677 677 682
rect 589 660 669 676
rect 681 668 717 689
rect 778 684 967 708
rect 1012 707 1059 708
rect 1025 702 1059 707
rect 793 681 967 684
rect 786 678 967 681
rect 995 701 1059 702
rect 589 658 608 660
rect 623 658 657 660
rect 589 642 669 658
rect 589 636 608 642
rect 305 610 408 620
rect 259 608 408 610
rect 429 608 464 620
rect 98 606 260 608
rect 110 586 129 606
rect 144 604 174 606
rect -7 578 34 586
rect 116 582 129 586
rect 181 590 260 606
rect 292 606 464 608
rect 292 590 371 606
rect 378 604 408 606
rect -1 568 28 578
rect 43 568 73 582
rect 116 568 159 582
rect 181 578 371 590
rect 436 586 442 606
rect 166 568 196 578
rect 197 568 355 578
rect 359 568 389 578
rect 393 568 423 582
rect 451 568 464 606
rect 536 620 565 636
rect 579 620 608 636
rect 623 626 653 642
rect 681 620 687 668
rect 690 662 709 668
rect 724 662 754 670
rect 690 654 754 662
rect 690 638 770 654
rect 786 647 848 678
rect 864 647 926 678
rect 995 676 1044 701
rect 1059 676 1089 692
rect 958 662 988 670
rect 995 668 1105 676
rect 958 654 1003 662
rect 690 636 709 638
rect 724 636 770 638
rect 690 620 770 636
rect 797 634 832 647
rect 873 644 910 647
rect 873 642 915 644
rect 802 631 832 634
rect 811 627 818 631
rect 818 626 819 627
rect 777 620 787 626
rect 536 612 571 620
rect 536 586 537 612
rect 544 586 571 612
rect 479 568 509 582
rect 536 578 571 586
rect 573 612 614 620
rect 573 586 588 612
rect 595 586 614 612
rect 678 608 709 620
rect 724 608 827 620
rect 839 610 865 636
rect 880 631 910 642
rect 942 638 1004 654
rect 942 636 988 638
rect 942 620 1004 636
rect 1016 620 1022 668
rect 1025 660 1105 668
rect 1025 658 1044 660
rect 1059 658 1093 660
rect 1025 642 1105 658
rect 1025 620 1044 642
rect 1059 626 1089 642
rect 1117 636 1123 710
rect 1126 636 1145 780
rect 1160 636 1166 780
rect 1175 710 1188 780
rect 1240 776 1262 780
rect 1233 754 1262 768
rect 1315 754 1331 768
rect 1369 764 1375 766
rect 1382 764 1490 780
rect 1497 764 1503 766
rect 1511 764 1526 780
rect 1592 774 1611 777
rect 1233 752 1331 754
rect 1358 752 1526 764
rect 1541 754 1557 768
rect 1592 755 1614 774
rect 1624 768 1640 769
rect 1623 766 1640 768
rect 1624 761 1640 766
rect 1614 754 1620 755
rect 1623 754 1652 761
rect 1541 753 1652 754
rect 1541 752 1658 753
rect 1217 744 1268 752
rect 1315 744 1349 752
rect 1217 732 1242 744
rect 1249 732 1268 744
rect 1322 742 1349 744
rect 1358 742 1579 752
rect 1614 749 1620 752
rect 1322 738 1579 742
rect 1217 724 1268 732
rect 1315 724 1579 738
rect 1623 744 1658 752
rect 1169 676 1188 710
rect 1233 716 1262 724
rect 1233 710 1250 716
rect 1233 708 1267 710
rect 1315 708 1331 724
rect 1332 714 1540 724
rect 1541 714 1557 724
rect 1605 720 1620 735
rect 1623 732 1624 744
rect 1631 732 1658 744
rect 1623 724 1658 732
rect 1623 723 1652 724
rect 1343 710 1557 714
rect 1358 708 1557 710
rect 1592 710 1605 720
rect 1623 710 1640 723
rect 1592 708 1640 710
rect 1234 704 1267 708
rect 1230 702 1267 704
rect 1230 701 1297 702
rect 1230 696 1261 701
rect 1267 696 1297 701
rect 1230 692 1297 696
rect 1203 689 1297 692
rect 1203 682 1252 689
rect 1203 676 1233 682
rect 1252 677 1257 682
rect 1169 660 1249 676
rect 1261 668 1297 689
rect 1358 684 1547 708
rect 1592 707 1639 708
rect 1605 702 1639 707
rect 1373 681 1547 684
rect 1366 678 1547 681
rect 1575 701 1639 702
rect 1169 658 1188 660
rect 1203 658 1237 660
rect 1169 642 1249 658
rect 1169 636 1188 642
rect 885 610 988 620
rect 839 608 988 610
rect 1009 608 1044 620
rect 678 606 840 608
rect 690 586 709 606
rect 724 604 754 606
rect 573 578 614 586
rect 696 582 709 586
rect 761 590 840 606
rect 872 606 1044 608
rect 872 590 951 606
rect 958 604 988 606
rect 536 568 565 578
rect 579 568 608 578
rect 623 568 653 582
rect 696 568 739 582
rect 761 578 951 590
rect 1016 586 1022 606
rect 746 568 776 578
rect 777 568 935 578
rect 939 568 969 578
rect 973 568 1003 582
rect 1031 568 1044 606
rect 1116 620 1145 636
rect 1159 620 1188 636
rect 1203 626 1233 642
rect 1261 620 1267 668
rect 1270 662 1289 668
rect 1304 662 1334 670
rect 1270 654 1334 662
rect 1270 638 1350 654
rect 1366 647 1428 678
rect 1444 647 1506 678
rect 1575 676 1624 701
rect 1639 676 1669 692
rect 1538 662 1568 670
rect 1575 668 1685 676
rect 1538 654 1583 662
rect 1270 636 1289 638
rect 1304 636 1350 638
rect 1270 620 1350 636
rect 1377 634 1412 647
rect 1453 644 1490 647
rect 1453 642 1495 644
rect 1382 631 1412 634
rect 1391 627 1398 631
rect 1398 626 1399 627
rect 1357 620 1367 626
rect 1116 612 1151 620
rect 1116 586 1117 612
rect 1124 586 1151 612
rect 1059 568 1089 582
rect 1116 578 1151 586
rect 1153 612 1194 620
rect 1153 586 1168 612
rect 1175 586 1194 612
rect 1258 608 1289 620
rect 1304 608 1407 620
rect 1419 610 1445 636
rect 1460 631 1490 642
rect 1522 638 1584 654
rect 1522 636 1568 638
rect 1522 620 1584 636
rect 1596 620 1602 668
rect 1605 660 1685 668
rect 1605 658 1624 660
rect 1639 658 1673 660
rect 1605 642 1685 658
rect 1605 620 1624 642
rect 1639 626 1669 642
rect 1697 636 1703 710
rect 1706 636 1725 780
rect 1740 636 1746 780
rect 1755 710 1768 780
rect 1820 776 1842 780
rect 1813 754 1842 768
rect 1895 754 1911 768
rect 1949 764 1955 766
rect 1962 764 2070 780
rect 2077 764 2083 766
rect 2091 764 2106 780
rect 2172 774 2191 777
rect 1813 752 1911 754
rect 1938 752 2106 764
rect 2121 754 2137 768
rect 2172 755 2194 774
rect 2204 768 2220 769
rect 2203 766 2220 768
rect 2204 761 2220 766
rect 2194 754 2200 755
rect 2203 754 2232 761
rect 2121 753 2232 754
rect 2121 752 2238 753
rect 1797 744 1848 752
rect 1895 744 1929 752
rect 1797 732 1822 744
rect 1829 732 1848 744
rect 1902 742 1929 744
rect 1938 742 2159 752
rect 2194 749 2200 752
rect 1902 738 2159 742
rect 1797 724 1848 732
rect 1895 724 2159 738
rect 2203 744 2238 752
rect 1749 676 1768 710
rect 1813 716 1842 724
rect 1813 710 1830 716
rect 1813 708 1847 710
rect 1895 708 1911 724
rect 1912 714 2120 724
rect 2121 714 2137 724
rect 2185 720 2200 735
rect 2203 732 2204 744
rect 2211 732 2238 744
rect 2203 724 2238 732
rect 2203 723 2232 724
rect 1923 710 2137 714
rect 1938 708 2137 710
rect 2172 710 2185 720
rect 2203 710 2220 723
rect 2172 708 2220 710
rect 1814 704 1847 708
rect 1810 702 1847 704
rect 1810 701 1877 702
rect 1810 696 1841 701
rect 1847 696 1877 701
rect 1810 692 1877 696
rect 1783 689 1877 692
rect 1783 682 1832 689
rect 1783 676 1813 682
rect 1832 677 1837 682
rect 1749 660 1829 676
rect 1841 668 1877 689
rect 1938 684 2127 708
rect 2172 707 2219 708
rect 2185 702 2219 707
rect 1953 681 2127 684
rect 1946 678 2127 681
rect 2155 701 2219 702
rect 1749 658 1768 660
rect 1783 658 1817 660
rect 1749 642 1829 658
rect 1749 636 1768 642
rect 1465 610 1568 620
rect 1419 608 1568 610
rect 1589 608 1624 620
rect 1258 606 1420 608
rect 1270 586 1289 606
rect 1304 604 1334 606
rect 1153 578 1194 586
rect 1276 582 1289 586
rect 1341 590 1420 606
rect 1452 606 1624 608
rect 1452 590 1531 606
rect 1538 604 1568 606
rect 1116 568 1145 578
rect 1159 568 1188 578
rect 1203 568 1233 582
rect 1276 568 1319 582
rect 1341 578 1531 590
rect 1596 586 1602 606
rect 1326 568 1356 578
rect 1357 568 1515 578
rect 1519 568 1549 578
rect 1553 568 1583 582
rect 1611 568 1624 606
rect 1696 620 1725 636
rect 1739 620 1768 636
rect 1783 626 1813 642
rect 1841 620 1847 668
rect 1850 662 1869 668
rect 1884 662 1914 670
rect 1850 654 1914 662
rect 1850 638 1930 654
rect 1946 647 2008 678
rect 2024 647 2086 678
rect 2155 676 2204 701
rect 2219 676 2249 692
rect 2118 662 2148 670
rect 2155 668 2265 676
rect 2118 654 2163 662
rect 1850 636 1869 638
rect 1884 636 1930 638
rect 1850 620 1930 636
rect 1957 634 1992 647
rect 2033 644 2070 647
rect 2033 642 2075 644
rect 1962 631 1992 634
rect 1971 627 1978 631
rect 1978 626 1979 627
rect 1937 620 1947 626
rect 1696 612 1731 620
rect 1696 586 1697 612
rect 1704 586 1731 612
rect 1639 568 1669 582
rect 1696 578 1731 586
rect 1733 612 1774 620
rect 1733 586 1748 612
rect 1755 586 1774 612
rect 1838 608 1869 620
rect 1884 608 1987 620
rect 1999 610 2025 636
rect 2040 631 2070 642
rect 2102 638 2164 654
rect 2102 636 2148 638
rect 2102 620 2164 636
rect 2176 620 2182 668
rect 2185 660 2265 668
rect 2185 658 2204 660
rect 2219 658 2253 660
rect 2185 642 2265 658
rect 2185 620 2204 642
rect 2219 626 2249 642
rect 2277 636 2283 710
rect 2286 636 2305 780
rect 2320 636 2326 780
rect 2335 710 2348 780
rect 2400 776 2422 780
rect 2393 754 2422 768
rect 2475 754 2491 768
rect 2529 764 2535 766
rect 2542 764 2650 780
rect 2657 764 2663 766
rect 2671 764 2686 780
rect 2752 774 2771 777
rect 2393 752 2491 754
rect 2518 752 2686 764
rect 2701 754 2717 768
rect 2752 755 2774 774
rect 2784 768 2800 769
rect 2783 766 2800 768
rect 2784 761 2800 766
rect 2774 754 2780 755
rect 2783 754 2812 761
rect 2701 753 2812 754
rect 2701 752 2818 753
rect 2377 744 2428 752
rect 2475 744 2509 752
rect 2377 732 2402 744
rect 2409 732 2428 744
rect 2482 742 2509 744
rect 2518 742 2739 752
rect 2774 749 2780 752
rect 2482 738 2739 742
rect 2377 724 2428 732
rect 2475 724 2739 738
rect 2783 744 2818 752
rect 2329 676 2348 710
rect 2393 716 2422 724
rect 2393 710 2410 716
rect 2393 708 2427 710
rect 2475 708 2491 724
rect 2492 714 2700 724
rect 2701 714 2717 724
rect 2765 720 2780 735
rect 2783 732 2784 744
rect 2791 732 2818 744
rect 2783 724 2818 732
rect 2783 723 2812 724
rect 2503 710 2717 714
rect 2518 708 2717 710
rect 2752 710 2765 720
rect 2783 710 2800 723
rect 2752 708 2800 710
rect 2394 704 2427 708
rect 2390 702 2427 704
rect 2390 701 2457 702
rect 2390 696 2421 701
rect 2427 696 2457 701
rect 2390 692 2457 696
rect 2363 689 2457 692
rect 2363 682 2412 689
rect 2363 676 2393 682
rect 2412 677 2417 682
rect 2329 660 2409 676
rect 2421 668 2457 689
rect 2518 684 2707 708
rect 2752 707 2799 708
rect 2765 702 2799 707
rect 2533 681 2707 684
rect 2526 678 2707 681
rect 2735 701 2799 702
rect 2329 658 2348 660
rect 2363 658 2397 660
rect 2329 642 2409 658
rect 2329 636 2348 642
rect 2045 610 2148 620
rect 1999 608 2148 610
rect 2169 608 2204 620
rect 1838 606 2000 608
rect 1850 586 1869 606
rect 1884 604 1914 606
rect 1733 578 1774 586
rect 1856 582 1869 586
rect 1921 590 2000 606
rect 2032 606 2204 608
rect 2032 590 2111 606
rect 2118 604 2148 606
rect 1696 568 1725 578
rect 1739 568 1768 578
rect 1783 568 1813 582
rect 1856 568 1899 582
rect 1921 578 2111 590
rect 2176 586 2182 606
rect 1906 568 1936 578
rect 1937 568 2095 578
rect 2099 568 2129 578
rect 2133 568 2163 582
rect 2191 568 2204 606
rect 2276 620 2305 636
rect 2319 620 2348 636
rect 2363 626 2393 642
rect 2421 620 2427 668
rect 2430 662 2449 668
rect 2464 662 2494 670
rect 2430 654 2494 662
rect 2430 638 2510 654
rect 2526 647 2588 678
rect 2604 647 2666 678
rect 2735 676 2784 701
rect 2799 676 2829 692
rect 2698 662 2728 670
rect 2735 668 2845 676
rect 2698 654 2743 662
rect 2430 636 2449 638
rect 2464 636 2510 638
rect 2430 620 2510 636
rect 2537 634 2572 647
rect 2613 644 2650 647
rect 2613 642 2655 644
rect 2542 631 2572 634
rect 2551 627 2558 631
rect 2558 626 2559 627
rect 2517 620 2527 626
rect 2276 612 2311 620
rect 2276 586 2277 612
rect 2284 586 2311 612
rect 2219 568 2249 582
rect 2276 578 2311 586
rect 2313 612 2354 620
rect 2313 586 2328 612
rect 2335 586 2354 612
rect 2418 608 2449 620
rect 2464 608 2567 620
rect 2579 610 2605 636
rect 2620 631 2650 642
rect 2682 638 2744 654
rect 2682 636 2728 638
rect 2682 620 2744 636
rect 2756 620 2762 668
rect 2765 660 2845 668
rect 2765 658 2784 660
rect 2799 658 2833 660
rect 2765 642 2845 658
rect 2765 620 2784 642
rect 2799 626 2829 642
rect 2857 636 2863 710
rect 2866 636 2885 780
rect 2900 636 2906 780
rect 2915 710 2928 780
rect 2980 776 3002 780
rect 2973 754 3002 768
rect 3055 754 3071 768
rect 3109 764 3115 766
rect 3122 764 3230 780
rect 3237 764 3243 766
rect 3251 764 3266 780
rect 3332 774 3351 777
rect 2973 752 3071 754
rect 3098 752 3266 764
rect 3281 754 3297 768
rect 3332 755 3354 774
rect 3364 768 3380 769
rect 3363 766 3380 768
rect 3364 761 3380 766
rect 3354 754 3360 755
rect 3363 754 3392 761
rect 3281 753 3392 754
rect 3281 752 3398 753
rect 2957 744 3008 752
rect 3055 744 3089 752
rect 2957 732 2982 744
rect 2989 732 3008 744
rect 3062 742 3089 744
rect 3098 742 3319 752
rect 3354 749 3360 752
rect 3062 738 3319 742
rect 2957 724 3008 732
rect 3055 724 3319 738
rect 3363 744 3398 752
rect 2909 676 2928 710
rect 2973 716 3002 724
rect 2973 710 2990 716
rect 2973 708 3007 710
rect 3055 708 3071 724
rect 3072 714 3280 724
rect 3281 714 3297 724
rect 3345 720 3360 735
rect 3363 732 3364 744
rect 3371 732 3398 744
rect 3363 724 3398 732
rect 3363 723 3392 724
rect 3083 710 3297 714
rect 3098 708 3297 710
rect 3332 710 3345 720
rect 3363 710 3380 723
rect 3332 708 3380 710
rect 2974 704 3007 708
rect 2970 702 3007 704
rect 2970 701 3037 702
rect 2970 696 3001 701
rect 3007 696 3037 701
rect 2970 692 3037 696
rect 2943 689 3037 692
rect 2943 682 2992 689
rect 2943 676 2973 682
rect 2992 677 2997 682
rect 2909 660 2989 676
rect 3001 668 3037 689
rect 3098 684 3287 708
rect 3332 707 3379 708
rect 3345 702 3379 707
rect 3113 681 3287 684
rect 3106 678 3287 681
rect 3315 701 3379 702
rect 2909 658 2928 660
rect 2943 658 2977 660
rect 2909 642 2989 658
rect 2909 636 2928 642
rect 2625 610 2728 620
rect 2579 608 2728 610
rect 2749 608 2784 620
rect 2418 606 2580 608
rect 2430 586 2449 606
rect 2464 604 2494 606
rect 2313 578 2354 586
rect 2436 582 2449 586
rect 2501 590 2580 606
rect 2612 606 2784 608
rect 2612 590 2691 606
rect 2698 604 2728 606
rect 2276 568 2305 578
rect 2319 568 2348 578
rect 2363 568 2393 582
rect 2436 568 2479 582
rect 2501 578 2691 590
rect 2756 586 2762 606
rect 2486 568 2516 578
rect 2517 568 2675 578
rect 2679 568 2709 578
rect 2713 568 2743 582
rect 2771 568 2784 606
rect 2856 620 2885 636
rect 2899 620 2928 636
rect 2943 626 2973 642
rect 3001 620 3007 668
rect 3010 662 3029 668
rect 3044 662 3074 670
rect 3010 654 3074 662
rect 3010 638 3090 654
rect 3106 647 3168 678
rect 3184 647 3246 678
rect 3315 676 3364 701
rect 3379 676 3409 692
rect 3278 662 3308 670
rect 3315 668 3425 676
rect 3278 654 3323 662
rect 3010 636 3029 638
rect 3044 636 3090 638
rect 3010 620 3090 636
rect 3117 634 3152 647
rect 3193 644 3230 647
rect 3193 642 3235 644
rect 3122 631 3152 634
rect 3131 627 3138 631
rect 3138 626 3139 627
rect 3097 620 3107 626
rect 2856 612 2891 620
rect 2856 586 2857 612
rect 2864 586 2891 612
rect 2799 568 2829 582
rect 2856 578 2891 586
rect 2893 612 2934 620
rect 2893 586 2908 612
rect 2915 586 2934 612
rect 2998 608 3029 620
rect 3044 608 3147 620
rect 3159 610 3185 636
rect 3200 631 3230 642
rect 3262 638 3324 654
rect 3262 636 3308 638
rect 3262 620 3324 636
rect 3336 620 3342 668
rect 3345 660 3425 668
rect 3345 658 3364 660
rect 3379 658 3413 660
rect 3345 642 3425 658
rect 3345 620 3364 642
rect 3379 626 3409 642
rect 3437 636 3443 710
rect 3446 636 3465 780
rect 3480 636 3486 780
rect 3495 710 3508 780
rect 3560 776 3582 780
rect 3553 754 3582 768
rect 3635 754 3651 768
rect 3689 764 3695 766
rect 3702 764 3810 780
rect 3817 764 3823 766
rect 3831 764 3846 780
rect 3912 774 3931 777
rect 3553 752 3651 754
rect 3678 752 3846 764
rect 3861 754 3877 768
rect 3912 755 3934 774
rect 3944 768 3960 769
rect 3943 766 3960 768
rect 3944 761 3960 766
rect 3934 754 3940 755
rect 3943 754 3972 761
rect 3861 753 3972 754
rect 3861 752 3978 753
rect 3537 744 3588 752
rect 3635 744 3669 752
rect 3537 732 3562 744
rect 3569 732 3588 744
rect 3642 742 3669 744
rect 3678 742 3899 752
rect 3934 749 3940 752
rect 3642 738 3899 742
rect 3537 724 3588 732
rect 3635 724 3899 738
rect 3943 744 3978 752
rect 3489 676 3508 710
rect 3553 716 3582 724
rect 3553 710 3570 716
rect 3553 708 3587 710
rect 3635 708 3651 724
rect 3652 714 3860 724
rect 3861 714 3877 724
rect 3925 720 3940 735
rect 3943 732 3944 744
rect 3951 732 3978 744
rect 3943 724 3978 732
rect 3943 723 3972 724
rect 3663 710 3877 714
rect 3678 708 3877 710
rect 3912 710 3925 720
rect 3943 710 3960 723
rect 3912 708 3960 710
rect 3554 704 3587 708
rect 3550 702 3587 704
rect 3550 701 3617 702
rect 3550 696 3581 701
rect 3587 696 3617 701
rect 3550 692 3617 696
rect 3523 689 3617 692
rect 3523 682 3572 689
rect 3523 676 3553 682
rect 3572 677 3577 682
rect 3489 660 3569 676
rect 3581 668 3617 689
rect 3678 684 3867 708
rect 3912 707 3959 708
rect 3925 702 3959 707
rect 3693 681 3867 684
rect 3686 678 3867 681
rect 3895 701 3959 702
rect 3489 658 3508 660
rect 3523 658 3557 660
rect 3489 642 3569 658
rect 3489 636 3508 642
rect 3205 610 3308 620
rect 3159 608 3308 610
rect 3329 608 3364 620
rect 2998 606 3160 608
rect 3010 586 3029 606
rect 3044 604 3074 606
rect 2893 578 2934 586
rect 3016 582 3029 586
rect 3081 590 3160 606
rect 3192 606 3364 608
rect 3192 590 3271 606
rect 3278 604 3308 606
rect 2856 568 2885 578
rect 2899 568 2928 578
rect 2943 568 2973 582
rect 3016 568 3059 582
rect 3081 578 3271 590
rect 3336 586 3342 606
rect 3066 568 3096 578
rect 3097 568 3255 578
rect 3259 568 3289 578
rect 3293 568 3323 582
rect 3351 568 3364 606
rect 3436 620 3465 636
rect 3479 620 3508 636
rect 3523 626 3553 642
rect 3581 620 3587 668
rect 3590 662 3609 668
rect 3624 662 3654 670
rect 3590 654 3654 662
rect 3590 638 3670 654
rect 3686 647 3748 678
rect 3764 647 3826 678
rect 3895 676 3944 701
rect 3959 676 3989 692
rect 3858 662 3888 670
rect 3895 668 4005 676
rect 3858 654 3903 662
rect 3590 636 3609 638
rect 3624 636 3670 638
rect 3590 620 3670 636
rect 3697 634 3732 647
rect 3773 644 3810 647
rect 3773 642 3815 644
rect 3702 631 3732 634
rect 3711 627 3718 631
rect 3718 626 3719 627
rect 3677 620 3687 626
rect 3436 612 3471 620
rect 3436 586 3437 612
rect 3444 586 3471 612
rect 3379 568 3409 582
rect 3436 578 3471 586
rect 3473 612 3514 620
rect 3473 586 3488 612
rect 3495 586 3514 612
rect 3578 608 3609 620
rect 3624 608 3727 620
rect 3739 610 3765 636
rect 3780 631 3810 642
rect 3842 638 3904 654
rect 3842 636 3888 638
rect 3842 620 3904 636
rect 3916 620 3922 668
rect 3925 660 4005 668
rect 3925 658 3944 660
rect 3959 658 3993 660
rect 3925 642 4005 658
rect 3925 620 3944 642
rect 3959 626 3989 642
rect 4017 636 4023 710
rect 4026 636 4045 780
rect 4060 636 4066 780
rect 4075 710 4088 780
rect 4140 776 4162 780
rect 4133 754 4162 768
rect 4215 754 4231 768
rect 4269 764 4275 766
rect 4282 764 4390 780
rect 4397 764 4403 766
rect 4411 764 4426 780
rect 4492 774 4511 777
rect 4133 752 4231 754
rect 4258 752 4426 764
rect 4441 754 4457 768
rect 4492 755 4514 774
rect 4524 768 4540 769
rect 4523 766 4540 768
rect 4524 761 4540 766
rect 4514 754 4520 755
rect 4523 754 4552 761
rect 4441 753 4552 754
rect 4441 752 4558 753
rect 4117 744 4168 752
rect 4215 744 4249 752
rect 4117 732 4142 744
rect 4149 732 4168 744
rect 4222 742 4249 744
rect 4258 742 4479 752
rect 4514 749 4520 752
rect 4222 738 4479 742
rect 4117 724 4168 732
rect 4215 724 4479 738
rect 4523 744 4558 752
rect 4069 676 4088 710
rect 4133 716 4162 724
rect 4133 710 4150 716
rect 4133 708 4167 710
rect 4215 708 4231 724
rect 4232 714 4440 724
rect 4441 714 4457 724
rect 4505 720 4520 735
rect 4523 732 4524 744
rect 4531 732 4558 744
rect 4523 724 4558 732
rect 4523 723 4552 724
rect 4243 710 4457 714
rect 4258 708 4457 710
rect 4492 710 4505 720
rect 4523 710 4540 723
rect 4492 708 4540 710
rect 4134 704 4167 708
rect 4130 702 4167 704
rect 4130 701 4197 702
rect 4130 696 4161 701
rect 4167 696 4197 701
rect 4130 692 4197 696
rect 4103 689 4197 692
rect 4103 682 4152 689
rect 4103 676 4133 682
rect 4152 677 4157 682
rect 4069 660 4149 676
rect 4161 668 4197 689
rect 4258 684 4447 708
rect 4492 707 4539 708
rect 4505 702 4539 707
rect 4273 681 4447 684
rect 4266 678 4447 681
rect 4475 701 4539 702
rect 4069 658 4088 660
rect 4103 658 4137 660
rect 4069 642 4149 658
rect 4069 636 4088 642
rect 3785 610 3888 620
rect 3739 608 3888 610
rect 3909 608 3944 620
rect 3578 606 3740 608
rect 3590 586 3609 606
rect 3624 604 3654 606
rect 3473 578 3514 586
rect 3596 582 3609 586
rect 3661 590 3740 606
rect 3772 606 3944 608
rect 3772 590 3851 606
rect 3858 604 3888 606
rect 3436 568 3465 578
rect 3479 568 3508 578
rect 3523 568 3553 582
rect 3596 568 3639 582
rect 3661 578 3851 590
rect 3916 586 3922 606
rect 3646 568 3676 578
rect 3677 568 3835 578
rect 3839 568 3869 578
rect 3873 568 3903 582
rect 3931 568 3944 606
rect 4016 620 4045 636
rect 4059 620 4088 636
rect 4103 626 4133 642
rect 4161 620 4167 668
rect 4170 662 4189 668
rect 4204 662 4234 670
rect 4170 654 4234 662
rect 4170 638 4250 654
rect 4266 647 4328 678
rect 4344 647 4406 678
rect 4475 676 4524 701
rect 4539 676 4569 692
rect 4438 662 4468 670
rect 4475 668 4585 676
rect 4438 654 4483 662
rect 4170 636 4189 638
rect 4204 636 4250 638
rect 4170 620 4250 636
rect 4277 634 4312 647
rect 4353 644 4390 647
rect 4353 642 4395 644
rect 4282 631 4312 634
rect 4291 627 4298 631
rect 4298 626 4299 627
rect 4257 620 4267 626
rect 4016 612 4051 620
rect 4016 586 4017 612
rect 4024 586 4051 612
rect 3959 568 3989 582
rect 4016 578 4051 586
rect 4053 612 4094 620
rect 4053 586 4068 612
rect 4075 586 4094 612
rect 4158 608 4189 620
rect 4204 608 4307 620
rect 4319 610 4345 636
rect 4360 631 4390 642
rect 4422 638 4484 654
rect 4422 636 4468 638
rect 4422 620 4484 636
rect 4496 620 4502 668
rect 4505 660 4585 668
rect 4505 658 4524 660
rect 4539 658 4573 660
rect 4505 642 4585 658
rect 4505 620 4524 642
rect 4539 626 4569 642
rect 4597 636 4603 710
rect 4606 636 4625 780
rect 4640 636 4646 780
rect 4655 710 4668 780
rect 4720 776 4742 780
rect 4713 754 4742 768
rect 4795 754 4811 768
rect 4849 765 4855 766
rect 4862 765 4970 780
rect 4977 765 4983 766
rect 4991 765 5006 780
rect 5072 774 5091 777
rect 4713 752 4811 754
rect 4838 752 5006 765
rect 5021 754 5037 768
rect 5072 755 5094 774
rect 5104 768 5120 769
rect 5103 766 5120 768
rect 5104 761 5120 766
rect 5094 754 5100 755
rect 5103 754 5132 761
rect 5021 753 5132 754
rect 5021 752 5138 753
rect 4697 744 4748 752
rect 4795 744 4829 752
rect 4697 732 4722 744
rect 4729 732 4748 744
rect 4802 742 4829 744
rect 4838 742 5059 752
rect 5094 749 5100 752
rect 4802 738 5059 742
rect 4697 724 4748 732
rect 4795 724 5059 738
rect 5103 744 5138 752
rect 4649 676 4668 710
rect 4713 716 4742 724
rect 4713 710 4730 716
rect 4713 708 4747 710
rect 4795 708 4811 724
rect 4812 714 5020 724
rect 5021 714 5037 724
rect 5085 720 5100 735
rect 5103 732 5104 744
rect 5111 732 5138 744
rect 5103 724 5138 732
rect 5103 723 5132 724
rect 4823 710 5037 714
rect 4838 708 5037 710
rect 5072 710 5085 720
rect 5103 710 5120 723
rect 5072 708 5120 710
rect 4714 704 4747 708
rect 4710 702 4747 704
rect 4710 701 4777 702
rect 4710 696 4741 701
rect 4747 696 4777 701
rect 4710 692 4777 696
rect 4683 689 4777 692
rect 4683 682 4732 689
rect 4683 676 4713 682
rect 4732 677 4737 682
rect 4649 660 4729 676
rect 4741 668 4777 689
rect 4838 684 5027 708
rect 5072 707 5119 708
rect 5085 702 5119 707
rect 4853 681 5027 684
rect 4846 678 5027 681
rect 5055 701 5119 702
rect 4649 658 4668 660
rect 4683 658 4717 660
rect 4649 642 4729 658
rect 4649 636 4668 642
rect 4365 610 4468 620
rect 4319 608 4468 610
rect 4489 608 4524 620
rect 4158 606 4320 608
rect 4170 586 4189 606
rect 4204 604 4234 606
rect 4053 578 4094 586
rect 4176 582 4189 586
rect 4241 590 4320 606
rect 4352 606 4524 608
rect 4352 590 4431 606
rect 4438 604 4468 606
rect 4016 568 4045 578
rect 4059 568 4088 578
rect 4103 568 4133 582
rect 4176 568 4219 582
rect 4241 578 4431 590
rect 4496 586 4502 606
rect 4226 568 4256 578
rect 4257 568 4415 578
rect 4419 568 4449 578
rect 4453 568 4483 582
rect 4511 568 4524 606
rect 4596 620 4625 636
rect 4639 620 4668 636
rect 4683 626 4713 642
rect 4741 620 4747 668
rect 4750 662 4769 668
rect 4784 662 4814 670
rect 4750 654 4814 662
rect 4750 638 4830 654
rect 4846 647 4908 678
rect 4924 647 4986 678
rect 5055 676 5104 701
rect 5119 676 5149 692
rect 5018 662 5048 670
rect 5055 668 5165 676
rect 5018 654 5063 662
rect 4750 636 4769 638
rect 4784 636 4830 638
rect 4750 620 4830 636
rect 4857 634 4892 647
rect 4933 644 4970 647
rect 4933 642 4975 644
rect 4862 631 4892 634
rect 4871 627 4878 631
rect 4878 626 4879 627
rect 4837 620 4847 626
rect 4596 612 4631 620
rect 4596 586 4597 612
rect 4604 586 4631 612
rect 4539 568 4569 582
rect 4596 578 4631 586
rect 4633 612 4674 620
rect 4633 586 4648 612
rect 4655 586 4674 612
rect 4738 608 4769 620
rect 4784 608 4887 620
rect 4899 610 4925 636
rect 4940 631 4970 642
rect 5002 638 5064 654
rect 5002 636 5048 638
rect 5002 620 5064 636
rect 5076 620 5082 668
rect 5085 660 5165 668
rect 5085 658 5104 660
rect 5119 658 5153 660
rect 5085 642 5165 658
rect 5085 620 5104 642
rect 5119 626 5149 642
rect 5177 636 5183 710
rect 5186 636 5205 780
rect 5220 636 5226 780
rect 5235 710 5248 780
rect 5300 776 5322 780
rect 5293 754 5322 768
rect 5375 754 5391 768
rect 5429 765 5435 766
rect 5442 765 5550 780
rect 5557 765 5563 766
rect 5571 765 5586 780
rect 5652 774 5671 777
rect 5293 752 5391 754
rect 5418 752 5586 765
rect 5601 754 5617 768
rect 5652 755 5674 774
rect 5684 768 5700 769
rect 5683 766 5700 768
rect 5684 761 5700 766
rect 5674 754 5680 755
rect 5683 754 5712 761
rect 5601 753 5712 754
rect 5601 752 5718 753
rect 5277 744 5328 752
rect 5375 744 5409 752
rect 5277 732 5302 744
rect 5309 732 5328 744
rect 5382 742 5409 744
rect 5418 742 5639 752
rect 5674 749 5680 752
rect 5382 738 5639 742
rect 5277 724 5328 732
rect 5375 724 5639 738
rect 5683 744 5718 752
rect 5229 676 5248 710
rect 5293 716 5322 724
rect 5293 710 5310 716
rect 5293 708 5327 710
rect 5375 708 5391 724
rect 5392 714 5600 724
rect 5601 714 5617 724
rect 5665 720 5680 735
rect 5683 732 5684 744
rect 5691 732 5718 744
rect 5683 724 5718 732
rect 5683 723 5712 724
rect 5403 710 5617 714
rect 5418 708 5617 710
rect 5652 710 5665 720
rect 5683 710 5700 723
rect 5652 708 5700 710
rect 5294 704 5327 708
rect 5290 702 5327 704
rect 5290 701 5357 702
rect 5290 696 5321 701
rect 5327 696 5357 701
rect 5290 692 5357 696
rect 5263 689 5357 692
rect 5263 682 5312 689
rect 5263 676 5293 682
rect 5312 677 5317 682
rect 5229 660 5309 676
rect 5321 668 5357 689
rect 5418 684 5607 708
rect 5652 707 5699 708
rect 5665 702 5699 707
rect 5433 681 5607 684
rect 5426 678 5607 681
rect 5635 701 5699 702
rect 5229 658 5248 660
rect 5263 658 5297 660
rect 5229 642 5309 658
rect 5229 636 5248 642
rect 4945 610 5048 620
rect 4899 608 5048 610
rect 5069 608 5104 620
rect 4738 606 4900 608
rect 4750 586 4769 606
rect 4784 604 4814 606
rect 4633 578 4674 586
rect 4756 583 4769 586
rect 4821 590 4900 606
rect 4932 606 5104 608
rect 4932 590 5011 606
rect 5018 604 5048 606
rect 4596 568 4625 578
rect 4639 568 4668 578
rect 4683 568 4713 583
rect 4756 579 4799 583
rect 4821 579 5011 590
rect 5076 586 5082 606
rect 5033 579 5063 583
rect 4756 578 5063 579
rect 4756 568 4799 578
rect 4806 568 4836 578
rect 4837 568 4995 578
rect 4999 568 5029 578
rect 5033 568 5063 578
rect 5091 568 5104 606
rect 5176 620 5205 636
rect 5219 620 5248 636
rect 5263 626 5293 642
rect 5321 620 5327 668
rect 5330 662 5349 668
rect 5364 662 5394 670
rect 5330 654 5394 662
rect 5330 638 5410 654
rect 5426 647 5488 678
rect 5504 647 5566 678
rect 5635 676 5684 701
rect 5699 676 5729 692
rect 5598 662 5628 670
rect 5635 668 5745 676
rect 5598 654 5643 662
rect 5330 636 5349 638
rect 5364 636 5410 638
rect 5330 620 5410 636
rect 5437 634 5472 647
rect 5513 644 5550 647
rect 5513 642 5555 644
rect 5442 631 5472 634
rect 5451 627 5458 631
rect 5458 626 5459 627
rect 5417 620 5427 626
rect 5176 612 5211 620
rect 5176 586 5177 612
rect 5184 586 5211 612
rect 5119 568 5149 583
rect 5176 578 5211 586
rect 5213 612 5254 620
rect 5213 586 5228 612
rect 5235 586 5254 612
rect 5318 608 5349 620
rect 5364 608 5467 620
rect 5479 610 5505 636
rect 5520 631 5550 642
rect 5582 638 5644 654
rect 5582 636 5628 638
rect 5582 620 5644 636
rect 5656 620 5662 668
rect 5665 660 5745 668
rect 5665 658 5684 660
rect 5699 658 5733 660
rect 5665 642 5745 658
rect 5665 620 5684 642
rect 5699 626 5729 642
rect 5757 636 5763 710
rect 5766 636 5785 780
rect 5800 636 5806 780
rect 5815 710 5828 780
rect 5880 776 5902 780
rect 5873 754 5902 768
rect 5955 754 5971 768
rect 6009 765 6015 766
rect 6022 765 6130 780
rect 6137 765 6143 766
rect 6151 765 6166 780
rect 6232 774 6251 777
rect 5873 752 5971 754
rect 5998 752 6166 765
rect 6181 754 6197 768
rect 6232 755 6254 774
rect 6264 768 6280 769
rect 6263 766 6280 768
rect 6264 761 6280 766
rect 6254 754 6260 755
rect 6263 754 6292 761
rect 6181 753 6292 754
rect 6181 752 6298 753
rect 5857 744 5908 752
rect 5955 744 5989 752
rect 5857 732 5882 744
rect 5889 732 5908 744
rect 5962 742 5989 744
rect 5998 742 6219 752
rect 6254 749 6260 752
rect 5962 738 6219 742
rect 5857 724 5908 732
rect 5955 724 6219 738
rect 6263 744 6298 752
rect 5809 676 5828 710
rect 5873 716 5902 724
rect 5873 710 5890 716
rect 5873 708 5907 710
rect 5955 708 5971 724
rect 5972 714 6180 724
rect 6181 714 6197 724
rect 6245 720 6260 735
rect 6263 732 6264 744
rect 6271 732 6298 744
rect 6263 724 6298 732
rect 6263 723 6292 724
rect 5983 710 6197 714
rect 5998 708 6197 710
rect 6232 710 6245 720
rect 6263 710 6280 723
rect 6232 708 6280 710
rect 5874 704 5907 708
rect 5870 702 5907 704
rect 5870 701 5937 702
rect 5870 696 5901 701
rect 5907 696 5937 701
rect 5870 692 5937 696
rect 5843 689 5937 692
rect 5843 682 5892 689
rect 5843 676 5873 682
rect 5892 677 5897 682
rect 5809 660 5889 676
rect 5901 668 5937 689
rect 5998 684 6187 708
rect 6232 707 6279 708
rect 6245 702 6279 707
rect 6013 681 6187 684
rect 6006 678 6187 681
rect 6215 701 6279 702
rect 5809 658 5828 660
rect 5843 658 5877 660
rect 5809 642 5889 658
rect 5809 636 5828 642
rect 5525 610 5628 620
rect 5479 608 5628 610
rect 5649 608 5684 620
rect 5318 606 5480 608
rect 5330 586 5349 606
rect 5364 604 5394 606
rect 5213 578 5254 586
rect 5336 583 5349 586
rect 5401 590 5480 606
rect 5512 606 5684 608
rect 5512 590 5591 606
rect 5598 604 5628 606
rect 5176 568 5205 578
rect 5219 568 5248 578
rect 5263 568 5293 583
rect 5336 579 5379 583
rect 5401 579 5591 590
rect 5656 586 5662 606
rect 5613 579 5643 583
rect 5336 578 5643 579
rect 5336 568 5379 578
rect 5386 568 5416 578
rect 5417 568 5575 578
rect 5579 568 5609 578
rect 5613 568 5643 578
rect 5671 568 5684 606
rect 5756 620 5785 636
rect 5799 620 5828 636
rect 5843 626 5873 642
rect 5901 620 5907 668
rect 5910 662 5929 668
rect 5944 662 5974 670
rect 5910 654 5974 662
rect 5910 638 5990 654
rect 6006 647 6068 678
rect 6084 647 6146 678
rect 6215 676 6264 701
rect 6279 676 6309 692
rect 6178 662 6208 670
rect 6215 668 6325 676
rect 6178 654 6223 662
rect 5910 636 5929 638
rect 5944 636 5990 638
rect 5910 620 5990 636
rect 6017 634 6052 647
rect 6093 644 6130 647
rect 6093 642 6135 644
rect 6022 631 6052 634
rect 6031 627 6038 631
rect 6038 626 6039 627
rect 5997 620 6007 626
rect 5756 612 5791 620
rect 5756 586 5757 612
rect 5764 586 5791 612
rect 5699 568 5729 583
rect 5756 578 5791 586
rect 5793 612 5834 620
rect 5793 586 5808 612
rect 5815 586 5834 612
rect 5898 608 5929 620
rect 5944 608 6047 620
rect 6059 610 6085 636
rect 6100 631 6130 642
rect 6162 638 6224 654
rect 6162 636 6208 638
rect 6162 620 6224 636
rect 6236 620 6242 668
rect 6245 660 6325 668
rect 6245 658 6264 660
rect 6279 658 6313 660
rect 6245 642 6325 658
rect 6245 620 6264 642
rect 6279 626 6309 642
rect 6337 636 6343 710
rect 6346 636 6365 780
rect 6380 636 6386 780
rect 6395 710 6408 780
rect 6460 776 6482 780
rect 6453 754 6482 768
rect 6535 754 6551 768
rect 6589 765 6595 766
rect 6602 765 6710 780
rect 6717 765 6723 766
rect 6731 765 6746 780
rect 6812 774 6831 777
rect 6453 752 6551 754
rect 6578 752 6746 765
rect 6761 754 6777 768
rect 6812 755 6834 774
rect 6844 768 6860 769
rect 6843 766 6860 768
rect 6844 761 6860 766
rect 6834 754 6840 755
rect 6843 754 6872 761
rect 6761 753 6872 754
rect 6761 752 6878 753
rect 6437 744 6488 752
rect 6535 744 6569 752
rect 6437 732 6462 744
rect 6469 732 6488 744
rect 6542 742 6569 744
rect 6578 742 6799 752
rect 6834 749 6840 752
rect 6542 738 6799 742
rect 6437 724 6488 732
rect 6535 724 6799 738
rect 6843 744 6878 752
rect 6389 676 6408 710
rect 6453 716 6482 724
rect 6453 710 6470 716
rect 6453 708 6487 710
rect 6535 708 6551 724
rect 6552 714 6760 724
rect 6761 714 6777 724
rect 6825 720 6840 735
rect 6843 732 6844 744
rect 6851 732 6878 744
rect 6843 724 6878 732
rect 6843 723 6872 724
rect 6563 710 6777 714
rect 6578 708 6777 710
rect 6812 710 6825 720
rect 6843 710 6860 723
rect 6812 708 6860 710
rect 6454 704 6487 708
rect 6450 702 6487 704
rect 6450 701 6517 702
rect 6450 696 6481 701
rect 6487 696 6517 701
rect 6450 692 6517 696
rect 6423 689 6517 692
rect 6423 682 6472 689
rect 6423 676 6453 682
rect 6472 677 6477 682
rect 6389 660 6469 676
rect 6481 668 6517 689
rect 6578 684 6767 708
rect 6812 707 6859 708
rect 6825 702 6859 707
rect 6593 681 6767 684
rect 6586 678 6767 681
rect 6795 701 6859 702
rect 6389 658 6408 660
rect 6423 658 6457 660
rect 6389 642 6469 658
rect 6389 636 6408 642
rect 6105 610 6208 620
rect 6059 608 6208 610
rect 6229 608 6264 620
rect 5898 606 6060 608
rect 5910 586 5929 606
rect 5944 604 5974 606
rect 5793 578 5834 586
rect 5916 583 5929 586
rect 5981 590 6060 606
rect 6092 606 6264 608
rect 6092 590 6171 606
rect 6178 604 6208 606
rect 5756 568 5785 578
rect 5799 568 5828 578
rect 5843 568 5873 583
rect 5916 579 5959 583
rect 5981 579 6171 590
rect 6236 586 6242 606
rect 6193 579 6223 583
rect 5916 578 6223 579
rect 5916 568 5959 578
rect 5966 568 5996 578
rect 5997 568 6155 578
rect 6159 568 6189 578
rect 6193 568 6223 578
rect 6251 568 6264 606
rect 6336 620 6365 636
rect 6379 620 6408 636
rect 6423 626 6453 642
rect 6481 620 6487 668
rect 6490 662 6509 668
rect 6524 662 6554 670
rect 6490 654 6554 662
rect 6490 638 6570 654
rect 6586 647 6648 678
rect 6664 647 6726 678
rect 6795 676 6844 701
rect 6859 676 6889 692
rect 6758 662 6788 670
rect 6795 668 6905 676
rect 6758 654 6803 662
rect 6490 636 6509 638
rect 6524 636 6570 638
rect 6490 620 6570 636
rect 6597 634 6632 647
rect 6673 644 6710 647
rect 6673 642 6715 644
rect 6602 631 6632 634
rect 6611 627 6618 631
rect 6618 626 6619 627
rect 6577 620 6587 626
rect 6336 612 6371 620
rect 6336 586 6337 612
rect 6344 586 6371 612
rect 6279 568 6309 583
rect 6336 578 6371 586
rect 6373 612 6414 620
rect 6373 586 6388 612
rect 6395 586 6414 612
rect 6478 608 6509 620
rect 6524 608 6627 620
rect 6639 610 6665 636
rect 6680 631 6710 642
rect 6742 638 6804 654
rect 6742 636 6788 638
rect 6742 620 6804 636
rect 6816 620 6822 668
rect 6825 660 6905 668
rect 6825 658 6844 660
rect 6859 658 6893 660
rect 6825 642 6905 658
rect 6825 620 6844 642
rect 6859 626 6889 642
rect 6917 636 6923 710
rect 6926 636 6945 780
rect 6960 636 6966 780
rect 6975 710 6988 780
rect 7040 776 7062 780
rect 7033 754 7062 768
rect 7115 754 7131 768
rect 7169 765 7175 766
rect 7182 765 7290 780
rect 7297 765 7303 766
rect 7311 765 7326 780
rect 7392 774 7411 777
rect 7033 752 7131 754
rect 7158 752 7326 765
rect 7341 754 7357 768
rect 7392 755 7414 774
rect 7424 768 7440 769
rect 7423 766 7440 768
rect 7424 761 7440 766
rect 7414 754 7420 755
rect 7423 754 7452 761
rect 7341 753 7452 754
rect 7341 752 7458 753
rect 7017 744 7068 752
rect 7115 744 7149 752
rect 7017 732 7042 744
rect 7049 732 7068 744
rect 7122 742 7149 744
rect 7158 742 7379 752
rect 7414 749 7420 752
rect 7122 738 7379 742
rect 7017 724 7068 732
rect 7115 724 7379 738
rect 7423 744 7458 752
rect 6969 676 6988 710
rect 7033 716 7062 724
rect 7033 710 7050 716
rect 7033 708 7067 710
rect 7115 708 7131 724
rect 7132 714 7340 724
rect 7341 714 7357 724
rect 7405 720 7420 735
rect 7423 732 7424 744
rect 7431 732 7458 744
rect 7423 724 7458 732
rect 7423 723 7452 724
rect 7151 710 7357 714
rect 7158 708 7357 710
rect 7392 710 7405 720
rect 7423 710 7440 723
rect 7392 708 7440 710
rect 7034 704 7067 708
rect 7030 702 7067 704
rect 7030 701 7097 702
rect 7030 696 7061 701
rect 7067 696 7097 701
rect 7030 692 7097 696
rect 7003 689 7097 692
rect 7003 682 7052 689
rect 7003 676 7033 682
rect 7052 677 7057 682
rect 6969 660 7049 676
rect 7061 668 7097 689
rect 7158 684 7347 708
rect 7392 707 7439 708
rect 7405 702 7439 707
rect 7173 681 7347 684
rect 7166 678 7347 681
rect 7375 701 7439 702
rect 6969 658 6988 660
rect 7003 658 7037 660
rect 6969 642 7049 658
rect 6969 636 6988 642
rect 6685 610 6788 620
rect 6639 608 6788 610
rect 6809 608 6844 620
rect 6478 606 6640 608
rect 6490 586 6509 606
rect 6524 604 6554 606
rect 6373 578 6414 586
rect 6496 583 6509 586
rect 6561 590 6640 606
rect 6672 606 6844 608
rect 6672 590 6751 606
rect 6758 604 6788 606
rect 6336 568 6365 578
rect 6379 568 6408 578
rect 6423 568 6453 583
rect 6496 579 6539 583
rect 6561 579 6751 590
rect 6816 586 6822 606
rect 6773 579 6803 583
rect 6496 578 6803 579
rect 6496 568 6539 578
rect 6546 568 6576 578
rect 6577 568 6735 578
rect 6739 568 6769 578
rect 6773 568 6803 578
rect 6831 568 6844 606
rect 6916 620 6945 636
rect 6959 620 6988 636
rect 7003 626 7033 642
rect 7061 620 7067 668
rect 7070 662 7089 668
rect 7104 662 7134 670
rect 7070 654 7134 662
rect 7070 638 7150 654
rect 7166 647 7228 678
rect 7244 647 7306 678
rect 7375 676 7424 701
rect 7439 676 7469 692
rect 7338 662 7368 670
rect 7375 668 7485 676
rect 7338 654 7383 662
rect 7070 636 7089 638
rect 7104 636 7150 638
rect 7070 620 7150 636
rect 7177 634 7212 647
rect 7253 644 7290 647
rect 7253 642 7295 644
rect 7182 631 7212 634
rect 7191 627 7198 631
rect 7198 626 7199 627
rect 7157 620 7167 626
rect 6916 612 6951 620
rect 6916 586 6917 612
rect 6924 586 6951 612
rect 6859 568 6889 583
rect 6916 578 6951 586
rect 6953 612 6994 620
rect 6953 586 6968 612
rect 6975 586 6994 612
rect 7058 608 7089 620
rect 7104 608 7207 620
rect 7219 610 7245 636
rect 7260 631 7290 642
rect 7322 638 7384 654
rect 7322 636 7368 638
rect 7322 620 7384 636
rect 7396 620 7402 668
rect 7405 660 7485 668
rect 7405 658 7424 660
rect 7439 658 7473 660
rect 7405 642 7485 658
rect 7405 620 7424 642
rect 7439 626 7469 642
rect 7497 636 7503 710
rect 7506 636 7525 780
rect 7540 636 7546 780
rect 7555 710 7568 780
rect 7620 776 7642 780
rect 7613 754 7642 768
rect 7695 754 7711 768
rect 7749 765 7755 766
rect 7762 765 7870 780
rect 7877 765 7883 766
rect 7891 765 7906 780
rect 7972 774 7991 777
rect 7613 752 7711 754
rect 7738 752 7906 765
rect 7921 754 7937 768
rect 7972 755 7994 774
rect 8004 768 8020 769
rect 8003 766 8020 768
rect 8004 761 8020 766
rect 7994 754 8000 755
rect 8003 754 8032 761
rect 7921 753 8032 754
rect 7921 752 8038 753
rect 7597 744 7648 752
rect 7695 744 7729 752
rect 7597 732 7622 744
rect 7629 732 7648 744
rect 7702 742 7729 744
rect 7738 742 7959 752
rect 7994 749 8000 752
rect 7702 738 7959 742
rect 7597 724 7648 732
rect 7695 724 7959 738
rect 8003 744 8038 752
rect 7549 676 7568 710
rect 7613 716 7642 724
rect 7613 710 7630 716
rect 7613 708 7647 710
rect 7695 708 7711 724
rect 7712 714 7920 724
rect 7921 714 7937 724
rect 7985 720 8000 735
rect 8003 732 8004 744
rect 8011 732 8038 744
rect 8003 724 8038 732
rect 8003 723 8032 724
rect 7723 710 7937 714
rect 7738 708 7937 710
rect 7972 710 7985 720
rect 8003 710 8020 723
rect 7972 708 8020 710
rect 7614 704 7647 708
rect 7610 702 7647 704
rect 7610 701 7677 702
rect 7610 696 7641 701
rect 7647 696 7677 701
rect 7610 692 7677 696
rect 7583 689 7677 692
rect 7583 682 7632 689
rect 7583 676 7613 682
rect 7632 677 7637 682
rect 7549 660 7629 676
rect 7641 668 7677 689
rect 7738 684 7927 708
rect 7972 707 8019 708
rect 7985 702 8019 707
rect 7753 681 7927 684
rect 7746 678 7927 681
rect 7955 701 8019 702
rect 7549 658 7568 660
rect 7583 658 7617 660
rect 7549 642 7629 658
rect 7549 636 7568 642
rect 7265 610 7368 620
rect 7219 608 7368 610
rect 7389 608 7424 620
rect 7058 606 7220 608
rect 7070 586 7089 606
rect 7104 604 7134 606
rect 6953 578 6994 586
rect 7076 583 7089 586
rect 7141 590 7220 606
rect 7252 606 7424 608
rect 7252 590 7331 606
rect 7338 604 7368 606
rect 6916 568 6945 578
rect 6959 568 6988 578
rect 7003 568 7033 583
rect 7076 579 7119 583
rect 7141 579 7331 590
rect 7396 586 7402 606
rect 7353 579 7383 583
rect 7076 578 7383 579
rect 7076 568 7119 578
rect 7126 568 7156 578
rect 7157 568 7315 578
rect 7319 568 7349 578
rect 7353 568 7383 578
rect 7411 568 7424 606
rect 7496 620 7525 636
rect 7539 620 7568 636
rect 7583 626 7613 642
rect 7641 620 7647 668
rect 7650 662 7669 668
rect 7684 662 7714 670
rect 7650 654 7714 662
rect 7650 638 7730 654
rect 7746 647 7808 678
rect 7824 647 7886 678
rect 7955 676 8004 701
rect 8019 676 8049 692
rect 7918 662 7948 670
rect 7955 668 8065 676
rect 7918 654 7963 662
rect 7650 636 7669 638
rect 7684 636 7730 638
rect 7650 620 7730 636
rect 7757 634 7792 647
rect 7833 644 7870 647
rect 7833 642 7875 644
rect 7762 631 7792 634
rect 7771 627 7778 631
rect 7778 626 7779 627
rect 7737 620 7747 626
rect 7496 612 7531 620
rect 7496 586 7497 612
rect 7504 586 7531 612
rect 7439 568 7469 583
rect 7496 578 7531 586
rect 7533 612 7574 620
rect 7533 586 7548 612
rect 7555 586 7574 612
rect 7638 608 7669 620
rect 7684 608 7787 620
rect 7799 610 7825 636
rect 7840 631 7870 642
rect 7902 638 7964 654
rect 7902 636 7948 638
rect 7902 620 7964 636
rect 7976 620 7982 668
rect 7985 660 8065 668
rect 7985 658 8004 660
rect 8019 658 8053 660
rect 7985 642 8065 658
rect 7985 620 8004 642
rect 8019 626 8049 642
rect 8077 636 8083 710
rect 8086 636 8105 780
rect 8120 636 8126 780
rect 8135 710 8148 780
rect 8200 776 8222 780
rect 8193 754 8222 768
rect 8275 754 8291 768
rect 8329 765 8335 766
rect 8342 765 8450 780
rect 8457 765 8463 766
rect 8471 765 8486 780
rect 8552 774 8571 777
rect 8193 752 8291 754
rect 8318 752 8486 765
rect 8501 754 8517 768
rect 8552 755 8574 774
rect 8584 768 8600 769
rect 8583 766 8600 768
rect 8584 761 8600 766
rect 8574 754 8580 755
rect 8583 754 8612 761
rect 8501 753 8612 754
rect 8501 752 8618 753
rect 8177 744 8228 752
rect 8275 744 8309 752
rect 8177 732 8202 744
rect 8209 732 8228 744
rect 8282 742 8309 744
rect 8318 742 8539 752
rect 8574 749 8580 752
rect 8282 738 8539 742
rect 8177 724 8228 732
rect 8275 724 8539 738
rect 8583 744 8618 752
rect 8129 676 8148 710
rect 8193 716 8222 724
rect 8193 710 8210 716
rect 8193 708 8227 710
rect 8275 708 8291 724
rect 8292 714 8500 724
rect 8501 714 8517 724
rect 8565 720 8580 735
rect 8583 732 8584 744
rect 8591 732 8618 744
rect 8583 724 8618 732
rect 8583 723 8612 724
rect 8303 710 8517 714
rect 8318 708 8517 710
rect 8552 710 8565 720
rect 8583 710 8600 723
rect 8552 708 8600 710
rect 8194 704 8227 708
rect 8190 702 8227 704
rect 8190 701 8257 702
rect 8190 696 8221 701
rect 8227 696 8257 701
rect 8190 692 8257 696
rect 8163 689 8257 692
rect 8163 682 8212 689
rect 8163 676 8193 682
rect 8212 677 8217 682
rect 8129 660 8209 676
rect 8221 668 8257 689
rect 8318 684 8507 708
rect 8552 707 8599 708
rect 8565 702 8599 707
rect 8333 681 8507 684
rect 8326 678 8507 681
rect 8535 701 8599 702
rect 8129 658 8148 660
rect 8163 658 8197 660
rect 8129 642 8209 658
rect 8129 636 8148 642
rect 7845 610 7948 620
rect 7799 608 7948 610
rect 7969 608 8004 620
rect 7638 606 7800 608
rect 7650 586 7669 606
rect 7684 604 7714 606
rect 7533 578 7574 586
rect 7656 583 7669 586
rect 7721 590 7800 606
rect 7832 606 8004 608
rect 7832 590 7911 606
rect 7918 604 7948 606
rect 7496 568 7525 578
rect 7539 568 7568 578
rect 7583 568 7613 583
rect 7656 579 7699 583
rect 7721 579 7911 590
rect 7976 586 7982 606
rect 7933 579 7963 583
rect 7656 578 7963 579
rect 7656 568 7699 578
rect 7706 568 7736 578
rect 7737 568 7895 578
rect 7899 568 7929 578
rect 7933 568 7963 578
rect 7991 568 8004 606
rect 8076 620 8105 636
rect 8119 620 8148 636
rect 8163 626 8193 642
rect 8221 620 8227 668
rect 8230 662 8249 668
rect 8264 662 8294 670
rect 8230 654 8294 662
rect 8230 638 8310 654
rect 8326 647 8388 678
rect 8404 647 8466 678
rect 8535 676 8584 701
rect 8599 676 8629 692
rect 8498 662 8528 670
rect 8535 668 8645 676
rect 8498 654 8543 662
rect 8230 636 8249 638
rect 8264 636 8310 638
rect 8230 620 8310 636
rect 8337 634 8372 647
rect 8413 644 8450 647
rect 8413 642 8455 644
rect 8342 631 8372 634
rect 8351 627 8358 631
rect 8358 626 8359 627
rect 8317 620 8327 626
rect 8076 612 8111 620
rect 8076 586 8077 612
rect 8084 586 8111 612
rect 8019 568 8049 583
rect 8076 578 8111 586
rect 8113 612 8154 620
rect 8113 586 8128 612
rect 8135 586 8154 612
rect 8218 608 8249 620
rect 8264 608 8367 620
rect 8379 610 8405 636
rect 8420 631 8450 642
rect 8482 638 8544 654
rect 8482 636 8528 638
rect 8482 620 8544 636
rect 8556 620 8562 668
rect 8565 660 8645 668
rect 8565 658 8584 660
rect 8599 658 8633 660
rect 8565 642 8645 658
rect 8565 620 8584 642
rect 8599 626 8629 642
rect 8657 636 8663 710
rect 8666 636 8685 780
rect 8700 636 8706 780
rect 8715 710 8728 780
rect 8780 776 8802 780
rect 8773 754 8802 768
rect 8855 754 8871 768
rect 8909 765 8915 766
rect 8922 765 9030 780
rect 9037 765 9043 766
rect 9051 765 9066 780
rect 9132 774 9151 777
rect 8773 752 8871 754
rect 8898 752 9066 765
rect 9081 754 9097 768
rect 9132 755 9154 774
rect 9164 768 9180 769
rect 9163 766 9180 768
rect 9164 761 9180 766
rect 9154 754 9160 755
rect 9163 754 9192 761
rect 9081 753 9192 754
rect 9081 752 9198 753
rect 8757 744 8808 752
rect 8855 744 8889 752
rect 8757 732 8782 744
rect 8789 732 8808 744
rect 8862 742 8889 744
rect 8898 742 9119 752
rect 9154 749 9160 752
rect 8862 738 9119 742
rect 8757 724 8808 732
rect 8855 724 9119 738
rect 9163 744 9198 752
rect 8709 676 8728 710
rect 8773 716 8802 724
rect 8773 710 8790 716
rect 8773 708 8807 710
rect 8855 708 8871 724
rect 8872 714 9080 724
rect 9081 714 9097 724
rect 9145 720 9160 735
rect 9163 732 9164 744
rect 9171 732 9198 744
rect 9163 724 9198 732
rect 9163 723 9192 724
rect 8883 710 9097 714
rect 8898 708 9097 710
rect 9132 710 9145 720
rect 9163 710 9180 723
rect 9132 708 9180 710
rect 8774 704 8807 708
rect 8770 702 8807 704
rect 8770 701 8837 702
rect 8770 696 8801 701
rect 8807 696 8837 701
rect 8770 692 8837 696
rect 8743 689 8837 692
rect 8743 682 8792 689
rect 8743 676 8773 682
rect 8792 677 8797 682
rect 8709 660 8789 676
rect 8801 668 8837 689
rect 8898 684 9087 708
rect 9132 707 9179 708
rect 9145 702 9179 707
rect 8913 681 9087 684
rect 8906 678 9087 681
rect 9115 701 9179 702
rect 8709 658 8728 660
rect 8743 658 8777 660
rect 8709 642 8789 658
rect 8709 636 8728 642
rect 8425 610 8528 620
rect 8379 608 8528 610
rect 8549 608 8584 620
rect 8218 606 8380 608
rect 8230 586 8249 606
rect 8264 604 8294 606
rect 8113 578 8154 586
rect 8236 583 8249 586
rect 8301 590 8380 606
rect 8412 606 8584 608
rect 8412 590 8491 606
rect 8498 604 8528 606
rect 8076 568 8105 578
rect 8119 568 8148 578
rect 8163 568 8193 583
rect 8236 579 8279 583
rect 8301 579 8491 590
rect 8556 586 8562 606
rect 8513 579 8543 583
rect 8236 578 8543 579
rect 8236 568 8279 578
rect 8286 568 8316 578
rect 8317 568 8475 578
rect 8479 568 8509 578
rect 8513 568 8543 578
rect 8571 568 8584 606
rect 8656 620 8685 636
rect 8699 620 8728 636
rect 8743 626 8773 642
rect 8801 620 8807 668
rect 8810 662 8829 668
rect 8844 662 8874 670
rect 8810 654 8874 662
rect 8810 638 8890 654
rect 8906 647 8968 678
rect 8984 647 9046 678
rect 9115 676 9164 701
rect 9179 676 9209 692
rect 9078 662 9108 670
rect 9115 668 9225 676
rect 9078 654 9123 662
rect 8810 636 8829 638
rect 8844 636 8890 638
rect 8810 620 8890 636
rect 8917 634 8952 647
rect 8993 644 9030 647
rect 8993 642 9035 644
rect 8922 631 8952 634
rect 8931 627 8938 631
rect 8938 626 8939 627
rect 8897 620 8907 626
rect 8656 612 8691 620
rect 8656 586 8657 612
rect 8664 586 8691 612
rect 8599 568 8629 583
rect 8656 578 8691 586
rect 8693 612 8734 620
rect 8693 586 8708 612
rect 8715 586 8734 612
rect 8798 608 8829 620
rect 8844 608 8947 620
rect 8959 610 8985 636
rect 9000 631 9030 642
rect 9062 638 9124 654
rect 9062 636 9108 638
rect 9062 620 9124 636
rect 9136 620 9142 668
rect 9145 660 9225 668
rect 9145 658 9164 660
rect 9179 658 9213 660
rect 9145 642 9225 658
rect 9145 620 9164 642
rect 9179 626 9209 642
rect 9237 636 9243 710
rect 9246 636 9265 780
rect 9280 636 9286 780
rect 9295 710 9308 780
rect 9360 776 9382 780
rect 9353 754 9382 768
rect 9435 754 9451 768
rect 9489 765 9495 766
rect 9502 765 9610 780
rect 9617 765 9623 766
rect 9631 765 9646 780
rect 9712 774 9731 777
rect 9353 752 9451 754
rect 9478 752 9646 765
rect 9661 754 9677 768
rect 9712 755 9734 774
rect 9744 768 9760 769
rect 9743 766 9760 768
rect 9744 761 9760 766
rect 9734 754 9740 755
rect 9743 754 9772 761
rect 9661 753 9772 754
rect 9661 752 9778 753
rect 9337 744 9388 752
rect 9435 744 9469 752
rect 9337 732 9362 744
rect 9369 732 9388 744
rect 9442 742 9469 744
rect 9478 742 9699 752
rect 9734 749 9740 752
rect 9442 738 9699 742
rect 9337 724 9388 732
rect 9435 724 9699 738
rect 9743 744 9778 752
rect 9289 676 9308 710
rect 9353 716 9382 724
rect 9353 710 9370 716
rect 9353 708 9387 710
rect 9435 708 9451 724
rect 9452 714 9660 724
rect 9661 714 9677 724
rect 9725 720 9740 735
rect 9743 732 9744 744
rect 9751 732 9778 744
rect 9743 724 9778 732
rect 9743 723 9772 724
rect 9463 710 9677 714
rect 9478 708 9677 710
rect 9712 710 9725 720
rect 9743 710 9760 723
rect 9712 708 9760 710
rect 9354 704 9387 708
rect 9350 702 9387 704
rect 9350 701 9417 702
rect 9350 696 9381 701
rect 9387 696 9417 701
rect 9350 692 9417 696
rect 9323 689 9417 692
rect 9323 682 9372 689
rect 9323 676 9353 682
rect 9372 677 9377 682
rect 9289 660 9369 676
rect 9381 668 9417 689
rect 9478 684 9667 708
rect 9712 707 9759 708
rect 9725 702 9759 707
rect 9493 681 9667 684
rect 9486 678 9667 681
rect 9695 701 9759 702
rect 9289 658 9308 660
rect 9323 658 9357 660
rect 9289 642 9369 658
rect 9289 636 9308 642
rect 9005 610 9108 620
rect 8959 608 9108 610
rect 9129 608 9164 620
rect 8798 606 8960 608
rect 8810 586 8829 606
rect 8844 604 8874 606
rect 8693 578 8734 586
rect 8816 583 8829 586
rect 8881 590 8960 606
rect 8992 606 9164 608
rect 8992 590 9071 606
rect 9078 604 9108 606
rect 8656 568 8685 578
rect 8699 568 8728 578
rect 8743 568 8773 583
rect 8816 579 8859 583
rect 8881 579 9071 590
rect 9136 586 9142 606
rect 9093 579 9123 583
rect 8816 578 9123 579
rect 8816 568 8859 578
rect 8866 568 8896 578
rect 8897 568 9055 578
rect 9059 568 9089 578
rect 9093 568 9123 578
rect 9151 568 9164 606
rect 9236 620 9265 636
rect 9279 620 9308 636
rect 9323 626 9353 642
rect 9381 620 9387 668
rect 9390 662 9409 668
rect 9424 662 9454 670
rect 9390 654 9454 662
rect 9390 638 9470 654
rect 9486 647 9548 678
rect 9564 647 9626 678
rect 9695 676 9744 701
rect 9759 676 9789 692
rect 9658 662 9688 670
rect 9695 668 9805 676
rect 9658 654 9703 662
rect 9390 636 9409 638
rect 9424 636 9470 638
rect 9390 620 9470 636
rect 9497 634 9532 647
rect 9573 644 9610 647
rect 9573 642 9615 644
rect 9502 631 9532 634
rect 9511 627 9518 631
rect 9518 626 9519 627
rect 9477 620 9487 626
rect 9236 612 9271 620
rect 9236 586 9237 612
rect 9244 586 9271 612
rect 9179 568 9209 583
rect 9236 578 9271 586
rect 9273 612 9314 620
rect 9273 586 9288 612
rect 9295 586 9314 612
rect 9378 608 9409 620
rect 9424 608 9527 620
rect 9539 610 9565 636
rect 9580 631 9610 642
rect 9642 638 9704 654
rect 9642 636 9688 638
rect 9642 620 9704 636
rect 9716 620 9722 668
rect 9725 660 9805 668
rect 9725 658 9744 660
rect 9759 658 9793 660
rect 9725 642 9805 658
rect 9725 620 9744 642
rect 9759 626 9789 642
rect 9817 636 9823 710
rect 9826 636 9845 780
rect 9860 636 9866 780
rect 9875 710 9888 780
rect 9940 776 9962 780
rect 9933 754 9962 768
rect 10015 754 10031 768
rect 10069 765 10075 766
rect 10082 765 10190 780
rect 10197 765 10203 766
rect 10211 765 10226 780
rect 10292 774 10311 777
rect 9933 752 10031 754
rect 10058 752 10226 765
rect 10241 754 10257 768
rect 10292 755 10314 774
rect 10324 768 10340 769
rect 10323 766 10340 768
rect 10324 761 10340 766
rect 10314 754 10320 755
rect 10323 754 10352 761
rect 10241 753 10352 754
rect 10241 752 10358 753
rect 9917 744 9968 752
rect 10015 744 10049 752
rect 9917 732 9942 744
rect 9949 732 9968 744
rect 10022 742 10049 744
rect 10058 742 10279 752
rect 10314 749 10320 752
rect 10022 738 10279 742
rect 9917 724 9968 732
rect 10015 724 10279 738
rect 10323 744 10358 752
rect 9869 676 9888 710
rect 9933 716 9962 724
rect 9933 710 9950 716
rect 9933 708 9967 710
rect 10015 708 10031 724
rect 10032 714 10240 724
rect 10241 714 10257 724
rect 10305 720 10320 735
rect 10323 732 10324 744
rect 10331 732 10358 744
rect 10323 724 10358 732
rect 10323 723 10352 724
rect 10043 710 10257 714
rect 10058 708 10257 710
rect 10292 710 10305 720
rect 10323 710 10340 723
rect 10292 708 10340 710
rect 9934 704 9967 708
rect 9930 702 9967 704
rect 9930 701 9997 702
rect 9930 696 9961 701
rect 9967 696 9997 701
rect 9930 692 9997 696
rect 9903 689 9997 692
rect 9903 682 9952 689
rect 9903 676 9933 682
rect 9952 677 9957 682
rect 9869 660 9949 676
rect 9961 668 9997 689
rect 10058 684 10247 708
rect 10292 707 10339 708
rect 10305 702 10339 707
rect 10073 681 10247 684
rect 10066 678 10247 681
rect 10275 701 10339 702
rect 9869 658 9888 660
rect 9903 658 9937 660
rect 9869 642 9949 658
rect 9869 636 9888 642
rect 9585 610 9688 620
rect 9539 608 9688 610
rect 9709 608 9744 620
rect 9378 606 9540 608
rect 9390 586 9409 606
rect 9424 604 9454 606
rect 9273 578 9314 586
rect 9396 583 9409 586
rect 9461 590 9540 606
rect 9572 606 9744 608
rect 9572 590 9651 606
rect 9658 604 9688 606
rect 9236 569 9265 578
rect 9279 569 9308 578
rect 9224 568 9308 569
rect 9323 568 9353 583
rect 9396 579 9439 583
rect 9461 579 9651 590
rect 9716 586 9722 606
rect 9673 579 9703 583
rect 9396 578 9703 579
rect 9396 568 9439 578
rect 9446 568 9476 578
rect 9477 568 9635 578
rect 9639 568 9669 578
rect 9673 568 9703 578
rect 9731 568 9744 606
rect 9816 620 9845 636
rect 9859 620 9888 636
rect 9903 626 9933 642
rect 9961 620 9967 668
rect 9970 662 9989 668
rect 10004 662 10034 670
rect 9970 654 10034 662
rect 9970 638 10050 654
rect 10066 647 10128 678
rect 10144 647 10206 678
rect 10275 676 10324 701
rect 10339 676 10369 692
rect 10238 662 10268 670
rect 10275 668 10385 676
rect 10238 654 10283 662
rect 9970 636 9989 638
rect 10004 636 10050 638
rect 9970 620 10050 636
rect 10077 634 10112 647
rect 10153 644 10190 647
rect 10153 642 10195 644
rect 10082 631 10112 634
rect 10091 627 10098 631
rect 10098 626 10099 627
rect 10057 620 10067 626
rect 9816 612 9851 620
rect 9816 586 9817 612
rect 9824 586 9851 612
rect 9759 568 9789 583
rect 9816 578 9851 586
rect 9853 612 9894 620
rect 9853 586 9868 612
rect 9875 586 9894 612
rect 9958 608 9989 620
rect 10004 608 10107 620
rect 10119 610 10145 636
rect 10160 631 10190 642
rect 10222 638 10284 654
rect 10222 636 10268 638
rect 10222 620 10284 636
rect 10296 620 10302 668
rect 10305 660 10385 668
rect 10305 658 10324 660
rect 10339 658 10373 660
rect 10305 642 10385 658
rect 10305 620 10324 642
rect 10339 626 10369 642
rect 10397 636 10403 710
rect 10406 636 10425 780
rect 10440 636 10446 780
rect 10455 710 10468 780
rect 10520 776 10542 780
rect 10513 754 10542 768
rect 10595 754 10611 768
rect 10649 765 10655 766
rect 10662 765 10770 780
rect 10777 765 10783 766
rect 10791 765 10806 780
rect 10872 774 10891 777
rect 10513 752 10611 754
rect 10638 752 10806 765
rect 10821 754 10837 768
rect 10872 755 10894 774
rect 10904 768 10920 769
rect 10903 766 10920 768
rect 10904 761 10920 766
rect 10894 754 10900 755
rect 10903 754 10932 761
rect 10821 753 10932 754
rect 10821 752 10938 753
rect 10497 744 10548 752
rect 10595 744 10629 752
rect 10497 732 10522 744
rect 10529 732 10548 744
rect 10602 742 10629 744
rect 10638 742 10859 752
rect 10894 749 10900 752
rect 10602 738 10859 742
rect 10497 724 10548 732
rect 10595 724 10859 738
rect 10903 744 10938 752
rect 10449 676 10468 710
rect 10513 716 10542 724
rect 10513 710 10530 716
rect 10513 708 10547 710
rect 10595 708 10611 724
rect 10612 714 10820 724
rect 10821 714 10837 724
rect 10885 720 10900 735
rect 10903 732 10904 744
rect 10911 732 10938 744
rect 10903 724 10938 732
rect 10903 723 10932 724
rect 10623 710 10837 714
rect 10638 708 10837 710
rect 10872 710 10885 720
rect 10903 710 10920 723
rect 10872 708 10920 710
rect 10514 704 10547 708
rect 10510 702 10547 704
rect 10510 701 10577 702
rect 10510 696 10541 701
rect 10547 696 10577 701
rect 10510 692 10577 696
rect 10483 689 10577 692
rect 10483 682 10532 689
rect 10483 676 10513 682
rect 10532 677 10537 682
rect 10449 660 10529 676
rect 10541 668 10577 689
rect 10638 684 10827 708
rect 10872 707 10919 708
rect 10885 702 10919 707
rect 10653 681 10827 684
rect 10646 678 10827 681
rect 10855 701 10919 702
rect 10449 658 10468 660
rect 10483 658 10517 660
rect 10449 642 10529 658
rect 10449 636 10468 642
rect 10165 610 10268 620
rect 10119 608 10268 610
rect 10289 608 10324 620
rect 9958 606 10120 608
rect 9970 586 9989 606
rect 10004 604 10034 606
rect 9853 578 9894 586
rect 9976 583 9989 586
rect 10041 590 10120 606
rect 10152 606 10324 608
rect 10152 590 10231 606
rect 10238 604 10268 606
rect 9816 568 9845 578
rect 9859 568 9888 578
rect 9903 568 9933 583
rect 9976 579 10019 583
rect 10041 579 10231 590
rect 10296 586 10302 606
rect 10253 579 10283 583
rect 9976 578 10283 579
rect 9976 568 10019 578
rect 10026 568 10056 578
rect 10057 568 10215 578
rect 10219 568 10249 578
rect 10253 568 10283 578
rect 10311 568 10324 606
rect 10396 620 10425 636
rect 10439 620 10468 636
rect 10483 626 10513 642
rect 10541 620 10547 668
rect 10550 662 10569 668
rect 10584 662 10614 670
rect 10550 654 10614 662
rect 10550 638 10630 654
rect 10646 647 10708 678
rect 10724 647 10786 678
rect 10855 676 10904 701
rect 10919 676 10949 692
rect 10818 662 10848 670
rect 10855 668 10965 676
rect 10818 654 10863 662
rect 10550 636 10569 638
rect 10584 636 10630 638
rect 10550 620 10630 636
rect 10657 634 10692 647
rect 10733 644 10770 647
rect 10733 642 10775 644
rect 10662 631 10692 634
rect 10671 627 10678 631
rect 10678 626 10679 627
rect 10637 620 10647 626
rect 10396 612 10431 620
rect 10396 586 10397 612
rect 10404 586 10431 612
rect 10339 568 10369 583
rect 10396 578 10431 586
rect 10433 612 10474 620
rect 10433 586 10448 612
rect 10455 586 10474 612
rect 10538 608 10569 620
rect 10584 608 10687 620
rect 10699 610 10725 636
rect 10740 631 10770 642
rect 10802 638 10864 654
rect 10802 636 10848 638
rect 10802 620 10864 636
rect 10876 620 10882 668
rect 10885 660 10965 668
rect 10885 658 10904 660
rect 10919 658 10953 660
rect 10885 642 10965 658
rect 10885 620 10904 642
rect 10919 626 10949 642
rect 10977 636 10983 710
rect 10986 636 11005 780
rect 11020 636 11026 780
rect 11035 710 11048 780
rect 11100 776 11122 780
rect 11093 754 11122 768
rect 11175 754 11191 768
rect 11229 765 11235 766
rect 11242 765 11350 780
rect 11357 765 11363 766
rect 11371 765 11386 780
rect 11452 774 11471 777
rect 11093 752 11191 754
rect 11218 752 11386 765
rect 11401 754 11417 768
rect 11452 755 11474 774
rect 11484 768 11500 769
rect 11483 766 11500 768
rect 11484 761 11500 766
rect 11474 754 11480 755
rect 11483 754 11512 761
rect 11401 753 11512 754
rect 11401 752 11518 753
rect 11077 744 11128 752
rect 11175 744 11209 752
rect 11077 732 11102 744
rect 11109 732 11128 744
rect 11182 742 11209 744
rect 11218 742 11439 752
rect 11474 749 11480 752
rect 11182 738 11439 742
rect 11077 724 11128 732
rect 11175 724 11439 738
rect 11483 744 11518 752
rect 11029 676 11048 710
rect 11093 716 11122 724
rect 11093 710 11110 716
rect 11093 708 11127 710
rect 11175 708 11191 724
rect 11192 714 11400 724
rect 11401 714 11417 724
rect 11465 720 11480 735
rect 11483 732 11484 744
rect 11491 732 11518 744
rect 11483 724 11518 732
rect 11483 723 11512 724
rect 11203 710 11417 714
rect 11218 708 11417 710
rect 11452 710 11465 720
rect 11483 710 11500 723
rect 11452 708 11500 710
rect 11094 704 11127 708
rect 11090 702 11127 704
rect 11090 701 11157 702
rect 11090 696 11121 701
rect 11127 696 11157 701
rect 11090 692 11157 696
rect 11063 689 11157 692
rect 11063 682 11112 689
rect 11063 676 11093 682
rect 11112 677 11117 682
rect 11029 660 11109 676
rect 11121 668 11157 689
rect 11218 684 11407 708
rect 11452 707 11499 708
rect 11465 702 11499 707
rect 11233 681 11407 684
rect 11226 678 11407 681
rect 11435 701 11499 702
rect 11029 658 11048 660
rect 11063 658 11097 660
rect 11029 642 11109 658
rect 11029 636 11048 642
rect 10745 610 10848 620
rect 10699 608 10848 610
rect 10869 608 10904 620
rect 10538 606 10700 608
rect 10550 586 10569 606
rect 10584 604 10614 606
rect 10433 578 10474 586
rect 10556 583 10569 586
rect 10621 590 10700 606
rect 10732 606 10904 608
rect 10732 590 10811 606
rect 10818 604 10848 606
rect 10396 568 10425 578
rect 10439 568 10468 578
rect 10483 568 10513 583
rect 10556 579 10599 583
rect 10621 579 10811 590
rect 10876 586 10882 606
rect 10833 579 10863 583
rect 10556 578 10863 579
rect 10556 568 10599 578
rect 10606 568 10636 578
rect 10637 568 10795 578
rect 10799 568 10829 578
rect 10833 568 10863 578
rect 10891 568 10904 606
rect 10976 620 11005 636
rect 11019 620 11048 636
rect 11063 626 11093 642
rect 11121 620 11127 668
rect 11130 662 11149 668
rect 11164 662 11194 670
rect 11130 654 11194 662
rect 11130 638 11210 654
rect 11226 647 11288 678
rect 11304 647 11366 678
rect 11435 676 11484 701
rect 11499 676 11529 692
rect 11398 662 11428 670
rect 11435 668 11545 676
rect 11398 654 11443 662
rect 11130 636 11149 638
rect 11164 636 11210 638
rect 11130 620 11210 636
rect 11237 634 11272 647
rect 11313 644 11350 647
rect 11313 642 11355 644
rect 11242 631 11272 634
rect 11251 627 11258 631
rect 11258 626 11259 627
rect 11217 620 11227 626
rect 10976 612 11011 620
rect 10976 586 10977 612
rect 10984 586 11011 612
rect 10919 568 10949 583
rect 10976 578 11011 586
rect 11013 612 11054 620
rect 11013 586 11028 612
rect 11035 586 11054 612
rect 11118 608 11149 620
rect 11164 608 11267 620
rect 11279 610 11305 636
rect 11320 631 11350 642
rect 11382 638 11444 654
rect 11382 636 11428 638
rect 11382 620 11444 636
rect 11456 620 11462 668
rect 11465 660 11545 668
rect 11465 658 11484 660
rect 11499 658 11533 660
rect 11465 642 11545 658
rect 11465 620 11484 642
rect 11499 626 11529 642
rect 11557 636 11563 710
rect 11566 636 11585 780
rect 11600 636 11606 780
rect 11615 710 11628 780
rect 11680 776 11702 780
rect 11673 754 11702 768
rect 11755 754 11771 768
rect 11809 765 11815 766
rect 11822 765 11930 780
rect 11937 765 11943 766
rect 11951 765 11966 780
rect 12032 774 12051 777
rect 11673 752 11771 754
rect 11798 752 11966 765
rect 11981 754 11997 768
rect 12032 755 12054 774
rect 12064 768 12080 769
rect 12063 766 12080 768
rect 12064 761 12080 766
rect 12054 754 12060 755
rect 12063 754 12092 761
rect 11981 753 12092 754
rect 11981 752 12098 753
rect 11657 744 11708 752
rect 11755 744 11789 752
rect 11657 732 11682 744
rect 11689 732 11708 744
rect 11762 742 11789 744
rect 11798 742 12019 752
rect 12054 749 12060 752
rect 11762 738 12019 742
rect 11657 724 11708 732
rect 11755 724 12019 738
rect 12063 744 12098 752
rect 11609 676 11628 710
rect 11673 716 11702 724
rect 11673 710 11690 716
rect 11673 708 11707 710
rect 11755 708 11771 724
rect 11772 714 11980 724
rect 11981 714 11997 724
rect 12045 720 12060 735
rect 12063 732 12064 744
rect 12071 732 12098 744
rect 12063 724 12098 732
rect 12063 723 12092 724
rect 11783 710 11997 714
rect 11798 708 11997 710
rect 12032 710 12045 720
rect 12063 710 12080 723
rect 12032 708 12080 710
rect 11674 704 11707 708
rect 11670 702 11707 704
rect 11670 701 11737 702
rect 11670 696 11701 701
rect 11707 696 11737 701
rect 11670 692 11737 696
rect 11643 689 11737 692
rect 11643 682 11692 689
rect 11643 676 11673 682
rect 11692 677 11697 682
rect 11609 660 11689 676
rect 11701 668 11737 689
rect 11798 684 11987 708
rect 12032 707 12079 708
rect 12045 702 12079 707
rect 11813 681 11987 684
rect 11806 678 11987 681
rect 12015 701 12079 702
rect 11609 658 11628 660
rect 11643 658 11677 660
rect 11609 642 11689 658
rect 11609 636 11628 642
rect 11325 610 11428 620
rect 11279 608 11428 610
rect 11449 608 11484 620
rect 11118 606 11280 608
rect 11130 586 11149 606
rect 11164 604 11194 606
rect 11013 578 11054 586
rect 11136 583 11149 586
rect 11201 590 11280 606
rect 11312 606 11484 608
rect 11312 590 11391 606
rect 11398 604 11428 606
rect 10976 568 11005 578
rect 11019 568 11048 578
rect 11063 568 11093 583
rect 11136 579 11179 583
rect 11201 579 11391 590
rect 11456 586 11462 606
rect 11413 579 11443 583
rect 11136 578 11443 579
rect 11136 568 11179 578
rect 11186 568 11216 578
rect 11217 568 11375 578
rect 11379 568 11409 578
rect 11413 568 11443 578
rect 11471 568 11484 606
rect 11556 620 11585 636
rect 11599 620 11628 636
rect 11643 626 11673 642
rect 11701 620 11707 668
rect 11710 662 11729 668
rect 11744 662 11774 670
rect 11710 654 11774 662
rect 11710 638 11790 654
rect 11806 647 11868 678
rect 11884 647 11946 678
rect 12015 676 12064 701
rect 12079 676 12109 692
rect 11978 662 12008 670
rect 12015 668 12125 676
rect 11978 654 12023 662
rect 11710 636 11729 638
rect 11744 636 11790 638
rect 11710 620 11790 636
rect 11817 634 11852 647
rect 11893 644 11930 647
rect 11893 642 11935 644
rect 11822 631 11852 634
rect 11831 627 11838 631
rect 11838 626 11839 627
rect 11797 620 11807 626
rect 11556 612 11591 620
rect 11556 586 11557 612
rect 11564 586 11591 612
rect 11499 568 11529 583
rect 11556 578 11591 586
rect 11593 612 11634 620
rect 11593 586 11608 612
rect 11615 586 11634 612
rect 11698 608 11729 620
rect 11744 608 11847 620
rect 11859 610 11885 636
rect 11900 631 11930 642
rect 11962 638 12024 654
rect 11962 636 12008 638
rect 11962 620 12024 636
rect 12036 620 12042 668
rect 12045 660 12125 668
rect 12045 658 12064 660
rect 12079 658 12113 660
rect 12045 642 12125 658
rect 12045 620 12064 642
rect 12079 626 12109 642
rect 12137 636 12143 710
rect 12146 636 12165 780
rect 12180 636 12186 780
rect 12195 710 12208 780
rect 12260 776 12282 780
rect 12253 754 12282 768
rect 12335 754 12351 768
rect 12389 765 12395 766
rect 12402 765 12510 780
rect 12517 765 12523 766
rect 12531 765 12546 780
rect 12612 774 12631 777
rect 12253 752 12351 754
rect 12378 752 12546 765
rect 12561 754 12577 768
rect 12612 755 12634 774
rect 12644 768 12660 769
rect 12643 766 12660 768
rect 12644 761 12660 766
rect 12634 754 12640 755
rect 12643 754 12672 761
rect 12561 753 12672 754
rect 12561 752 12678 753
rect 12237 744 12288 752
rect 12335 744 12369 752
rect 12237 732 12262 744
rect 12269 732 12288 744
rect 12342 742 12369 744
rect 12378 742 12599 752
rect 12634 749 12640 752
rect 12342 738 12599 742
rect 12237 724 12288 732
rect 12335 724 12599 738
rect 12643 744 12678 752
rect 12189 676 12208 710
rect 12253 716 12282 724
rect 12253 710 12270 716
rect 12253 708 12287 710
rect 12335 708 12351 724
rect 12352 714 12560 724
rect 12561 714 12577 724
rect 12625 720 12640 735
rect 12643 732 12644 744
rect 12651 732 12678 744
rect 12643 724 12678 732
rect 12643 723 12672 724
rect 12363 710 12577 714
rect 12378 708 12577 710
rect 12612 710 12625 720
rect 12643 710 12660 723
rect 12612 708 12660 710
rect 12254 704 12287 708
rect 12250 702 12287 704
rect 12250 701 12317 702
rect 12250 696 12281 701
rect 12287 696 12317 701
rect 12250 692 12317 696
rect 12223 689 12317 692
rect 12223 682 12272 689
rect 12223 676 12253 682
rect 12272 677 12277 682
rect 12189 660 12269 676
rect 12281 668 12317 689
rect 12378 684 12567 708
rect 12612 707 12659 708
rect 12625 702 12659 707
rect 12393 681 12567 684
rect 12386 678 12567 681
rect 12595 701 12659 702
rect 12189 658 12208 660
rect 12223 658 12257 660
rect 12189 642 12269 658
rect 12189 636 12208 642
rect 11905 610 12008 620
rect 11859 608 12008 610
rect 12029 608 12064 620
rect 11698 606 11860 608
rect 11710 586 11729 606
rect 11744 604 11774 606
rect 11593 578 11634 586
rect 11716 583 11729 586
rect 11781 590 11860 606
rect 11892 606 12064 608
rect 11892 590 11971 606
rect 11978 604 12008 606
rect 11556 568 11585 578
rect 11599 568 11628 578
rect 11643 568 11673 583
rect 11716 568 11759 583
rect 11781 579 11971 590
rect 12036 586 12042 606
rect 11993 579 12023 583
rect 11776 578 12023 579
rect 11766 568 11796 578
rect 11797 568 11955 578
rect 11959 568 11989 578
rect 11993 568 12023 578
rect 12051 568 12064 606
rect 12136 620 12165 636
rect 12179 620 12208 636
rect 12223 626 12253 642
rect 12281 620 12287 668
rect 12290 662 12309 668
rect 12324 662 12354 670
rect 12290 654 12354 662
rect 12290 638 12370 654
rect 12386 647 12448 678
rect 12464 647 12526 678
rect 12595 676 12644 701
rect 12659 676 12689 692
rect 12558 662 12588 670
rect 12595 668 12705 676
rect 12558 654 12603 662
rect 12290 636 12309 638
rect 12324 636 12370 638
rect 12290 620 12370 636
rect 12397 634 12432 647
rect 12473 644 12510 647
rect 12473 642 12515 644
rect 12402 631 12432 634
rect 12411 627 12418 631
rect 12418 626 12419 627
rect 12377 620 12387 626
rect 12136 612 12171 620
rect 12136 586 12137 612
rect 12144 586 12171 612
rect 12079 568 12109 583
rect 12136 578 12171 586
rect 12173 612 12214 620
rect 12173 586 12188 612
rect 12195 586 12214 612
rect 12278 608 12309 620
rect 12324 608 12427 620
rect 12439 610 12465 636
rect 12480 631 12510 642
rect 12542 638 12604 654
rect 12542 636 12588 638
rect 12542 620 12604 636
rect 12616 620 12622 668
rect 12625 660 12705 668
rect 12625 658 12644 660
rect 12659 658 12693 660
rect 12625 642 12705 658
rect 12625 620 12644 642
rect 12659 626 12689 642
rect 12717 636 12723 710
rect 12726 636 12745 780
rect 12760 636 12766 780
rect 12775 710 12788 780
rect 12840 776 12862 780
rect 12833 754 12862 768
rect 12915 754 12931 768
rect 12969 765 12975 766
rect 12982 765 13090 780
rect 13097 765 13103 766
rect 13111 765 13126 780
rect 13192 774 13211 777
rect 12833 752 12931 754
rect 12958 752 13126 765
rect 13141 754 13157 768
rect 13192 755 13214 774
rect 13224 768 13240 769
rect 13223 766 13240 768
rect 13224 761 13240 766
rect 13214 754 13220 755
rect 13223 754 13252 761
rect 13141 753 13252 754
rect 13141 752 13258 753
rect 12817 744 12868 752
rect 12915 744 12949 752
rect 12817 732 12842 744
rect 12849 732 12868 744
rect 12922 742 12949 744
rect 12958 742 13179 752
rect 13214 749 13220 752
rect 12922 738 13179 742
rect 12817 724 12868 732
rect 12915 724 13179 738
rect 13223 744 13258 752
rect 12769 676 12788 710
rect 12833 716 12862 724
rect 12833 710 12850 716
rect 12833 708 12867 710
rect 12915 708 12931 724
rect 12932 714 13140 724
rect 13141 714 13157 724
rect 13205 720 13220 735
rect 13223 732 13224 744
rect 13231 732 13258 744
rect 13223 724 13258 732
rect 13223 723 13252 724
rect 12943 710 13157 714
rect 12958 708 13157 710
rect 13192 710 13205 720
rect 13223 710 13240 723
rect 13192 708 13240 710
rect 12834 704 12867 708
rect 12830 702 12867 704
rect 12830 701 12897 702
rect 12830 696 12861 701
rect 12867 696 12897 701
rect 12830 692 12897 696
rect 12803 689 12897 692
rect 12803 682 12852 689
rect 12803 676 12833 682
rect 12852 677 12857 682
rect 12769 660 12849 676
rect 12861 668 12897 689
rect 12958 684 13147 708
rect 13192 707 13239 708
rect 13205 702 13239 707
rect 12973 681 13147 684
rect 12966 678 13147 681
rect 13175 701 13239 702
rect 12769 658 12788 660
rect 12803 658 12837 660
rect 12769 642 12849 658
rect 12769 636 12788 642
rect 12485 610 12588 620
rect 12439 608 12588 610
rect 12609 608 12644 620
rect 12278 606 12440 608
rect 12290 586 12309 606
rect 12324 604 12354 606
rect 12173 578 12214 586
rect 12296 583 12309 586
rect 12361 590 12440 606
rect 12472 606 12644 608
rect 12472 590 12551 606
rect 12558 604 12588 606
rect 12136 568 12165 578
rect 12179 568 12208 578
rect 12223 568 12253 583
rect 12296 579 12339 583
rect 12361 579 12551 590
rect 12616 586 12622 606
rect 12573 579 12603 583
rect 12296 578 12603 579
rect 12296 568 12339 578
rect 12346 568 12376 578
rect 12377 568 12535 578
rect 12539 568 12569 578
rect 12573 568 12603 578
rect 12631 568 12644 606
rect 12716 620 12745 636
rect 12759 620 12788 636
rect 12803 626 12833 642
rect 12861 620 12867 668
rect 12870 662 12889 668
rect 12904 662 12934 670
rect 12870 654 12934 662
rect 12870 638 12950 654
rect 12966 647 13028 678
rect 13044 647 13106 678
rect 13175 676 13224 701
rect 13239 676 13269 692
rect 13138 662 13168 670
rect 13175 668 13285 676
rect 13138 654 13183 662
rect 12870 636 12889 638
rect 12904 636 12950 638
rect 12870 620 12950 636
rect 12977 634 13012 647
rect 13053 644 13090 647
rect 13053 642 13095 644
rect 12982 631 13012 634
rect 12991 627 12998 631
rect 12998 626 12999 627
rect 12957 620 12967 626
rect 12716 612 12751 620
rect 12716 586 12717 612
rect 12724 586 12751 612
rect 12659 568 12689 583
rect 12716 578 12751 586
rect 12753 612 12794 620
rect 12753 586 12768 612
rect 12775 586 12794 612
rect 12858 608 12889 620
rect 12904 608 13007 620
rect 13019 610 13045 636
rect 13060 631 13090 642
rect 13122 638 13184 654
rect 13122 636 13168 638
rect 13122 620 13184 636
rect 13196 620 13202 668
rect 13205 660 13285 668
rect 13205 658 13224 660
rect 13239 658 13273 660
rect 13205 642 13285 658
rect 13205 620 13224 642
rect 13239 626 13269 642
rect 13297 636 13303 710
rect 13306 636 13325 780
rect 13340 636 13346 780
rect 13355 710 13368 780
rect 13420 776 13442 780
rect 13413 754 13442 768
rect 13495 754 13511 768
rect 13549 765 13555 766
rect 13562 765 13670 780
rect 13677 765 13683 766
rect 13691 765 13706 780
rect 13772 774 13791 777
rect 13413 752 13511 754
rect 13538 752 13706 765
rect 13721 754 13737 768
rect 13772 755 13794 774
rect 13804 768 13820 769
rect 13803 766 13820 768
rect 13804 761 13820 766
rect 13794 754 13800 755
rect 13803 754 13832 761
rect 13721 753 13832 754
rect 13721 752 13838 753
rect 13397 744 13448 752
rect 13495 744 13529 752
rect 13397 732 13422 744
rect 13429 732 13448 744
rect 13502 742 13529 744
rect 13538 742 13759 752
rect 13794 749 13800 752
rect 13502 738 13759 742
rect 13397 724 13448 732
rect 13495 724 13759 738
rect 13803 744 13838 752
rect 13349 676 13368 710
rect 13413 716 13442 724
rect 13413 710 13430 716
rect 13413 708 13447 710
rect 13495 708 13511 724
rect 13512 714 13720 724
rect 13721 714 13737 724
rect 13785 720 13800 735
rect 13803 732 13804 744
rect 13811 732 13838 744
rect 13803 724 13838 732
rect 13803 723 13832 724
rect 13523 710 13737 714
rect 13538 708 13737 710
rect 13772 710 13785 720
rect 13803 710 13820 723
rect 13772 708 13820 710
rect 13414 704 13447 708
rect 13410 702 13447 704
rect 13410 701 13477 702
rect 13410 696 13441 701
rect 13447 696 13477 701
rect 13410 692 13477 696
rect 13383 689 13477 692
rect 13383 682 13432 689
rect 13383 676 13413 682
rect 13432 677 13437 682
rect 13349 660 13429 676
rect 13441 668 13477 689
rect 13538 684 13727 708
rect 13772 707 13819 708
rect 13785 702 13819 707
rect 13553 681 13727 684
rect 13546 678 13727 681
rect 13755 701 13819 702
rect 13349 658 13368 660
rect 13383 658 13417 660
rect 13349 642 13429 658
rect 13349 636 13368 642
rect 13065 610 13168 620
rect 13019 608 13168 610
rect 13189 608 13224 620
rect 12858 606 13020 608
rect 12870 586 12889 606
rect 12904 604 12934 606
rect 12753 578 12794 586
rect 12876 583 12889 586
rect 12941 590 13020 606
rect 13052 606 13224 608
rect 13052 590 13131 606
rect 13138 604 13168 606
rect 12716 568 12745 578
rect 12759 568 12788 578
rect 12803 568 12833 583
rect 12876 579 12919 583
rect 12941 579 13131 590
rect 13196 586 13202 606
rect 13153 579 13183 583
rect 12876 578 13183 579
rect 12876 568 12919 578
rect 12926 568 12956 578
rect 12957 568 13115 578
rect 13119 568 13149 578
rect 13153 568 13183 578
rect 13211 568 13224 606
rect 13296 620 13325 636
rect 13339 620 13368 636
rect 13383 626 13413 642
rect 13441 620 13447 668
rect 13450 662 13469 668
rect 13484 662 13514 670
rect 13450 654 13514 662
rect 13450 638 13530 654
rect 13546 647 13608 678
rect 13624 647 13686 678
rect 13755 676 13804 701
rect 13819 676 13849 692
rect 13718 662 13748 670
rect 13755 668 13865 676
rect 13718 654 13763 662
rect 13450 636 13469 638
rect 13484 636 13530 638
rect 13450 620 13530 636
rect 13557 634 13592 647
rect 13633 644 13670 647
rect 13633 642 13675 644
rect 13562 631 13592 634
rect 13571 627 13578 631
rect 13578 626 13579 627
rect 13537 620 13547 626
rect 13296 612 13331 620
rect 13296 586 13297 612
rect 13304 586 13331 612
rect 13239 568 13269 583
rect 13296 578 13331 586
rect 13333 612 13374 620
rect 13333 586 13348 612
rect 13355 586 13374 612
rect 13438 608 13469 620
rect 13484 608 13587 620
rect 13599 610 13625 636
rect 13640 631 13670 642
rect 13702 638 13764 654
rect 13702 636 13748 638
rect 13702 620 13764 636
rect 13776 620 13782 668
rect 13785 660 13865 668
rect 13785 658 13804 660
rect 13819 658 13853 660
rect 13785 642 13865 658
rect 13785 620 13804 642
rect 13819 626 13849 642
rect 13877 636 13883 710
rect 13886 636 13905 780
rect 13920 636 13926 780
rect 13935 710 13948 780
rect 14000 776 14022 780
rect 13993 754 14022 768
rect 14075 754 14091 768
rect 14129 765 14135 766
rect 14142 765 14250 780
rect 14257 765 14263 766
rect 14271 765 14286 780
rect 14352 774 14371 777
rect 13993 752 14091 754
rect 14118 752 14286 765
rect 14301 754 14317 768
rect 14352 755 14374 774
rect 14384 768 14400 769
rect 14383 766 14400 768
rect 14384 761 14400 766
rect 14374 754 14380 755
rect 14383 754 14412 761
rect 14301 753 14412 754
rect 14301 752 14418 753
rect 13977 744 14028 752
rect 14075 744 14109 752
rect 13977 732 14002 744
rect 14009 732 14028 744
rect 14082 742 14109 744
rect 14118 742 14339 752
rect 14374 749 14380 752
rect 14082 738 14339 742
rect 13977 724 14028 732
rect 14075 724 14339 738
rect 14383 744 14418 752
rect 13929 676 13948 710
rect 13993 716 14022 724
rect 13993 710 14010 716
rect 13993 708 14027 710
rect 14075 708 14091 724
rect 14092 714 14300 724
rect 14301 714 14317 724
rect 14365 720 14380 735
rect 14383 732 14384 744
rect 14391 732 14418 744
rect 14383 724 14418 732
rect 14383 723 14412 724
rect 14103 710 14317 714
rect 14118 708 14317 710
rect 14352 710 14365 720
rect 14383 710 14400 723
rect 14352 708 14400 710
rect 13994 704 14027 708
rect 13990 702 14027 704
rect 13990 701 14057 702
rect 13990 696 14021 701
rect 14027 696 14057 701
rect 13990 692 14057 696
rect 13963 689 14057 692
rect 13963 682 14012 689
rect 13963 676 13993 682
rect 14012 677 14017 682
rect 13929 660 14009 676
rect 14021 668 14057 689
rect 14118 684 14307 708
rect 14352 707 14399 708
rect 14365 702 14399 707
rect 14133 681 14307 684
rect 14126 678 14307 681
rect 14335 701 14399 702
rect 13929 658 13948 660
rect 13963 658 13997 660
rect 13929 642 14009 658
rect 13929 636 13948 642
rect 13645 610 13748 620
rect 13599 608 13748 610
rect 13769 608 13804 620
rect 13438 606 13600 608
rect 13450 586 13469 606
rect 13484 604 13514 606
rect 13333 578 13374 586
rect 13456 583 13469 586
rect 13521 590 13600 606
rect 13632 606 13804 608
rect 13632 590 13711 606
rect 13718 604 13748 606
rect 13296 568 13325 578
rect 13339 568 13368 578
rect 13383 568 13413 583
rect 13456 579 13499 583
rect 13521 579 13711 590
rect 13776 586 13782 606
rect 13733 579 13763 583
rect 13456 578 13763 579
rect 13456 568 13499 578
rect 13506 568 13536 578
rect 13537 568 13695 578
rect 13699 568 13729 578
rect 13733 568 13763 578
rect 13791 568 13804 606
rect 13876 620 13905 636
rect 13919 620 13948 636
rect 13963 626 13993 642
rect 14021 620 14027 668
rect 14030 662 14049 668
rect 14064 662 14094 670
rect 14030 654 14094 662
rect 14030 638 14110 654
rect 14126 647 14188 678
rect 14204 647 14266 678
rect 14335 676 14384 701
rect 14399 676 14429 692
rect 14298 662 14328 670
rect 14335 668 14445 676
rect 14298 654 14343 662
rect 14030 636 14049 638
rect 14064 636 14110 638
rect 14030 620 14110 636
rect 14137 634 14172 647
rect 14213 644 14250 647
rect 14213 642 14255 644
rect 14142 631 14172 634
rect 14151 627 14158 631
rect 14158 626 14159 627
rect 14117 620 14127 626
rect 13876 612 13911 620
rect 13876 586 13877 612
rect 13884 586 13911 612
rect 13819 568 13849 583
rect 13876 578 13911 586
rect 13913 612 13954 620
rect 13913 586 13928 612
rect 13935 586 13954 612
rect 14018 608 14049 620
rect 14064 608 14167 620
rect 14179 610 14205 636
rect 14220 631 14250 642
rect 14282 638 14344 654
rect 14282 636 14328 638
rect 14282 620 14344 636
rect 14356 620 14362 668
rect 14365 660 14445 668
rect 14365 658 14384 660
rect 14399 658 14433 660
rect 14365 642 14445 658
rect 14365 620 14384 642
rect 14399 626 14429 642
rect 14457 636 14463 710
rect 14466 636 14485 780
rect 14500 636 14506 780
rect 14515 710 14528 780
rect 14580 776 14602 780
rect 14573 754 14602 768
rect 14655 754 14671 768
rect 14709 765 14715 766
rect 14722 765 14830 780
rect 14837 765 14843 766
rect 14851 765 14866 780
rect 14932 774 14951 777
rect 14573 752 14671 754
rect 14698 752 14866 765
rect 14881 754 14897 768
rect 14932 755 14954 774
rect 14964 768 14980 769
rect 14963 766 14980 768
rect 14964 761 14980 766
rect 14954 754 14960 755
rect 14963 754 14992 761
rect 14881 753 14992 754
rect 14881 752 14998 753
rect 14557 744 14608 752
rect 14655 744 14689 752
rect 14557 732 14582 744
rect 14589 732 14608 744
rect 14662 742 14689 744
rect 14698 742 14919 752
rect 14954 749 14960 752
rect 14662 738 14919 742
rect 14557 724 14608 732
rect 14655 724 14919 738
rect 14963 744 14998 752
rect 14509 676 14528 710
rect 14573 716 14602 724
rect 14573 710 14590 716
rect 14573 708 14607 710
rect 14655 708 14671 724
rect 14672 714 14880 724
rect 14881 714 14897 724
rect 14945 720 14960 735
rect 14963 732 14964 744
rect 14971 732 14998 744
rect 14963 724 14998 732
rect 14963 723 14992 724
rect 14683 710 14897 714
rect 14698 708 14897 710
rect 14932 710 14945 720
rect 14963 710 14980 723
rect 14932 708 14980 710
rect 14574 704 14607 708
rect 14570 702 14607 704
rect 14570 701 14637 702
rect 14570 696 14601 701
rect 14607 696 14637 701
rect 14570 692 14637 696
rect 14543 689 14637 692
rect 14543 682 14592 689
rect 14543 676 14573 682
rect 14592 677 14597 682
rect 14509 660 14589 676
rect 14601 668 14637 689
rect 14698 684 14887 708
rect 14932 707 14979 708
rect 14945 702 14979 707
rect 14713 681 14887 684
rect 14706 678 14887 681
rect 14915 701 14979 702
rect 14509 658 14528 660
rect 14543 658 14577 660
rect 14509 642 14589 658
rect 14509 636 14528 642
rect 14225 610 14328 620
rect 14179 608 14328 610
rect 14349 608 14384 620
rect 14018 606 14180 608
rect 14030 586 14049 606
rect 14064 604 14094 606
rect 13913 578 13954 586
rect 14036 583 14049 586
rect 14101 590 14180 606
rect 14212 606 14384 608
rect 14212 590 14291 606
rect 14298 604 14328 606
rect 13876 568 13905 578
rect 13919 568 13948 578
rect 13963 568 13993 583
rect 14036 579 14079 583
rect 14101 579 14291 590
rect 14356 586 14362 606
rect 14313 579 14343 583
rect 14036 578 14343 579
rect 14036 568 14079 578
rect 14086 568 14116 578
rect 14117 568 14275 578
rect 14279 568 14309 578
rect 14313 568 14343 578
rect 14371 568 14384 606
rect 14456 620 14485 636
rect 14499 620 14528 636
rect 14543 626 14573 642
rect 14601 620 14607 668
rect 14610 662 14629 668
rect 14644 662 14674 670
rect 14610 654 14674 662
rect 14610 638 14690 654
rect 14706 647 14768 678
rect 14784 647 14846 678
rect 14915 676 14964 701
rect 14979 676 15009 692
rect 14878 662 14908 670
rect 14915 668 15025 676
rect 14878 654 14923 662
rect 14610 636 14629 638
rect 14644 636 14690 638
rect 14610 620 14690 636
rect 14717 634 14752 647
rect 14793 644 14830 647
rect 14793 642 14835 644
rect 14722 631 14752 634
rect 14731 627 14738 631
rect 14738 626 14739 627
rect 14697 620 14707 626
rect 14456 612 14491 620
rect 14456 586 14457 612
rect 14464 586 14491 612
rect 14399 568 14429 583
rect 14456 578 14491 586
rect 14493 612 14534 620
rect 14493 586 14508 612
rect 14515 586 14534 612
rect 14598 608 14629 620
rect 14644 608 14747 620
rect 14759 610 14785 636
rect 14800 631 14830 642
rect 14862 638 14924 654
rect 14862 636 14908 638
rect 14862 620 14924 636
rect 14936 620 14942 668
rect 14945 660 15025 668
rect 14945 658 14964 660
rect 14979 658 15013 660
rect 14945 642 15025 658
rect 14945 620 14964 642
rect 14979 626 15009 642
rect 15037 636 15043 710
rect 15046 636 15065 780
rect 15080 636 15086 780
rect 15095 710 15108 780
rect 15160 776 15182 780
rect 15153 754 15182 768
rect 15235 754 15251 768
rect 15289 765 15295 766
rect 15302 765 15410 780
rect 15417 765 15423 766
rect 15431 765 15446 780
rect 15512 774 15531 777
rect 15153 752 15251 754
rect 15278 752 15446 765
rect 15461 754 15477 768
rect 15512 755 15534 774
rect 15544 768 15560 769
rect 15543 766 15560 768
rect 15544 761 15560 766
rect 15534 754 15540 755
rect 15543 754 15572 761
rect 15461 753 15572 754
rect 15461 752 15578 753
rect 15137 744 15188 752
rect 15235 744 15269 752
rect 15137 732 15162 744
rect 15169 732 15188 744
rect 15242 742 15269 744
rect 15278 742 15499 752
rect 15534 749 15540 752
rect 15242 738 15499 742
rect 15137 724 15188 732
rect 15235 724 15499 738
rect 15543 744 15578 752
rect 15089 676 15108 710
rect 15153 716 15182 724
rect 15153 710 15170 716
rect 15153 708 15187 710
rect 15235 708 15251 724
rect 15252 714 15460 724
rect 15461 714 15477 724
rect 15525 720 15540 735
rect 15543 732 15544 744
rect 15551 732 15578 744
rect 15543 724 15578 732
rect 15543 723 15572 724
rect 15263 710 15477 714
rect 15278 708 15477 710
rect 15512 710 15525 720
rect 15543 710 15560 723
rect 15512 708 15560 710
rect 15154 704 15187 708
rect 15150 702 15187 704
rect 15150 701 15217 702
rect 15150 696 15181 701
rect 15187 696 15217 701
rect 15150 692 15217 696
rect 15123 689 15217 692
rect 15123 682 15172 689
rect 15123 676 15153 682
rect 15172 677 15177 682
rect 15089 660 15169 676
rect 15181 668 15217 689
rect 15278 684 15467 708
rect 15512 707 15559 708
rect 15525 702 15559 707
rect 15293 681 15467 684
rect 15286 678 15467 681
rect 15495 701 15559 702
rect 15089 658 15108 660
rect 15123 658 15157 660
rect 15089 642 15169 658
rect 15089 636 15108 642
rect 14805 610 14908 620
rect 14759 608 14908 610
rect 14929 608 14964 620
rect 14598 606 14760 608
rect 14610 586 14629 606
rect 14644 604 14674 606
rect 14493 578 14534 586
rect 14616 583 14629 586
rect 14681 590 14760 606
rect 14792 606 14964 608
rect 14792 590 14871 606
rect 14878 604 14908 606
rect 14456 568 14485 578
rect 14499 568 14528 578
rect 14543 568 14573 583
rect 14616 579 14659 583
rect 14681 579 14871 590
rect 14936 586 14942 606
rect 14893 579 14923 583
rect 14616 578 14923 579
rect 14616 568 14659 578
rect 14666 568 14696 578
rect 14697 568 14855 578
rect 14859 568 14889 578
rect 14893 568 14923 578
rect 14951 568 14964 606
rect 15036 620 15065 636
rect 15079 620 15108 636
rect 15123 626 15153 642
rect 15181 620 15187 668
rect 15190 662 15209 668
rect 15224 662 15254 670
rect 15190 654 15254 662
rect 15190 638 15270 654
rect 15286 647 15348 678
rect 15364 647 15426 678
rect 15495 676 15544 701
rect 15559 676 15589 692
rect 15458 662 15488 670
rect 15495 668 15605 676
rect 15458 654 15503 662
rect 15190 636 15209 638
rect 15224 636 15270 638
rect 15190 620 15270 636
rect 15297 634 15332 647
rect 15373 644 15410 647
rect 15373 642 15415 644
rect 15302 631 15332 634
rect 15311 627 15318 631
rect 15318 626 15319 627
rect 15277 620 15287 626
rect 15036 612 15071 620
rect 15036 586 15037 612
rect 15044 586 15071 612
rect 14979 568 15009 583
rect 15036 578 15071 586
rect 15073 612 15114 620
rect 15073 586 15088 612
rect 15095 586 15114 612
rect 15178 608 15209 620
rect 15224 608 15327 620
rect 15339 610 15365 636
rect 15380 631 15410 642
rect 15442 638 15504 654
rect 15442 636 15488 638
rect 15442 620 15504 636
rect 15516 620 15522 668
rect 15525 660 15605 668
rect 15525 658 15544 660
rect 15559 658 15593 660
rect 15525 642 15605 658
rect 15525 620 15544 642
rect 15559 626 15589 642
rect 15617 636 15623 710
rect 15626 636 15645 780
rect 15660 636 15666 780
rect 15675 710 15688 780
rect 15740 776 15762 780
rect 15733 754 15762 768
rect 15815 754 15831 768
rect 15869 765 15875 766
rect 15882 765 15990 780
rect 15997 765 16003 766
rect 16011 765 16026 780
rect 16092 774 16111 777
rect 15733 752 15831 754
rect 15858 752 16026 765
rect 16041 754 16057 768
rect 16092 755 16114 774
rect 16124 768 16140 769
rect 16123 766 16140 768
rect 16124 761 16140 766
rect 16114 754 16120 755
rect 16123 754 16152 761
rect 16041 753 16152 754
rect 16041 752 16158 753
rect 15717 744 15768 752
rect 15815 744 15849 752
rect 15717 732 15742 744
rect 15749 732 15768 744
rect 15822 742 15849 744
rect 15858 742 16079 752
rect 16114 749 16120 752
rect 15822 738 16079 742
rect 15717 724 15768 732
rect 15815 724 16079 738
rect 16123 744 16158 752
rect 15669 676 15688 710
rect 15733 716 15762 724
rect 15733 710 15750 716
rect 15733 708 15767 710
rect 15815 708 15831 724
rect 15832 714 16040 724
rect 16041 714 16057 724
rect 16105 720 16120 735
rect 16123 732 16124 744
rect 16131 732 16158 744
rect 16123 724 16158 732
rect 16123 723 16152 724
rect 15843 710 16057 714
rect 15858 708 16057 710
rect 16092 710 16105 720
rect 16123 710 16140 723
rect 16092 708 16140 710
rect 15734 704 15767 708
rect 15730 702 15767 704
rect 15730 701 15797 702
rect 15730 696 15761 701
rect 15767 696 15797 701
rect 15730 692 15797 696
rect 15703 689 15797 692
rect 15703 682 15752 689
rect 15703 676 15733 682
rect 15752 677 15757 682
rect 15669 660 15749 676
rect 15761 668 15797 689
rect 15858 684 16047 708
rect 16092 707 16139 708
rect 16105 702 16139 707
rect 15873 681 16047 684
rect 15866 678 16047 681
rect 16075 701 16139 702
rect 15669 658 15688 660
rect 15703 658 15737 660
rect 15669 642 15749 658
rect 15669 636 15688 642
rect 15385 610 15488 620
rect 15339 608 15488 610
rect 15509 608 15544 620
rect 15178 606 15340 608
rect 15190 586 15209 606
rect 15224 604 15254 606
rect 15073 578 15114 586
rect 15196 583 15209 586
rect 15261 590 15340 606
rect 15372 606 15544 608
rect 15372 590 15451 606
rect 15458 604 15488 606
rect 15036 568 15065 578
rect 15079 568 15108 578
rect 15123 568 15153 583
rect 15196 579 15239 583
rect 15261 579 15451 590
rect 15516 586 15522 606
rect 15473 579 15503 583
rect 15196 578 15503 579
rect 15196 568 15239 578
rect 15246 568 15276 578
rect 15277 568 15435 578
rect 15439 568 15469 578
rect 15473 568 15503 578
rect 15531 568 15544 606
rect 15616 620 15645 636
rect 15659 620 15688 636
rect 15703 626 15733 642
rect 15761 620 15767 668
rect 15770 662 15789 668
rect 15804 662 15834 670
rect 15770 654 15834 662
rect 15770 638 15850 654
rect 15866 647 15928 678
rect 15944 647 16006 678
rect 16075 676 16124 701
rect 16139 676 16169 692
rect 16038 662 16068 670
rect 16075 668 16185 676
rect 16038 654 16083 662
rect 15770 636 15789 638
rect 15804 636 15850 638
rect 15770 620 15850 636
rect 15877 634 15912 647
rect 15953 644 15990 647
rect 15953 642 15995 644
rect 15882 631 15912 634
rect 15891 627 15898 631
rect 15898 626 15899 627
rect 15857 620 15867 626
rect 15616 612 15651 620
rect 15616 586 15617 612
rect 15624 586 15651 612
rect 15559 568 15589 583
rect 15616 578 15651 586
rect 15653 612 15694 620
rect 15653 586 15668 612
rect 15675 586 15694 612
rect 15758 608 15789 620
rect 15804 608 15907 620
rect 15919 610 15945 636
rect 15960 631 15990 642
rect 16022 638 16084 654
rect 16022 636 16068 638
rect 16022 620 16084 636
rect 16096 620 16102 668
rect 16105 660 16185 668
rect 16105 658 16124 660
rect 16139 658 16173 660
rect 16105 642 16185 658
rect 16105 620 16124 642
rect 16139 626 16169 642
rect 16197 636 16203 710
rect 16206 636 16225 780
rect 16240 636 16246 780
rect 16255 710 16268 780
rect 16320 776 16342 780
rect 16313 754 16342 768
rect 16395 754 16411 768
rect 16449 765 16455 766
rect 16462 765 16570 780
rect 16577 765 16583 766
rect 16591 765 16606 780
rect 16672 774 16691 777
rect 16313 752 16411 754
rect 16438 752 16606 765
rect 16621 754 16637 768
rect 16672 755 16694 774
rect 16704 768 16720 769
rect 16703 766 16720 768
rect 16704 761 16720 766
rect 16694 754 16700 755
rect 16703 754 16732 761
rect 16621 753 16732 754
rect 16621 752 16738 753
rect 16297 744 16348 752
rect 16395 744 16429 752
rect 16297 732 16322 744
rect 16329 732 16348 744
rect 16402 742 16429 744
rect 16438 742 16659 752
rect 16694 749 16700 752
rect 16402 738 16659 742
rect 16297 724 16348 732
rect 16395 724 16659 738
rect 16703 744 16738 752
rect 16249 676 16268 710
rect 16313 716 16342 724
rect 16313 710 16330 716
rect 16313 708 16347 710
rect 16395 708 16411 724
rect 16412 714 16620 724
rect 16621 714 16637 724
rect 16685 720 16700 735
rect 16703 732 16704 744
rect 16711 732 16738 744
rect 16703 724 16738 732
rect 16703 723 16732 724
rect 16423 710 16637 714
rect 16438 708 16637 710
rect 16672 710 16685 720
rect 16703 710 16720 723
rect 16672 708 16720 710
rect 16314 704 16347 708
rect 16310 702 16347 704
rect 16310 701 16377 702
rect 16310 696 16341 701
rect 16347 696 16377 701
rect 16310 692 16377 696
rect 16283 689 16377 692
rect 16283 682 16332 689
rect 16283 676 16313 682
rect 16332 677 16337 682
rect 16249 660 16329 676
rect 16341 668 16377 689
rect 16438 684 16627 708
rect 16672 707 16719 708
rect 16685 702 16719 707
rect 16453 681 16627 684
rect 16446 678 16627 681
rect 16655 701 16719 702
rect 16249 658 16268 660
rect 16283 658 16317 660
rect 16249 642 16329 658
rect 16249 636 16268 642
rect 15965 610 16068 620
rect 15919 608 16068 610
rect 16089 608 16124 620
rect 15758 606 15920 608
rect 15770 586 15789 606
rect 15804 604 15834 606
rect 15653 578 15694 586
rect 15776 583 15789 586
rect 15841 590 15920 606
rect 15952 606 16124 608
rect 15952 590 16031 606
rect 16038 604 16068 606
rect 15616 568 15645 578
rect 15659 568 15688 578
rect 15703 568 15733 583
rect 15776 579 15819 583
rect 15841 579 16031 590
rect 16096 586 16102 606
rect 16053 579 16083 583
rect 15776 578 16083 579
rect 15776 568 15819 578
rect 15826 568 15856 578
rect 15857 568 16015 578
rect 16019 568 16049 578
rect 16053 568 16083 578
rect 16111 568 16124 606
rect 16196 620 16225 636
rect 16239 620 16268 636
rect 16283 626 16313 642
rect 16341 620 16347 668
rect 16350 662 16369 668
rect 16384 662 16414 670
rect 16350 654 16414 662
rect 16350 638 16430 654
rect 16446 647 16508 678
rect 16524 647 16586 678
rect 16655 676 16704 701
rect 16719 676 16749 692
rect 16618 662 16648 670
rect 16655 668 16765 676
rect 16618 654 16663 662
rect 16350 636 16369 638
rect 16384 636 16430 638
rect 16350 620 16430 636
rect 16457 634 16492 647
rect 16533 644 16570 647
rect 16533 642 16575 644
rect 16462 631 16492 634
rect 16471 627 16478 631
rect 16478 626 16479 627
rect 16437 620 16447 626
rect 16196 612 16231 620
rect 16196 586 16197 612
rect 16204 586 16231 612
rect 16139 568 16169 583
rect 16196 578 16231 586
rect 16233 612 16274 620
rect 16233 586 16248 612
rect 16255 586 16274 612
rect 16338 608 16369 620
rect 16384 608 16487 620
rect 16499 610 16525 636
rect 16540 631 16570 642
rect 16602 638 16664 654
rect 16602 636 16648 638
rect 16602 620 16664 636
rect 16676 620 16682 668
rect 16685 660 16765 668
rect 16685 658 16704 660
rect 16719 658 16753 660
rect 16685 642 16765 658
rect 16685 620 16704 642
rect 16719 626 16749 642
rect 16777 636 16783 710
rect 16786 636 16805 780
rect 16820 636 16826 780
rect 16835 710 16848 780
rect 16900 776 16922 780
rect 16893 754 16922 768
rect 16975 754 16991 768
rect 17029 765 17035 766
rect 17042 765 17150 780
rect 17157 765 17163 766
rect 17171 765 17186 780
rect 17252 774 17271 777
rect 16893 752 16991 754
rect 17018 752 17186 765
rect 17201 754 17217 768
rect 17252 755 17274 774
rect 17284 768 17300 769
rect 17283 766 17300 768
rect 17284 761 17300 766
rect 17274 754 17280 755
rect 17283 754 17312 761
rect 17201 753 17312 754
rect 17201 752 17318 753
rect 16877 744 16928 752
rect 16975 744 17009 752
rect 16877 732 16902 744
rect 16909 732 16928 744
rect 16982 742 17009 744
rect 17018 742 17239 752
rect 17274 749 17280 752
rect 16982 738 17239 742
rect 16877 724 16928 732
rect 16975 724 17239 738
rect 17283 744 17318 752
rect 16829 676 16848 710
rect 16893 716 16922 724
rect 16893 710 16910 716
rect 16893 708 16927 710
rect 16975 708 16991 724
rect 16992 714 17200 724
rect 17201 714 17217 724
rect 17265 720 17280 735
rect 17283 732 17284 744
rect 17291 732 17318 744
rect 17283 724 17318 732
rect 17283 723 17312 724
rect 17003 710 17217 714
rect 17018 708 17217 710
rect 17252 710 17265 720
rect 17283 710 17300 723
rect 17252 708 17300 710
rect 16894 704 16927 708
rect 16890 702 16927 704
rect 16890 701 16957 702
rect 16890 696 16921 701
rect 16927 696 16957 701
rect 16890 692 16957 696
rect 16863 689 16957 692
rect 16863 682 16912 689
rect 16863 676 16893 682
rect 16912 677 16917 682
rect 16829 660 16909 676
rect 16921 668 16957 689
rect 17018 684 17207 708
rect 17252 707 17299 708
rect 17265 702 17299 707
rect 17033 681 17207 684
rect 17026 678 17207 681
rect 17235 701 17299 702
rect 16829 658 16848 660
rect 16863 658 16897 660
rect 16829 642 16909 658
rect 16829 636 16848 642
rect 16545 610 16648 620
rect 16499 608 16648 610
rect 16669 608 16704 620
rect 16338 606 16500 608
rect 16350 586 16369 606
rect 16384 604 16414 606
rect 16233 578 16274 586
rect 16356 583 16369 586
rect 16421 590 16500 606
rect 16532 606 16704 608
rect 16532 590 16611 606
rect 16618 604 16648 606
rect 16196 568 16225 578
rect 16239 568 16268 578
rect 16283 568 16313 583
rect 16356 579 16399 583
rect 16421 579 16611 590
rect 16676 586 16682 606
rect 16633 579 16663 583
rect 16356 578 16663 579
rect 16356 568 16399 578
rect 16406 568 16436 578
rect 16437 568 16595 578
rect 16599 568 16629 578
rect 16633 568 16663 578
rect 16691 568 16704 606
rect 16776 620 16805 636
rect 16819 620 16848 636
rect 16863 626 16893 642
rect 16921 620 16927 668
rect 16930 662 16949 668
rect 16964 662 16994 670
rect 16930 654 16994 662
rect 16930 638 17010 654
rect 17026 647 17088 678
rect 17104 647 17166 678
rect 17235 676 17284 701
rect 17299 676 17329 692
rect 17198 662 17228 670
rect 17235 668 17345 676
rect 17198 654 17243 662
rect 16930 636 16949 638
rect 16964 636 17010 638
rect 16930 620 17010 636
rect 17037 634 17072 647
rect 17113 644 17150 647
rect 17113 642 17155 644
rect 17042 631 17072 634
rect 17051 627 17058 631
rect 17058 626 17059 627
rect 17017 620 17027 626
rect 16776 612 16811 620
rect 16776 586 16777 612
rect 16784 586 16811 612
rect 16719 568 16749 583
rect 16776 578 16811 586
rect 16813 612 16854 620
rect 16813 586 16828 612
rect 16835 586 16854 612
rect 16918 608 16949 620
rect 16964 608 17067 620
rect 17079 610 17105 636
rect 17120 631 17150 642
rect 17182 638 17244 654
rect 17182 636 17228 638
rect 17182 620 17244 636
rect 17256 620 17262 668
rect 17265 660 17345 668
rect 17265 658 17284 660
rect 17299 658 17333 660
rect 17265 642 17345 658
rect 17265 620 17284 642
rect 17299 626 17329 642
rect 17357 636 17363 710
rect 17366 636 17385 780
rect 17400 636 17406 780
rect 17415 710 17428 780
rect 17480 776 17502 780
rect 17473 754 17502 768
rect 17555 754 17571 768
rect 17609 765 17615 766
rect 17622 765 17730 780
rect 17737 765 17743 766
rect 17751 765 17766 780
rect 17832 774 17851 777
rect 17473 752 17571 754
rect 17598 752 17766 765
rect 17781 754 17797 768
rect 17832 755 17854 774
rect 17864 768 17880 769
rect 17863 766 17880 768
rect 17864 761 17880 766
rect 17854 754 17860 755
rect 17863 754 17892 761
rect 17781 753 17892 754
rect 17781 752 17898 753
rect 17457 744 17508 752
rect 17555 744 17589 752
rect 17457 732 17482 744
rect 17489 732 17508 744
rect 17562 742 17589 744
rect 17598 742 17819 752
rect 17854 749 17860 752
rect 17562 738 17819 742
rect 17457 724 17508 732
rect 17555 724 17819 738
rect 17863 744 17898 752
rect 17409 676 17428 710
rect 17473 716 17502 724
rect 17473 710 17490 716
rect 17473 708 17507 710
rect 17555 708 17571 724
rect 17572 714 17780 724
rect 17781 714 17797 724
rect 17845 720 17860 735
rect 17863 732 17864 744
rect 17871 732 17898 744
rect 17863 724 17898 732
rect 17863 723 17892 724
rect 17583 710 17797 714
rect 17598 708 17797 710
rect 17832 710 17845 720
rect 17863 710 17880 723
rect 17832 708 17880 710
rect 17474 704 17507 708
rect 17470 702 17507 704
rect 17470 701 17537 702
rect 17470 696 17501 701
rect 17507 696 17537 701
rect 17470 692 17537 696
rect 17443 689 17537 692
rect 17443 682 17492 689
rect 17443 676 17473 682
rect 17492 677 17497 682
rect 17409 660 17489 676
rect 17501 668 17537 689
rect 17598 684 17787 708
rect 17832 707 17879 708
rect 17845 702 17879 707
rect 17613 681 17787 684
rect 17606 678 17787 681
rect 17815 701 17879 702
rect 17409 658 17428 660
rect 17443 658 17477 660
rect 17409 642 17489 658
rect 17409 636 17428 642
rect 17125 610 17228 620
rect 17079 608 17228 610
rect 17249 608 17284 620
rect 16918 606 17080 608
rect 16930 586 16949 606
rect 16964 604 16994 606
rect 16813 578 16854 586
rect 16936 583 16949 586
rect 17001 590 17080 606
rect 17112 606 17284 608
rect 17112 590 17191 606
rect 17198 604 17228 606
rect 16776 568 16805 578
rect 16819 568 16848 578
rect 16863 568 16893 583
rect 16936 579 16979 583
rect 17001 579 17191 590
rect 17256 586 17262 606
rect 17213 579 17243 583
rect 16936 578 17243 579
rect 16936 568 16979 578
rect 16986 568 17016 578
rect 17017 568 17175 578
rect 17179 568 17209 578
rect 17213 568 17243 578
rect 17271 568 17284 606
rect 17356 620 17385 636
rect 17399 620 17428 636
rect 17443 626 17473 642
rect 17501 620 17507 668
rect 17510 662 17529 668
rect 17544 662 17574 670
rect 17510 654 17574 662
rect 17510 638 17590 654
rect 17606 647 17668 678
rect 17684 647 17746 678
rect 17815 676 17864 701
rect 17879 676 17909 692
rect 17778 662 17808 670
rect 17815 668 17925 676
rect 17778 654 17823 662
rect 17510 636 17529 638
rect 17544 636 17590 638
rect 17510 620 17590 636
rect 17617 634 17652 647
rect 17693 644 17730 647
rect 17693 642 17735 644
rect 17622 631 17652 634
rect 17631 627 17638 631
rect 17638 626 17639 627
rect 17597 620 17607 626
rect 17356 612 17391 620
rect 17356 586 17357 612
rect 17364 586 17391 612
rect 17299 568 17329 583
rect 17356 578 17391 586
rect 17393 612 17434 620
rect 17393 586 17408 612
rect 17415 586 17434 612
rect 17498 608 17529 620
rect 17544 608 17647 620
rect 17659 610 17685 636
rect 17700 631 17730 642
rect 17762 638 17824 654
rect 17762 636 17808 638
rect 17762 620 17824 636
rect 17836 620 17842 668
rect 17845 660 17925 668
rect 17845 658 17864 660
rect 17879 658 17913 660
rect 17845 642 17925 658
rect 17845 620 17864 642
rect 17879 626 17909 642
rect 17937 636 17943 710
rect 17946 636 17965 780
rect 17980 636 17986 780
rect 17995 710 18008 780
rect 18060 776 18082 780
rect 18053 754 18082 768
rect 18135 754 18151 768
rect 18189 765 18195 766
rect 18202 765 18310 780
rect 18317 765 18323 766
rect 18331 765 18346 780
rect 18412 774 18431 777
rect 18053 752 18151 754
rect 18178 752 18346 765
rect 18361 754 18377 768
rect 18412 755 18434 774
rect 18444 768 18460 769
rect 18443 766 18460 768
rect 18444 761 18460 766
rect 18434 754 18440 755
rect 18443 754 18472 761
rect 18361 753 18472 754
rect 18361 752 18478 753
rect 18037 744 18088 752
rect 18135 744 18169 752
rect 18037 732 18062 744
rect 18069 732 18088 744
rect 18142 742 18169 744
rect 18178 742 18399 752
rect 18434 749 18440 752
rect 18142 738 18399 742
rect 18037 724 18088 732
rect 18135 724 18399 738
rect 18443 744 18478 752
rect 17989 676 18008 710
rect 18053 716 18082 724
rect 18053 710 18070 716
rect 18053 708 18087 710
rect 18135 708 18151 724
rect 18152 714 18360 724
rect 18361 714 18377 724
rect 18425 720 18440 735
rect 18443 732 18444 744
rect 18451 732 18478 744
rect 18443 724 18478 732
rect 18443 723 18472 724
rect 18163 710 18377 714
rect 18178 708 18377 710
rect 18412 710 18425 720
rect 18443 710 18460 723
rect 18412 708 18460 710
rect 18054 704 18087 708
rect 18050 702 18087 704
rect 18050 701 18117 702
rect 18050 696 18081 701
rect 18087 696 18117 701
rect 18050 692 18117 696
rect 18023 689 18117 692
rect 18023 682 18072 689
rect 18023 676 18053 682
rect 18072 677 18077 682
rect 17989 660 18069 676
rect 18081 668 18117 689
rect 18178 684 18367 708
rect 18412 707 18459 708
rect 18425 702 18459 707
rect 18193 681 18367 684
rect 18186 678 18367 681
rect 18395 701 18459 702
rect 17989 658 18008 660
rect 18023 658 18057 660
rect 17989 642 18069 658
rect 17989 636 18008 642
rect 17705 610 17808 620
rect 17659 608 17808 610
rect 17829 608 17864 620
rect 17498 606 17660 608
rect 17510 586 17529 606
rect 17544 604 17574 606
rect 17393 578 17434 586
rect 17516 583 17529 586
rect 17581 590 17660 606
rect 17692 606 17864 608
rect 17692 590 17771 606
rect 17778 604 17808 606
rect 17356 568 17385 578
rect 17399 568 17428 578
rect 17443 568 17473 583
rect 17516 579 17559 583
rect 17581 579 17771 590
rect 17836 586 17842 606
rect 17793 579 17823 583
rect 17516 578 17823 579
rect 17516 568 17559 578
rect 17566 568 17596 578
rect 17597 568 17755 578
rect 17759 568 17789 578
rect 17793 568 17823 578
rect 17851 568 17864 606
rect 17936 620 17965 636
rect 17979 620 18008 636
rect 18023 626 18053 642
rect 18081 620 18087 668
rect 18090 662 18109 668
rect 18124 662 18154 670
rect 18090 654 18154 662
rect 18090 638 18170 654
rect 18186 647 18248 678
rect 18264 647 18326 678
rect 18395 676 18444 701
rect 18459 676 18489 692
rect 18358 662 18388 670
rect 18395 668 18505 676
rect 18358 654 18403 662
rect 18090 636 18109 638
rect 18124 636 18170 638
rect 18090 620 18170 636
rect 18197 634 18232 647
rect 18273 644 18310 647
rect 18273 642 18315 644
rect 18202 631 18232 634
rect 18211 627 18218 631
rect 18218 626 18219 627
rect 18177 620 18187 626
rect 17936 612 17971 620
rect 17936 586 17937 612
rect 17944 586 17971 612
rect 17879 568 17909 583
rect 17936 578 17971 586
rect 17973 612 18014 620
rect 17973 586 17988 612
rect 17995 586 18014 612
rect 18078 608 18109 620
rect 18124 608 18227 620
rect 18239 610 18265 636
rect 18280 631 18310 642
rect 18342 638 18404 654
rect 18342 636 18388 638
rect 18342 620 18404 636
rect 18416 620 18422 668
rect 18425 660 18505 668
rect 18425 658 18444 660
rect 18459 658 18493 660
rect 18425 642 18505 658
rect 18425 620 18444 642
rect 18459 626 18489 642
rect 18517 636 18523 710
rect 18532 636 18545 780
rect 18285 610 18388 620
rect 18239 608 18388 610
rect 18409 608 18444 620
rect 18078 606 18240 608
rect 18090 586 18109 606
rect 18124 604 18154 606
rect 17973 578 18014 586
rect 18096 583 18109 586
rect 18161 590 18240 606
rect 18272 606 18444 608
rect 18272 590 18351 606
rect 18358 604 18388 606
rect 17936 568 17965 578
rect 17979 568 18008 578
rect 18023 568 18053 583
rect 18096 579 18139 583
rect 18161 579 18351 590
rect 18416 586 18422 606
rect 18373 579 18403 583
rect 18096 578 18403 579
rect 18096 568 18139 578
rect 18146 568 18176 578
rect 18177 568 18335 578
rect 18339 568 18369 578
rect 18373 568 18403 578
rect 18431 568 18444 606
rect 18516 620 18545 636
rect 18516 612 18551 620
rect 18516 586 18517 612
rect 18524 586 18551 612
rect 18459 568 18489 583
rect 18516 578 18551 586
rect 18516 568 18545 578
rect -1 562 18545 568
rect 0 555 18545 562
rect 0 554 9211 555
rect 15 524 28 554
rect 43 540 73 554
rect 116 540 159 554
rect 166 540 386 554
rect 393 540 423 554
rect 83 526 98 538
rect 117 526 130 540
rect 198 536 351 540
rect 80 524 102 526
rect 180 524 372 536
rect 451 524 464 554
rect 479 540 509 554
rect 546 524 565 554
rect 580 524 586 554
rect 595 524 608 554
rect 623 540 653 554
rect 696 540 739 554
rect 746 540 966 554
rect 973 540 1003 554
rect 663 526 678 538
rect 697 526 710 540
rect 778 536 931 540
rect 660 524 682 526
rect 760 524 952 536
rect 1031 524 1044 554
rect 1059 540 1089 554
rect 1126 524 1145 554
rect 1160 524 1166 554
rect 1175 524 1188 554
rect 1203 540 1233 554
rect 1276 540 1319 554
rect 1326 540 1546 554
rect 1553 540 1583 554
rect 1243 526 1258 538
rect 1277 526 1290 540
rect 1358 536 1511 540
rect 1240 524 1262 526
rect 1340 524 1532 536
rect 1611 524 1624 554
rect 1639 540 1669 554
rect 1706 524 1725 554
rect 1740 524 1746 554
rect 1755 524 1768 554
rect 1783 540 1813 554
rect 1856 540 1899 554
rect 1906 540 2126 554
rect 2133 540 2163 554
rect 1823 526 1838 538
rect 1857 526 1870 540
rect 1938 536 2091 540
rect 1820 524 1842 526
rect 1920 524 2112 536
rect 2191 524 2204 554
rect 2219 540 2249 554
rect 2286 524 2305 554
rect 2320 524 2326 554
rect 2335 524 2348 554
rect 2363 540 2393 554
rect 2436 540 2479 554
rect 2486 540 2706 554
rect 2713 540 2743 554
rect 2403 526 2418 538
rect 2437 526 2450 540
rect 2518 536 2671 540
rect 2400 524 2422 526
rect 2500 524 2692 536
rect 2771 524 2784 554
rect 2799 540 2829 554
rect 2866 524 2885 554
rect 2900 524 2906 554
rect 2915 524 2928 554
rect 2943 540 2973 554
rect 3016 540 3059 554
rect 3066 540 3286 554
rect 3293 540 3323 554
rect 2983 526 2998 538
rect 3017 526 3030 540
rect 3098 536 3251 540
rect 2980 524 3002 526
rect 3080 524 3272 536
rect 3351 524 3364 554
rect 3379 540 3409 554
rect 3446 524 3465 554
rect 3480 524 3486 554
rect 3495 524 3508 554
rect 3523 540 3553 554
rect 3596 540 3639 554
rect 3646 540 3866 554
rect 3873 540 3903 554
rect 3563 526 3578 538
rect 3597 526 3610 540
rect 3678 536 3831 540
rect 3560 524 3582 526
rect 3660 524 3852 536
rect 3931 524 3944 554
rect 3959 540 3989 554
rect 4026 524 4045 554
rect 4060 524 4066 554
rect 4075 524 4088 554
rect 4103 540 4133 554
rect 4176 540 4219 554
rect 4226 540 4446 554
rect 4453 540 4483 554
rect 4143 526 4158 538
rect 4177 526 4190 540
rect 4258 536 4411 540
rect 4140 524 4162 526
rect 4240 524 4432 536
rect 4511 524 4524 554
rect 4539 540 4569 554
rect 4606 524 4625 554
rect 4640 525 4646 554
rect 4655 525 4668 554
rect 4683 541 4713 554
rect 4756 541 4799 554
rect 4723 527 4738 539
rect 4757 527 4770 541
rect 4806 540 5026 554
rect 5033 541 5063 554
rect 4838 537 4991 540
rect 4720 525 4742 527
rect 4820 525 5012 537
rect 5091 525 5104 554
rect 5119 541 5149 554
rect 5186 525 5205 554
rect 5220 525 5226 554
rect 5235 525 5248 554
rect 5263 541 5293 554
rect 5336 541 5379 554
rect 5303 527 5318 539
rect 5337 527 5350 541
rect 5386 540 5606 554
rect 5613 541 5643 554
rect 5418 537 5571 540
rect 5300 525 5322 527
rect 5400 525 5592 537
rect 5671 525 5684 554
rect 5699 541 5729 554
rect 5766 525 5785 554
rect 5800 525 5806 554
rect 5815 525 5828 554
rect 5843 541 5873 554
rect 5916 541 5959 554
rect 5883 527 5898 539
rect 5917 527 5930 541
rect 5966 540 6186 554
rect 6193 541 6223 554
rect 5998 537 6151 540
rect 5880 525 5902 527
rect 5980 525 6172 537
rect 6251 525 6264 554
rect 6279 541 6309 554
rect 6346 525 6365 554
rect 6380 525 6386 554
rect 6395 525 6408 554
rect 6423 541 6453 554
rect 6496 541 6539 554
rect 6463 527 6478 539
rect 6497 527 6510 541
rect 6546 540 6766 554
rect 6773 541 6803 554
rect 6578 537 6731 540
rect 6460 525 6482 527
rect 6560 525 6752 537
rect 6831 525 6844 554
rect 6859 541 6889 554
rect 6926 525 6945 554
rect 6960 525 6966 554
rect 6975 525 6988 554
rect 7003 541 7033 554
rect 7076 541 7119 554
rect 7043 527 7058 539
rect 7077 527 7090 541
rect 7126 540 7346 554
rect 7353 541 7383 554
rect 7158 537 7311 540
rect 7040 525 7062 527
rect 7140 525 7332 537
rect 7411 525 7424 554
rect 7439 541 7469 554
rect 7506 525 7525 554
rect 7540 525 7546 554
rect 7555 525 7568 554
rect 7583 541 7613 554
rect 7656 541 7699 554
rect 7623 527 7638 539
rect 7657 527 7670 541
rect 7706 540 7926 554
rect 7933 541 7963 554
rect 7738 537 7891 540
rect 7620 525 7642 527
rect 7720 525 7912 537
rect 7991 525 8004 554
rect 8019 541 8049 554
rect 8086 525 8105 554
rect 8120 525 8126 554
rect 8135 525 8148 554
rect 8163 541 8193 554
rect 8236 541 8279 554
rect 8203 527 8218 539
rect 8237 527 8250 541
rect 8286 540 8506 554
rect 8513 541 8543 554
rect 8318 537 8471 540
rect 8200 525 8222 527
rect 8300 525 8492 537
rect 8571 525 8584 554
rect 8599 541 8629 554
rect 8666 525 8685 554
rect 8700 525 8706 554
rect 8715 525 8728 554
rect 8743 541 8773 554
rect 8816 541 8859 554
rect 8783 527 8798 539
rect 8817 527 8830 541
rect 8866 540 9086 554
rect 9093 541 9123 554
rect 8898 537 9051 540
rect 8780 525 8802 527
rect 8880 525 9072 537
rect 9151 525 9164 554
rect 9179 541 9209 554
rect 9246 525 9265 555
rect 9280 525 9286 555
rect 9295 525 9308 555
rect 9323 554 18545 555
rect 9323 541 9353 554
rect 9396 541 9439 554
rect 9363 527 9378 539
rect 9397 527 9410 541
rect 9446 540 9666 554
rect 9673 541 9703 554
rect 9478 537 9631 540
rect 9360 525 9382 527
rect 9460 525 9652 537
rect 9731 525 9744 554
rect 9759 541 9789 554
rect 9826 525 9845 554
rect 9860 525 9866 554
rect 9875 525 9888 554
rect 9903 541 9933 554
rect 9976 541 10019 554
rect 9943 527 9958 539
rect 9977 527 9990 541
rect 10026 540 10246 554
rect 10253 541 10283 554
rect 10058 537 10211 540
rect 9940 525 9962 527
rect 10040 525 10232 537
rect 10311 525 10324 554
rect 10339 541 10369 554
rect 10406 525 10425 554
rect 10440 525 10446 554
rect 10455 525 10468 554
rect 10483 541 10513 554
rect 10556 541 10599 554
rect 10523 527 10538 539
rect 10557 527 10570 541
rect 10606 540 10826 554
rect 10833 541 10863 554
rect 10638 537 10791 540
rect 10520 525 10542 527
rect 10620 525 10812 537
rect 10891 525 10904 554
rect 10919 541 10949 554
rect 10986 525 11005 554
rect 11020 525 11026 554
rect 11035 525 11048 554
rect 11063 541 11093 554
rect 11136 541 11179 554
rect 11103 527 11118 539
rect 11137 527 11150 541
rect 11186 540 11406 554
rect 11413 541 11443 554
rect 11218 537 11371 540
rect 11100 525 11122 527
rect 11200 525 11392 537
rect 11471 525 11484 554
rect 11499 541 11529 554
rect 11566 525 11585 554
rect 11600 525 11606 554
rect 11615 525 11628 554
rect 11643 541 11673 554
rect 11716 541 11759 554
rect 11683 527 11698 539
rect 11717 527 11730 541
rect 11766 540 11986 554
rect 11993 541 12023 554
rect 11798 537 11951 540
rect 11680 525 11702 527
rect 11780 525 11972 537
rect 12051 525 12064 554
rect 12079 541 12109 554
rect 12146 525 12165 554
rect 12180 525 12186 554
rect 12195 525 12208 554
rect 12223 541 12253 554
rect 12296 541 12339 554
rect 12263 527 12278 539
rect 12297 527 12310 541
rect 12346 540 12566 554
rect 12573 541 12603 554
rect 12378 537 12531 540
rect 12260 525 12282 527
rect 12360 525 12552 537
rect 12631 525 12644 554
rect 12659 541 12689 554
rect 12726 525 12745 554
rect 12760 525 12766 554
rect 12775 525 12788 554
rect 12803 541 12833 554
rect 12876 541 12919 554
rect 12843 527 12858 539
rect 12877 527 12890 541
rect 12926 540 13146 554
rect 13153 541 13183 554
rect 12958 537 13111 540
rect 12840 525 12862 527
rect 12940 525 13132 537
rect 13211 525 13224 554
rect 13239 541 13269 554
rect 13306 525 13325 554
rect 13340 525 13346 554
rect 13355 525 13368 554
rect 13383 541 13413 554
rect 13456 541 13499 554
rect 13423 527 13438 539
rect 13457 527 13470 541
rect 13506 540 13726 554
rect 13733 541 13763 554
rect 13538 537 13691 540
rect 13420 525 13442 527
rect 13520 525 13712 537
rect 13791 525 13804 554
rect 13819 541 13849 554
rect 13886 525 13905 554
rect 13920 541 13926 554
rect 13920 540 13934 541
rect 13920 525 13926 540
rect 13935 525 13948 554
rect 13963 541 13993 554
rect 14036 541 14079 554
rect 14003 527 14018 539
rect 14037 527 14050 541
rect 14086 540 14306 554
rect 14313 541 14343 554
rect 14118 537 14271 540
rect 14000 525 14022 527
rect 14100 525 14292 537
rect 14371 525 14384 554
rect 14399 541 14429 554
rect 14466 525 14485 554
rect 14500 525 14506 554
rect 14515 525 14528 554
rect 14543 541 14573 554
rect 14616 541 14659 554
rect 14583 527 14598 539
rect 14617 527 14630 541
rect 14666 540 14886 554
rect 14893 541 14923 554
rect 14698 537 14851 540
rect 14580 525 14602 527
rect 14680 525 14872 537
rect 14951 525 14964 554
rect 14979 541 15009 554
rect 15046 525 15065 554
rect 15080 525 15086 554
rect 15095 525 15108 554
rect 15123 541 15153 554
rect 15196 541 15239 554
rect 15163 527 15178 539
rect 15197 527 15210 541
rect 15246 540 15466 554
rect 15473 541 15503 554
rect 15278 537 15431 540
rect 15160 525 15182 527
rect 15260 525 15452 537
rect 15531 525 15544 554
rect 15559 541 15589 554
rect 15626 525 15645 554
rect 15660 525 15666 554
rect 15675 525 15688 554
rect 15703 541 15733 554
rect 15776 541 15819 554
rect 15743 527 15758 539
rect 15777 527 15790 541
rect 15826 540 16046 554
rect 16053 541 16083 554
rect 15858 537 16011 540
rect 15740 525 15762 527
rect 15840 525 16032 537
rect 16111 525 16124 554
rect 16139 541 16169 554
rect 16206 525 16225 554
rect 16240 525 16246 554
rect 16255 525 16268 554
rect 16283 541 16313 554
rect 16356 541 16399 554
rect 16323 527 16338 539
rect 16357 527 16370 541
rect 16406 540 16626 554
rect 16633 541 16663 554
rect 16438 537 16591 540
rect 16320 525 16342 527
rect 16420 525 16612 537
rect 16691 525 16704 554
rect 16719 541 16749 554
rect 16786 525 16805 554
rect 16820 525 16826 554
rect 16835 525 16848 554
rect 16863 541 16893 554
rect 16936 541 16979 554
rect 16903 527 16918 539
rect 16937 527 16950 541
rect 16986 540 17206 554
rect 17213 541 17243 554
rect 17018 537 17171 540
rect 16900 525 16922 527
rect 17000 525 17192 537
rect 17271 525 17284 554
rect 17299 541 17329 554
rect 17366 525 17385 554
rect 17400 525 17406 554
rect 17415 525 17428 554
rect 17443 541 17473 554
rect 17516 541 17559 554
rect 17483 527 17498 539
rect 17517 527 17530 541
rect 17566 540 17786 554
rect 17793 541 17823 554
rect 17598 537 17751 540
rect 17480 525 17502 527
rect 17580 525 17772 537
rect 17851 525 17864 554
rect 17879 541 17909 554
rect 17946 525 17965 554
rect 17980 525 17986 554
rect 17995 525 18008 554
rect 18023 541 18053 554
rect 18096 541 18139 554
rect 18063 527 18078 539
rect 18097 527 18110 541
rect 18146 540 18366 554
rect 18373 541 18403 554
rect 18178 537 18331 540
rect 18060 525 18082 527
rect 18160 525 18352 537
rect 18431 525 18444 554
rect 18459 541 18489 554
rect 18532 525 18545 554
rect 4627 524 18545 525
rect -13 511 18545 524
rect -13 510 4646 511
rect -13 496 0 510
rect 15 440 28 510
rect 80 506 102 510
rect 73 484 102 498
rect 155 484 171 498
rect 209 494 215 496
rect 222 494 330 510
rect 337 494 343 496
rect 351 494 366 510
rect 432 504 451 507
rect 73 482 171 484
rect 198 482 366 494
rect 381 484 397 498
rect 432 485 454 504
rect 464 498 480 499
rect 463 496 480 498
rect 464 491 480 496
rect 454 484 460 485
rect 463 484 492 491
rect 381 483 492 484
rect 381 482 498 483
rect 57 474 108 482
rect 155 474 189 482
rect 57 462 82 474
rect 89 462 108 474
rect 162 472 189 474
rect 198 472 419 482
rect 454 479 460 482
rect 162 468 419 472
rect 57 454 108 462
rect 155 454 419 468
rect 463 474 498 482
rect 9 406 28 440
rect 73 446 102 454
rect 73 440 90 446
rect 73 438 107 440
rect 155 438 171 454
rect 172 444 380 454
rect 381 444 397 454
rect 445 450 460 465
rect 463 462 464 474
rect 471 462 498 474
rect 463 454 498 462
rect 463 453 492 454
rect 183 440 397 444
rect 198 438 397 440
rect 432 440 445 450
rect 463 440 480 453
rect 432 438 480 440
rect 74 434 107 438
rect 70 432 107 434
rect 70 431 137 432
rect 70 426 101 431
rect 107 426 137 431
rect 70 422 137 426
rect 43 419 137 422
rect 43 412 92 419
rect 43 406 73 412
rect 92 407 97 412
rect -13 372 0 400
rect 9 390 89 406
rect 101 398 137 419
rect 198 414 387 438
rect 432 437 479 438
rect 445 432 479 437
rect 213 411 387 414
rect 206 408 387 411
rect 415 431 479 432
rect 9 388 28 390
rect 43 388 77 390
rect 9 372 89 388
rect 9 366 28 372
rect -1 350 28 366
rect 43 356 73 372
rect 101 350 107 398
rect 110 392 129 398
rect 144 392 174 400
rect 110 384 174 392
rect 110 368 190 384
rect 206 377 268 408
rect 284 377 346 408
rect 415 406 464 431
rect 479 406 509 422
rect 378 392 408 400
rect 415 398 525 406
rect 378 384 423 392
rect 110 366 129 368
rect 144 366 190 368
rect 110 350 190 366
rect 217 364 252 377
rect 293 374 330 377
rect 293 372 335 374
rect 222 361 252 364
rect 231 357 238 361
rect 238 356 239 357
rect 197 350 207 356
rect -7 342 34 350
rect -7 316 8 342
rect 15 316 34 342
rect 98 338 129 350
rect 144 338 247 350
rect 259 340 285 366
rect 300 361 330 372
rect 362 368 424 384
rect 362 366 408 368
rect 362 350 424 366
rect 436 350 442 398
rect 445 390 525 398
rect 445 388 464 390
rect 479 388 513 390
rect 445 372 525 388
rect 445 350 464 372
rect 479 356 509 372
rect 537 366 543 440
rect 546 366 565 510
rect 580 366 586 510
rect 595 440 608 510
rect 660 506 682 510
rect 653 484 682 498
rect 735 484 751 498
rect 789 494 795 496
rect 802 494 910 510
rect 917 494 923 496
rect 931 494 946 510
rect 1012 504 1031 507
rect 653 482 751 484
rect 778 482 946 494
rect 961 484 977 498
rect 1012 485 1034 504
rect 1044 498 1060 499
rect 1043 496 1060 498
rect 1044 491 1060 496
rect 1034 484 1040 485
rect 1043 484 1072 491
rect 961 483 1072 484
rect 961 482 1078 483
rect 637 474 688 482
rect 735 474 769 482
rect 637 462 662 474
rect 669 462 688 474
rect 742 472 769 474
rect 778 472 999 482
rect 1034 479 1040 482
rect 742 468 999 472
rect 637 454 688 462
rect 735 454 999 468
rect 1043 474 1078 482
rect 589 406 608 440
rect 653 446 682 454
rect 653 440 670 446
rect 653 438 687 440
rect 735 438 751 454
rect 752 444 960 454
rect 961 444 977 454
rect 1025 450 1040 465
rect 1043 462 1044 474
rect 1051 462 1078 474
rect 1043 454 1078 462
rect 1043 453 1072 454
rect 763 440 977 444
rect 778 438 977 440
rect 1012 440 1025 450
rect 1043 440 1060 453
rect 1012 438 1060 440
rect 654 434 687 438
rect 650 432 687 434
rect 650 431 717 432
rect 650 426 681 431
rect 687 426 717 431
rect 650 422 717 426
rect 623 419 717 422
rect 623 412 672 419
rect 623 406 653 412
rect 672 407 677 412
rect 589 390 669 406
rect 681 398 717 419
rect 778 414 967 438
rect 1012 437 1059 438
rect 1025 432 1059 437
rect 793 411 967 414
rect 786 408 967 411
rect 995 431 1059 432
rect 589 388 608 390
rect 623 388 657 390
rect 589 372 669 388
rect 589 366 608 372
rect 305 340 408 350
rect 259 338 408 340
rect 429 338 464 350
rect 98 336 260 338
rect 110 316 129 336
rect 144 334 174 336
rect -7 308 34 316
rect 116 312 129 316
rect 181 320 260 336
rect 292 336 464 338
rect 292 320 371 336
rect 378 334 408 336
rect -1 298 28 308
rect 43 298 73 312
rect 116 298 159 312
rect 181 308 371 320
rect 436 316 442 336
rect 166 298 196 308
rect 197 298 355 308
rect 359 298 389 308
rect 393 298 423 312
rect 451 298 464 336
rect 536 350 565 366
rect 579 350 608 366
rect 623 356 653 372
rect 681 350 687 398
rect 690 392 709 398
rect 724 392 754 400
rect 690 384 754 392
rect 690 368 770 384
rect 786 377 848 408
rect 864 377 926 408
rect 995 406 1044 431
rect 1059 406 1089 422
rect 958 392 988 400
rect 995 398 1105 406
rect 958 384 1003 392
rect 690 366 709 368
rect 724 366 770 368
rect 690 350 770 366
rect 797 364 832 377
rect 873 374 910 377
rect 873 372 915 374
rect 802 361 832 364
rect 811 357 818 361
rect 818 356 819 357
rect 777 350 787 356
rect 536 342 571 350
rect 536 316 537 342
rect 544 316 571 342
rect 479 298 509 312
rect 536 308 571 316
rect 573 342 614 350
rect 573 316 588 342
rect 595 316 614 342
rect 678 338 709 350
rect 724 338 827 350
rect 839 340 865 366
rect 880 361 910 372
rect 942 368 1004 384
rect 942 366 988 368
rect 942 350 1004 366
rect 1016 350 1022 398
rect 1025 390 1105 398
rect 1025 388 1044 390
rect 1059 388 1093 390
rect 1025 372 1105 388
rect 1025 350 1044 372
rect 1059 356 1089 372
rect 1117 366 1123 440
rect 1126 366 1145 510
rect 1160 366 1166 510
rect 1175 440 1188 510
rect 1240 506 1262 510
rect 1233 484 1262 498
rect 1315 484 1331 498
rect 1369 494 1375 496
rect 1382 494 1490 510
rect 1497 494 1503 496
rect 1511 494 1526 510
rect 1592 504 1611 507
rect 1233 482 1331 484
rect 1358 482 1526 494
rect 1541 484 1557 498
rect 1592 485 1614 504
rect 1624 498 1640 499
rect 1623 496 1640 498
rect 1624 491 1640 496
rect 1614 484 1620 485
rect 1623 484 1652 491
rect 1541 483 1652 484
rect 1541 482 1658 483
rect 1217 474 1268 482
rect 1315 474 1349 482
rect 1217 462 1242 474
rect 1249 462 1268 474
rect 1322 472 1349 474
rect 1358 472 1579 482
rect 1614 479 1620 482
rect 1322 468 1579 472
rect 1217 454 1268 462
rect 1315 454 1579 468
rect 1623 474 1658 482
rect 1169 406 1188 440
rect 1233 446 1262 454
rect 1233 440 1250 446
rect 1233 438 1267 440
rect 1315 438 1331 454
rect 1332 444 1540 454
rect 1541 444 1557 454
rect 1605 450 1620 465
rect 1623 462 1624 474
rect 1631 462 1658 474
rect 1623 454 1658 462
rect 1623 453 1652 454
rect 1343 440 1557 444
rect 1358 438 1557 440
rect 1592 440 1605 450
rect 1623 440 1640 453
rect 1592 438 1640 440
rect 1234 434 1267 438
rect 1230 432 1267 434
rect 1230 431 1297 432
rect 1230 426 1261 431
rect 1267 426 1297 431
rect 1230 422 1297 426
rect 1203 419 1297 422
rect 1203 412 1252 419
rect 1203 406 1233 412
rect 1252 407 1257 412
rect 1169 390 1249 406
rect 1261 398 1297 419
rect 1358 414 1547 438
rect 1592 437 1639 438
rect 1605 432 1639 437
rect 1373 411 1547 414
rect 1366 408 1547 411
rect 1575 431 1639 432
rect 1169 388 1188 390
rect 1203 388 1237 390
rect 1169 372 1249 388
rect 1169 366 1188 372
rect 885 340 988 350
rect 839 338 988 340
rect 1009 338 1044 350
rect 678 336 840 338
rect 690 316 709 336
rect 724 334 754 336
rect 573 308 614 316
rect 696 312 709 316
rect 761 320 840 336
rect 872 336 1044 338
rect 872 320 951 336
rect 958 334 988 336
rect 536 298 565 308
rect 579 298 608 308
rect 623 298 653 312
rect 696 298 739 312
rect 761 308 951 320
rect 1016 316 1022 336
rect 746 298 776 308
rect 777 298 935 308
rect 939 298 969 308
rect 973 298 1003 312
rect 1031 298 1044 336
rect 1116 350 1145 366
rect 1159 350 1188 366
rect 1203 356 1233 372
rect 1261 350 1267 398
rect 1270 392 1289 398
rect 1304 392 1334 400
rect 1270 384 1334 392
rect 1270 368 1350 384
rect 1366 377 1428 408
rect 1444 377 1506 408
rect 1575 406 1624 431
rect 1639 406 1669 422
rect 1538 392 1568 400
rect 1575 398 1685 406
rect 1538 384 1583 392
rect 1270 366 1289 368
rect 1304 366 1350 368
rect 1270 350 1350 366
rect 1377 364 1412 377
rect 1453 374 1490 377
rect 1453 372 1495 374
rect 1382 361 1412 364
rect 1391 357 1398 361
rect 1398 356 1399 357
rect 1357 350 1367 356
rect 1116 342 1151 350
rect 1116 316 1117 342
rect 1124 316 1151 342
rect 1059 298 1089 312
rect 1116 308 1151 316
rect 1153 342 1194 350
rect 1153 316 1168 342
rect 1175 316 1194 342
rect 1258 338 1289 350
rect 1304 338 1407 350
rect 1419 340 1445 366
rect 1460 361 1490 372
rect 1522 368 1584 384
rect 1522 366 1568 368
rect 1522 350 1584 366
rect 1596 350 1602 398
rect 1605 390 1685 398
rect 1605 388 1624 390
rect 1639 388 1673 390
rect 1605 372 1685 388
rect 1605 350 1624 372
rect 1639 356 1669 372
rect 1697 366 1703 440
rect 1706 366 1725 510
rect 1740 366 1746 510
rect 1755 440 1768 510
rect 1820 506 1842 510
rect 1813 484 1842 498
rect 1895 484 1911 498
rect 1949 494 1955 496
rect 1962 494 2070 510
rect 2077 494 2083 496
rect 2091 494 2106 510
rect 2172 504 2191 507
rect 1813 482 1911 484
rect 1938 482 2106 494
rect 2121 484 2137 498
rect 2172 485 2194 504
rect 2204 498 2220 499
rect 2203 496 2220 498
rect 2204 491 2220 496
rect 2194 484 2200 485
rect 2203 484 2232 491
rect 2121 483 2232 484
rect 2121 482 2238 483
rect 1797 474 1848 482
rect 1895 474 1929 482
rect 1797 462 1822 474
rect 1829 462 1848 474
rect 1902 472 1929 474
rect 1938 472 2159 482
rect 2194 479 2200 482
rect 1902 468 2159 472
rect 1797 454 1848 462
rect 1895 454 2159 468
rect 2203 474 2238 482
rect 1749 406 1768 440
rect 1813 446 1842 454
rect 1813 440 1830 446
rect 1813 438 1847 440
rect 1895 438 1911 454
rect 1912 444 2120 454
rect 2121 444 2137 454
rect 2185 450 2200 465
rect 2203 462 2204 474
rect 2211 462 2238 474
rect 2203 454 2238 462
rect 2203 453 2232 454
rect 1923 440 2137 444
rect 1938 438 2137 440
rect 2172 440 2185 450
rect 2203 440 2220 453
rect 2172 438 2220 440
rect 1814 434 1847 438
rect 1810 432 1847 434
rect 1810 431 1877 432
rect 1810 426 1841 431
rect 1847 426 1877 431
rect 1810 422 1877 426
rect 1783 419 1877 422
rect 1783 412 1832 419
rect 1783 406 1813 412
rect 1832 407 1837 412
rect 1749 390 1829 406
rect 1841 398 1877 419
rect 1938 414 2127 438
rect 2172 437 2219 438
rect 2185 432 2219 437
rect 1953 411 2127 414
rect 1946 408 2127 411
rect 2155 431 2219 432
rect 1749 388 1768 390
rect 1783 388 1817 390
rect 1749 372 1829 388
rect 1749 366 1768 372
rect 1465 340 1568 350
rect 1419 338 1568 340
rect 1589 338 1624 350
rect 1258 336 1420 338
rect 1270 316 1289 336
rect 1304 334 1334 336
rect 1153 308 1194 316
rect 1276 312 1289 316
rect 1341 320 1420 336
rect 1452 336 1624 338
rect 1452 320 1531 336
rect 1538 334 1568 336
rect 1116 298 1145 308
rect 1159 298 1188 308
rect 1203 298 1233 312
rect 1276 298 1319 312
rect 1341 308 1531 320
rect 1596 316 1602 336
rect 1326 298 1356 308
rect 1357 298 1515 308
rect 1519 298 1549 308
rect 1553 298 1583 312
rect 1611 298 1624 336
rect 1696 350 1725 366
rect 1739 350 1768 366
rect 1783 356 1813 372
rect 1841 350 1847 398
rect 1850 392 1869 398
rect 1884 392 1914 400
rect 1850 384 1914 392
rect 1850 368 1930 384
rect 1946 377 2008 408
rect 2024 377 2086 408
rect 2155 406 2204 431
rect 2219 406 2249 422
rect 2118 392 2148 400
rect 2155 398 2265 406
rect 2118 384 2163 392
rect 1850 366 1869 368
rect 1884 366 1930 368
rect 1850 350 1930 366
rect 1957 364 1992 377
rect 2033 374 2070 377
rect 2033 372 2075 374
rect 1962 361 1992 364
rect 1971 357 1978 361
rect 1978 356 1979 357
rect 1937 350 1947 356
rect 1696 342 1731 350
rect 1696 316 1697 342
rect 1704 316 1731 342
rect 1639 298 1669 312
rect 1696 308 1731 316
rect 1733 342 1774 350
rect 1733 316 1748 342
rect 1755 316 1774 342
rect 1838 338 1869 350
rect 1884 338 1987 350
rect 1999 340 2025 366
rect 2040 361 2070 372
rect 2102 368 2164 384
rect 2102 366 2148 368
rect 2102 350 2164 366
rect 2176 350 2182 398
rect 2185 390 2265 398
rect 2185 388 2204 390
rect 2219 388 2253 390
rect 2185 372 2265 388
rect 2185 350 2204 372
rect 2219 356 2249 372
rect 2277 366 2283 440
rect 2286 366 2305 510
rect 2320 366 2326 510
rect 2335 440 2348 510
rect 2400 506 2422 510
rect 2393 484 2422 498
rect 2475 484 2491 498
rect 2529 494 2535 496
rect 2542 494 2650 510
rect 2657 494 2663 496
rect 2671 494 2686 510
rect 2752 504 2771 507
rect 2393 482 2491 484
rect 2518 482 2686 494
rect 2701 484 2717 498
rect 2752 485 2774 504
rect 2784 498 2800 499
rect 2783 496 2800 498
rect 2784 491 2800 496
rect 2774 484 2780 485
rect 2783 484 2812 491
rect 2701 483 2812 484
rect 2701 482 2818 483
rect 2377 474 2428 482
rect 2475 474 2509 482
rect 2377 462 2402 474
rect 2409 462 2428 474
rect 2482 472 2509 474
rect 2518 472 2739 482
rect 2774 479 2780 482
rect 2482 468 2739 472
rect 2377 454 2428 462
rect 2475 454 2739 468
rect 2783 474 2818 482
rect 2329 406 2348 440
rect 2393 446 2422 454
rect 2393 440 2410 446
rect 2393 438 2427 440
rect 2475 438 2491 454
rect 2492 444 2700 454
rect 2701 444 2717 454
rect 2765 450 2780 465
rect 2783 462 2784 474
rect 2791 462 2818 474
rect 2783 454 2818 462
rect 2783 453 2812 454
rect 2503 440 2717 444
rect 2518 438 2717 440
rect 2752 440 2765 450
rect 2783 440 2800 453
rect 2752 438 2800 440
rect 2394 434 2427 438
rect 2390 432 2427 434
rect 2390 431 2457 432
rect 2390 426 2421 431
rect 2427 426 2457 431
rect 2390 422 2457 426
rect 2363 419 2457 422
rect 2363 412 2412 419
rect 2363 406 2393 412
rect 2412 407 2417 412
rect 2329 390 2409 406
rect 2421 398 2457 419
rect 2518 414 2707 438
rect 2752 437 2799 438
rect 2765 432 2799 437
rect 2533 411 2707 414
rect 2526 408 2707 411
rect 2735 431 2799 432
rect 2329 388 2348 390
rect 2363 388 2397 390
rect 2329 372 2409 388
rect 2329 366 2348 372
rect 2045 340 2148 350
rect 1999 338 2148 340
rect 2169 338 2204 350
rect 1838 336 2000 338
rect 1850 316 1869 336
rect 1884 334 1914 336
rect 1733 308 1774 316
rect 1856 312 1869 316
rect 1921 320 2000 336
rect 2032 336 2204 338
rect 2032 320 2111 336
rect 2118 334 2148 336
rect 1696 298 1725 308
rect 1739 298 1768 308
rect 1783 298 1813 312
rect 1856 298 1899 312
rect 1921 308 2111 320
rect 2176 316 2182 336
rect 1906 298 1936 308
rect 1937 298 2095 308
rect 2099 298 2129 308
rect 2133 298 2163 312
rect 2191 298 2204 336
rect 2276 350 2305 366
rect 2319 350 2348 366
rect 2363 356 2393 372
rect 2421 350 2427 398
rect 2430 392 2449 398
rect 2464 392 2494 400
rect 2430 384 2494 392
rect 2430 368 2510 384
rect 2526 377 2588 408
rect 2604 377 2666 408
rect 2735 406 2784 431
rect 2799 406 2829 422
rect 2698 392 2728 400
rect 2735 398 2845 406
rect 2698 384 2743 392
rect 2430 366 2449 368
rect 2464 366 2510 368
rect 2430 350 2510 366
rect 2537 364 2572 377
rect 2613 374 2650 377
rect 2613 372 2655 374
rect 2542 361 2572 364
rect 2551 357 2558 361
rect 2558 356 2559 357
rect 2517 350 2527 356
rect 2276 342 2311 350
rect 2276 316 2277 342
rect 2284 316 2311 342
rect 2219 298 2249 312
rect 2276 308 2311 316
rect 2313 342 2354 350
rect 2313 316 2328 342
rect 2335 316 2354 342
rect 2418 338 2449 350
rect 2464 338 2567 350
rect 2579 340 2605 366
rect 2620 361 2650 372
rect 2682 368 2744 384
rect 2682 366 2728 368
rect 2682 350 2744 366
rect 2756 350 2762 398
rect 2765 390 2845 398
rect 2765 388 2784 390
rect 2799 388 2833 390
rect 2765 372 2845 388
rect 2765 350 2784 372
rect 2799 356 2829 372
rect 2857 366 2863 440
rect 2866 366 2885 510
rect 2900 366 2906 510
rect 2915 440 2928 510
rect 2980 506 3002 510
rect 2973 484 3002 498
rect 3055 484 3071 498
rect 3109 494 3115 496
rect 3122 494 3230 510
rect 3237 494 3243 496
rect 3251 494 3266 510
rect 3332 504 3351 507
rect 2973 482 3071 484
rect 3098 482 3266 494
rect 3281 484 3297 498
rect 3332 485 3354 504
rect 3364 498 3380 499
rect 3363 496 3380 498
rect 3364 491 3380 496
rect 3354 484 3360 485
rect 3363 484 3392 491
rect 3281 483 3392 484
rect 3281 482 3398 483
rect 2957 474 3008 482
rect 3055 474 3089 482
rect 2957 462 2982 474
rect 2989 462 3008 474
rect 3062 472 3089 474
rect 3098 472 3319 482
rect 3354 479 3360 482
rect 3062 468 3319 472
rect 2957 454 3008 462
rect 3055 454 3319 468
rect 3363 474 3398 482
rect 2909 406 2928 440
rect 2973 446 3002 454
rect 2973 440 2990 446
rect 2973 438 3007 440
rect 3055 438 3071 454
rect 3072 444 3280 454
rect 3281 444 3297 454
rect 3345 450 3360 465
rect 3363 462 3364 474
rect 3371 462 3398 474
rect 3363 454 3398 462
rect 3363 453 3392 454
rect 3083 440 3297 444
rect 3098 438 3297 440
rect 3332 440 3345 450
rect 3363 440 3380 453
rect 3332 438 3380 440
rect 2974 434 3007 438
rect 2970 432 3007 434
rect 2970 431 3037 432
rect 2970 426 3001 431
rect 3007 426 3037 431
rect 2970 422 3037 426
rect 2943 419 3037 422
rect 2943 412 2992 419
rect 2943 406 2973 412
rect 2992 407 2997 412
rect 2909 390 2989 406
rect 3001 398 3037 419
rect 3098 414 3287 438
rect 3332 437 3379 438
rect 3345 432 3379 437
rect 3113 411 3287 414
rect 3106 408 3287 411
rect 3315 431 3379 432
rect 2909 388 2928 390
rect 2943 388 2977 390
rect 2909 372 2989 388
rect 2909 366 2928 372
rect 2625 340 2728 350
rect 2579 338 2728 340
rect 2749 338 2784 350
rect 2418 336 2580 338
rect 2430 316 2449 336
rect 2464 334 2494 336
rect 2313 308 2354 316
rect 2436 312 2449 316
rect 2501 320 2580 336
rect 2612 336 2784 338
rect 2612 320 2691 336
rect 2698 334 2728 336
rect 2276 298 2305 308
rect 2319 298 2348 308
rect 2363 298 2393 312
rect 2436 298 2479 312
rect 2501 308 2691 320
rect 2756 316 2762 336
rect 2486 298 2516 308
rect 2517 298 2675 308
rect 2679 298 2709 308
rect 2713 298 2743 312
rect 2771 298 2784 336
rect 2856 350 2885 366
rect 2899 350 2928 366
rect 2943 356 2973 372
rect 3001 350 3007 398
rect 3010 392 3029 398
rect 3044 392 3074 400
rect 3010 384 3074 392
rect 3010 368 3090 384
rect 3106 377 3168 408
rect 3184 377 3246 408
rect 3315 406 3364 431
rect 3379 406 3409 422
rect 3278 392 3308 400
rect 3315 398 3425 406
rect 3278 384 3323 392
rect 3010 366 3029 368
rect 3044 366 3090 368
rect 3010 350 3090 366
rect 3117 364 3152 377
rect 3193 374 3230 377
rect 3193 372 3235 374
rect 3122 361 3152 364
rect 3131 357 3138 361
rect 3138 356 3139 357
rect 3097 350 3107 356
rect 2856 342 2891 350
rect 2856 316 2857 342
rect 2864 316 2891 342
rect 2799 298 2829 312
rect 2856 308 2891 316
rect 2893 342 2934 350
rect 2893 316 2908 342
rect 2915 316 2934 342
rect 2998 338 3029 350
rect 3044 338 3147 350
rect 3159 340 3185 366
rect 3200 361 3230 372
rect 3262 368 3324 384
rect 3262 366 3308 368
rect 3262 350 3324 366
rect 3336 350 3342 398
rect 3345 390 3425 398
rect 3345 388 3364 390
rect 3379 388 3413 390
rect 3345 372 3425 388
rect 3345 350 3364 372
rect 3379 356 3409 372
rect 3437 366 3443 440
rect 3446 366 3465 510
rect 3480 366 3486 510
rect 3495 440 3508 510
rect 3560 506 3582 510
rect 3553 484 3582 498
rect 3635 484 3651 498
rect 3689 494 3695 496
rect 3702 494 3810 510
rect 3817 494 3823 496
rect 3831 494 3846 510
rect 3912 504 3931 507
rect 3553 482 3651 484
rect 3678 482 3846 494
rect 3861 484 3877 498
rect 3912 485 3934 504
rect 3944 498 3960 499
rect 3943 496 3960 498
rect 3944 491 3960 496
rect 3934 484 3940 485
rect 3943 484 3972 491
rect 3861 483 3972 484
rect 3861 482 3978 483
rect 3537 474 3588 482
rect 3635 474 3669 482
rect 3537 462 3562 474
rect 3569 462 3588 474
rect 3642 472 3669 474
rect 3678 472 3899 482
rect 3934 479 3940 482
rect 3642 468 3899 472
rect 3537 454 3588 462
rect 3635 454 3899 468
rect 3943 474 3978 482
rect 3489 406 3508 440
rect 3553 446 3582 454
rect 3553 440 3570 446
rect 3553 438 3587 440
rect 3635 438 3651 454
rect 3652 444 3860 454
rect 3861 444 3877 454
rect 3925 450 3940 465
rect 3943 462 3944 474
rect 3951 462 3978 474
rect 3943 454 3978 462
rect 3943 453 3972 454
rect 3663 440 3877 444
rect 3678 438 3877 440
rect 3912 440 3925 450
rect 3943 440 3960 453
rect 3912 438 3960 440
rect 3554 434 3587 438
rect 3550 432 3587 434
rect 3550 431 3617 432
rect 3550 426 3581 431
rect 3587 426 3617 431
rect 3550 422 3617 426
rect 3523 419 3617 422
rect 3523 412 3572 419
rect 3523 406 3553 412
rect 3572 407 3577 412
rect 3489 390 3569 406
rect 3581 398 3617 419
rect 3678 414 3867 438
rect 3912 437 3959 438
rect 3925 432 3959 437
rect 3693 411 3867 414
rect 3686 408 3867 411
rect 3895 431 3959 432
rect 3489 388 3508 390
rect 3523 388 3557 390
rect 3489 372 3569 388
rect 3489 366 3508 372
rect 3205 340 3308 350
rect 3159 338 3308 340
rect 3329 338 3364 350
rect 2998 336 3160 338
rect 3010 316 3029 336
rect 3044 334 3074 336
rect 2893 308 2934 316
rect 3016 312 3029 316
rect 3081 320 3160 336
rect 3192 336 3364 338
rect 3192 320 3271 336
rect 3278 334 3308 336
rect 2856 298 2885 308
rect 2899 298 2928 308
rect 2943 298 2973 312
rect 3016 298 3059 312
rect 3081 308 3271 320
rect 3336 316 3342 336
rect 3066 298 3096 308
rect 3097 298 3255 308
rect 3259 298 3289 308
rect 3293 298 3323 312
rect 3351 298 3364 336
rect 3436 350 3465 366
rect 3479 350 3508 366
rect 3523 356 3553 372
rect 3581 350 3587 398
rect 3590 392 3609 398
rect 3624 392 3654 400
rect 3590 384 3654 392
rect 3590 368 3670 384
rect 3686 377 3748 408
rect 3764 377 3826 408
rect 3895 406 3944 431
rect 3959 406 3989 422
rect 3858 392 3888 400
rect 3895 398 4005 406
rect 3858 384 3903 392
rect 3590 366 3609 368
rect 3624 366 3670 368
rect 3590 350 3670 366
rect 3697 364 3732 377
rect 3773 374 3810 377
rect 3773 372 3815 374
rect 3702 361 3732 364
rect 3711 357 3718 361
rect 3718 356 3719 357
rect 3677 350 3687 356
rect 3436 342 3471 350
rect 3436 316 3437 342
rect 3444 316 3471 342
rect 3379 298 3409 312
rect 3436 308 3471 316
rect 3473 342 3514 350
rect 3473 316 3488 342
rect 3495 316 3514 342
rect 3578 338 3609 350
rect 3624 338 3727 350
rect 3739 340 3765 366
rect 3780 361 3810 372
rect 3842 368 3904 384
rect 3842 366 3888 368
rect 3842 350 3904 366
rect 3916 350 3922 398
rect 3925 390 4005 398
rect 3925 388 3944 390
rect 3959 388 3993 390
rect 3925 372 4005 388
rect 3925 350 3944 372
rect 3959 356 3989 372
rect 4017 366 4023 440
rect 4026 366 4045 510
rect 4060 366 4066 510
rect 4075 440 4088 510
rect 4140 506 4162 510
rect 4133 484 4162 498
rect 4215 484 4231 498
rect 4269 494 4275 496
rect 4282 494 4390 510
rect 4397 494 4403 496
rect 4411 494 4426 510
rect 4492 504 4511 507
rect 4133 482 4231 484
rect 4258 482 4426 494
rect 4441 484 4457 498
rect 4492 485 4514 504
rect 4524 498 4540 499
rect 4523 496 4540 498
rect 4524 491 4540 496
rect 4514 484 4520 485
rect 4523 484 4552 491
rect 4441 483 4552 484
rect 4441 482 4558 483
rect 4117 474 4168 482
rect 4215 474 4249 482
rect 4117 462 4142 474
rect 4149 462 4168 474
rect 4222 472 4249 474
rect 4258 472 4479 482
rect 4514 479 4520 482
rect 4222 468 4479 472
rect 4117 454 4168 462
rect 4215 454 4479 468
rect 4523 474 4558 482
rect 4069 406 4088 440
rect 4133 446 4162 454
rect 4133 440 4150 446
rect 4133 438 4167 440
rect 4215 438 4231 454
rect 4232 444 4440 454
rect 4441 444 4457 454
rect 4505 450 4520 465
rect 4523 462 4524 474
rect 4531 462 4558 474
rect 4523 454 4558 462
rect 4523 453 4552 454
rect 4243 440 4457 444
rect 4258 438 4457 440
rect 4492 440 4505 450
rect 4523 440 4540 453
rect 4492 438 4540 440
rect 4134 434 4167 438
rect 4130 432 4167 434
rect 4130 431 4197 432
rect 4130 426 4161 431
rect 4167 426 4197 431
rect 4130 422 4197 426
rect 4103 419 4197 422
rect 4103 412 4152 419
rect 4103 406 4133 412
rect 4152 407 4157 412
rect 4069 390 4149 406
rect 4161 398 4197 419
rect 4258 414 4447 438
rect 4492 437 4539 438
rect 4505 432 4539 437
rect 4273 411 4447 414
rect 4266 408 4447 411
rect 4475 431 4539 432
rect 4069 388 4088 390
rect 4103 388 4137 390
rect 4069 372 4149 388
rect 4069 366 4088 372
rect 3785 340 3888 350
rect 3739 338 3888 340
rect 3909 338 3944 350
rect 3578 336 3740 338
rect 3590 316 3609 336
rect 3624 334 3654 336
rect 3473 308 3514 316
rect 3596 312 3609 316
rect 3661 320 3740 336
rect 3772 336 3944 338
rect 3772 320 3851 336
rect 3858 334 3888 336
rect 3436 298 3465 308
rect 3479 298 3508 308
rect 3523 298 3553 312
rect 3596 298 3639 312
rect 3661 308 3851 320
rect 3916 316 3922 336
rect 3646 298 3676 308
rect 3677 298 3835 308
rect 3839 298 3869 308
rect 3873 298 3903 312
rect 3931 298 3944 336
rect 4016 350 4045 366
rect 4059 350 4088 366
rect 4103 356 4133 372
rect 4161 350 4167 398
rect 4170 392 4189 398
rect 4204 392 4234 400
rect 4170 384 4234 392
rect 4170 368 4250 384
rect 4266 377 4328 408
rect 4344 377 4406 408
rect 4475 406 4524 431
rect 4539 406 4569 422
rect 4438 392 4468 400
rect 4475 398 4585 406
rect 4438 384 4483 392
rect 4170 366 4189 368
rect 4204 366 4250 368
rect 4170 350 4250 366
rect 4277 364 4312 377
rect 4353 374 4390 377
rect 4353 372 4395 374
rect 4282 361 4312 364
rect 4291 357 4298 361
rect 4298 356 4299 357
rect 4257 350 4267 356
rect 4016 342 4051 350
rect 4016 316 4017 342
rect 4024 316 4051 342
rect 3959 298 3989 312
rect 4016 308 4051 316
rect 4053 342 4094 350
rect 4053 316 4068 342
rect 4075 316 4094 342
rect 4158 338 4189 350
rect 4204 338 4307 350
rect 4319 340 4345 366
rect 4360 361 4390 372
rect 4422 368 4484 384
rect 4422 366 4468 368
rect 4422 350 4484 366
rect 4496 350 4502 398
rect 4505 390 4585 398
rect 4505 388 4524 390
rect 4539 388 4573 390
rect 4505 372 4585 388
rect 4505 350 4524 372
rect 4539 356 4569 372
rect 4597 366 4603 440
rect 4606 366 4625 510
rect 4640 367 4646 510
rect 4655 441 4668 511
rect 4720 506 4742 511
rect 4713 485 4742 499
rect 4795 485 4811 499
rect 4849 495 4855 497
rect 4862 495 4970 511
rect 4977 495 4983 497
rect 4991 495 5006 511
rect 5072 505 5091 508
rect 4713 483 4811 485
rect 4838 483 5006 495
rect 5021 485 5037 499
rect 5072 486 5094 505
rect 5104 499 5120 500
rect 5103 497 5120 499
rect 5104 492 5120 497
rect 5094 485 5100 486
rect 5103 485 5132 492
rect 5021 484 5132 485
rect 5021 483 5138 484
rect 4697 475 4748 483
rect 4795 475 4829 483
rect 4697 463 4722 475
rect 4729 463 4748 475
rect 4802 473 4829 475
rect 4838 473 5059 483
rect 5094 480 5100 483
rect 4802 469 5059 473
rect 4697 455 4748 463
rect 4795 455 5059 469
rect 5103 475 5138 483
rect 4649 407 4668 441
rect 4713 447 4742 455
rect 4713 441 4730 447
rect 4713 439 4747 441
rect 4795 439 4811 455
rect 4812 445 5020 455
rect 5021 445 5037 455
rect 5085 451 5100 466
rect 5103 463 5104 475
rect 5111 463 5138 475
rect 5103 455 5138 463
rect 5103 454 5132 455
rect 4823 441 5037 445
rect 4838 439 5037 441
rect 5072 441 5085 451
rect 5103 441 5120 454
rect 5072 439 5120 441
rect 4714 435 4747 439
rect 4710 433 4747 435
rect 4710 432 4777 433
rect 4710 427 4741 432
rect 4747 427 4777 432
rect 4710 423 4777 427
rect 4683 420 4777 423
rect 4683 413 4732 420
rect 4683 407 4713 413
rect 4732 408 4737 413
rect 4649 391 4729 407
rect 4741 399 4777 420
rect 4838 415 5027 439
rect 5072 438 5119 439
rect 5085 433 5119 438
rect 4853 412 5027 415
rect 4846 409 5027 412
rect 5055 432 5119 433
rect 4649 389 4668 391
rect 4683 389 4717 391
rect 4649 373 4729 389
rect 4649 367 4668 373
rect 4365 340 4468 350
rect 4319 338 4468 340
rect 4489 338 4524 350
rect 4158 336 4320 338
rect 4170 316 4189 336
rect 4204 334 4234 336
rect 4053 308 4094 316
rect 4176 312 4189 316
rect 4241 320 4320 336
rect 4352 336 4524 338
rect 4352 320 4431 336
rect 4438 334 4468 336
rect 4016 298 4045 308
rect 4059 298 4088 308
rect 4103 298 4133 312
rect 4176 298 4219 312
rect 4241 308 4431 320
rect 4496 316 4502 336
rect 4226 298 4256 308
rect 4257 298 4415 308
rect 4419 298 4449 308
rect 4453 298 4483 312
rect 4511 298 4524 336
rect 4596 350 4625 366
rect 4639 351 4668 367
rect 4683 357 4713 373
rect 4741 351 4747 399
rect 4750 393 4769 399
rect 4784 393 4814 401
rect 4750 385 4814 393
rect 4750 369 4830 385
rect 4846 378 4908 409
rect 4924 378 4986 409
rect 5055 407 5104 432
rect 5119 407 5149 423
rect 5018 393 5048 401
rect 5055 399 5165 407
rect 5018 385 5063 393
rect 4750 367 4769 369
rect 4784 367 4830 369
rect 4750 351 4830 367
rect 4857 365 4892 378
rect 4933 375 4970 378
rect 4933 373 4975 375
rect 4862 362 4892 365
rect 4871 358 4878 362
rect 4878 357 4879 358
rect 4837 351 4847 357
rect 4596 342 4631 350
rect 4596 316 4597 342
rect 4604 316 4631 342
rect 4539 298 4569 312
rect 4596 308 4631 316
rect 4633 343 4674 351
rect 4633 317 4648 343
rect 4655 317 4674 343
rect 4738 339 4769 351
rect 4784 339 4887 351
rect 4899 341 4925 367
rect 4940 362 4970 373
rect 5002 369 5064 385
rect 5002 367 5048 369
rect 5002 351 5064 367
rect 5076 351 5082 399
rect 5085 391 5165 399
rect 5085 389 5104 391
rect 5119 389 5153 391
rect 5085 373 5165 389
rect 5085 351 5104 373
rect 5119 357 5149 373
rect 5177 367 5183 441
rect 5186 367 5205 511
rect 5220 367 5226 511
rect 5235 441 5248 511
rect 5300 506 5322 511
rect 5293 485 5322 499
rect 5375 485 5391 499
rect 5429 495 5435 497
rect 5442 495 5550 511
rect 5557 495 5563 497
rect 5571 495 5586 511
rect 5652 505 5671 508
rect 5293 483 5391 485
rect 5418 483 5586 495
rect 5601 485 5617 499
rect 5652 486 5674 505
rect 5684 499 5700 500
rect 5683 497 5700 499
rect 5684 492 5700 497
rect 5674 485 5680 486
rect 5683 485 5712 492
rect 5601 484 5712 485
rect 5601 483 5718 484
rect 5277 475 5328 483
rect 5375 475 5409 483
rect 5277 463 5302 475
rect 5309 463 5328 475
rect 5382 473 5409 475
rect 5418 473 5639 483
rect 5674 480 5680 483
rect 5382 469 5639 473
rect 5277 455 5328 463
rect 5375 455 5639 469
rect 5683 475 5718 483
rect 5229 407 5248 441
rect 5293 447 5322 455
rect 5293 441 5310 447
rect 5293 439 5327 441
rect 5375 439 5391 455
rect 5392 445 5600 455
rect 5601 445 5617 455
rect 5665 451 5680 466
rect 5683 463 5684 475
rect 5691 463 5718 475
rect 5683 455 5718 463
rect 5683 454 5712 455
rect 5403 441 5617 445
rect 5418 439 5617 441
rect 5652 441 5665 451
rect 5683 441 5700 454
rect 5652 439 5700 441
rect 5294 435 5327 439
rect 5290 433 5327 435
rect 5290 432 5357 433
rect 5290 427 5321 432
rect 5327 427 5357 432
rect 5290 423 5357 427
rect 5263 420 5357 423
rect 5263 413 5312 420
rect 5263 407 5293 413
rect 5312 408 5317 413
rect 5229 391 5309 407
rect 5321 399 5357 420
rect 5418 415 5607 439
rect 5652 438 5699 439
rect 5665 433 5699 438
rect 5433 412 5607 415
rect 5426 409 5607 412
rect 5635 432 5699 433
rect 5229 389 5248 391
rect 5263 389 5297 391
rect 5229 373 5309 389
rect 5229 367 5248 373
rect 4945 341 5048 351
rect 4899 339 5048 341
rect 5069 339 5104 351
rect 4738 337 4900 339
rect 4750 317 4769 337
rect 4784 335 4814 337
rect 4633 309 4674 317
rect 4756 313 4769 317
rect 4821 321 4900 337
rect 4932 337 5104 339
rect 4932 321 5011 337
rect 5018 335 5048 337
rect 4596 299 4625 308
rect 4639 299 4668 309
rect 4683 299 4713 313
rect 4756 299 4799 313
rect 4821 309 5011 321
rect 5076 317 5082 337
rect 4806 299 4836 309
rect 4837 299 4995 309
rect 4999 299 5029 309
rect 5033 299 5063 313
rect 5091 299 5104 337
rect 5176 351 5205 367
rect 5219 351 5248 367
rect 5263 357 5293 373
rect 5321 351 5327 399
rect 5330 393 5349 399
rect 5364 393 5394 401
rect 5330 385 5394 393
rect 5330 369 5410 385
rect 5426 378 5488 409
rect 5504 378 5566 409
rect 5635 407 5684 432
rect 5699 407 5729 423
rect 5598 393 5628 401
rect 5635 399 5745 407
rect 5598 385 5643 393
rect 5330 367 5349 369
rect 5364 367 5410 369
rect 5330 351 5410 367
rect 5437 365 5472 378
rect 5513 375 5550 378
rect 5513 373 5555 375
rect 5442 362 5472 365
rect 5451 358 5458 362
rect 5458 357 5459 358
rect 5417 351 5427 357
rect 5176 343 5211 351
rect 5176 317 5177 343
rect 5184 317 5211 343
rect 5119 299 5149 313
rect 5176 309 5211 317
rect 5213 343 5254 351
rect 5213 317 5228 343
rect 5235 317 5254 343
rect 5318 339 5349 351
rect 5364 339 5467 351
rect 5479 341 5505 367
rect 5520 362 5550 373
rect 5582 369 5644 385
rect 5582 367 5628 369
rect 5582 351 5644 367
rect 5656 351 5662 399
rect 5665 391 5745 399
rect 5665 389 5684 391
rect 5699 389 5733 391
rect 5665 373 5745 389
rect 5665 351 5684 373
rect 5699 357 5729 373
rect 5757 367 5763 441
rect 5766 367 5785 511
rect 5800 367 5806 511
rect 5815 441 5828 511
rect 5880 506 5902 511
rect 5873 485 5902 499
rect 5955 485 5971 499
rect 6009 495 6015 497
rect 6022 495 6130 511
rect 6137 495 6143 497
rect 6151 495 6166 511
rect 6232 505 6251 508
rect 5873 483 5971 485
rect 5998 483 6166 495
rect 6181 485 6197 499
rect 6232 486 6254 505
rect 6264 499 6280 500
rect 6263 497 6280 499
rect 6264 492 6280 497
rect 6254 485 6260 486
rect 6263 485 6292 492
rect 6181 484 6292 485
rect 6181 483 6298 484
rect 5857 475 5908 483
rect 5955 475 5989 483
rect 5857 463 5882 475
rect 5889 463 5908 475
rect 5962 473 5989 475
rect 5998 473 6219 483
rect 6254 480 6260 483
rect 5962 469 6219 473
rect 5857 455 5908 463
rect 5955 455 6219 469
rect 6263 475 6298 483
rect 5809 407 5828 441
rect 5873 447 5902 455
rect 5873 441 5890 447
rect 5873 439 5907 441
rect 5955 439 5971 455
rect 5972 445 6180 455
rect 6181 445 6197 455
rect 6245 451 6260 466
rect 6263 463 6264 475
rect 6271 463 6298 475
rect 6263 455 6298 463
rect 6263 454 6292 455
rect 5983 441 6197 445
rect 5998 439 6197 441
rect 6232 441 6245 451
rect 6263 441 6280 454
rect 6232 439 6280 441
rect 5874 435 5907 439
rect 5870 433 5907 435
rect 5870 432 5937 433
rect 5870 427 5901 432
rect 5907 427 5937 432
rect 5870 423 5937 427
rect 5843 420 5937 423
rect 5843 413 5892 420
rect 5843 407 5873 413
rect 5892 408 5897 413
rect 5809 391 5889 407
rect 5901 399 5937 420
rect 5998 415 6187 439
rect 6232 438 6279 439
rect 6245 433 6279 438
rect 6013 412 6187 415
rect 6006 409 6187 412
rect 6215 432 6279 433
rect 5809 389 5828 391
rect 5843 389 5877 391
rect 5809 373 5889 389
rect 5809 367 5828 373
rect 5525 341 5628 351
rect 5479 339 5628 341
rect 5649 339 5684 351
rect 5318 337 5480 339
rect 5330 317 5349 337
rect 5364 335 5394 337
rect 5213 309 5254 317
rect 5336 313 5349 317
rect 5401 321 5480 337
rect 5512 337 5684 339
rect 5512 321 5591 337
rect 5598 335 5628 337
rect 5176 299 5205 309
rect 5219 299 5248 309
rect 5263 299 5293 313
rect 5336 299 5379 313
rect 5401 309 5591 321
rect 5656 317 5662 337
rect 5386 299 5416 309
rect 5417 299 5575 309
rect 5579 299 5609 309
rect 5613 299 5643 313
rect 5671 299 5684 337
rect 5756 351 5785 367
rect 5799 351 5828 367
rect 5843 357 5873 373
rect 5901 351 5907 399
rect 5910 393 5929 399
rect 5944 393 5974 401
rect 5910 385 5974 393
rect 5910 369 5990 385
rect 6006 378 6068 409
rect 6084 378 6146 409
rect 6215 407 6264 432
rect 6279 407 6309 423
rect 6178 393 6208 401
rect 6215 399 6325 407
rect 6178 385 6223 393
rect 5910 367 5929 369
rect 5944 367 5990 369
rect 5910 351 5990 367
rect 6017 365 6052 378
rect 6093 375 6130 378
rect 6093 373 6135 375
rect 6022 362 6052 365
rect 6031 358 6038 362
rect 6038 357 6039 358
rect 5997 351 6007 357
rect 5756 343 5791 351
rect 5756 317 5757 343
rect 5764 317 5791 343
rect 5699 299 5729 313
rect 5756 309 5791 317
rect 5793 343 5834 351
rect 5793 317 5808 343
rect 5815 317 5834 343
rect 5898 339 5929 351
rect 5944 339 6047 351
rect 6059 341 6085 367
rect 6100 362 6130 373
rect 6162 369 6224 385
rect 6162 367 6208 369
rect 6162 351 6224 367
rect 6236 351 6242 399
rect 6245 391 6325 399
rect 6245 389 6264 391
rect 6279 389 6313 391
rect 6245 373 6325 389
rect 6245 351 6264 373
rect 6279 357 6309 373
rect 6337 367 6343 441
rect 6346 367 6365 511
rect 6380 367 6386 511
rect 6395 441 6408 511
rect 6460 506 6482 511
rect 6453 485 6482 499
rect 6535 485 6551 499
rect 6589 495 6595 497
rect 6602 495 6710 511
rect 6717 495 6723 497
rect 6731 495 6746 511
rect 6812 505 6831 508
rect 6453 483 6551 485
rect 6578 483 6746 495
rect 6761 485 6777 499
rect 6812 486 6834 505
rect 6844 499 6860 500
rect 6843 497 6860 499
rect 6844 492 6860 497
rect 6834 485 6840 486
rect 6843 485 6872 492
rect 6761 484 6872 485
rect 6761 483 6878 484
rect 6437 475 6488 483
rect 6535 475 6569 483
rect 6437 463 6462 475
rect 6469 463 6488 475
rect 6542 473 6569 475
rect 6578 473 6799 483
rect 6834 480 6840 483
rect 6542 469 6799 473
rect 6437 455 6488 463
rect 6535 455 6799 469
rect 6843 475 6878 483
rect 6389 407 6408 441
rect 6453 447 6482 455
rect 6453 441 6470 447
rect 6453 439 6487 441
rect 6535 439 6551 455
rect 6552 445 6760 455
rect 6761 445 6777 455
rect 6825 451 6840 466
rect 6843 463 6844 475
rect 6851 463 6878 475
rect 6843 455 6878 463
rect 6843 454 6872 455
rect 6563 441 6777 445
rect 6578 439 6777 441
rect 6812 441 6825 451
rect 6843 441 6860 454
rect 6812 439 6860 441
rect 6454 435 6487 439
rect 6450 433 6487 435
rect 6450 432 6517 433
rect 6450 427 6481 432
rect 6487 427 6517 432
rect 6450 423 6517 427
rect 6423 420 6517 423
rect 6423 413 6472 420
rect 6423 407 6453 413
rect 6472 408 6477 413
rect 6389 391 6469 407
rect 6481 399 6517 420
rect 6578 415 6767 439
rect 6812 438 6859 439
rect 6825 433 6859 438
rect 6593 412 6767 415
rect 6586 409 6767 412
rect 6795 432 6859 433
rect 6389 389 6408 391
rect 6423 389 6457 391
rect 6389 373 6469 389
rect 6389 367 6408 373
rect 6105 341 6208 351
rect 6059 339 6208 341
rect 6229 339 6264 351
rect 5898 337 6060 339
rect 5910 317 5929 337
rect 5944 335 5974 337
rect 5793 309 5834 317
rect 5916 313 5929 317
rect 5981 321 6060 337
rect 6092 337 6264 339
rect 6092 321 6171 337
rect 6178 335 6208 337
rect 5756 299 5785 309
rect 5799 299 5828 309
rect 5843 299 5873 313
rect 5916 299 5959 313
rect 5981 309 6171 321
rect 6236 317 6242 337
rect 5966 299 5996 309
rect 5997 299 6155 309
rect 6159 299 6189 309
rect 6193 299 6223 313
rect 6251 299 6264 337
rect 6336 351 6365 367
rect 6379 351 6408 367
rect 6423 357 6453 373
rect 6481 351 6487 399
rect 6490 393 6509 399
rect 6524 393 6554 401
rect 6490 385 6554 393
rect 6490 369 6570 385
rect 6586 378 6648 409
rect 6664 378 6726 409
rect 6795 407 6844 432
rect 6859 407 6889 423
rect 6758 393 6788 401
rect 6795 399 6905 407
rect 6758 385 6803 393
rect 6490 367 6509 369
rect 6524 367 6570 369
rect 6490 351 6570 367
rect 6597 365 6632 378
rect 6673 375 6710 378
rect 6673 373 6715 375
rect 6602 362 6632 365
rect 6611 358 6618 362
rect 6618 357 6619 358
rect 6577 351 6587 357
rect 6336 343 6371 351
rect 6336 317 6337 343
rect 6344 317 6371 343
rect 6279 299 6309 313
rect 6336 309 6371 317
rect 6373 343 6414 351
rect 6373 317 6388 343
rect 6395 317 6414 343
rect 6478 339 6509 351
rect 6524 339 6627 351
rect 6639 341 6665 367
rect 6680 362 6710 373
rect 6742 369 6804 385
rect 6742 367 6788 369
rect 6742 351 6804 367
rect 6816 351 6822 399
rect 6825 391 6905 399
rect 6825 389 6844 391
rect 6859 389 6893 391
rect 6825 373 6905 389
rect 6825 351 6844 373
rect 6859 357 6889 373
rect 6917 367 6923 441
rect 6926 367 6945 511
rect 6960 367 6966 511
rect 6975 441 6988 511
rect 7040 506 7062 511
rect 7033 485 7062 499
rect 7115 485 7131 499
rect 7169 495 7175 497
rect 7182 495 7290 511
rect 7297 495 7303 497
rect 7311 495 7326 511
rect 7392 505 7411 508
rect 7033 483 7131 485
rect 7158 483 7326 495
rect 7341 485 7357 499
rect 7392 486 7414 505
rect 7424 499 7440 500
rect 7423 497 7440 499
rect 7424 492 7440 497
rect 7414 485 7420 486
rect 7423 485 7452 492
rect 7341 484 7452 485
rect 7341 483 7458 484
rect 7017 475 7068 483
rect 7115 475 7149 483
rect 7017 463 7042 475
rect 7049 463 7068 475
rect 7122 473 7149 475
rect 7158 473 7379 483
rect 7414 480 7420 483
rect 7122 469 7379 473
rect 7017 455 7068 463
rect 7115 455 7379 469
rect 7423 475 7458 483
rect 6969 407 6988 441
rect 7033 447 7062 455
rect 7033 441 7050 447
rect 7033 439 7067 441
rect 7115 439 7131 455
rect 7132 445 7340 455
rect 7341 445 7357 455
rect 7405 451 7420 466
rect 7423 463 7424 475
rect 7431 463 7458 475
rect 7423 455 7458 463
rect 7423 454 7452 455
rect 7151 441 7357 445
rect 7158 439 7357 441
rect 7392 441 7405 451
rect 7423 441 7440 454
rect 7392 439 7440 441
rect 7034 435 7067 439
rect 7030 433 7067 435
rect 7030 432 7097 433
rect 7030 427 7061 432
rect 7067 427 7097 432
rect 7030 423 7097 427
rect 7003 420 7097 423
rect 7003 413 7052 420
rect 7003 407 7033 413
rect 7052 408 7057 413
rect 6969 391 7049 407
rect 7061 399 7097 420
rect 7158 415 7347 439
rect 7392 438 7439 439
rect 7405 433 7439 438
rect 7173 412 7347 415
rect 7166 409 7347 412
rect 7375 432 7439 433
rect 6969 389 6988 391
rect 7003 389 7037 391
rect 6969 373 7049 389
rect 6969 367 6988 373
rect 6685 341 6788 351
rect 6639 339 6788 341
rect 6809 339 6844 351
rect 6478 337 6640 339
rect 6490 317 6509 337
rect 6524 335 6554 337
rect 6373 309 6414 317
rect 6496 313 6509 317
rect 6561 321 6640 337
rect 6672 337 6844 339
rect 6672 321 6751 337
rect 6758 335 6788 337
rect 6336 299 6365 309
rect 6379 299 6408 309
rect 6423 299 6453 313
rect 6496 299 6539 313
rect 6561 309 6751 321
rect 6816 317 6822 337
rect 6546 299 6576 309
rect 6577 299 6735 309
rect 6739 299 6769 309
rect 6773 299 6803 313
rect 6831 299 6844 337
rect 6916 351 6945 367
rect 6959 351 6988 367
rect 7003 357 7033 373
rect 7061 351 7067 399
rect 7070 393 7089 399
rect 7104 393 7134 401
rect 7070 385 7134 393
rect 7070 369 7150 385
rect 7166 378 7228 409
rect 7244 378 7306 409
rect 7375 407 7424 432
rect 7439 407 7469 423
rect 7338 393 7368 401
rect 7375 399 7485 407
rect 7338 385 7383 393
rect 7070 367 7089 369
rect 7104 367 7150 369
rect 7070 351 7150 367
rect 7177 365 7212 378
rect 7253 375 7290 378
rect 7253 373 7295 375
rect 7182 362 7212 365
rect 7191 358 7198 362
rect 7198 357 7199 358
rect 7157 351 7167 357
rect 6916 343 6951 351
rect 6916 317 6917 343
rect 6924 317 6951 343
rect 6859 299 6889 313
rect 6916 309 6951 317
rect 6953 343 6994 351
rect 6953 317 6968 343
rect 6975 317 6994 343
rect 7058 339 7089 351
rect 7104 339 7207 351
rect 7219 341 7245 367
rect 7260 362 7290 373
rect 7322 369 7384 385
rect 7322 367 7368 369
rect 7322 351 7384 367
rect 7396 351 7402 399
rect 7405 391 7485 399
rect 7405 389 7424 391
rect 7439 389 7473 391
rect 7405 373 7485 389
rect 7405 351 7424 373
rect 7439 357 7469 373
rect 7497 367 7503 441
rect 7506 367 7525 511
rect 7540 367 7546 511
rect 7555 441 7568 511
rect 7620 506 7642 511
rect 7613 485 7642 499
rect 7695 485 7711 499
rect 7749 495 7755 497
rect 7762 495 7870 511
rect 7877 495 7883 497
rect 7891 495 7906 511
rect 7972 505 7991 508
rect 7613 483 7711 485
rect 7738 483 7906 495
rect 7921 485 7937 499
rect 7972 486 7994 505
rect 8004 499 8020 500
rect 8003 497 8020 499
rect 8004 492 8020 497
rect 7994 485 8000 486
rect 8003 485 8032 492
rect 7921 484 8032 485
rect 7921 483 8038 484
rect 7597 475 7648 483
rect 7695 475 7729 483
rect 7597 463 7622 475
rect 7629 463 7648 475
rect 7702 473 7729 475
rect 7738 473 7959 483
rect 7994 480 8000 483
rect 7702 469 7959 473
rect 7597 455 7648 463
rect 7695 455 7959 469
rect 8003 475 8038 483
rect 7549 407 7568 441
rect 7613 447 7642 455
rect 7613 441 7630 447
rect 7613 439 7647 441
rect 7695 439 7711 455
rect 7712 445 7920 455
rect 7921 445 7937 455
rect 7985 451 8000 466
rect 8003 463 8004 475
rect 8011 463 8038 475
rect 8003 455 8038 463
rect 8003 454 8032 455
rect 7723 441 7937 445
rect 7738 439 7937 441
rect 7972 441 7985 451
rect 8003 441 8020 454
rect 7972 439 8020 441
rect 7614 435 7647 439
rect 7610 433 7647 435
rect 7610 432 7677 433
rect 7610 427 7641 432
rect 7647 427 7677 432
rect 7610 423 7677 427
rect 7583 420 7677 423
rect 7583 413 7632 420
rect 7583 407 7613 413
rect 7632 408 7637 413
rect 7549 391 7629 407
rect 7641 399 7677 420
rect 7738 415 7927 439
rect 7972 438 8019 439
rect 7985 433 8019 438
rect 7753 412 7927 415
rect 7746 409 7927 412
rect 7955 432 8019 433
rect 7549 389 7568 391
rect 7583 389 7617 391
rect 7549 373 7629 389
rect 7549 367 7568 373
rect 7265 341 7368 351
rect 7219 339 7368 341
rect 7389 339 7424 351
rect 7058 337 7220 339
rect 7070 317 7089 337
rect 7104 335 7134 337
rect 6953 309 6994 317
rect 7076 313 7089 317
rect 7141 321 7220 337
rect 7252 337 7424 339
rect 7252 321 7331 337
rect 7338 335 7368 337
rect 6916 299 6945 309
rect 6959 299 6988 309
rect 7003 299 7033 313
rect 7076 299 7119 313
rect 7141 309 7331 321
rect 7396 317 7402 337
rect 7126 299 7156 309
rect 7157 299 7315 309
rect 7319 299 7349 309
rect 7353 299 7383 313
rect 7411 299 7424 337
rect 7496 351 7525 367
rect 7539 351 7568 367
rect 7583 357 7613 373
rect 7641 351 7647 399
rect 7650 393 7669 399
rect 7684 393 7714 401
rect 7650 385 7714 393
rect 7650 369 7730 385
rect 7746 378 7808 409
rect 7824 378 7886 409
rect 7955 407 8004 432
rect 8019 407 8049 423
rect 7918 393 7948 401
rect 7955 399 8065 407
rect 7918 385 7963 393
rect 7650 367 7669 369
rect 7684 367 7730 369
rect 7650 351 7730 367
rect 7757 365 7792 378
rect 7833 375 7870 378
rect 7833 373 7875 375
rect 7762 362 7792 365
rect 7771 358 7778 362
rect 7778 357 7779 358
rect 7737 351 7747 357
rect 7496 343 7531 351
rect 7496 317 7497 343
rect 7504 317 7531 343
rect 7439 299 7469 313
rect 7496 309 7531 317
rect 7533 343 7574 351
rect 7533 317 7548 343
rect 7555 317 7574 343
rect 7638 339 7669 351
rect 7684 339 7787 351
rect 7799 341 7825 367
rect 7840 362 7870 373
rect 7902 369 7964 385
rect 7902 367 7948 369
rect 7902 351 7964 367
rect 7976 351 7982 399
rect 7985 391 8065 399
rect 7985 389 8004 391
rect 8019 389 8053 391
rect 7985 373 8065 389
rect 7985 351 8004 373
rect 8019 357 8049 373
rect 8077 367 8083 441
rect 8086 367 8105 511
rect 8120 367 8126 511
rect 8135 441 8148 511
rect 8200 506 8222 511
rect 8193 485 8222 499
rect 8275 485 8291 499
rect 8329 495 8335 497
rect 8342 495 8450 511
rect 8457 495 8463 497
rect 8471 495 8486 511
rect 8552 505 8571 508
rect 8193 483 8291 485
rect 8318 483 8486 495
rect 8501 485 8517 499
rect 8552 486 8574 505
rect 8584 499 8600 500
rect 8583 497 8600 499
rect 8584 492 8600 497
rect 8574 485 8580 486
rect 8583 485 8612 492
rect 8501 484 8612 485
rect 8501 483 8618 484
rect 8177 475 8228 483
rect 8275 475 8309 483
rect 8177 463 8202 475
rect 8209 463 8228 475
rect 8282 473 8309 475
rect 8318 473 8539 483
rect 8574 480 8580 483
rect 8282 469 8539 473
rect 8177 455 8228 463
rect 8275 455 8539 469
rect 8583 475 8618 483
rect 8129 407 8148 441
rect 8193 447 8222 455
rect 8193 441 8210 447
rect 8193 439 8227 441
rect 8275 439 8291 455
rect 8292 445 8500 455
rect 8501 445 8517 455
rect 8565 451 8580 466
rect 8583 463 8584 475
rect 8591 463 8618 475
rect 8583 455 8618 463
rect 8583 454 8612 455
rect 8303 441 8517 445
rect 8318 439 8517 441
rect 8552 441 8565 451
rect 8583 441 8600 454
rect 8552 439 8600 441
rect 8194 435 8227 439
rect 8190 433 8227 435
rect 8190 432 8257 433
rect 8190 427 8221 432
rect 8227 427 8257 432
rect 8190 423 8257 427
rect 8163 420 8257 423
rect 8163 413 8212 420
rect 8163 407 8193 413
rect 8212 408 8217 413
rect 8129 391 8209 407
rect 8221 399 8257 420
rect 8318 415 8507 439
rect 8552 438 8599 439
rect 8565 433 8599 438
rect 8333 412 8507 415
rect 8326 409 8507 412
rect 8535 432 8599 433
rect 8129 389 8148 391
rect 8163 389 8197 391
rect 8129 373 8209 389
rect 8129 367 8148 373
rect 7845 341 7948 351
rect 7799 339 7948 341
rect 7969 339 8004 351
rect 7638 337 7800 339
rect 7650 317 7669 337
rect 7684 335 7714 337
rect 7533 309 7574 317
rect 7656 313 7669 317
rect 7721 321 7800 337
rect 7832 337 8004 339
rect 7832 321 7911 337
rect 7918 335 7948 337
rect 7496 299 7525 309
rect 7539 299 7568 309
rect 7583 299 7613 313
rect 7656 299 7699 313
rect 7721 309 7911 321
rect 7976 317 7982 337
rect 7706 299 7736 309
rect 7737 299 7895 309
rect 7899 299 7929 309
rect 7933 299 7963 313
rect 7991 299 8004 337
rect 8076 351 8105 367
rect 8119 351 8148 367
rect 8163 357 8193 373
rect 8221 351 8227 399
rect 8230 393 8249 399
rect 8264 393 8294 401
rect 8230 385 8294 393
rect 8230 369 8310 385
rect 8326 378 8388 409
rect 8404 378 8466 409
rect 8535 407 8584 432
rect 8599 407 8629 423
rect 8498 393 8528 401
rect 8535 399 8645 407
rect 8498 385 8543 393
rect 8230 367 8249 369
rect 8264 367 8310 369
rect 8230 351 8310 367
rect 8337 365 8372 378
rect 8413 375 8450 378
rect 8413 373 8455 375
rect 8342 362 8372 365
rect 8351 358 8358 362
rect 8358 357 8359 358
rect 8317 351 8327 357
rect 8076 343 8111 351
rect 8076 317 8077 343
rect 8084 317 8111 343
rect 8019 299 8049 313
rect 8076 309 8111 317
rect 8113 343 8154 351
rect 8113 317 8128 343
rect 8135 317 8154 343
rect 8218 339 8249 351
rect 8264 339 8367 351
rect 8379 341 8405 367
rect 8420 362 8450 373
rect 8482 369 8544 385
rect 8482 367 8528 369
rect 8482 351 8544 367
rect 8556 351 8562 399
rect 8565 391 8645 399
rect 8565 389 8584 391
rect 8599 389 8633 391
rect 8565 373 8645 389
rect 8565 351 8584 373
rect 8599 357 8629 373
rect 8657 367 8663 441
rect 8666 367 8685 511
rect 8700 367 8706 511
rect 8715 441 8728 511
rect 8780 506 8802 511
rect 8773 485 8802 499
rect 8855 485 8871 499
rect 8909 495 8915 497
rect 8922 495 9030 511
rect 9037 495 9043 497
rect 9051 495 9066 511
rect 9132 505 9151 508
rect 8773 483 8871 485
rect 8898 483 9066 495
rect 9081 485 9097 499
rect 9132 486 9154 505
rect 9164 499 9180 500
rect 9163 497 9180 499
rect 9164 492 9180 497
rect 9154 485 9160 486
rect 9163 485 9192 492
rect 9081 484 9192 485
rect 9081 483 9198 484
rect 8757 475 8808 483
rect 8855 475 8889 483
rect 8757 463 8782 475
rect 8789 463 8808 475
rect 8862 473 8889 475
rect 8898 473 9119 483
rect 9154 480 9160 483
rect 8862 469 9119 473
rect 8757 455 8808 463
rect 8855 455 9119 469
rect 9163 475 9198 483
rect 8709 407 8728 441
rect 8773 447 8802 455
rect 8773 441 8790 447
rect 8773 439 8807 441
rect 8855 439 8871 455
rect 8872 445 9080 455
rect 9081 445 9097 455
rect 9145 451 9160 466
rect 9163 463 9164 475
rect 9171 463 9198 475
rect 9163 455 9198 463
rect 9163 454 9192 455
rect 8883 441 9097 445
rect 8898 439 9097 441
rect 9132 441 9145 451
rect 9163 441 9180 454
rect 9132 439 9180 441
rect 8774 435 8807 439
rect 8770 433 8807 435
rect 8770 432 8837 433
rect 8770 427 8801 432
rect 8807 427 8837 432
rect 8770 423 8837 427
rect 8743 420 8837 423
rect 8743 413 8792 420
rect 8743 407 8773 413
rect 8792 408 8797 413
rect 8709 391 8789 407
rect 8801 399 8837 420
rect 8898 415 9087 439
rect 9132 438 9179 439
rect 9145 433 9179 438
rect 8913 412 9087 415
rect 8906 409 9087 412
rect 9115 432 9179 433
rect 8709 389 8728 391
rect 8743 389 8777 391
rect 8709 373 8789 389
rect 8709 367 8728 373
rect 8425 341 8528 351
rect 8379 339 8528 341
rect 8549 339 8584 351
rect 8218 337 8380 339
rect 8230 317 8249 337
rect 8264 335 8294 337
rect 8113 309 8154 317
rect 8236 313 8249 317
rect 8301 321 8380 337
rect 8412 337 8584 339
rect 8412 321 8491 337
rect 8498 335 8528 337
rect 8076 299 8105 309
rect 8119 299 8148 309
rect 8163 299 8193 313
rect 8236 299 8279 313
rect 8301 309 8491 321
rect 8556 317 8562 337
rect 8286 299 8316 309
rect 8317 299 8475 309
rect 8479 299 8509 309
rect 8513 299 8543 313
rect 8571 299 8584 337
rect 8656 351 8685 367
rect 8699 351 8728 367
rect 8743 357 8773 373
rect 8801 351 8807 399
rect 8810 393 8829 399
rect 8844 393 8874 401
rect 8810 385 8874 393
rect 8810 369 8890 385
rect 8906 378 8968 409
rect 8984 378 9046 409
rect 9115 407 9164 432
rect 9179 407 9209 423
rect 9078 393 9108 401
rect 9115 399 9225 407
rect 9078 385 9123 393
rect 8810 367 8829 369
rect 8844 367 8890 369
rect 8810 351 8890 367
rect 8917 365 8952 378
rect 8993 375 9030 378
rect 8993 373 9035 375
rect 8922 362 8952 365
rect 8931 358 8938 362
rect 8938 357 8939 358
rect 8897 351 8907 357
rect 8656 343 8691 351
rect 8656 317 8657 343
rect 8664 317 8691 343
rect 8599 299 8629 313
rect 8656 309 8691 317
rect 8693 343 8734 351
rect 8693 317 8708 343
rect 8715 317 8734 343
rect 8798 339 8829 351
rect 8844 339 8947 351
rect 8959 341 8985 367
rect 9000 362 9030 373
rect 9062 369 9124 385
rect 9062 367 9108 369
rect 9062 351 9124 367
rect 9136 351 9142 399
rect 9145 391 9225 399
rect 9145 389 9164 391
rect 9179 389 9213 391
rect 9145 373 9225 389
rect 9145 351 9164 373
rect 9179 357 9209 373
rect 9237 367 9243 441
rect 9246 367 9265 511
rect 9280 367 9286 511
rect 9295 441 9308 511
rect 9360 506 9382 511
rect 9353 485 9382 499
rect 9435 485 9451 499
rect 9489 495 9495 497
rect 9502 495 9610 511
rect 9617 495 9623 497
rect 9631 495 9646 511
rect 9712 505 9731 508
rect 9353 483 9451 485
rect 9478 483 9646 495
rect 9661 485 9677 499
rect 9712 486 9734 505
rect 9744 499 9760 500
rect 9743 497 9760 499
rect 9744 492 9760 497
rect 9734 485 9740 486
rect 9743 485 9772 492
rect 9661 484 9772 485
rect 9661 483 9778 484
rect 9337 475 9388 483
rect 9435 475 9469 483
rect 9337 463 9362 475
rect 9369 463 9388 475
rect 9442 473 9469 475
rect 9478 473 9699 483
rect 9734 480 9740 483
rect 9442 469 9699 473
rect 9337 455 9388 463
rect 9435 455 9699 469
rect 9743 475 9778 483
rect 9289 407 9308 441
rect 9353 447 9382 455
rect 9353 441 9370 447
rect 9353 439 9387 441
rect 9435 439 9451 455
rect 9452 445 9660 455
rect 9661 445 9677 455
rect 9725 451 9740 466
rect 9743 463 9744 475
rect 9751 463 9778 475
rect 9743 455 9778 463
rect 9743 454 9772 455
rect 9463 441 9677 445
rect 9478 439 9677 441
rect 9712 441 9725 451
rect 9743 441 9760 454
rect 9712 439 9760 441
rect 9354 435 9387 439
rect 9350 433 9387 435
rect 9350 432 9417 433
rect 9350 427 9381 432
rect 9387 427 9417 432
rect 9350 423 9417 427
rect 9323 420 9417 423
rect 9323 413 9372 420
rect 9323 407 9353 413
rect 9372 408 9377 413
rect 9289 391 9369 407
rect 9381 399 9417 420
rect 9478 415 9667 439
rect 9712 438 9759 439
rect 9725 433 9759 438
rect 9493 412 9667 415
rect 9486 409 9667 412
rect 9695 432 9759 433
rect 9289 389 9308 391
rect 9323 389 9357 391
rect 9289 373 9369 389
rect 9289 367 9308 373
rect 9005 341 9108 351
rect 8959 339 9108 341
rect 9129 339 9164 351
rect 8798 337 8960 339
rect 8810 317 8829 337
rect 8844 335 8874 337
rect 8693 309 8734 317
rect 8816 313 8829 317
rect 8881 321 8960 337
rect 8992 337 9164 339
rect 8992 321 9071 337
rect 9078 335 9108 337
rect 8656 299 8685 309
rect 8699 299 8728 309
rect 8743 299 8773 313
rect 8816 299 8859 313
rect 8881 309 9071 321
rect 9136 317 9142 337
rect 8866 299 8896 309
rect 8897 299 9055 309
rect 9059 299 9089 309
rect 9093 299 9123 313
rect 9151 299 9164 337
rect 9236 351 9265 367
rect 9279 351 9308 367
rect 9323 357 9353 373
rect 9381 351 9387 399
rect 9390 393 9409 399
rect 9424 393 9454 401
rect 9390 385 9454 393
rect 9390 369 9470 385
rect 9486 378 9548 409
rect 9564 378 9626 409
rect 9695 407 9744 432
rect 9759 407 9789 423
rect 9658 393 9688 401
rect 9695 399 9805 407
rect 9658 385 9703 393
rect 9390 367 9409 369
rect 9424 367 9470 369
rect 9390 351 9470 367
rect 9497 365 9532 378
rect 9573 375 9610 378
rect 9573 373 9615 375
rect 9502 362 9532 365
rect 9511 358 9518 362
rect 9518 357 9519 358
rect 9477 351 9487 357
rect 9236 343 9271 351
rect 9236 317 9237 343
rect 9244 317 9271 343
rect 9179 299 9209 313
rect 9236 309 9271 317
rect 9273 343 9314 351
rect 9273 317 9288 343
rect 9295 317 9314 343
rect 9378 339 9409 351
rect 9424 339 9527 351
rect 9539 341 9565 367
rect 9580 362 9610 373
rect 9642 369 9704 385
rect 9642 367 9688 369
rect 9642 351 9704 367
rect 9716 351 9722 399
rect 9725 391 9805 399
rect 9725 389 9744 391
rect 9759 389 9793 391
rect 9725 373 9805 389
rect 9725 351 9744 373
rect 9759 357 9789 373
rect 9817 367 9823 441
rect 9826 367 9845 511
rect 9860 367 9866 511
rect 9875 441 9888 511
rect 9940 506 9962 511
rect 9933 485 9962 499
rect 10015 485 10031 499
rect 10069 495 10075 497
rect 10082 495 10190 511
rect 10197 495 10203 497
rect 10211 495 10226 511
rect 10292 505 10311 508
rect 9933 483 10031 485
rect 10058 483 10226 495
rect 10241 485 10257 499
rect 10292 486 10314 505
rect 10324 499 10340 500
rect 10323 497 10340 499
rect 10324 492 10340 497
rect 10314 485 10320 486
rect 10323 485 10352 492
rect 10241 484 10352 485
rect 10241 483 10358 484
rect 9917 475 9968 483
rect 10015 475 10049 483
rect 9917 463 9942 475
rect 9949 463 9968 475
rect 10022 473 10049 475
rect 10058 473 10279 483
rect 10314 480 10320 483
rect 10022 469 10279 473
rect 9917 455 9968 463
rect 10015 455 10279 469
rect 10323 475 10358 483
rect 9869 407 9888 441
rect 9933 447 9962 455
rect 9933 441 9950 447
rect 9933 439 9967 441
rect 10015 439 10031 455
rect 10032 445 10240 455
rect 10241 445 10257 455
rect 10305 451 10320 466
rect 10323 463 10324 475
rect 10331 463 10358 475
rect 10323 455 10358 463
rect 10323 454 10352 455
rect 10043 441 10257 445
rect 10058 439 10257 441
rect 10292 441 10305 451
rect 10323 441 10340 454
rect 10292 439 10340 441
rect 9934 435 9967 439
rect 9930 433 9967 435
rect 9930 432 9997 433
rect 9930 427 9961 432
rect 9967 427 9997 432
rect 9930 423 9997 427
rect 9903 420 9997 423
rect 9903 413 9952 420
rect 9903 407 9933 413
rect 9952 408 9957 413
rect 9869 391 9949 407
rect 9961 399 9997 420
rect 10058 415 10247 439
rect 10292 438 10339 439
rect 10305 433 10339 438
rect 10073 412 10247 415
rect 10066 409 10247 412
rect 10275 432 10339 433
rect 9869 389 9888 391
rect 9903 389 9937 391
rect 9869 373 9949 389
rect 9869 367 9888 373
rect 9585 341 9688 351
rect 9539 339 9688 341
rect 9709 339 9744 351
rect 9378 337 9540 339
rect 9390 317 9409 337
rect 9424 335 9454 337
rect 9273 309 9314 317
rect 9396 313 9409 317
rect 9461 321 9540 337
rect 9572 337 9744 339
rect 9572 321 9651 337
rect 9658 335 9688 337
rect 9236 299 9265 309
rect 9279 299 9308 309
rect 9323 299 9353 313
rect 9396 299 9439 313
rect 9461 309 9651 321
rect 9716 317 9722 337
rect 9446 299 9476 309
rect 9477 299 9635 309
rect 9639 299 9669 309
rect 9673 299 9703 313
rect 9731 299 9744 337
rect 9816 351 9845 367
rect 9859 351 9888 367
rect 9903 357 9933 373
rect 9961 351 9967 399
rect 9970 393 9989 399
rect 10004 393 10034 401
rect 9970 385 10034 393
rect 9970 369 10050 385
rect 10066 378 10128 409
rect 10144 378 10206 409
rect 10275 407 10324 432
rect 10339 407 10369 423
rect 10238 393 10268 401
rect 10275 399 10385 407
rect 10238 385 10283 393
rect 9970 367 9989 369
rect 10004 367 10050 369
rect 9970 351 10050 367
rect 10077 365 10112 378
rect 10153 375 10190 378
rect 10153 373 10195 375
rect 10082 362 10112 365
rect 10091 358 10098 362
rect 10098 357 10099 358
rect 10057 351 10067 357
rect 9816 343 9851 351
rect 9816 317 9817 343
rect 9824 317 9851 343
rect 9759 299 9789 313
rect 9816 309 9851 317
rect 9853 343 9894 351
rect 9853 317 9868 343
rect 9875 317 9894 343
rect 9958 339 9989 351
rect 10004 339 10107 351
rect 10119 341 10145 367
rect 10160 362 10190 373
rect 10222 369 10284 385
rect 10222 367 10268 369
rect 10222 351 10284 367
rect 10296 351 10302 399
rect 10305 391 10385 399
rect 10305 389 10324 391
rect 10339 389 10373 391
rect 10305 373 10385 389
rect 10305 351 10324 373
rect 10339 357 10369 373
rect 10397 367 10403 441
rect 10406 367 10425 511
rect 10440 367 10446 511
rect 10455 441 10468 511
rect 10520 506 10542 511
rect 10513 485 10542 499
rect 10595 485 10611 499
rect 10649 495 10655 497
rect 10662 495 10770 511
rect 10777 495 10783 497
rect 10791 495 10806 511
rect 10872 505 10891 508
rect 10513 483 10611 485
rect 10638 483 10806 495
rect 10821 485 10837 499
rect 10872 486 10894 505
rect 10904 499 10920 500
rect 10903 497 10920 499
rect 10904 492 10920 497
rect 10894 485 10900 486
rect 10903 485 10932 492
rect 10821 484 10932 485
rect 10821 483 10938 484
rect 10497 475 10548 483
rect 10595 475 10629 483
rect 10497 463 10522 475
rect 10529 463 10548 475
rect 10602 473 10629 475
rect 10638 473 10859 483
rect 10894 480 10900 483
rect 10602 469 10859 473
rect 10497 455 10548 463
rect 10595 455 10859 469
rect 10903 475 10938 483
rect 10449 407 10468 441
rect 10513 447 10542 455
rect 10513 441 10530 447
rect 10513 439 10547 441
rect 10595 439 10611 455
rect 10612 445 10820 455
rect 10821 445 10837 455
rect 10885 451 10900 466
rect 10903 463 10904 475
rect 10911 463 10938 475
rect 10903 455 10938 463
rect 10903 454 10932 455
rect 10623 441 10837 445
rect 10638 439 10837 441
rect 10872 441 10885 451
rect 10903 441 10920 454
rect 10872 439 10920 441
rect 10514 435 10547 439
rect 10510 433 10547 435
rect 10510 432 10577 433
rect 10510 427 10541 432
rect 10547 427 10577 432
rect 10510 423 10577 427
rect 10483 420 10577 423
rect 10483 413 10532 420
rect 10483 407 10513 413
rect 10532 408 10537 413
rect 10449 391 10529 407
rect 10541 399 10577 420
rect 10638 415 10827 439
rect 10872 438 10919 439
rect 10885 433 10919 438
rect 10653 412 10827 415
rect 10646 409 10827 412
rect 10855 432 10919 433
rect 10449 389 10468 391
rect 10483 389 10517 391
rect 10449 373 10529 389
rect 10449 367 10468 373
rect 10165 341 10268 351
rect 10119 339 10268 341
rect 10289 339 10324 351
rect 9958 337 10120 339
rect 9970 317 9989 337
rect 10004 335 10034 337
rect 9853 309 9894 317
rect 9976 313 9989 317
rect 10041 321 10120 337
rect 10152 337 10324 339
rect 10152 321 10231 337
rect 10238 335 10268 337
rect 9816 299 9845 309
rect 9859 299 9888 309
rect 9903 299 9933 313
rect 9976 299 10019 313
rect 10041 309 10231 321
rect 10296 317 10302 337
rect 10026 299 10056 309
rect 10057 299 10215 309
rect 10219 299 10249 309
rect 10253 299 10283 313
rect 10311 299 10324 337
rect 10396 351 10425 367
rect 10439 351 10468 367
rect 10483 357 10513 373
rect 10541 351 10547 399
rect 10550 393 10569 399
rect 10584 393 10614 401
rect 10550 385 10614 393
rect 10550 369 10630 385
rect 10646 378 10708 409
rect 10724 378 10786 409
rect 10855 407 10904 432
rect 10919 407 10949 423
rect 10818 393 10848 401
rect 10855 399 10965 407
rect 10818 385 10863 393
rect 10550 367 10569 369
rect 10584 367 10630 369
rect 10550 351 10630 367
rect 10657 365 10692 378
rect 10733 375 10770 378
rect 10733 373 10775 375
rect 10662 362 10692 365
rect 10671 358 10678 362
rect 10678 357 10679 358
rect 10637 351 10647 357
rect 10396 343 10431 351
rect 10396 317 10397 343
rect 10404 317 10431 343
rect 10339 299 10369 313
rect 10396 309 10431 317
rect 10433 343 10474 351
rect 10433 317 10448 343
rect 10455 317 10474 343
rect 10538 339 10569 351
rect 10584 339 10687 351
rect 10699 341 10725 367
rect 10740 362 10770 373
rect 10802 369 10864 385
rect 10802 367 10848 369
rect 10802 351 10864 367
rect 10876 351 10882 399
rect 10885 391 10965 399
rect 10885 389 10904 391
rect 10919 389 10953 391
rect 10885 373 10965 389
rect 10885 351 10904 373
rect 10919 357 10949 373
rect 10977 367 10983 441
rect 10986 367 11005 511
rect 11020 367 11026 511
rect 11035 441 11048 511
rect 11100 506 11122 511
rect 11093 485 11122 499
rect 11175 485 11191 499
rect 11229 495 11235 497
rect 11242 495 11350 511
rect 11357 495 11363 497
rect 11371 495 11386 511
rect 11452 505 11471 508
rect 11093 483 11191 485
rect 11218 483 11386 495
rect 11401 485 11417 499
rect 11452 486 11474 505
rect 11484 499 11500 500
rect 11483 497 11500 499
rect 11484 492 11500 497
rect 11474 485 11480 486
rect 11483 485 11512 492
rect 11401 484 11512 485
rect 11401 483 11518 484
rect 11077 475 11128 483
rect 11175 475 11209 483
rect 11077 463 11102 475
rect 11109 463 11128 475
rect 11182 473 11209 475
rect 11218 473 11439 483
rect 11474 480 11480 483
rect 11182 469 11439 473
rect 11077 455 11128 463
rect 11175 455 11439 469
rect 11483 475 11518 483
rect 11029 407 11048 441
rect 11093 447 11122 455
rect 11093 441 11110 447
rect 11093 439 11127 441
rect 11175 439 11191 455
rect 11192 445 11400 455
rect 11401 445 11417 455
rect 11465 451 11480 466
rect 11483 463 11484 475
rect 11491 463 11518 475
rect 11483 455 11518 463
rect 11483 454 11512 455
rect 11203 441 11417 445
rect 11218 439 11417 441
rect 11452 441 11465 451
rect 11483 441 11500 454
rect 11452 439 11500 441
rect 11094 435 11127 439
rect 11090 433 11127 435
rect 11090 432 11157 433
rect 11090 427 11121 432
rect 11127 427 11157 432
rect 11090 423 11157 427
rect 11063 420 11157 423
rect 11063 413 11112 420
rect 11063 407 11093 413
rect 11112 408 11117 413
rect 11029 391 11109 407
rect 11121 399 11157 420
rect 11218 415 11407 439
rect 11452 438 11499 439
rect 11465 433 11499 438
rect 11233 412 11407 415
rect 11226 409 11407 412
rect 11435 432 11499 433
rect 11029 389 11048 391
rect 11063 389 11097 391
rect 11029 373 11109 389
rect 11029 367 11048 373
rect 10745 341 10848 351
rect 10699 339 10848 341
rect 10869 339 10904 351
rect 10538 337 10700 339
rect 10550 317 10569 337
rect 10584 335 10614 337
rect 10433 309 10474 317
rect 10556 313 10569 317
rect 10621 321 10700 337
rect 10732 337 10904 339
rect 10732 321 10811 337
rect 10818 335 10848 337
rect 10396 299 10425 309
rect 10439 299 10468 309
rect 10483 299 10513 313
rect 10556 299 10599 313
rect 10621 309 10811 321
rect 10876 317 10882 337
rect 10606 299 10636 309
rect 10637 299 10795 309
rect 10799 299 10829 309
rect 10833 299 10863 313
rect 10891 299 10904 337
rect 10976 351 11005 367
rect 11019 351 11048 367
rect 11063 357 11093 373
rect 11121 351 11127 399
rect 11130 393 11149 399
rect 11164 393 11194 401
rect 11130 385 11194 393
rect 11130 369 11210 385
rect 11226 378 11288 409
rect 11304 378 11366 409
rect 11435 407 11484 432
rect 11499 407 11529 423
rect 11398 393 11428 401
rect 11435 399 11545 407
rect 11398 385 11443 393
rect 11130 367 11149 369
rect 11164 367 11210 369
rect 11130 351 11210 367
rect 11237 365 11272 378
rect 11313 375 11350 378
rect 11313 373 11355 375
rect 11242 362 11272 365
rect 11251 358 11258 362
rect 11258 357 11259 358
rect 11217 351 11227 357
rect 10976 343 11011 351
rect 10976 317 10977 343
rect 10984 317 11011 343
rect 10919 299 10949 313
rect 10976 309 11011 317
rect 11013 343 11054 351
rect 11013 317 11028 343
rect 11035 317 11054 343
rect 11118 339 11149 351
rect 11164 339 11267 351
rect 11279 341 11305 367
rect 11320 362 11350 373
rect 11382 369 11444 385
rect 11382 367 11428 369
rect 11382 351 11444 367
rect 11456 351 11462 399
rect 11465 391 11545 399
rect 11465 389 11484 391
rect 11499 389 11533 391
rect 11465 373 11545 389
rect 11465 351 11484 373
rect 11499 357 11529 373
rect 11557 367 11563 441
rect 11566 367 11585 511
rect 11600 367 11606 511
rect 11615 441 11628 511
rect 11680 506 11702 511
rect 11673 485 11702 499
rect 11755 485 11771 499
rect 11809 495 11815 497
rect 11822 495 11930 511
rect 11937 495 11943 497
rect 11951 495 11966 511
rect 12032 505 12051 508
rect 11673 483 11771 485
rect 11798 483 11966 495
rect 11981 485 11997 499
rect 12032 486 12054 505
rect 12064 499 12080 500
rect 12063 497 12080 499
rect 12064 492 12080 497
rect 12054 485 12060 486
rect 12063 485 12092 492
rect 11981 484 12092 485
rect 11981 483 12098 484
rect 11657 475 11708 483
rect 11755 475 11789 483
rect 11657 463 11682 475
rect 11689 463 11708 475
rect 11762 473 11789 475
rect 11798 473 12019 483
rect 12054 480 12060 483
rect 11762 469 12019 473
rect 11657 455 11708 463
rect 11755 455 12019 469
rect 12063 475 12098 483
rect 11609 407 11628 441
rect 11673 447 11702 455
rect 11673 441 11690 447
rect 11673 439 11707 441
rect 11755 439 11771 455
rect 11772 445 11980 455
rect 11981 445 11997 455
rect 12045 451 12060 466
rect 12063 463 12064 475
rect 12071 463 12098 475
rect 12063 455 12098 463
rect 12063 454 12092 455
rect 11783 441 11997 445
rect 11798 439 11997 441
rect 12032 441 12045 451
rect 12063 441 12080 454
rect 12032 439 12080 441
rect 11674 435 11707 439
rect 11670 433 11707 435
rect 11670 432 11737 433
rect 11670 427 11701 432
rect 11707 427 11737 432
rect 11670 423 11737 427
rect 11643 420 11737 423
rect 11643 413 11692 420
rect 11643 407 11673 413
rect 11692 408 11697 413
rect 11609 391 11689 407
rect 11701 399 11737 420
rect 11798 415 11987 439
rect 12032 438 12079 439
rect 12045 433 12079 438
rect 11813 412 11987 415
rect 11806 409 11987 412
rect 12015 432 12079 433
rect 11609 389 11628 391
rect 11643 389 11677 391
rect 11609 373 11689 389
rect 11609 367 11628 373
rect 11325 341 11428 351
rect 11279 339 11428 341
rect 11449 339 11484 351
rect 11118 337 11280 339
rect 11130 317 11149 337
rect 11164 335 11194 337
rect 11013 309 11054 317
rect 11136 313 11149 317
rect 11201 321 11280 337
rect 11312 337 11484 339
rect 11312 321 11391 337
rect 11398 335 11428 337
rect 10976 299 11005 309
rect 11019 299 11048 309
rect 11063 299 11093 313
rect 11136 299 11179 313
rect 11201 309 11391 321
rect 11456 317 11462 337
rect 11186 299 11216 309
rect 11217 299 11375 309
rect 11379 299 11409 309
rect 11413 299 11443 313
rect 11471 299 11484 337
rect 11556 351 11585 367
rect 11599 351 11628 367
rect 11643 357 11673 373
rect 11701 351 11707 399
rect 11710 393 11729 399
rect 11744 393 11774 401
rect 11710 385 11774 393
rect 11710 369 11790 385
rect 11806 378 11868 409
rect 11884 378 11946 409
rect 12015 407 12064 432
rect 12079 407 12109 423
rect 11978 393 12008 401
rect 12015 399 12125 407
rect 11978 385 12023 393
rect 11710 367 11729 369
rect 11744 367 11790 369
rect 11710 351 11790 367
rect 11817 365 11852 378
rect 11893 375 11930 378
rect 11893 373 11935 375
rect 11822 362 11852 365
rect 11831 358 11838 362
rect 11838 357 11839 358
rect 11797 351 11807 357
rect 11556 343 11591 351
rect 11556 317 11557 343
rect 11564 317 11591 343
rect 11499 299 11529 313
rect 11556 309 11591 317
rect 11593 343 11634 351
rect 11593 317 11608 343
rect 11615 317 11634 343
rect 11698 339 11729 351
rect 11744 339 11847 351
rect 11859 341 11885 367
rect 11900 362 11930 373
rect 11962 369 12024 385
rect 11962 367 12008 369
rect 11962 351 12024 367
rect 12036 351 12042 399
rect 12045 391 12125 399
rect 12045 389 12064 391
rect 12079 389 12113 391
rect 12045 373 12125 389
rect 12045 351 12064 373
rect 12079 357 12109 373
rect 12137 367 12143 441
rect 12146 367 12165 511
rect 12180 367 12186 511
rect 12195 441 12208 511
rect 12260 506 12282 511
rect 12253 485 12282 499
rect 12335 485 12351 499
rect 12389 495 12395 497
rect 12402 495 12510 511
rect 12517 495 12523 497
rect 12531 495 12546 511
rect 12612 505 12631 508
rect 12253 483 12351 485
rect 12378 483 12546 495
rect 12561 485 12577 499
rect 12612 486 12634 505
rect 12644 499 12660 500
rect 12643 497 12660 499
rect 12644 492 12660 497
rect 12634 485 12640 486
rect 12643 485 12672 492
rect 12561 484 12672 485
rect 12561 483 12678 484
rect 12237 475 12288 483
rect 12335 475 12369 483
rect 12237 463 12262 475
rect 12269 463 12288 475
rect 12342 473 12369 475
rect 12378 473 12599 483
rect 12634 480 12640 483
rect 12342 469 12599 473
rect 12237 455 12288 463
rect 12335 455 12599 469
rect 12643 475 12678 483
rect 12189 407 12208 441
rect 12253 447 12282 455
rect 12253 441 12270 447
rect 12253 439 12287 441
rect 12335 439 12351 455
rect 12352 445 12560 455
rect 12561 445 12577 455
rect 12625 451 12640 466
rect 12643 463 12644 475
rect 12651 463 12678 475
rect 12643 455 12678 463
rect 12643 454 12672 455
rect 12363 441 12577 445
rect 12378 439 12577 441
rect 12612 441 12625 451
rect 12643 441 12660 454
rect 12612 439 12660 441
rect 12254 435 12287 439
rect 12250 433 12287 435
rect 12250 432 12317 433
rect 12250 427 12281 432
rect 12287 427 12317 432
rect 12250 423 12317 427
rect 12223 420 12317 423
rect 12223 413 12272 420
rect 12223 407 12253 413
rect 12272 408 12277 413
rect 12189 391 12269 407
rect 12281 399 12317 420
rect 12378 415 12567 439
rect 12612 438 12659 439
rect 12625 433 12659 438
rect 12393 412 12567 415
rect 12386 409 12567 412
rect 12595 432 12659 433
rect 12189 389 12208 391
rect 12223 389 12257 391
rect 12189 373 12269 389
rect 12189 367 12208 373
rect 11905 341 12008 351
rect 11859 339 12008 341
rect 12029 339 12064 351
rect 11698 337 11860 339
rect 11710 317 11729 337
rect 11744 335 11774 337
rect 11593 309 11634 317
rect 11716 313 11729 317
rect 11781 321 11860 337
rect 11892 337 12064 339
rect 11892 321 11971 337
rect 11978 335 12008 337
rect 11556 299 11585 309
rect 11599 299 11628 309
rect 11643 299 11673 313
rect 11716 299 11759 313
rect 11781 309 11971 321
rect 12036 317 12042 337
rect 11766 299 11796 309
rect 11797 299 11955 309
rect 11959 299 11989 309
rect 11993 299 12023 313
rect 12051 299 12064 337
rect 12136 351 12165 367
rect 12179 351 12208 367
rect 12223 357 12253 373
rect 12281 351 12287 399
rect 12290 393 12309 399
rect 12324 393 12354 401
rect 12290 385 12354 393
rect 12290 369 12370 385
rect 12386 378 12448 409
rect 12464 378 12526 409
rect 12595 407 12644 432
rect 12659 407 12689 423
rect 12558 393 12588 401
rect 12595 399 12705 407
rect 12558 385 12603 393
rect 12290 367 12309 369
rect 12324 367 12370 369
rect 12290 351 12370 367
rect 12397 365 12432 378
rect 12473 375 12510 378
rect 12473 373 12515 375
rect 12402 362 12432 365
rect 12411 358 12418 362
rect 12418 357 12419 358
rect 12377 351 12387 357
rect 12136 343 12171 351
rect 12136 317 12137 343
rect 12144 317 12171 343
rect 12079 299 12109 313
rect 12136 309 12171 317
rect 12173 343 12214 351
rect 12173 317 12188 343
rect 12195 317 12214 343
rect 12278 339 12309 351
rect 12324 339 12427 351
rect 12439 341 12465 367
rect 12480 362 12510 373
rect 12542 369 12604 385
rect 12542 367 12588 369
rect 12542 351 12604 367
rect 12616 351 12622 399
rect 12625 391 12705 399
rect 12625 389 12644 391
rect 12659 389 12693 391
rect 12625 373 12705 389
rect 12625 351 12644 373
rect 12659 357 12689 373
rect 12717 367 12723 441
rect 12726 367 12745 511
rect 12760 367 12766 511
rect 12775 441 12788 511
rect 12840 506 12862 511
rect 12833 485 12862 499
rect 12915 485 12931 499
rect 12969 495 12975 497
rect 12982 495 13090 511
rect 13097 495 13103 497
rect 13111 495 13126 511
rect 13192 505 13211 508
rect 12833 483 12931 485
rect 12958 483 13126 495
rect 13141 485 13157 499
rect 13192 486 13214 505
rect 13224 499 13240 500
rect 13223 497 13240 499
rect 13224 492 13240 497
rect 13214 485 13220 486
rect 13223 485 13252 492
rect 13141 484 13252 485
rect 13141 483 13258 484
rect 12817 475 12868 483
rect 12915 475 12949 483
rect 12817 463 12842 475
rect 12849 463 12868 475
rect 12922 473 12949 475
rect 12958 473 13179 483
rect 13214 480 13220 483
rect 12922 469 13179 473
rect 12817 455 12868 463
rect 12915 455 13179 469
rect 13223 475 13258 483
rect 12769 407 12788 441
rect 12833 447 12862 455
rect 12833 441 12850 447
rect 12833 439 12867 441
rect 12915 439 12931 455
rect 12932 445 13140 455
rect 13141 445 13157 455
rect 13205 451 13220 466
rect 13223 463 13224 475
rect 13231 463 13258 475
rect 13223 455 13258 463
rect 13223 454 13252 455
rect 12943 441 13157 445
rect 12958 439 13157 441
rect 13192 441 13205 451
rect 13223 441 13240 454
rect 13192 439 13240 441
rect 12834 435 12867 439
rect 12830 433 12867 435
rect 12830 432 12897 433
rect 12830 427 12861 432
rect 12867 427 12897 432
rect 12830 423 12897 427
rect 12803 420 12897 423
rect 12803 413 12852 420
rect 12803 407 12833 413
rect 12852 408 12857 413
rect 12769 391 12849 407
rect 12861 399 12897 420
rect 12958 415 13147 439
rect 13192 438 13239 439
rect 13205 433 13239 438
rect 12973 412 13147 415
rect 12966 409 13147 412
rect 13175 432 13239 433
rect 12769 389 12788 391
rect 12803 389 12837 391
rect 12769 373 12849 389
rect 12769 367 12788 373
rect 12485 341 12588 351
rect 12439 339 12588 341
rect 12609 339 12644 351
rect 12278 337 12440 339
rect 12290 317 12309 337
rect 12324 335 12354 337
rect 12173 309 12214 317
rect 12296 313 12309 317
rect 12361 321 12440 337
rect 12472 337 12644 339
rect 12472 321 12551 337
rect 12558 335 12588 337
rect 12136 299 12165 309
rect 12179 299 12208 309
rect 12223 299 12253 313
rect 12296 299 12339 313
rect 12361 309 12551 321
rect 12616 317 12622 337
rect 12346 299 12376 309
rect 12377 299 12535 309
rect 12539 299 12569 309
rect 12573 299 12603 313
rect 12631 299 12644 337
rect 12716 351 12745 367
rect 12759 351 12788 367
rect 12803 357 12833 373
rect 12861 351 12867 399
rect 12870 393 12889 399
rect 12904 393 12934 401
rect 12870 385 12934 393
rect 12870 369 12950 385
rect 12966 378 13028 409
rect 13044 378 13106 409
rect 13175 407 13224 432
rect 13239 407 13269 423
rect 13138 393 13168 401
rect 13175 399 13285 407
rect 13138 385 13183 393
rect 12870 367 12889 369
rect 12904 367 12950 369
rect 12870 351 12950 367
rect 12977 365 13012 378
rect 13053 375 13090 378
rect 13053 373 13095 375
rect 12982 362 13012 365
rect 12991 358 12998 362
rect 12998 357 12999 358
rect 12957 351 12967 357
rect 12716 343 12751 351
rect 12716 317 12717 343
rect 12724 317 12751 343
rect 12659 299 12689 313
rect 12716 309 12751 317
rect 12753 343 12794 351
rect 12753 317 12768 343
rect 12775 317 12794 343
rect 12858 339 12889 351
rect 12904 339 13007 351
rect 13019 341 13045 367
rect 13060 362 13090 373
rect 13122 369 13184 385
rect 13122 367 13168 369
rect 13122 351 13184 367
rect 13196 351 13202 399
rect 13205 391 13285 399
rect 13205 389 13224 391
rect 13239 389 13273 391
rect 13205 373 13285 389
rect 13205 351 13224 373
rect 13239 357 13269 373
rect 13297 367 13303 441
rect 13306 367 13325 511
rect 13340 367 13346 511
rect 13355 441 13368 511
rect 13420 506 13442 511
rect 13413 485 13442 499
rect 13495 485 13511 499
rect 13549 495 13555 497
rect 13562 495 13670 511
rect 13677 495 13683 497
rect 13691 495 13706 511
rect 13886 510 13926 511
rect 13772 505 13791 508
rect 13413 483 13511 485
rect 13538 483 13706 495
rect 13721 485 13737 499
rect 13772 486 13794 505
rect 13804 499 13820 500
rect 13803 497 13820 499
rect 13804 492 13820 497
rect 13794 485 13800 486
rect 13803 485 13832 492
rect 13721 484 13832 485
rect 13721 483 13838 484
rect 13397 475 13448 483
rect 13495 475 13529 483
rect 13397 463 13422 475
rect 13429 463 13448 475
rect 13502 473 13529 475
rect 13538 473 13759 483
rect 13794 480 13800 483
rect 13502 469 13759 473
rect 13397 455 13448 463
rect 13495 455 13759 469
rect 13803 475 13838 483
rect 13349 407 13368 441
rect 13413 447 13442 455
rect 13413 441 13430 447
rect 13413 439 13447 441
rect 13495 439 13511 455
rect 13512 445 13720 455
rect 13721 445 13737 455
rect 13785 451 13800 466
rect 13803 463 13804 475
rect 13811 463 13838 475
rect 13803 455 13838 463
rect 13803 454 13832 455
rect 13523 441 13737 445
rect 13538 439 13737 441
rect 13772 441 13785 451
rect 13803 441 13820 454
rect 13772 439 13820 441
rect 13414 435 13447 439
rect 13410 433 13447 435
rect 13410 432 13477 433
rect 13410 427 13441 432
rect 13447 427 13477 432
rect 13410 423 13477 427
rect 13383 420 13477 423
rect 13383 413 13432 420
rect 13383 407 13413 413
rect 13432 408 13437 413
rect 13349 391 13429 407
rect 13441 399 13477 420
rect 13538 415 13727 439
rect 13772 438 13819 439
rect 13785 433 13819 438
rect 13553 412 13727 415
rect 13546 409 13727 412
rect 13755 432 13819 433
rect 13349 389 13368 391
rect 13383 389 13417 391
rect 13349 373 13429 389
rect 13349 367 13368 373
rect 13065 341 13168 351
rect 13019 339 13168 341
rect 13189 339 13224 351
rect 12858 337 13020 339
rect 12870 317 12889 337
rect 12904 335 12934 337
rect 12753 309 12794 317
rect 12876 313 12889 317
rect 12941 321 13020 337
rect 13052 337 13224 339
rect 13052 321 13131 337
rect 13138 335 13168 337
rect 12716 299 12745 309
rect 12759 299 12788 309
rect 12803 299 12833 313
rect 12876 299 12919 313
rect 12941 309 13131 321
rect 13196 317 13202 337
rect 12926 299 12956 309
rect 12957 299 13115 309
rect 13119 299 13149 309
rect 13153 299 13183 313
rect 13211 299 13224 337
rect 13296 351 13325 367
rect 13339 351 13368 367
rect 13383 357 13413 373
rect 13441 351 13447 399
rect 13450 393 13469 399
rect 13484 393 13514 401
rect 13450 385 13514 393
rect 13450 369 13530 385
rect 13546 378 13608 409
rect 13624 378 13686 409
rect 13755 407 13804 432
rect 13819 407 13849 423
rect 13718 393 13748 401
rect 13755 399 13865 407
rect 13718 385 13763 393
rect 13450 367 13469 369
rect 13484 367 13530 369
rect 13450 351 13530 367
rect 13557 365 13592 378
rect 13633 375 13670 378
rect 13633 373 13675 375
rect 13562 362 13592 365
rect 13571 358 13578 362
rect 13578 357 13579 358
rect 13537 351 13547 357
rect 13296 343 13331 351
rect 13296 317 13297 343
rect 13304 317 13331 343
rect 13239 299 13269 313
rect 13296 309 13331 317
rect 13333 343 13374 351
rect 13333 317 13348 343
rect 13355 317 13374 343
rect 13438 339 13469 351
rect 13484 339 13587 351
rect 13599 341 13625 367
rect 13640 362 13670 373
rect 13702 369 13764 385
rect 13702 367 13748 369
rect 13702 351 13764 367
rect 13776 351 13782 399
rect 13785 391 13865 399
rect 13785 389 13804 391
rect 13819 389 13853 391
rect 13785 373 13865 389
rect 13785 351 13804 373
rect 13819 357 13849 373
rect 13877 367 13883 441
rect 13886 367 13905 510
rect 13920 367 13926 510
rect 13935 441 13948 511
rect 14000 506 14022 511
rect 13993 485 14022 499
rect 14075 485 14091 499
rect 14129 495 14135 497
rect 14142 495 14250 511
rect 14257 495 14263 497
rect 14271 495 14286 511
rect 14352 505 14371 508
rect 13993 483 14091 485
rect 14118 483 14286 495
rect 14301 485 14317 499
rect 14352 486 14374 505
rect 14384 499 14400 500
rect 14383 497 14400 499
rect 14384 492 14400 497
rect 14374 485 14380 486
rect 14383 485 14412 492
rect 14301 484 14412 485
rect 14301 483 14418 484
rect 13977 475 14028 483
rect 14075 475 14109 483
rect 13977 463 14002 475
rect 14009 463 14028 475
rect 14082 473 14109 475
rect 14118 473 14339 483
rect 14374 480 14380 483
rect 14082 469 14339 473
rect 13977 455 14028 463
rect 14075 455 14339 469
rect 14383 475 14418 483
rect 13929 407 13948 441
rect 13993 447 14022 455
rect 13993 441 14010 447
rect 13993 439 14027 441
rect 14075 439 14091 455
rect 14092 445 14300 455
rect 14301 445 14317 455
rect 14365 451 14380 466
rect 14383 463 14384 475
rect 14391 463 14418 475
rect 14383 455 14418 463
rect 14383 454 14412 455
rect 14103 441 14317 445
rect 14118 439 14317 441
rect 14352 441 14365 451
rect 14383 441 14400 454
rect 14352 439 14400 441
rect 13994 435 14027 439
rect 13990 433 14027 435
rect 13990 432 14057 433
rect 13990 427 14021 432
rect 14027 427 14057 432
rect 13990 423 14057 427
rect 13963 420 14057 423
rect 13963 413 14012 420
rect 13963 407 13993 413
rect 14012 408 14017 413
rect 13929 391 14009 407
rect 14021 399 14057 420
rect 14118 415 14307 439
rect 14352 438 14399 439
rect 14365 433 14399 438
rect 14133 412 14307 415
rect 14126 409 14307 412
rect 14335 432 14399 433
rect 13929 389 13948 391
rect 13963 389 13997 391
rect 13929 373 14009 389
rect 13929 367 13948 373
rect 13645 341 13748 351
rect 13599 339 13748 341
rect 13769 339 13804 351
rect 13438 337 13600 339
rect 13450 317 13469 337
rect 13484 335 13514 337
rect 13333 309 13374 317
rect 13456 313 13469 317
rect 13521 321 13600 337
rect 13632 337 13804 339
rect 13632 321 13711 337
rect 13718 335 13748 337
rect 13296 299 13325 309
rect 13339 299 13368 309
rect 13383 299 13413 313
rect 13456 299 13499 313
rect 13521 309 13711 321
rect 13776 317 13782 337
rect 13506 299 13536 309
rect 13537 299 13695 309
rect 13699 299 13729 309
rect 13733 299 13763 313
rect 13791 299 13804 337
rect 13876 351 13905 367
rect 13919 351 13948 367
rect 13963 357 13993 373
rect 14021 351 14027 399
rect 14030 393 14049 399
rect 14064 393 14094 401
rect 14030 385 14094 393
rect 14030 369 14110 385
rect 14126 378 14188 409
rect 14204 378 14266 409
rect 14335 407 14384 432
rect 14399 407 14429 423
rect 14298 393 14328 401
rect 14335 399 14445 407
rect 14298 385 14343 393
rect 14030 367 14049 369
rect 14064 367 14110 369
rect 14030 351 14110 367
rect 14137 365 14172 378
rect 14213 375 14250 378
rect 14213 373 14255 375
rect 14142 362 14172 365
rect 14151 358 14158 362
rect 14158 357 14159 358
rect 14117 351 14127 357
rect 13876 343 13911 351
rect 13876 317 13877 343
rect 13884 317 13911 343
rect 13819 299 13849 313
rect 13876 309 13911 317
rect 13913 343 13954 351
rect 13913 317 13928 343
rect 13935 317 13954 343
rect 14018 339 14049 351
rect 14064 339 14167 351
rect 14179 341 14205 367
rect 14220 362 14250 373
rect 14282 369 14344 385
rect 14282 367 14328 369
rect 14282 351 14344 367
rect 14356 351 14362 399
rect 14365 391 14445 399
rect 14365 389 14384 391
rect 14399 389 14433 391
rect 14365 373 14445 389
rect 14365 351 14384 373
rect 14399 357 14429 373
rect 14457 367 14463 441
rect 14466 367 14485 511
rect 14500 367 14506 511
rect 14515 441 14528 511
rect 14580 506 14602 511
rect 14573 485 14602 499
rect 14655 485 14671 499
rect 14709 495 14715 497
rect 14722 495 14830 511
rect 14837 495 14843 497
rect 14851 495 14866 511
rect 14932 505 14951 508
rect 14573 483 14671 485
rect 14698 483 14866 495
rect 14881 485 14897 499
rect 14932 486 14954 505
rect 14964 499 14980 500
rect 14963 497 14980 499
rect 14964 492 14980 497
rect 14954 485 14960 486
rect 14963 485 14992 492
rect 14881 484 14992 485
rect 14881 483 14998 484
rect 14557 475 14608 483
rect 14655 475 14689 483
rect 14557 463 14582 475
rect 14589 463 14608 475
rect 14662 473 14689 475
rect 14698 473 14919 483
rect 14954 480 14960 483
rect 14662 469 14919 473
rect 14557 455 14608 463
rect 14655 455 14919 469
rect 14963 475 14998 483
rect 14509 407 14528 441
rect 14573 447 14602 455
rect 14573 441 14590 447
rect 14573 439 14607 441
rect 14655 439 14671 455
rect 14672 445 14880 455
rect 14881 445 14897 455
rect 14945 451 14960 466
rect 14963 463 14964 475
rect 14971 463 14998 475
rect 14963 455 14998 463
rect 14963 454 14992 455
rect 14683 441 14897 445
rect 14698 439 14897 441
rect 14932 441 14945 451
rect 14963 441 14980 454
rect 14932 439 14980 441
rect 14574 435 14607 439
rect 14570 433 14607 435
rect 14570 432 14637 433
rect 14570 427 14601 432
rect 14607 427 14637 432
rect 14570 423 14637 427
rect 14543 420 14637 423
rect 14543 413 14592 420
rect 14543 407 14573 413
rect 14592 408 14597 413
rect 14509 391 14589 407
rect 14601 399 14637 420
rect 14698 415 14887 439
rect 14932 438 14979 439
rect 14945 433 14979 438
rect 14713 412 14887 415
rect 14706 409 14887 412
rect 14915 432 14979 433
rect 14509 389 14528 391
rect 14543 389 14577 391
rect 14509 373 14589 389
rect 14509 367 14528 373
rect 14225 341 14328 351
rect 14179 339 14328 341
rect 14349 339 14384 351
rect 14018 337 14180 339
rect 14030 317 14049 337
rect 14064 335 14094 337
rect 13913 309 13954 317
rect 14036 313 14049 317
rect 14101 321 14180 337
rect 14212 337 14384 339
rect 14212 321 14291 337
rect 14298 335 14328 337
rect 13876 299 13905 309
rect 13919 299 13948 309
rect 13963 299 13993 313
rect 14036 299 14079 313
rect 14101 309 14291 321
rect 14356 317 14362 337
rect 14086 299 14116 309
rect 14117 299 14275 309
rect 14279 299 14309 309
rect 14313 299 14343 313
rect 14371 299 14384 337
rect 14456 351 14485 367
rect 14499 351 14528 367
rect 14543 357 14573 373
rect 14601 351 14607 399
rect 14610 393 14629 399
rect 14644 393 14674 401
rect 14610 385 14674 393
rect 14610 369 14690 385
rect 14706 378 14768 409
rect 14784 378 14846 409
rect 14915 407 14964 432
rect 14979 407 15009 423
rect 14878 393 14908 401
rect 14915 399 15025 407
rect 14878 385 14923 393
rect 14610 367 14629 369
rect 14644 367 14690 369
rect 14610 351 14690 367
rect 14717 365 14752 378
rect 14793 375 14830 378
rect 14793 373 14835 375
rect 14722 362 14752 365
rect 14731 358 14738 362
rect 14738 357 14739 358
rect 14697 351 14707 357
rect 14456 343 14491 351
rect 14456 317 14457 343
rect 14464 317 14491 343
rect 14399 299 14429 313
rect 14456 309 14491 317
rect 14493 343 14534 351
rect 14493 317 14508 343
rect 14515 317 14534 343
rect 14598 339 14629 351
rect 14644 339 14747 351
rect 14759 341 14785 367
rect 14800 362 14830 373
rect 14862 369 14924 385
rect 14862 367 14908 369
rect 14862 351 14924 367
rect 14936 351 14942 399
rect 14945 391 15025 399
rect 14945 389 14964 391
rect 14979 389 15013 391
rect 14945 373 15025 389
rect 14945 351 14964 373
rect 14979 357 15009 373
rect 15037 367 15043 441
rect 15046 367 15065 511
rect 15080 367 15086 511
rect 15095 441 15108 511
rect 15160 506 15182 511
rect 15153 485 15182 499
rect 15235 485 15251 499
rect 15289 495 15295 497
rect 15302 495 15410 511
rect 15417 495 15423 497
rect 15431 495 15446 511
rect 15512 505 15531 508
rect 15153 483 15251 485
rect 15278 483 15446 495
rect 15461 485 15477 499
rect 15512 486 15534 505
rect 15544 499 15560 500
rect 15543 497 15560 499
rect 15544 492 15560 497
rect 15534 485 15540 486
rect 15543 485 15572 492
rect 15461 484 15572 485
rect 15461 483 15578 484
rect 15137 475 15188 483
rect 15235 475 15269 483
rect 15137 463 15162 475
rect 15169 463 15188 475
rect 15242 473 15269 475
rect 15278 473 15499 483
rect 15534 480 15540 483
rect 15242 469 15499 473
rect 15137 455 15188 463
rect 15235 455 15499 469
rect 15543 475 15578 483
rect 15089 407 15108 441
rect 15153 447 15182 455
rect 15153 441 15170 447
rect 15153 439 15187 441
rect 15235 439 15251 455
rect 15252 445 15460 455
rect 15461 445 15477 455
rect 15525 451 15540 466
rect 15543 463 15544 475
rect 15551 463 15578 475
rect 15543 455 15578 463
rect 15543 454 15572 455
rect 15263 441 15477 445
rect 15278 439 15477 441
rect 15512 441 15525 451
rect 15543 441 15560 454
rect 15512 439 15560 441
rect 15154 435 15187 439
rect 15150 433 15187 435
rect 15150 432 15217 433
rect 15150 427 15181 432
rect 15187 427 15217 432
rect 15150 423 15217 427
rect 15123 420 15217 423
rect 15123 413 15172 420
rect 15123 407 15153 413
rect 15172 408 15177 413
rect 15089 391 15169 407
rect 15181 399 15217 420
rect 15278 415 15467 439
rect 15512 438 15559 439
rect 15525 433 15559 438
rect 15293 412 15467 415
rect 15286 409 15467 412
rect 15495 432 15559 433
rect 15089 389 15108 391
rect 15123 389 15157 391
rect 15089 373 15169 389
rect 15089 367 15108 373
rect 14805 341 14908 351
rect 14759 339 14908 341
rect 14929 339 14964 351
rect 14598 337 14760 339
rect 14610 317 14629 337
rect 14644 335 14674 337
rect 14493 309 14534 317
rect 14616 313 14629 317
rect 14681 321 14760 337
rect 14792 337 14964 339
rect 14792 321 14871 337
rect 14878 335 14908 337
rect 14456 299 14485 309
rect 14499 299 14528 309
rect 14543 299 14573 313
rect 14616 299 14659 313
rect 14681 309 14871 321
rect 14936 317 14942 337
rect 14666 299 14696 309
rect 14697 299 14855 309
rect 14859 299 14889 309
rect 14893 299 14923 313
rect 14951 299 14964 337
rect 15036 351 15065 367
rect 15079 351 15108 367
rect 15123 357 15153 373
rect 15181 351 15187 399
rect 15190 393 15209 399
rect 15224 393 15254 401
rect 15190 385 15254 393
rect 15190 369 15270 385
rect 15286 378 15348 409
rect 15364 378 15426 409
rect 15495 407 15544 432
rect 15559 407 15589 423
rect 15458 393 15488 401
rect 15495 399 15605 407
rect 15458 385 15503 393
rect 15190 367 15209 369
rect 15224 367 15270 369
rect 15190 351 15270 367
rect 15297 365 15332 378
rect 15373 375 15410 378
rect 15373 373 15415 375
rect 15302 362 15332 365
rect 15311 358 15318 362
rect 15318 357 15319 358
rect 15277 351 15287 357
rect 15036 343 15071 351
rect 15036 317 15037 343
rect 15044 317 15071 343
rect 14979 299 15009 313
rect 15036 309 15071 317
rect 15073 343 15114 351
rect 15073 317 15088 343
rect 15095 317 15114 343
rect 15178 339 15209 351
rect 15224 339 15327 351
rect 15339 341 15365 367
rect 15380 362 15410 373
rect 15442 369 15504 385
rect 15442 367 15488 369
rect 15442 351 15504 367
rect 15516 351 15522 399
rect 15525 391 15605 399
rect 15525 389 15544 391
rect 15559 389 15593 391
rect 15525 373 15605 389
rect 15525 351 15544 373
rect 15559 357 15589 373
rect 15617 367 15623 441
rect 15626 367 15645 511
rect 15660 367 15666 511
rect 15675 441 15688 511
rect 15740 506 15762 511
rect 15733 485 15762 499
rect 15815 485 15831 499
rect 15869 495 15875 497
rect 15882 495 15990 511
rect 15997 495 16003 497
rect 16011 495 16026 511
rect 16092 505 16111 508
rect 15733 483 15831 485
rect 15858 483 16026 495
rect 16041 485 16057 499
rect 16092 486 16114 505
rect 16124 499 16140 500
rect 16123 497 16140 499
rect 16124 492 16140 497
rect 16114 485 16120 486
rect 16123 485 16152 492
rect 16041 484 16152 485
rect 16041 483 16158 484
rect 15717 475 15768 483
rect 15815 475 15849 483
rect 15717 463 15742 475
rect 15749 463 15768 475
rect 15822 473 15849 475
rect 15858 473 16079 483
rect 16114 480 16120 483
rect 15822 469 16079 473
rect 15717 455 15768 463
rect 15815 455 16079 469
rect 16123 475 16158 483
rect 15669 407 15688 441
rect 15733 447 15762 455
rect 15733 441 15750 447
rect 15733 439 15767 441
rect 15815 439 15831 455
rect 15832 445 16040 455
rect 16041 445 16057 455
rect 16105 451 16120 466
rect 16123 463 16124 475
rect 16131 463 16158 475
rect 16123 455 16158 463
rect 16123 454 16152 455
rect 15843 441 16057 445
rect 15858 439 16057 441
rect 16092 441 16105 451
rect 16123 441 16140 454
rect 16092 439 16140 441
rect 15734 435 15767 439
rect 15730 433 15767 435
rect 15730 432 15797 433
rect 15730 427 15761 432
rect 15767 427 15797 432
rect 15730 423 15797 427
rect 15703 420 15797 423
rect 15703 413 15752 420
rect 15703 407 15733 413
rect 15752 408 15757 413
rect 15669 391 15749 407
rect 15761 399 15797 420
rect 15858 415 16047 439
rect 16092 438 16139 439
rect 16105 433 16139 438
rect 15873 412 16047 415
rect 15866 409 16047 412
rect 16075 432 16139 433
rect 15669 389 15688 391
rect 15703 389 15737 391
rect 15669 373 15749 389
rect 15669 367 15688 373
rect 15385 341 15488 351
rect 15339 339 15488 341
rect 15509 339 15544 351
rect 15178 337 15340 339
rect 15190 317 15209 337
rect 15224 335 15254 337
rect 15073 309 15114 317
rect 15196 313 15209 317
rect 15261 321 15340 337
rect 15372 337 15544 339
rect 15372 321 15451 337
rect 15458 335 15488 337
rect 15036 299 15065 309
rect 15079 299 15108 309
rect 15123 299 15153 313
rect 15196 299 15239 313
rect 15261 309 15451 321
rect 15516 317 15522 337
rect 15246 299 15276 309
rect 15277 299 15435 309
rect 15439 299 15469 309
rect 15473 299 15503 313
rect 15531 299 15544 337
rect 15616 351 15645 367
rect 15659 351 15688 367
rect 15703 357 15733 373
rect 15761 351 15767 399
rect 15770 393 15789 399
rect 15804 393 15834 401
rect 15770 385 15834 393
rect 15770 369 15850 385
rect 15866 378 15928 409
rect 15944 378 16006 409
rect 16075 407 16124 432
rect 16139 407 16169 423
rect 16038 393 16068 401
rect 16075 399 16185 407
rect 16038 385 16083 393
rect 15770 367 15789 369
rect 15804 367 15850 369
rect 15770 351 15850 367
rect 15877 365 15912 378
rect 15953 375 15990 378
rect 15953 373 15995 375
rect 15882 362 15912 365
rect 15891 358 15898 362
rect 15898 357 15899 358
rect 15857 351 15867 357
rect 15616 343 15651 351
rect 15616 317 15617 343
rect 15624 317 15651 343
rect 15559 299 15589 313
rect 15616 309 15651 317
rect 15653 343 15694 351
rect 15653 317 15668 343
rect 15675 317 15694 343
rect 15758 339 15789 351
rect 15804 339 15907 351
rect 15919 341 15945 367
rect 15960 362 15990 373
rect 16022 369 16084 385
rect 16022 367 16068 369
rect 16022 351 16084 367
rect 16096 351 16102 399
rect 16105 391 16185 399
rect 16105 389 16124 391
rect 16139 389 16173 391
rect 16105 373 16185 389
rect 16105 351 16124 373
rect 16139 357 16169 373
rect 16197 367 16203 441
rect 16206 367 16225 511
rect 16240 367 16246 511
rect 16255 441 16268 511
rect 16320 506 16342 511
rect 16313 485 16342 499
rect 16395 485 16411 499
rect 16449 495 16455 497
rect 16462 495 16570 511
rect 16577 495 16583 497
rect 16591 495 16606 511
rect 16672 505 16691 508
rect 16313 483 16411 485
rect 16438 483 16606 495
rect 16621 485 16637 499
rect 16672 486 16694 505
rect 16704 499 16720 500
rect 16703 497 16720 499
rect 16704 492 16720 497
rect 16694 485 16700 486
rect 16703 485 16732 492
rect 16621 484 16732 485
rect 16621 483 16738 484
rect 16297 475 16348 483
rect 16395 475 16429 483
rect 16297 463 16322 475
rect 16329 463 16348 475
rect 16402 473 16429 475
rect 16438 473 16659 483
rect 16694 480 16700 483
rect 16402 469 16659 473
rect 16297 455 16348 463
rect 16395 455 16659 469
rect 16703 475 16738 483
rect 16249 407 16268 441
rect 16313 447 16342 455
rect 16313 441 16330 447
rect 16313 439 16347 441
rect 16395 439 16411 455
rect 16412 445 16620 455
rect 16621 445 16637 455
rect 16685 451 16700 466
rect 16703 463 16704 475
rect 16711 463 16738 475
rect 16703 455 16738 463
rect 16703 454 16732 455
rect 16423 441 16637 445
rect 16438 439 16637 441
rect 16672 441 16685 451
rect 16703 441 16720 454
rect 16672 439 16720 441
rect 16314 435 16347 439
rect 16310 433 16347 435
rect 16310 432 16377 433
rect 16310 427 16341 432
rect 16347 427 16377 432
rect 16310 423 16377 427
rect 16283 420 16377 423
rect 16283 413 16332 420
rect 16283 407 16313 413
rect 16332 408 16337 413
rect 16249 391 16329 407
rect 16341 399 16377 420
rect 16438 415 16627 439
rect 16672 438 16719 439
rect 16685 433 16719 438
rect 16453 412 16627 415
rect 16446 409 16627 412
rect 16655 432 16719 433
rect 16249 389 16268 391
rect 16283 389 16317 391
rect 16249 373 16329 389
rect 16249 367 16268 373
rect 15965 341 16068 351
rect 15919 339 16068 341
rect 16089 339 16124 351
rect 15758 337 15920 339
rect 15770 317 15789 337
rect 15804 335 15834 337
rect 15653 309 15694 317
rect 15776 313 15789 317
rect 15841 321 15920 337
rect 15952 337 16124 339
rect 15952 321 16031 337
rect 16038 335 16068 337
rect 15616 299 15645 309
rect 15659 299 15688 309
rect 15703 299 15733 313
rect 15776 299 15819 313
rect 15841 309 16031 321
rect 16096 317 16102 337
rect 15826 299 15856 309
rect 15857 299 16015 309
rect 16019 299 16049 309
rect 16053 299 16083 313
rect 16111 299 16124 337
rect 16196 351 16225 367
rect 16239 351 16268 367
rect 16283 357 16313 373
rect 16341 351 16347 399
rect 16350 393 16369 399
rect 16384 393 16414 401
rect 16350 385 16414 393
rect 16350 369 16430 385
rect 16446 378 16508 409
rect 16524 378 16586 409
rect 16655 407 16704 432
rect 16719 407 16749 423
rect 16618 393 16648 401
rect 16655 399 16765 407
rect 16618 385 16663 393
rect 16350 367 16369 369
rect 16384 367 16430 369
rect 16350 351 16430 367
rect 16457 365 16492 378
rect 16533 375 16570 378
rect 16533 373 16575 375
rect 16462 362 16492 365
rect 16471 358 16478 362
rect 16478 357 16479 358
rect 16437 351 16447 357
rect 16196 343 16231 351
rect 16196 317 16197 343
rect 16204 317 16231 343
rect 16139 299 16169 313
rect 16196 309 16231 317
rect 16233 343 16274 351
rect 16233 317 16248 343
rect 16255 317 16274 343
rect 16338 339 16369 351
rect 16384 339 16487 351
rect 16499 341 16525 367
rect 16540 362 16570 373
rect 16602 369 16664 385
rect 16602 367 16648 369
rect 16602 351 16664 367
rect 16676 351 16682 399
rect 16685 391 16765 399
rect 16685 389 16704 391
rect 16719 389 16753 391
rect 16685 373 16765 389
rect 16685 351 16704 373
rect 16719 357 16749 373
rect 16777 367 16783 441
rect 16786 367 16805 511
rect 16820 367 16826 511
rect 16835 441 16848 511
rect 16900 506 16922 511
rect 16893 485 16922 499
rect 16975 485 16991 499
rect 17029 495 17035 497
rect 17042 495 17150 511
rect 17157 495 17163 497
rect 17171 495 17186 511
rect 17252 505 17271 508
rect 16893 483 16991 485
rect 17018 483 17186 495
rect 17201 485 17217 499
rect 17252 486 17274 505
rect 17284 499 17300 500
rect 17283 497 17300 499
rect 17284 492 17300 497
rect 17274 485 17280 486
rect 17283 485 17312 492
rect 17201 484 17312 485
rect 17201 483 17318 484
rect 16877 475 16928 483
rect 16975 475 17009 483
rect 16877 463 16902 475
rect 16909 463 16928 475
rect 16982 473 17009 475
rect 17018 473 17239 483
rect 17274 480 17280 483
rect 16982 469 17239 473
rect 16877 455 16928 463
rect 16975 455 17239 469
rect 17283 475 17318 483
rect 16829 407 16848 441
rect 16893 447 16922 455
rect 16893 441 16910 447
rect 16893 439 16927 441
rect 16975 439 16991 455
rect 16992 445 17200 455
rect 17201 445 17217 455
rect 17265 451 17280 466
rect 17283 463 17284 475
rect 17291 463 17318 475
rect 17283 455 17318 463
rect 17283 454 17312 455
rect 17003 441 17217 445
rect 17018 439 17217 441
rect 17252 441 17265 451
rect 17283 441 17300 454
rect 17252 439 17300 441
rect 16894 435 16927 439
rect 16890 433 16927 435
rect 16890 432 16957 433
rect 16890 427 16921 432
rect 16927 427 16957 432
rect 16890 423 16957 427
rect 16863 420 16957 423
rect 16863 413 16912 420
rect 16863 407 16893 413
rect 16912 408 16917 413
rect 16829 391 16909 407
rect 16921 399 16957 420
rect 17018 415 17207 439
rect 17252 438 17299 439
rect 17265 433 17299 438
rect 17033 412 17207 415
rect 17026 409 17207 412
rect 17235 432 17299 433
rect 16829 389 16848 391
rect 16863 389 16897 391
rect 16829 373 16909 389
rect 16829 367 16848 373
rect 16545 341 16648 351
rect 16499 339 16648 341
rect 16669 339 16704 351
rect 16338 337 16500 339
rect 16350 317 16369 337
rect 16384 335 16414 337
rect 16233 309 16274 317
rect 16356 313 16369 317
rect 16421 321 16500 337
rect 16532 337 16704 339
rect 16532 321 16611 337
rect 16618 335 16648 337
rect 16196 299 16225 309
rect 16239 299 16268 309
rect 16283 299 16313 313
rect 16356 299 16399 313
rect 16421 309 16611 321
rect 16676 317 16682 337
rect 16406 299 16436 309
rect 16437 299 16595 309
rect 16599 299 16629 309
rect 16633 299 16663 313
rect 16691 299 16704 337
rect 16776 351 16805 367
rect 16819 351 16848 367
rect 16863 357 16893 373
rect 16921 351 16927 399
rect 16930 393 16949 399
rect 16964 393 16994 401
rect 16930 385 16994 393
rect 16930 369 17010 385
rect 17026 378 17088 409
rect 17104 378 17166 409
rect 17235 407 17284 432
rect 17299 407 17329 423
rect 17198 393 17228 401
rect 17235 399 17345 407
rect 17198 385 17243 393
rect 16930 367 16949 369
rect 16964 367 17010 369
rect 16930 351 17010 367
rect 17037 365 17072 378
rect 17113 375 17150 378
rect 17113 373 17155 375
rect 17042 362 17072 365
rect 17051 358 17058 362
rect 17058 357 17059 358
rect 17017 351 17027 357
rect 16776 343 16811 351
rect 16776 317 16777 343
rect 16784 317 16811 343
rect 16719 299 16749 313
rect 16776 309 16811 317
rect 16813 343 16854 351
rect 16813 317 16828 343
rect 16835 317 16854 343
rect 16918 339 16949 351
rect 16964 339 17067 351
rect 17079 341 17105 367
rect 17120 362 17150 373
rect 17182 369 17244 385
rect 17182 367 17228 369
rect 17182 351 17244 367
rect 17256 351 17262 399
rect 17265 391 17345 399
rect 17265 389 17284 391
rect 17299 389 17333 391
rect 17265 373 17345 389
rect 17265 351 17284 373
rect 17299 357 17329 373
rect 17357 367 17363 441
rect 17366 367 17385 511
rect 17400 367 17406 511
rect 17415 441 17428 511
rect 17480 506 17502 511
rect 17473 485 17502 499
rect 17555 485 17571 499
rect 17609 495 17615 497
rect 17622 495 17730 511
rect 17737 495 17743 497
rect 17751 495 17766 511
rect 17832 505 17851 508
rect 17473 483 17571 485
rect 17598 483 17766 495
rect 17781 485 17797 499
rect 17832 486 17854 505
rect 17864 499 17880 500
rect 17863 497 17880 499
rect 17864 492 17880 497
rect 17854 485 17860 486
rect 17863 485 17892 492
rect 17781 484 17892 485
rect 17781 483 17898 484
rect 17457 475 17508 483
rect 17555 475 17589 483
rect 17457 463 17482 475
rect 17489 463 17508 475
rect 17562 473 17589 475
rect 17598 473 17819 483
rect 17854 480 17860 483
rect 17562 469 17819 473
rect 17457 455 17508 463
rect 17555 455 17819 469
rect 17863 475 17898 483
rect 17409 407 17428 441
rect 17473 447 17502 455
rect 17473 441 17490 447
rect 17473 439 17507 441
rect 17555 439 17571 455
rect 17572 445 17780 455
rect 17781 445 17797 455
rect 17845 451 17860 466
rect 17863 463 17864 475
rect 17871 463 17898 475
rect 17863 455 17898 463
rect 17863 454 17892 455
rect 17583 441 17797 445
rect 17598 439 17797 441
rect 17832 441 17845 451
rect 17863 441 17880 454
rect 17832 439 17880 441
rect 17474 435 17507 439
rect 17470 433 17507 435
rect 17470 432 17537 433
rect 17470 427 17501 432
rect 17507 427 17537 432
rect 17470 423 17537 427
rect 17443 420 17537 423
rect 17443 413 17492 420
rect 17443 407 17473 413
rect 17492 408 17497 413
rect 17409 391 17489 407
rect 17501 399 17537 420
rect 17598 415 17787 439
rect 17832 438 17879 439
rect 17845 433 17879 438
rect 17613 412 17787 415
rect 17606 409 17787 412
rect 17815 432 17879 433
rect 17409 389 17428 391
rect 17443 389 17477 391
rect 17409 373 17489 389
rect 17409 367 17428 373
rect 17125 341 17228 351
rect 17079 339 17228 341
rect 17249 339 17284 351
rect 16918 337 17080 339
rect 16930 317 16949 337
rect 16964 335 16994 337
rect 16813 309 16854 317
rect 16936 313 16949 317
rect 17001 321 17080 337
rect 17112 337 17284 339
rect 17112 321 17191 337
rect 17198 335 17228 337
rect 16776 299 16805 309
rect 16819 299 16848 309
rect 16863 299 16893 313
rect 16936 299 16979 313
rect 17001 309 17191 321
rect 17256 317 17262 337
rect 16986 299 17016 309
rect 17017 299 17175 309
rect 17179 299 17209 309
rect 17213 299 17243 313
rect 17271 299 17284 337
rect 17356 351 17385 367
rect 17399 351 17428 367
rect 17443 357 17473 373
rect 17501 351 17507 399
rect 17510 393 17529 399
rect 17544 393 17574 401
rect 17510 385 17574 393
rect 17510 369 17590 385
rect 17606 378 17668 409
rect 17684 378 17746 409
rect 17815 407 17864 432
rect 17879 407 17909 423
rect 17778 393 17808 401
rect 17815 399 17925 407
rect 17778 385 17823 393
rect 17510 367 17529 369
rect 17544 367 17590 369
rect 17510 351 17590 367
rect 17617 365 17652 378
rect 17693 375 17730 378
rect 17693 373 17735 375
rect 17622 362 17652 365
rect 17631 358 17638 362
rect 17638 357 17639 358
rect 17597 351 17607 357
rect 17356 343 17391 351
rect 17356 317 17357 343
rect 17364 317 17391 343
rect 17299 299 17329 313
rect 17356 309 17391 317
rect 17393 343 17434 351
rect 17393 317 17408 343
rect 17415 317 17434 343
rect 17498 339 17529 351
rect 17544 339 17647 351
rect 17659 341 17685 367
rect 17700 362 17730 373
rect 17762 369 17824 385
rect 17762 367 17808 369
rect 17762 351 17824 367
rect 17836 351 17842 399
rect 17845 391 17925 399
rect 17845 389 17864 391
rect 17879 389 17913 391
rect 17845 373 17925 389
rect 17845 351 17864 373
rect 17879 357 17909 373
rect 17937 367 17943 441
rect 17946 367 17965 511
rect 17980 367 17986 511
rect 17995 441 18008 511
rect 18060 506 18082 511
rect 18053 485 18082 499
rect 18135 485 18151 499
rect 18189 495 18195 497
rect 18202 495 18310 511
rect 18317 495 18323 497
rect 18331 495 18346 511
rect 18412 505 18431 508
rect 18053 483 18151 485
rect 18178 483 18346 495
rect 18361 485 18377 499
rect 18412 486 18434 505
rect 18444 499 18460 500
rect 18443 497 18460 499
rect 18444 492 18460 497
rect 18434 485 18440 486
rect 18443 485 18472 492
rect 18361 484 18472 485
rect 18361 483 18478 484
rect 18037 475 18088 483
rect 18135 475 18169 483
rect 18037 463 18062 475
rect 18069 463 18088 475
rect 18142 473 18169 475
rect 18178 473 18399 483
rect 18434 480 18440 483
rect 18142 469 18399 473
rect 18037 455 18088 463
rect 18135 455 18399 469
rect 18443 475 18478 483
rect 17989 407 18008 441
rect 18053 447 18082 455
rect 18053 441 18070 447
rect 18053 439 18087 441
rect 18135 439 18151 455
rect 18152 445 18360 455
rect 18361 445 18377 455
rect 18425 451 18440 466
rect 18443 463 18444 475
rect 18451 463 18478 475
rect 18443 455 18478 463
rect 18443 454 18472 455
rect 18163 441 18377 445
rect 18178 439 18377 441
rect 18412 441 18425 451
rect 18443 441 18460 454
rect 18412 439 18460 441
rect 18054 435 18087 439
rect 18050 433 18087 435
rect 18050 432 18117 433
rect 18050 427 18081 432
rect 18087 427 18117 432
rect 18050 423 18117 427
rect 18023 420 18117 423
rect 18023 413 18072 420
rect 18023 407 18053 413
rect 18072 408 18077 413
rect 17989 391 18069 407
rect 18081 399 18117 420
rect 18178 415 18367 439
rect 18412 438 18459 439
rect 18425 433 18459 438
rect 18193 412 18367 415
rect 18186 409 18367 412
rect 18395 432 18459 433
rect 17989 389 18008 391
rect 18023 389 18057 391
rect 17989 373 18069 389
rect 17989 367 18008 373
rect 17705 341 17808 351
rect 17659 339 17808 341
rect 17829 339 17864 351
rect 17498 337 17660 339
rect 17510 317 17529 337
rect 17544 335 17574 337
rect 17393 309 17434 317
rect 17516 313 17529 317
rect 17581 321 17660 337
rect 17692 337 17864 339
rect 17692 321 17771 337
rect 17778 335 17808 337
rect 17356 299 17385 309
rect 17399 299 17428 309
rect 17443 299 17473 313
rect 17516 299 17559 313
rect 17581 309 17771 321
rect 17836 317 17842 337
rect 17566 299 17596 309
rect 17597 299 17755 309
rect 17759 299 17789 309
rect 17793 299 17823 313
rect 17851 299 17864 337
rect 17936 351 17965 367
rect 17979 351 18008 367
rect 18023 357 18053 373
rect 18081 351 18087 399
rect 18090 393 18109 399
rect 18124 393 18154 401
rect 18090 385 18154 393
rect 18090 369 18170 385
rect 18186 378 18248 409
rect 18264 378 18326 409
rect 18395 407 18444 432
rect 18459 407 18489 423
rect 18358 393 18388 401
rect 18395 399 18505 407
rect 18358 385 18403 393
rect 18090 367 18109 369
rect 18124 367 18170 369
rect 18090 351 18170 367
rect 18197 365 18232 378
rect 18273 375 18310 378
rect 18273 373 18315 375
rect 18202 362 18232 365
rect 18211 358 18218 362
rect 18218 357 18219 358
rect 18177 351 18187 357
rect 17936 343 17971 351
rect 17936 317 17937 343
rect 17944 317 17971 343
rect 17879 299 17909 313
rect 17936 309 17971 317
rect 17973 343 18014 351
rect 17973 317 17988 343
rect 17995 317 18014 343
rect 18078 339 18109 351
rect 18124 339 18227 351
rect 18239 341 18265 367
rect 18280 362 18310 373
rect 18342 369 18404 385
rect 18342 367 18388 369
rect 18342 351 18404 367
rect 18416 351 18422 399
rect 18425 391 18505 399
rect 18425 389 18444 391
rect 18459 389 18493 391
rect 18425 373 18505 389
rect 18425 351 18444 373
rect 18459 357 18489 373
rect 18517 367 18523 441
rect 18532 367 18545 511
rect 18285 341 18388 351
rect 18239 339 18388 341
rect 18409 339 18444 351
rect 18078 337 18240 339
rect 18090 317 18109 337
rect 18124 335 18154 337
rect 17973 309 18014 317
rect 18096 313 18109 317
rect 18161 321 18240 337
rect 18272 337 18444 339
rect 18272 321 18351 337
rect 18358 335 18388 337
rect 17936 299 17965 309
rect 17979 299 18008 309
rect 18023 299 18053 313
rect 18096 299 18139 313
rect 18161 309 18351 321
rect 18416 317 18422 337
rect 18146 299 18176 309
rect 18177 299 18335 309
rect 18339 299 18369 309
rect 18373 299 18403 313
rect 18431 299 18444 337
rect 18516 351 18545 367
rect 18516 343 18551 351
rect 18516 317 18517 343
rect 18524 317 18551 343
rect 18459 299 18489 313
rect 18516 309 18551 317
rect 18516 299 18545 309
rect 4596 298 18545 299
rect -1 292 18545 298
rect 0 285 18545 292
rect 0 284 4631 285
rect 15 254 28 284
rect 43 270 73 284
rect 116 270 159 284
rect 166 270 386 284
rect 393 270 423 284
rect 83 256 98 268
rect 117 256 130 270
rect 198 266 351 270
rect 80 254 102 256
rect 180 254 372 266
rect 451 254 464 284
rect 479 270 509 284
rect 546 254 565 284
rect 580 254 586 284
rect 595 254 608 284
rect 623 270 653 284
rect 696 270 739 284
rect 746 270 966 284
rect 973 270 1003 284
rect 663 256 678 268
rect 697 256 710 270
rect 778 266 931 270
rect 660 254 682 256
rect 760 254 952 266
rect 1031 254 1044 284
rect 1059 270 1089 284
rect 1126 254 1145 284
rect 1160 254 1166 284
rect 1175 254 1188 284
rect 1203 270 1233 284
rect 1276 270 1319 284
rect 1326 270 1546 284
rect 1553 270 1583 284
rect 1243 256 1258 268
rect 1277 256 1290 270
rect 1358 266 1511 270
rect 1240 254 1262 256
rect 1340 254 1532 266
rect 1611 254 1624 284
rect 1639 270 1669 284
rect 1706 254 1725 284
rect 1740 254 1746 284
rect 1755 254 1768 284
rect 1783 270 1813 284
rect 1856 270 1899 284
rect 1906 270 2126 284
rect 2133 270 2163 284
rect 1823 256 1838 268
rect 1857 256 1870 270
rect 1938 266 2091 270
rect 1820 254 1842 256
rect 1920 254 2112 266
rect 2191 254 2204 284
rect 2219 270 2249 284
rect 2286 254 2305 284
rect 2320 254 2326 284
rect 2335 254 2348 284
rect 2363 270 2393 284
rect 2436 270 2479 284
rect 2486 270 2706 284
rect 2713 270 2743 284
rect 2403 256 2418 268
rect 2437 256 2450 270
rect 2518 266 2671 270
rect 2400 254 2422 256
rect 2500 254 2692 266
rect 2771 254 2784 284
rect 2799 270 2829 284
rect 2866 254 2885 284
rect 2900 254 2906 284
rect 2915 254 2928 284
rect 2943 270 2973 284
rect 3016 270 3059 284
rect 3066 270 3286 284
rect 3293 270 3323 284
rect 2983 256 2998 268
rect 3017 256 3030 270
rect 3098 266 3251 270
rect 2980 254 3002 256
rect 3080 254 3272 266
rect 3351 254 3364 284
rect 3379 270 3409 284
rect 3446 254 3465 284
rect 3480 254 3486 284
rect 3495 254 3508 284
rect 3523 270 3553 284
rect 3596 270 3639 284
rect 3646 270 3866 284
rect 3873 270 3903 284
rect 3563 256 3578 268
rect 3597 256 3610 270
rect 3678 266 3831 270
rect 3560 254 3582 256
rect 3660 254 3852 266
rect 3931 254 3944 284
rect 3959 270 3989 284
rect 4026 254 4045 284
rect 4060 254 4066 284
rect 4075 254 4088 284
rect 4103 270 4133 284
rect 4176 270 4219 284
rect 4226 270 4446 284
rect 4453 270 4483 284
rect 4143 256 4158 268
rect 4177 256 4190 270
rect 4258 266 4411 270
rect 4140 254 4162 256
rect 4240 254 4432 266
rect 4511 254 4524 284
rect 4539 270 4569 284
rect 4606 271 4625 284
rect 4601 270 4631 271
rect 4606 255 4625 270
rect 4640 255 4646 285
rect 4655 255 4668 285
rect 4683 271 4713 285
rect 4756 271 4799 285
rect 4806 271 5026 285
rect 5033 271 5063 285
rect 4723 257 4738 269
rect 4757 257 4770 271
rect 4838 267 4991 271
rect 4720 255 4742 257
rect 4820 255 5012 267
rect 5091 255 5104 285
rect 5119 271 5149 285
rect 5186 255 5205 285
rect 5220 255 5226 285
rect 5235 255 5248 285
rect 5263 271 5293 285
rect 5336 271 5379 285
rect 5386 271 5606 285
rect 5613 271 5643 285
rect 5303 257 5318 269
rect 5337 257 5350 271
rect 5418 267 5571 271
rect 5300 255 5322 257
rect 5400 255 5592 267
rect 5671 255 5684 285
rect 5699 271 5729 285
rect 5766 255 5785 285
rect 5800 255 5806 285
rect 5815 255 5828 285
rect 5843 271 5873 285
rect 5916 271 5959 285
rect 5966 271 6186 285
rect 6193 271 6223 285
rect 5883 257 5898 269
rect 5917 257 5930 271
rect 5998 267 6151 271
rect 5880 255 5902 257
rect 5980 255 6172 267
rect 6251 255 6264 285
rect 6279 271 6309 285
rect 6346 255 6365 285
rect 6380 255 6386 285
rect 6395 255 6408 285
rect 6423 271 6453 285
rect 6496 271 6539 285
rect 6546 271 6766 285
rect 6773 271 6803 285
rect 6463 257 6478 269
rect 6497 257 6510 271
rect 6578 267 6731 271
rect 6460 255 6482 257
rect 6560 255 6752 267
rect 6831 255 6844 285
rect 6859 271 6889 285
rect 6926 255 6945 285
rect 6960 255 6966 285
rect 6975 255 6988 285
rect 7003 271 7033 285
rect 7076 271 7119 285
rect 7126 271 7346 285
rect 7353 271 7383 285
rect 7043 257 7058 269
rect 7077 257 7090 271
rect 7158 267 7311 271
rect 7040 255 7062 257
rect 7140 255 7332 267
rect 7411 255 7424 285
rect 7439 271 7469 285
rect 7506 255 7525 285
rect 7540 255 7546 285
rect 7555 255 7568 285
rect 7583 271 7613 285
rect 7656 271 7699 285
rect 7706 271 7926 285
rect 7933 271 7963 285
rect 7623 257 7638 269
rect 7657 257 7670 271
rect 7738 267 7891 271
rect 7620 255 7642 257
rect 7720 255 7912 267
rect 7991 255 8004 285
rect 8019 271 8049 285
rect 8086 255 8105 285
rect 8120 255 8126 285
rect 8135 255 8148 285
rect 8163 271 8193 285
rect 8236 271 8279 285
rect 8286 271 8506 285
rect 8513 271 8543 285
rect 8203 257 8218 269
rect 8237 257 8250 271
rect 8318 267 8471 271
rect 8200 255 8222 257
rect 8300 255 8492 267
rect 8571 255 8584 285
rect 8599 271 8629 285
rect 8666 255 8685 285
rect 8700 255 8706 285
rect 8715 255 8728 285
rect 8743 271 8773 285
rect 8816 271 8859 285
rect 8866 271 9086 285
rect 9093 271 9123 285
rect 8783 257 8798 269
rect 8817 257 8830 271
rect 8898 267 9051 271
rect 8780 255 8802 257
rect 8880 255 9072 267
rect 9151 255 9164 285
rect 9179 271 9209 285
rect 9246 255 9265 285
rect 9280 255 9286 285
rect 9295 255 9308 285
rect 9323 271 9353 285
rect 9396 271 9439 285
rect 9446 271 9666 285
rect 9673 271 9703 285
rect 9363 257 9378 269
rect 9397 257 9410 271
rect 9478 267 9631 271
rect 9360 255 9382 257
rect 9460 255 9652 267
rect 9731 255 9744 285
rect 9759 271 9789 285
rect 9826 255 9845 285
rect 9860 255 9866 285
rect 9875 255 9888 285
rect 9903 271 9933 285
rect 9976 271 10019 285
rect 10026 271 10246 285
rect 10253 271 10283 285
rect 9943 257 9958 269
rect 9977 257 9990 271
rect 10058 267 10211 271
rect 9940 255 9962 257
rect 10040 255 10232 267
rect 10311 255 10324 285
rect 10339 271 10369 285
rect 10406 255 10425 285
rect 10440 255 10446 285
rect 10455 255 10468 285
rect 10483 271 10513 285
rect 10556 271 10599 285
rect 10606 271 10826 285
rect 10833 271 10863 285
rect 10523 257 10538 269
rect 10557 257 10570 271
rect 10638 267 10791 271
rect 10520 255 10542 257
rect 10620 255 10812 267
rect 10891 255 10904 285
rect 10919 271 10949 285
rect 10986 255 11005 285
rect 11020 255 11026 285
rect 11035 255 11048 285
rect 11063 271 11093 285
rect 11136 271 11179 285
rect 11186 271 11406 285
rect 11413 271 11443 285
rect 11103 257 11118 269
rect 11137 257 11150 271
rect 11218 267 11371 271
rect 11100 255 11122 257
rect 11200 255 11392 267
rect 11471 255 11484 285
rect 11499 271 11529 285
rect 11566 255 11585 285
rect 11600 255 11606 285
rect 11615 255 11628 285
rect 11643 271 11673 285
rect 11716 271 11759 285
rect 11766 271 11986 285
rect 11993 271 12023 285
rect 11683 257 11698 269
rect 11717 257 11730 271
rect 11798 267 11951 271
rect 11680 255 11702 257
rect 11780 255 11972 267
rect 12051 255 12064 285
rect 12079 271 12109 285
rect 12146 255 12165 285
rect 12180 255 12186 285
rect 12195 255 12208 285
rect 12223 271 12253 285
rect 12296 271 12339 285
rect 12346 271 12566 285
rect 12573 271 12603 285
rect 12263 257 12278 269
rect 12297 257 12310 271
rect 12378 267 12531 271
rect 12260 255 12282 257
rect 12360 255 12552 267
rect 12631 255 12644 285
rect 12659 271 12689 285
rect 12726 255 12745 285
rect 12760 255 12766 285
rect 12775 255 12788 285
rect 12803 271 12833 285
rect 12876 271 12919 285
rect 12926 271 13146 285
rect 13153 271 13183 285
rect 12843 257 12858 269
rect 12877 257 12890 271
rect 12958 267 13111 271
rect 12840 255 12862 257
rect 12940 255 13132 267
rect 13211 255 13224 285
rect 13239 271 13269 285
rect 13306 255 13325 285
rect 13340 255 13346 285
rect 13355 255 13368 285
rect 13383 271 13413 285
rect 13456 271 13499 285
rect 13506 271 13726 285
rect 13733 271 13763 285
rect 13423 257 13438 269
rect 13457 257 13470 271
rect 13538 267 13691 271
rect 13420 255 13442 257
rect 13520 255 13712 267
rect 13791 255 13804 285
rect 13819 271 13849 285
rect 13886 284 13926 285
rect 13886 255 13905 284
rect 13920 255 13926 284
rect 13935 255 13948 285
rect 13963 271 13993 285
rect 14036 271 14079 285
rect 14086 271 14306 285
rect 14313 271 14343 285
rect 14003 257 14018 269
rect 14037 257 14050 271
rect 14118 267 14271 271
rect 14000 255 14022 257
rect 14100 255 14292 267
rect 14371 255 14384 285
rect 14399 271 14429 285
rect 14466 255 14485 285
rect 14500 255 14506 285
rect 14515 255 14528 285
rect 14543 271 14573 285
rect 14616 271 14659 285
rect 14666 271 14886 285
rect 14893 271 14923 285
rect 14583 257 14598 269
rect 14617 257 14630 271
rect 14698 267 14851 271
rect 14580 255 14602 257
rect 14680 255 14872 267
rect 14951 255 14964 285
rect 14979 271 15009 285
rect 15046 255 15065 285
rect 15080 255 15086 285
rect 15095 255 15108 285
rect 15123 271 15153 285
rect 15196 271 15239 285
rect 15246 271 15466 285
rect 15473 271 15503 285
rect 15163 257 15178 269
rect 15197 257 15210 271
rect 15278 267 15431 271
rect 15160 255 15182 257
rect 15260 255 15452 267
rect 15531 255 15544 285
rect 15559 271 15589 285
rect 15626 255 15645 285
rect 15660 255 15666 285
rect 15675 255 15688 285
rect 15703 271 15733 285
rect 15776 271 15819 285
rect 15826 271 16046 285
rect 16053 271 16083 285
rect 15743 257 15758 269
rect 15777 257 15790 271
rect 15858 267 16011 271
rect 15740 255 15762 257
rect 15840 255 16032 267
rect 16111 255 16124 285
rect 16139 271 16169 285
rect 16206 255 16225 285
rect 16240 255 16246 285
rect 16255 255 16268 285
rect 16283 271 16313 285
rect 16356 271 16399 285
rect 16406 271 16626 285
rect 16633 271 16663 285
rect 16323 257 16338 269
rect 16357 257 16370 271
rect 16438 267 16591 271
rect 16320 255 16342 257
rect 16420 255 16612 267
rect 16691 255 16704 285
rect 16719 271 16749 285
rect 16786 255 16805 285
rect 16820 255 16826 285
rect 16835 255 16848 285
rect 16863 271 16893 285
rect 16936 271 16979 285
rect 16986 271 17206 285
rect 17213 271 17243 285
rect 16903 257 16918 269
rect 16937 257 16950 271
rect 17018 267 17171 271
rect 16900 255 16922 257
rect 17000 255 17192 267
rect 17271 255 17284 285
rect 17299 271 17329 285
rect 17366 255 17385 285
rect 17400 255 17406 285
rect 17415 255 17428 285
rect 17443 271 17473 285
rect 17516 271 17559 285
rect 17566 271 17786 285
rect 17793 271 17823 285
rect 17483 257 17498 269
rect 17517 257 17530 271
rect 17598 267 17751 271
rect 17480 255 17502 257
rect 17580 255 17772 267
rect 17851 255 17864 285
rect 17879 271 17909 285
rect 17946 255 17965 285
rect 17980 255 17986 285
rect 17995 255 18008 285
rect 18023 271 18053 285
rect 18096 271 18139 285
rect 18146 271 18366 285
rect 18373 271 18403 285
rect 18063 257 18078 269
rect 18097 257 18110 271
rect 18178 267 18331 271
rect 18060 255 18082 257
rect 18160 255 18352 267
rect 18431 255 18444 285
rect 18459 271 18489 285
rect 18532 255 18545 285
rect 4603 254 18545 255
rect 0 241 18545 254
rect 0 240 4631 241
rect 15 170 28 240
rect 80 236 102 240
rect 73 214 102 228
rect 155 214 171 228
rect 209 218 215 226
rect 222 224 330 240
rect 73 212 171 214
rect 57 204 108 212
rect 155 204 189 212
rect 57 192 82 204
rect 89 192 108 204
rect 162 202 189 204
rect 198 204 215 218
rect 260 204 292 224
rect 337 218 343 226
rect 351 218 366 240
rect 432 234 451 237
rect 337 212 366 218
rect 381 214 397 228
rect 432 215 454 234
rect 464 228 480 229
rect 463 226 480 228
rect 464 221 480 226
rect 454 214 460 215
rect 463 214 492 221
rect 381 213 492 214
rect 381 212 498 213
rect 337 204 419 212
rect 454 209 460 212
rect 198 202 419 204
rect 162 198 234 202
rect 262 200 290 202
rect 57 184 108 192
rect 155 190 287 198
rect 290 190 301 198
rect 155 188 234 190
rect 315 188 419 202
rect 463 204 498 212
rect 155 184 252 188
rect 9 136 28 170
rect 73 176 102 184
rect 73 170 90 176
rect 73 168 107 170
rect 155 168 171 184
rect 172 180 252 184
rect 300 184 419 188
rect 300 180 380 184
rect 172 174 380 180
rect 381 174 397 184
rect 445 180 460 195
rect 463 192 464 204
rect 471 192 498 204
rect 463 184 498 192
rect 463 183 492 184
rect 183 170 293 174
rect 74 164 107 168
rect 70 162 107 164
rect 70 161 137 162
rect 70 156 101 161
rect 107 156 137 161
rect 198 158 213 170
rect 70 152 137 156
rect 43 149 137 152
rect 43 142 92 149
rect 43 136 73 142
rect 92 137 97 142
rect 9 120 89 136
rect 101 128 137 149
rect 222 148 252 157
rect 275 152 293 170
rect 351 168 397 174
rect 432 170 445 180
rect 463 170 480 183
rect 432 168 480 170
rect 313 162 315 164
rect 315 160 317 162
rect 317 157 327 160
rect 300 150 330 157
rect 300 148 331 150
rect 351 148 387 168
rect 432 167 479 168
rect 445 162 479 167
rect 198 144 387 148
rect 213 141 387 144
rect 206 138 387 141
rect 415 161 479 162
rect 9 118 28 120
rect 43 118 77 120
rect 9 102 89 118
rect 9 96 28 102
rect -1 80 28 96
rect 43 86 73 102
rect 101 80 107 128
rect 110 122 129 128
rect 144 122 174 130
rect 110 114 174 122
rect 110 98 190 114
rect 206 107 268 138
rect 284 107 346 138
rect 415 136 464 161
rect 479 136 509 152
rect 378 122 408 130
rect 415 128 525 136
rect 378 114 423 122
rect 217 104 221 107
rect 222 104 252 107
rect 110 96 129 98
rect 144 96 190 98
rect 110 80 190 96
rect 221 94 252 104
rect 293 104 299 107
rect 300 104 330 107
rect 293 102 335 104
rect 222 91 252 94
rect 231 87 238 91
rect 238 86 239 87
rect 197 80 207 86
rect 259 80 275 96
rect 300 91 330 102
rect 362 98 424 114
rect 362 96 408 98
rect 362 80 424 96
rect 436 80 442 128
rect 445 120 525 128
rect 445 118 464 120
rect 479 118 513 120
rect 445 102 525 118
rect 445 80 464 102
rect 479 86 509 102
rect 537 96 543 170
rect 546 96 565 240
rect 580 96 586 240
rect 595 170 608 240
rect 660 236 682 240
rect 653 214 682 228
rect 735 214 751 228
rect 789 218 795 226
rect 802 224 910 240
rect 653 212 751 214
rect 637 204 688 212
rect 735 204 769 212
rect 637 192 662 204
rect 669 192 688 204
rect 742 202 769 204
rect 778 204 795 218
rect 840 204 872 224
rect 917 218 923 226
rect 931 218 946 240
rect 1012 234 1031 237
rect 917 212 946 218
rect 961 214 977 228
rect 1012 215 1034 234
rect 1044 228 1060 229
rect 1043 226 1060 228
rect 1044 221 1060 226
rect 1034 214 1040 215
rect 1043 214 1072 221
rect 961 213 1072 214
rect 961 212 1078 213
rect 917 204 999 212
rect 1034 209 1040 212
rect 778 202 999 204
rect 742 198 814 202
rect 842 200 870 202
rect 637 184 688 192
rect 735 190 867 198
rect 870 190 881 198
rect 735 188 814 190
rect 895 188 999 202
rect 1043 204 1078 212
rect 735 184 832 188
rect 589 136 608 170
rect 653 176 682 184
rect 653 170 670 176
rect 653 168 687 170
rect 735 168 751 184
rect 752 180 832 184
rect 880 184 999 188
rect 880 180 960 184
rect 752 174 960 180
rect 961 174 977 184
rect 1025 180 1040 195
rect 1043 192 1044 204
rect 1051 192 1078 204
rect 1043 184 1078 192
rect 1043 183 1072 184
rect 763 170 873 174
rect 654 164 687 168
rect 650 162 687 164
rect 650 161 717 162
rect 650 156 681 161
rect 687 156 717 161
rect 778 158 793 170
rect 650 152 717 156
rect 623 149 717 152
rect 623 142 672 149
rect 623 136 653 142
rect 672 137 677 142
rect 589 120 669 136
rect 681 128 717 149
rect 802 148 832 157
rect 855 152 873 170
rect 931 168 977 174
rect 1012 170 1025 180
rect 1043 170 1060 183
rect 1012 168 1060 170
rect 893 162 895 164
rect 895 160 897 162
rect 897 157 907 160
rect 880 150 910 157
rect 880 148 911 150
rect 931 148 967 168
rect 1012 167 1059 168
rect 1025 162 1059 167
rect 778 144 967 148
rect 793 141 967 144
rect 786 138 967 141
rect 995 161 1059 162
rect 589 118 608 120
rect 623 118 657 120
rect 589 102 669 118
rect 589 96 608 102
rect -7 72 34 80
rect -7 46 8 72
rect 15 46 34 72
rect 98 68 129 80
rect 144 68 247 80
rect 259 70 285 80
rect 305 70 408 80
rect 259 68 408 70
rect 429 68 464 80
rect 98 66 260 68
rect 110 46 129 66
rect 144 64 174 66
rect -7 38 34 46
rect -1 28 28 38
rect 116 28 129 46
rect 181 50 260 66
rect 292 66 464 68
rect 292 50 371 66
rect 378 64 408 66
rect 181 42 371 50
rect 436 46 442 66
rect 181 38 260 42
rect 262 38 290 42
rect 292 38 371 42
rect 166 28 174 38
rect 193 30 196 38
rect 197 30 215 38
rect 260 30 292 38
rect 337 30 355 38
rect 193 28 359 30
rect 378 28 389 38
rect 451 28 464 66
rect 536 80 565 96
rect 579 80 608 96
rect 623 86 653 102
rect 681 80 687 128
rect 690 122 709 128
rect 724 122 754 130
rect 690 114 754 122
rect 690 98 770 114
rect 786 107 848 138
rect 864 107 926 138
rect 995 136 1044 161
rect 1059 136 1089 152
rect 958 122 988 130
rect 995 128 1105 136
rect 958 114 1003 122
rect 797 104 801 107
rect 802 104 832 107
rect 690 96 709 98
rect 724 96 770 98
rect 690 80 770 96
rect 801 94 832 104
rect 873 104 879 107
rect 880 104 910 107
rect 873 102 915 104
rect 802 91 832 94
rect 811 87 818 91
rect 818 86 819 87
rect 777 80 787 86
rect 839 80 855 96
rect 880 91 910 102
rect 942 98 1004 114
rect 942 96 988 98
rect 942 80 1004 96
rect 1016 80 1022 128
rect 1025 120 1105 128
rect 1025 118 1044 120
rect 1059 118 1093 120
rect 1025 102 1105 118
rect 1025 80 1044 102
rect 1059 86 1089 102
rect 1117 96 1123 170
rect 1126 96 1145 240
rect 1160 96 1166 240
rect 1175 170 1188 240
rect 1240 236 1262 240
rect 1233 214 1262 228
rect 1315 214 1331 228
rect 1369 218 1375 226
rect 1382 224 1490 240
rect 1233 212 1331 214
rect 1217 204 1268 212
rect 1315 204 1349 212
rect 1217 192 1242 204
rect 1249 192 1268 204
rect 1322 202 1349 204
rect 1358 204 1375 218
rect 1420 204 1452 224
rect 1497 218 1503 226
rect 1511 218 1526 240
rect 1592 234 1611 237
rect 1497 212 1526 218
rect 1541 214 1557 228
rect 1592 215 1614 234
rect 1624 228 1640 229
rect 1623 226 1640 228
rect 1624 221 1640 226
rect 1614 214 1620 215
rect 1623 214 1652 221
rect 1541 213 1652 214
rect 1541 212 1658 213
rect 1497 204 1579 212
rect 1614 209 1620 212
rect 1358 202 1579 204
rect 1322 198 1394 202
rect 1422 200 1450 202
rect 1217 184 1268 192
rect 1315 190 1447 198
rect 1450 190 1461 198
rect 1315 188 1394 190
rect 1475 188 1579 202
rect 1623 204 1658 212
rect 1315 184 1412 188
rect 1169 136 1188 170
rect 1233 176 1262 184
rect 1233 170 1250 176
rect 1233 168 1267 170
rect 1315 168 1331 184
rect 1332 180 1412 184
rect 1460 184 1579 188
rect 1460 180 1540 184
rect 1332 174 1540 180
rect 1541 174 1557 184
rect 1605 180 1620 195
rect 1623 192 1624 204
rect 1631 192 1658 204
rect 1623 184 1658 192
rect 1623 183 1652 184
rect 1343 170 1453 174
rect 1234 164 1267 168
rect 1230 162 1267 164
rect 1230 161 1297 162
rect 1230 156 1261 161
rect 1267 156 1297 161
rect 1358 158 1373 170
rect 1230 152 1297 156
rect 1203 149 1297 152
rect 1203 142 1252 149
rect 1203 136 1233 142
rect 1252 137 1257 142
rect 1169 120 1249 136
rect 1261 128 1297 149
rect 1382 148 1412 157
rect 1435 152 1453 170
rect 1511 168 1557 174
rect 1592 170 1605 180
rect 1623 170 1640 183
rect 1592 168 1640 170
rect 1473 162 1475 164
rect 1475 160 1477 162
rect 1477 157 1487 160
rect 1460 150 1490 157
rect 1460 148 1491 150
rect 1511 148 1547 168
rect 1592 167 1639 168
rect 1605 162 1639 167
rect 1358 144 1547 148
rect 1373 141 1547 144
rect 1366 138 1547 141
rect 1575 161 1639 162
rect 1169 118 1188 120
rect 1203 118 1237 120
rect 1169 102 1249 118
rect 1169 96 1188 102
rect 536 72 571 80
rect 536 46 537 72
rect 544 46 571 72
rect 536 38 571 46
rect 573 72 614 80
rect 573 46 588 72
rect 595 46 614 72
rect 678 68 709 80
rect 724 68 827 80
rect 839 70 865 80
rect 885 70 988 80
rect 839 68 988 70
rect 1009 68 1044 80
rect 678 66 840 68
rect 690 46 709 66
rect 724 64 754 66
rect 573 38 614 46
rect 536 28 565 38
rect 579 28 608 38
rect 696 28 709 46
rect 761 50 840 66
rect 872 66 1044 68
rect 872 50 951 66
rect 958 64 988 66
rect 761 42 951 50
rect 1016 46 1022 66
rect 761 38 840 42
rect 842 38 870 42
rect 872 38 951 42
rect 746 28 754 38
rect 773 30 776 38
rect 777 30 795 38
rect 840 30 872 38
rect 917 30 935 38
rect 773 28 939 30
rect 958 28 969 38
rect 1031 28 1044 66
rect 1116 80 1145 96
rect 1159 80 1188 96
rect 1203 86 1233 102
rect 1261 80 1267 128
rect 1270 122 1289 128
rect 1304 122 1334 130
rect 1270 114 1334 122
rect 1270 98 1350 114
rect 1366 107 1428 138
rect 1444 107 1506 138
rect 1575 136 1624 161
rect 1639 136 1669 152
rect 1538 122 1568 130
rect 1575 128 1685 136
rect 1538 114 1583 122
rect 1377 104 1381 107
rect 1382 104 1412 107
rect 1270 96 1289 98
rect 1304 96 1350 98
rect 1270 80 1350 96
rect 1381 94 1412 104
rect 1453 104 1459 107
rect 1460 104 1490 107
rect 1453 102 1495 104
rect 1382 91 1412 94
rect 1391 87 1398 91
rect 1398 86 1399 87
rect 1357 80 1367 86
rect 1419 80 1435 96
rect 1460 91 1490 102
rect 1522 98 1584 114
rect 1522 96 1568 98
rect 1522 80 1584 96
rect 1596 80 1602 128
rect 1605 120 1685 128
rect 1605 118 1624 120
rect 1639 118 1673 120
rect 1605 102 1685 118
rect 1605 80 1624 102
rect 1639 86 1669 102
rect 1697 96 1703 170
rect 1706 96 1725 240
rect 1740 96 1746 240
rect 1755 170 1768 240
rect 1820 236 1842 240
rect 1813 214 1842 228
rect 1895 214 1911 228
rect 1949 218 1955 226
rect 1962 224 2070 240
rect 1813 212 1911 214
rect 1797 204 1848 212
rect 1895 204 1929 212
rect 1797 192 1822 204
rect 1829 192 1848 204
rect 1902 202 1929 204
rect 1938 204 1955 218
rect 2000 204 2032 224
rect 2077 218 2083 226
rect 2091 218 2106 240
rect 2172 234 2191 237
rect 2077 212 2106 218
rect 2121 214 2137 228
rect 2172 215 2194 234
rect 2204 228 2220 229
rect 2203 226 2220 228
rect 2204 221 2220 226
rect 2194 214 2200 215
rect 2203 214 2232 221
rect 2121 213 2232 214
rect 2121 212 2238 213
rect 2077 204 2159 212
rect 2194 209 2200 212
rect 1938 202 2159 204
rect 1902 198 1974 202
rect 2002 200 2030 202
rect 1797 184 1848 192
rect 1895 190 2027 198
rect 2030 190 2041 198
rect 1895 188 1974 190
rect 2055 188 2159 202
rect 2203 204 2238 212
rect 1895 184 1992 188
rect 1749 136 1768 170
rect 1813 176 1842 184
rect 1813 170 1830 176
rect 1813 168 1847 170
rect 1895 168 1911 184
rect 1912 180 1992 184
rect 2040 184 2159 188
rect 2040 180 2120 184
rect 1912 174 2120 180
rect 2121 174 2137 184
rect 2185 180 2200 195
rect 2203 192 2204 204
rect 2211 192 2238 204
rect 2203 184 2238 192
rect 2203 183 2232 184
rect 1923 170 2033 174
rect 1814 164 1847 168
rect 1810 162 1847 164
rect 1810 161 1877 162
rect 1810 156 1841 161
rect 1847 156 1877 161
rect 1938 158 1953 170
rect 1810 152 1877 156
rect 1783 149 1877 152
rect 1783 142 1832 149
rect 1783 136 1813 142
rect 1832 137 1837 142
rect 1749 120 1829 136
rect 1841 128 1877 149
rect 1962 148 1992 157
rect 2015 152 2033 170
rect 2091 168 2137 174
rect 2172 170 2185 180
rect 2203 170 2220 183
rect 2172 168 2220 170
rect 2053 162 2055 164
rect 2055 160 2057 162
rect 2057 157 2067 160
rect 2040 150 2070 157
rect 2040 148 2071 150
rect 2091 148 2127 168
rect 2172 167 2219 168
rect 2185 162 2219 167
rect 1938 144 2127 148
rect 1953 141 2127 144
rect 1946 138 2127 141
rect 2155 161 2219 162
rect 1749 118 1768 120
rect 1783 118 1817 120
rect 1749 102 1829 118
rect 1749 96 1768 102
rect 1116 72 1151 80
rect 1116 46 1117 72
rect 1124 46 1151 72
rect 1116 38 1151 46
rect 1153 72 1194 80
rect 1153 46 1168 72
rect 1175 46 1194 72
rect 1258 68 1289 80
rect 1304 68 1407 80
rect 1419 70 1445 80
rect 1465 70 1568 80
rect 1419 68 1568 70
rect 1589 68 1624 80
rect 1258 66 1420 68
rect 1270 46 1289 66
rect 1304 64 1334 66
rect 1153 38 1194 46
rect 1116 28 1145 38
rect 1159 28 1188 38
rect 1276 28 1289 46
rect 1341 50 1420 66
rect 1452 66 1624 68
rect 1452 50 1531 66
rect 1538 64 1568 66
rect 1341 42 1531 50
rect 1596 46 1602 66
rect 1341 38 1420 42
rect 1422 38 1450 42
rect 1452 38 1531 42
rect 1326 28 1334 38
rect 1353 30 1356 38
rect 1357 30 1375 38
rect 1420 30 1452 38
rect 1497 30 1515 38
rect 1353 28 1519 30
rect 1538 28 1549 38
rect 1611 28 1624 66
rect 1696 80 1725 96
rect 1739 80 1768 96
rect 1783 86 1813 102
rect 1841 80 1847 128
rect 1850 122 1869 128
rect 1884 122 1914 130
rect 1850 114 1914 122
rect 1850 98 1930 114
rect 1946 107 2008 138
rect 2024 107 2086 138
rect 2155 136 2204 161
rect 2219 136 2249 152
rect 2118 122 2148 130
rect 2155 128 2265 136
rect 2118 114 2163 122
rect 1957 104 1961 107
rect 1962 104 1992 107
rect 1850 96 1869 98
rect 1884 96 1930 98
rect 1850 80 1930 96
rect 1961 94 1992 104
rect 2033 104 2039 107
rect 2040 104 2070 107
rect 2033 102 2075 104
rect 1962 91 1992 94
rect 1971 87 1978 91
rect 1978 86 1979 87
rect 1937 80 1947 86
rect 1999 80 2015 96
rect 2040 91 2070 102
rect 2102 98 2164 114
rect 2102 96 2148 98
rect 2102 80 2164 96
rect 2176 80 2182 128
rect 2185 120 2265 128
rect 2185 118 2204 120
rect 2219 118 2253 120
rect 2185 102 2265 118
rect 2185 80 2204 102
rect 2219 86 2249 102
rect 2277 96 2283 170
rect 2286 96 2305 240
rect 2320 96 2326 240
rect 2335 170 2348 240
rect 2400 236 2422 240
rect 2393 214 2422 228
rect 2475 214 2491 228
rect 2529 218 2535 226
rect 2542 224 2650 240
rect 2393 212 2491 214
rect 2377 204 2428 212
rect 2475 204 2509 212
rect 2377 192 2402 204
rect 2409 192 2428 204
rect 2482 202 2509 204
rect 2518 204 2535 218
rect 2580 204 2612 224
rect 2657 218 2663 226
rect 2671 218 2686 240
rect 2752 234 2771 237
rect 2657 212 2686 218
rect 2701 214 2717 228
rect 2752 215 2774 234
rect 2784 228 2800 229
rect 2783 226 2800 228
rect 2784 221 2800 226
rect 2774 214 2780 215
rect 2783 214 2812 221
rect 2701 213 2812 214
rect 2701 212 2818 213
rect 2657 204 2739 212
rect 2774 209 2780 212
rect 2518 202 2739 204
rect 2482 198 2554 202
rect 2582 200 2610 202
rect 2377 184 2428 192
rect 2475 190 2607 198
rect 2610 190 2621 198
rect 2475 188 2554 190
rect 2635 188 2739 202
rect 2783 204 2818 212
rect 2475 184 2572 188
rect 2329 136 2348 170
rect 2393 176 2422 184
rect 2393 170 2410 176
rect 2393 168 2427 170
rect 2475 168 2491 184
rect 2492 180 2572 184
rect 2620 184 2739 188
rect 2620 180 2700 184
rect 2492 174 2700 180
rect 2701 174 2717 184
rect 2765 180 2780 195
rect 2783 192 2784 204
rect 2791 192 2818 204
rect 2783 184 2818 192
rect 2783 183 2812 184
rect 2503 170 2613 174
rect 2394 164 2427 168
rect 2390 162 2427 164
rect 2390 161 2457 162
rect 2390 156 2421 161
rect 2427 156 2457 161
rect 2518 158 2533 170
rect 2390 152 2457 156
rect 2363 149 2457 152
rect 2363 142 2412 149
rect 2363 136 2393 142
rect 2412 137 2417 142
rect 2329 120 2409 136
rect 2421 128 2457 149
rect 2542 148 2572 157
rect 2595 152 2613 170
rect 2671 168 2717 174
rect 2752 170 2765 180
rect 2783 170 2800 183
rect 2752 168 2800 170
rect 2633 162 2635 164
rect 2635 160 2637 162
rect 2637 157 2647 160
rect 2620 150 2650 157
rect 2620 148 2651 150
rect 2671 148 2707 168
rect 2752 167 2799 168
rect 2765 162 2799 167
rect 2518 144 2707 148
rect 2533 141 2707 144
rect 2526 138 2707 141
rect 2735 161 2799 162
rect 2329 118 2348 120
rect 2363 118 2397 120
rect 2329 102 2409 118
rect 2329 96 2348 102
rect 1696 72 1731 80
rect 1696 46 1697 72
rect 1704 46 1731 72
rect 1696 38 1731 46
rect 1733 72 1774 80
rect 1733 46 1748 72
rect 1755 46 1774 72
rect 1838 68 1869 80
rect 1884 68 1987 80
rect 1999 70 2025 80
rect 2045 70 2148 80
rect 1999 68 2148 70
rect 2169 68 2204 80
rect 1838 66 2000 68
rect 1850 46 1869 66
rect 1884 64 1914 66
rect 1733 38 1774 46
rect 1696 28 1725 38
rect 1739 28 1768 38
rect 1856 28 1869 46
rect 1921 50 2000 66
rect 2032 66 2204 68
rect 2032 50 2111 66
rect 2118 64 2148 66
rect 1921 42 2111 50
rect 2176 46 2182 66
rect 1921 38 2000 42
rect 2002 38 2030 42
rect 2032 38 2111 42
rect 1906 28 1914 38
rect 1933 30 1936 38
rect 1937 30 1955 38
rect 2000 30 2032 38
rect 2077 30 2095 38
rect 1933 28 2099 30
rect 2118 28 2129 38
rect 2191 28 2204 66
rect 2276 80 2305 96
rect 2319 80 2348 96
rect 2363 86 2393 102
rect 2421 80 2427 128
rect 2430 122 2449 128
rect 2464 122 2494 130
rect 2430 114 2494 122
rect 2430 98 2510 114
rect 2526 107 2588 138
rect 2604 107 2666 138
rect 2735 136 2784 161
rect 2799 136 2829 152
rect 2698 122 2728 130
rect 2735 128 2845 136
rect 2698 114 2743 122
rect 2537 104 2541 107
rect 2542 104 2572 107
rect 2430 96 2449 98
rect 2464 96 2510 98
rect 2430 80 2510 96
rect 2541 94 2572 104
rect 2613 104 2619 107
rect 2620 104 2650 107
rect 2613 102 2655 104
rect 2542 91 2572 94
rect 2551 87 2558 91
rect 2558 86 2559 87
rect 2517 80 2527 86
rect 2579 80 2595 96
rect 2620 91 2650 102
rect 2682 98 2744 114
rect 2682 96 2728 98
rect 2682 80 2744 96
rect 2756 80 2762 128
rect 2765 120 2845 128
rect 2765 118 2784 120
rect 2799 118 2833 120
rect 2765 102 2845 118
rect 2765 80 2784 102
rect 2799 86 2829 102
rect 2857 96 2863 170
rect 2866 96 2885 240
rect 2900 96 2906 240
rect 2915 170 2928 240
rect 2980 236 3002 240
rect 2973 214 3002 228
rect 3055 214 3071 228
rect 3109 218 3115 226
rect 3122 224 3230 240
rect 2973 212 3071 214
rect 2957 204 3008 212
rect 3055 204 3089 212
rect 2957 192 2982 204
rect 2989 192 3008 204
rect 3062 202 3089 204
rect 3098 204 3115 218
rect 3160 204 3192 224
rect 3237 218 3243 226
rect 3251 218 3266 240
rect 3332 234 3351 237
rect 3237 212 3266 218
rect 3281 214 3297 228
rect 3332 215 3354 234
rect 3364 228 3380 229
rect 3363 226 3380 228
rect 3364 221 3380 226
rect 3354 214 3360 215
rect 3363 214 3392 221
rect 3281 213 3392 214
rect 3281 212 3398 213
rect 3237 204 3319 212
rect 3354 209 3360 212
rect 3098 202 3319 204
rect 3062 198 3134 202
rect 3162 200 3190 202
rect 2957 184 3008 192
rect 3055 190 3187 198
rect 3190 190 3201 198
rect 3055 188 3134 190
rect 3215 188 3319 202
rect 3363 204 3398 212
rect 3055 184 3152 188
rect 2909 136 2928 170
rect 2973 176 3002 184
rect 2973 170 2990 176
rect 2973 168 3007 170
rect 3055 168 3071 184
rect 3072 180 3152 184
rect 3200 184 3319 188
rect 3200 180 3280 184
rect 3072 174 3280 180
rect 3281 174 3297 184
rect 3345 180 3360 195
rect 3363 192 3364 204
rect 3371 192 3398 204
rect 3363 184 3398 192
rect 3363 183 3392 184
rect 3083 170 3193 174
rect 2974 164 3007 168
rect 2970 162 3007 164
rect 2970 161 3037 162
rect 2970 156 3001 161
rect 3007 156 3037 161
rect 3098 158 3113 170
rect 2970 152 3037 156
rect 2943 149 3037 152
rect 2943 142 2992 149
rect 2943 136 2973 142
rect 2992 137 2997 142
rect 2909 120 2989 136
rect 3001 128 3037 149
rect 3122 148 3152 157
rect 3175 152 3193 170
rect 3251 168 3297 174
rect 3332 170 3345 180
rect 3363 170 3380 183
rect 3332 168 3380 170
rect 3213 162 3215 164
rect 3215 160 3217 162
rect 3217 157 3227 160
rect 3200 150 3230 157
rect 3200 148 3231 150
rect 3251 148 3287 168
rect 3332 167 3379 168
rect 3345 162 3379 167
rect 3098 144 3287 148
rect 3113 141 3287 144
rect 3106 138 3287 141
rect 3315 161 3379 162
rect 2909 118 2928 120
rect 2943 118 2977 120
rect 2909 102 2989 118
rect 2909 96 2928 102
rect 2276 72 2311 80
rect 2276 46 2277 72
rect 2284 46 2311 72
rect 2276 38 2311 46
rect 2313 72 2354 80
rect 2313 46 2328 72
rect 2335 46 2354 72
rect 2418 68 2449 80
rect 2464 68 2567 80
rect 2579 70 2605 80
rect 2625 70 2728 80
rect 2579 68 2728 70
rect 2749 68 2784 80
rect 2418 66 2580 68
rect 2430 46 2449 66
rect 2464 64 2494 66
rect 2313 38 2354 46
rect 2276 28 2305 38
rect 2319 28 2348 38
rect 2436 28 2449 46
rect 2501 50 2580 66
rect 2612 66 2784 68
rect 2612 50 2691 66
rect 2698 64 2728 66
rect 2501 42 2691 50
rect 2756 46 2762 66
rect 2501 38 2580 42
rect 2582 38 2610 42
rect 2612 38 2691 42
rect 2486 28 2494 38
rect 2513 30 2516 38
rect 2517 30 2535 38
rect 2580 30 2612 38
rect 2657 30 2675 38
rect 2513 28 2679 30
rect 2698 28 2709 38
rect 2771 28 2784 66
rect 2856 80 2885 96
rect 2899 80 2928 96
rect 2943 86 2973 102
rect 3001 80 3007 128
rect 3010 122 3029 128
rect 3044 122 3074 130
rect 3010 114 3074 122
rect 3010 98 3090 114
rect 3106 107 3168 138
rect 3184 107 3246 138
rect 3315 136 3364 161
rect 3379 136 3409 152
rect 3278 122 3308 130
rect 3315 128 3425 136
rect 3278 114 3323 122
rect 3117 104 3121 107
rect 3122 104 3152 107
rect 3010 96 3029 98
rect 3044 96 3090 98
rect 3010 80 3090 96
rect 3121 94 3152 104
rect 3193 104 3199 107
rect 3200 104 3230 107
rect 3193 102 3235 104
rect 3122 91 3152 94
rect 3131 87 3138 91
rect 3138 86 3139 87
rect 3097 80 3107 86
rect 3159 80 3175 96
rect 3200 91 3230 102
rect 3262 98 3324 114
rect 3262 96 3308 98
rect 3262 80 3324 96
rect 3336 80 3342 128
rect 3345 120 3425 128
rect 3345 118 3364 120
rect 3379 118 3413 120
rect 3345 102 3425 118
rect 3345 80 3364 102
rect 3379 86 3409 102
rect 3437 96 3443 170
rect 3446 96 3465 240
rect 3480 96 3486 240
rect 3495 170 3508 240
rect 3560 236 3582 240
rect 3553 214 3582 228
rect 3635 214 3651 228
rect 3689 218 3695 226
rect 3702 224 3810 240
rect 3553 212 3651 214
rect 3537 204 3588 212
rect 3635 204 3669 212
rect 3537 192 3562 204
rect 3569 192 3588 204
rect 3642 202 3669 204
rect 3678 204 3695 218
rect 3740 204 3772 224
rect 3817 218 3823 226
rect 3831 218 3846 240
rect 3912 234 3931 237
rect 3817 212 3846 218
rect 3861 214 3877 228
rect 3912 215 3934 234
rect 3944 228 3960 229
rect 3943 226 3960 228
rect 3944 221 3960 226
rect 3934 214 3940 215
rect 3943 214 3972 221
rect 3861 213 3972 214
rect 3861 212 3978 213
rect 3817 204 3899 212
rect 3934 209 3940 212
rect 3678 202 3899 204
rect 3642 198 3714 202
rect 3742 200 3770 202
rect 3537 184 3588 192
rect 3635 190 3767 198
rect 3770 190 3781 198
rect 3635 188 3714 190
rect 3795 188 3899 202
rect 3943 204 3978 212
rect 3635 184 3732 188
rect 3489 136 3508 170
rect 3553 176 3582 184
rect 3553 170 3570 176
rect 3553 168 3587 170
rect 3635 168 3651 184
rect 3652 180 3732 184
rect 3780 184 3899 188
rect 3780 180 3860 184
rect 3652 174 3860 180
rect 3861 174 3877 184
rect 3925 180 3940 195
rect 3943 192 3944 204
rect 3951 192 3978 204
rect 3943 184 3978 192
rect 3943 183 3972 184
rect 3663 170 3773 174
rect 3554 164 3587 168
rect 3550 162 3587 164
rect 3550 161 3617 162
rect 3550 156 3581 161
rect 3587 156 3617 161
rect 3678 158 3693 170
rect 3550 152 3617 156
rect 3523 149 3617 152
rect 3523 142 3572 149
rect 3523 136 3553 142
rect 3572 137 3577 142
rect 3489 120 3569 136
rect 3581 128 3617 149
rect 3702 148 3732 157
rect 3755 152 3773 170
rect 3831 168 3877 174
rect 3912 170 3925 180
rect 3943 170 3960 183
rect 3912 168 3960 170
rect 3793 162 3795 164
rect 3795 160 3797 162
rect 3797 157 3807 160
rect 3780 150 3810 157
rect 3780 148 3811 150
rect 3831 148 3867 168
rect 3912 167 3959 168
rect 3925 162 3959 167
rect 3678 144 3867 148
rect 3693 141 3867 144
rect 3686 138 3867 141
rect 3895 161 3959 162
rect 3489 118 3508 120
rect 3523 118 3557 120
rect 3489 102 3569 118
rect 3489 96 3508 102
rect 2856 72 2891 80
rect 2856 46 2857 72
rect 2864 46 2891 72
rect 2856 38 2891 46
rect 2893 72 2934 80
rect 2893 46 2908 72
rect 2915 46 2934 72
rect 2998 68 3029 80
rect 3044 68 3147 80
rect 3159 70 3185 80
rect 3205 70 3308 80
rect 3159 68 3308 70
rect 3329 68 3364 80
rect 2998 66 3160 68
rect 3010 46 3029 66
rect 3044 64 3074 66
rect 2893 38 2934 46
rect 2856 28 2885 38
rect 2899 28 2928 38
rect 3016 28 3029 46
rect 3081 50 3160 66
rect 3192 66 3364 68
rect 3192 50 3271 66
rect 3278 64 3308 66
rect 3081 42 3271 50
rect 3336 46 3342 66
rect 3081 38 3160 42
rect 3162 38 3190 42
rect 3192 38 3271 42
rect 3066 28 3074 38
rect 3093 30 3096 38
rect 3097 30 3115 38
rect 3160 30 3192 38
rect 3237 30 3255 38
rect 3093 28 3259 30
rect 3278 28 3289 38
rect 3351 28 3364 66
rect 3436 80 3465 96
rect 3479 80 3508 96
rect 3523 86 3553 102
rect 3581 80 3587 128
rect 3590 122 3609 128
rect 3624 122 3654 130
rect 3590 114 3654 122
rect 3590 98 3670 114
rect 3686 107 3748 138
rect 3764 107 3826 138
rect 3895 136 3944 161
rect 3959 136 3989 152
rect 3858 122 3888 130
rect 3895 128 4005 136
rect 3858 114 3903 122
rect 3697 104 3701 107
rect 3702 104 3732 107
rect 3590 96 3609 98
rect 3624 96 3670 98
rect 3590 80 3670 96
rect 3701 94 3732 104
rect 3773 104 3779 107
rect 3780 104 3810 107
rect 3773 102 3815 104
rect 3702 91 3732 94
rect 3711 87 3718 91
rect 3718 86 3719 87
rect 3677 80 3687 86
rect 3739 80 3755 96
rect 3780 91 3810 102
rect 3842 98 3904 114
rect 3842 96 3888 98
rect 3842 80 3904 96
rect 3916 80 3922 128
rect 3925 120 4005 128
rect 3925 118 3944 120
rect 3959 118 3993 120
rect 3925 102 4005 118
rect 3925 80 3944 102
rect 3959 86 3989 102
rect 4017 96 4023 170
rect 4026 96 4045 240
rect 4060 96 4066 240
rect 4075 170 4088 240
rect 4140 236 4162 240
rect 4133 214 4162 228
rect 4215 214 4231 228
rect 4269 218 4275 226
rect 4282 224 4390 240
rect 4133 212 4231 214
rect 4117 204 4168 212
rect 4215 204 4249 212
rect 4117 192 4142 204
rect 4149 192 4168 204
rect 4222 202 4249 204
rect 4258 204 4275 218
rect 4320 204 4352 224
rect 4397 218 4403 226
rect 4411 218 4426 240
rect 4492 234 4511 237
rect 4397 212 4426 218
rect 4441 214 4457 228
rect 4492 215 4514 234
rect 4524 228 4540 229
rect 4523 226 4540 228
rect 4524 221 4540 226
rect 4514 214 4520 215
rect 4523 214 4552 221
rect 4441 213 4552 214
rect 4441 212 4558 213
rect 4397 204 4479 212
rect 4514 209 4520 212
rect 4258 202 4479 204
rect 4222 198 4294 202
rect 4322 200 4350 202
rect 4117 184 4168 192
rect 4215 190 4347 198
rect 4350 190 4361 198
rect 4215 188 4294 190
rect 4375 188 4479 202
rect 4523 204 4558 212
rect 4215 184 4312 188
rect 4069 136 4088 170
rect 4133 176 4162 184
rect 4133 170 4150 176
rect 4133 168 4167 170
rect 4215 168 4231 184
rect 4232 180 4312 184
rect 4360 184 4479 188
rect 4360 180 4440 184
rect 4232 174 4440 180
rect 4441 174 4457 184
rect 4505 180 4520 195
rect 4523 192 4524 204
rect 4531 192 4558 204
rect 4523 184 4558 192
rect 4523 183 4552 184
rect 4243 170 4353 174
rect 4134 164 4167 168
rect 4130 162 4167 164
rect 4130 161 4197 162
rect 4130 156 4161 161
rect 4167 156 4197 161
rect 4258 158 4273 170
rect 4130 152 4197 156
rect 4103 149 4197 152
rect 4103 142 4152 149
rect 4103 136 4133 142
rect 4152 137 4157 142
rect 4069 120 4149 136
rect 4161 128 4197 149
rect 4282 148 4312 157
rect 4335 152 4353 170
rect 4411 168 4457 174
rect 4492 170 4505 180
rect 4523 170 4540 183
rect 4492 168 4540 170
rect 4373 162 4375 164
rect 4375 160 4377 162
rect 4377 157 4387 160
rect 4360 150 4390 157
rect 4360 148 4391 150
rect 4411 148 4447 168
rect 4492 167 4539 168
rect 4505 162 4539 167
rect 4258 144 4447 148
rect 4273 141 4447 144
rect 4266 138 4447 141
rect 4475 161 4539 162
rect 4069 118 4088 120
rect 4103 118 4137 120
rect 4069 102 4149 118
rect 4069 96 4088 102
rect 3436 72 3471 80
rect 3436 46 3437 72
rect 3444 46 3471 72
rect 3436 38 3471 46
rect 3473 72 3514 80
rect 3473 46 3488 72
rect 3495 46 3514 72
rect 3578 68 3609 80
rect 3624 68 3727 80
rect 3739 70 3765 80
rect 3785 70 3888 80
rect 3739 68 3888 70
rect 3909 68 3944 80
rect 3578 66 3740 68
rect 3590 46 3609 66
rect 3624 64 3654 66
rect 3473 38 3514 46
rect 3436 28 3465 38
rect 3479 28 3508 38
rect 3596 28 3609 46
rect 3661 50 3740 66
rect 3772 66 3944 68
rect 3772 50 3851 66
rect 3858 64 3888 66
rect 3661 42 3851 50
rect 3916 46 3922 66
rect 3661 38 3740 42
rect 3742 38 3770 42
rect 3772 38 3851 42
rect 3646 28 3654 38
rect 3673 30 3676 38
rect 3677 30 3695 38
rect 3740 30 3772 38
rect 3817 30 3835 38
rect 3673 28 3839 30
rect 3858 28 3869 38
rect 3931 28 3944 66
rect 4016 80 4045 96
rect 4059 80 4088 96
rect 4103 86 4133 102
rect 4161 80 4167 128
rect 4170 122 4189 128
rect 4204 122 4234 130
rect 4170 114 4234 122
rect 4170 98 4250 114
rect 4266 107 4328 138
rect 4344 107 4406 138
rect 4475 136 4524 161
rect 4539 136 4569 152
rect 4438 122 4468 130
rect 4475 128 4585 136
rect 4438 114 4483 122
rect 4277 104 4281 107
rect 4282 104 4312 107
rect 4170 96 4189 98
rect 4204 96 4250 98
rect 4170 80 4250 96
rect 4281 94 4312 104
rect 4353 104 4359 107
rect 4360 104 4390 107
rect 4353 102 4395 104
rect 4282 91 4312 94
rect 4291 87 4298 91
rect 4298 86 4299 87
rect 4257 80 4267 86
rect 4319 80 4335 96
rect 4360 91 4390 102
rect 4422 98 4484 114
rect 4422 96 4468 98
rect 4422 80 4484 96
rect 4496 80 4502 128
rect 4505 120 4585 128
rect 4505 118 4524 120
rect 4539 118 4573 120
rect 4505 102 4585 118
rect 4505 80 4524 102
rect 4539 86 4569 102
rect 4597 96 4603 170
rect 4606 96 4625 240
rect 4640 97 4646 241
rect 4655 171 4668 241
rect 4720 237 4742 241
rect 4713 215 4742 229
rect 4795 215 4811 229
rect 4849 219 4855 227
rect 4862 225 4970 241
rect 4713 213 4811 215
rect 4697 205 4748 213
rect 4795 205 4829 213
rect 4697 193 4722 205
rect 4729 193 4748 205
rect 4802 203 4829 205
rect 4838 205 4855 219
rect 4900 205 4932 225
rect 4977 219 4983 227
rect 4991 219 5006 241
rect 5072 235 5091 238
rect 4977 213 5006 219
rect 5021 215 5037 229
rect 5072 216 5094 235
rect 5104 229 5120 230
rect 5103 227 5120 229
rect 5104 222 5120 227
rect 5094 215 5100 216
rect 5103 215 5132 222
rect 5021 214 5132 215
rect 5021 213 5138 214
rect 4977 205 5059 213
rect 5094 210 5100 213
rect 4838 203 5059 205
rect 4802 199 4874 203
rect 4902 201 4930 203
rect 4697 185 4748 193
rect 4795 191 4927 199
rect 4930 191 4942 199
rect 4795 189 4874 191
rect 4955 189 5059 203
rect 4795 185 4892 189
rect 4649 137 4668 171
rect 4713 177 4742 185
rect 4713 171 4730 177
rect 4713 169 4747 171
rect 4795 169 4811 185
rect 4812 181 4892 185
rect 4940 185 5059 189
rect 4940 181 5020 185
rect 4812 175 5020 181
rect 5021 175 5037 185
rect 5085 181 5100 196
rect 5103 184 5138 213
rect 4823 171 4933 175
rect 4714 165 4747 169
rect 4710 163 4747 165
rect 4710 162 4777 163
rect 4710 157 4741 162
rect 4747 157 4777 162
rect 4838 159 4853 171
rect 4710 153 4777 157
rect 4683 150 4777 153
rect 4683 143 4732 150
rect 4683 137 4713 143
rect 4732 138 4737 143
rect 4649 121 4729 137
rect 4741 129 4777 150
rect 4862 149 4892 158
rect 4915 153 4933 171
rect 4991 169 5037 175
rect 5072 171 5085 181
rect 5103 171 5120 184
rect 4953 163 4955 165
rect 4955 160 4958 163
rect 4958 158 4967 160
rect 4940 151 4970 158
rect 4940 149 4971 151
rect 4991 149 5027 169
rect 5072 168 5120 171
rect 5085 163 5119 168
rect 4838 145 5027 149
rect 4853 142 5027 145
rect 4846 139 5027 142
rect 5055 162 5119 163
rect 4649 119 4668 121
rect 4683 119 4717 121
rect 4649 103 4729 119
rect 4649 97 4668 103
rect 4016 72 4051 80
rect 4016 46 4017 72
rect 4024 46 4051 72
rect 4016 38 4051 46
rect 4053 72 4094 80
rect 4053 46 4068 72
rect 4075 46 4094 72
rect 4158 68 4189 80
rect 4204 68 4307 80
rect 4319 70 4345 80
rect 4365 70 4468 80
rect 4319 68 4468 70
rect 4489 68 4524 80
rect 4158 66 4320 68
rect 4170 46 4189 66
rect 4204 64 4234 66
rect 4053 38 4094 46
rect 4016 28 4045 38
rect 4059 28 4088 38
rect 4176 28 4189 46
rect 4241 50 4320 66
rect 4352 66 4524 68
rect 4352 50 4431 66
rect 4438 64 4468 66
rect 4241 42 4431 50
rect 4496 46 4502 66
rect 4241 38 4320 42
rect 4322 38 4350 42
rect 4352 38 4431 42
rect 4226 28 4234 38
rect 4253 30 4256 38
rect 4257 30 4275 38
rect 4320 30 4352 38
rect 4397 30 4415 38
rect 4253 28 4419 30
rect 4438 28 4449 38
rect 4511 28 4524 66
rect 4596 80 4625 96
rect 4639 81 4668 97
rect 4683 87 4713 103
rect 4741 81 4747 129
rect 4750 123 4769 129
rect 4784 123 4814 131
rect 4750 115 4814 123
rect 4750 99 4830 115
rect 4846 108 4908 139
rect 4924 108 4986 139
rect 5055 137 5104 162
rect 5119 137 5149 153
rect 5018 123 5048 131
rect 5055 129 5165 137
rect 5018 115 5063 123
rect 4857 104 4892 108
rect 4750 97 4769 99
rect 4784 97 4830 99
rect 4750 81 4830 97
rect 4862 92 4892 104
rect 4933 105 4970 108
rect 4933 103 4975 105
rect 4871 88 4878 92
rect 4878 87 4879 88
rect 4837 81 4847 87
rect 4596 72 4631 80
rect 4596 46 4597 72
rect 4604 46 4631 72
rect 4596 38 4631 46
rect 4633 73 4674 81
rect 4633 47 4648 73
rect 4655 47 4674 73
rect 4738 69 4769 81
rect 4784 69 4887 81
rect 4899 80 4916 97
rect 4940 92 4970 103
rect 5002 99 5064 115
rect 5002 97 5048 99
rect 5002 81 5064 97
rect 5076 81 5082 129
rect 5085 121 5165 129
rect 5085 119 5104 121
rect 5119 119 5153 121
rect 5085 103 5165 119
rect 5085 81 5104 103
rect 5119 87 5149 103
rect 5177 97 5183 171
rect 5186 97 5205 241
rect 5220 97 5226 241
rect 5235 171 5248 241
rect 5300 237 5322 241
rect 5293 215 5322 229
rect 5375 215 5391 229
rect 5429 219 5435 227
rect 5442 225 5550 241
rect 5279 213 5391 215
rect 5277 185 5328 213
rect 5375 205 5409 213
rect 5382 203 5409 205
rect 5418 205 5435 219
rect 5480 205 5512 225
rect 5557 219 5563 227
rect 5571 219 5586 241
rect 5652 235 5671 238
rect 5557 213 5586 219
rect 5601 215 5617 229
rect 5652 216 5674 235
rect 5684 229 5700 230
rect 5683 227 5700 229
rect 5684 222 5700 227
rect 5674 215 5680 216
rect 5683 215 5712 222
rect 5601 214 5712 215
rect 5601 213 5718 214
rect 5557 205 5639 213
rect 5674 210 5680 213
rect 5418 203 5639 205
rect 5382 199 5454 203
rect 5482 201 5510 203
rect 5229 137 5248 171
rect 5293 184 5328 185
rect 5375 191 5507 199
rect 5510 191 5522 199
rect 5375 189 5454 191
rect 5535 189 5639 203
rect 5375 185 5472 189
rect 5293 177 5322 184
rect 5293 171 5310 177
rect 5293 168 5327 171
rect 5375 169 5391 185
rect 5392 181 5472 185
rect 5520 185 5639 189
rect 5520 181 5600 185
rect 5392 175 5600 181
rect 5601 175 5617 185
rect 5665 181 5680 196
rect 5683 184 5718 213
rect 5403 171 5513 175
rect 5294 165 5327 168
rect 5290 163 5327 165
rect 5290 162 5357 163
rect 5290 157 5321 162
rect 5327 157 5357 162
rect 5418 159 5433 171
rect 5290 153 5357 157
rect 5263 150 5357 153
rect 5263 143 5312 150
rect 5263 137 5293 143
rect 5312 138 5317 143
rect 5229 121 5309 137
rect 5321 129 5357 150
rect 5442 149 5472 158
rect 5495 153 5513 171
rect 5571 169 5617 175
rect 5652 171 5665 181
rect 5683 171 5700 184
rect 5533 163 5535 165
rect 5535 160 5538 163
rect 5538 158 5547 160
rect 5520 151 5550 158
rect 5520 149 5551 151
rect 5571 149 5607 169
rect 5652 168 5700 171
rect 5665 163 5699 168
rect 5418 145 5607 149
rect 5433 142 5607 145
rect 5426 139 5607 142
rect 5635 162 5699 163
rect 5229 119 5248 121
rect 5263 119 5297 121
rect 5229 103 5309 119
rect 5229 97 5248 103
rect 4899 71 4925 80
rect 4945 71 5048 81
rect 4899 69 5048 71
rect 5069 69 5104 81
rect 4738 67 4900 69
rect 4750 47 4769 67
rect 4784 65 4814 67
rect 4633 39 4674 47
rect 4596 29 4625 38
rect 4639 29 4668 39
rect 4756 29 4769 47
rect 4821 51 4900 67
rect 4932 67 5104 69
rect 4932 51 5011 67
rect 5018 65 5048 67
rect 4821 43 5011 51
rect 5076 47 5082 67
rect 4821 39 4900 43
rect 4902 39 4930 43
rect 4932 39 5011 43
rect 4806 29 4814 39
rect 4833 31 4836 39
rect 4837 31 4855 39
rect 4900 31 4932 39
rect 4977 31 4995 39
rect 4833 29 4999 31
rect 5018 29 5029 39
rect 5091 29 5104 67
rect 5176 81 5205 97
rect 5219 81 5248 97
rect 5263 87 5293 103
rect 5321 81 5327 129
rect 5330 123 5349 129
rect 5364 123 5394 131
rect 5330 115 5394 123
rect 5330 99 5410 115
rect 5426 108 5488 139
rect 5504 108 5566 139
rect 5635 137 5684 162
rect 5699 137 5729 153
rect 5598 123 5628 131
rect 5635 129 5745 137
rect 5598 115 5643 123
rect 5437 104 5472 108
rect 5330 97 5349 99
rect 5364 97 5410 99
rect 5330 81 5410 97
rect 5442 92 5472 104
rect 5513 105 5550 108
rect 5513 103 5555 105
rect 5451 88 5458 92
rect 5458 87 5459 88
rect 5417 81 5427 87
rect 5176 69 5211 81
rect 5213 69 5254 81
rect 5176 39 5254 69
rect 5318 69 5349 81
rect 5364 69 5467 81
rect 5479 80 5496 97
rect 5520 92 5550 103
rect 5582 99 5644 115
rect 5582 97 5628 99
rect 5582 81 5644 97
rect 5656 81 5662 129
rect 5665 121 5745 129
rect 5665 119 5684 121
rect 5699 119 5733 121
rect 5665 103 5745 119
rect 5665 81 5684 103
rect 5699 87 5729 103
rect 5757 97 5763 171
rect 5766 97 5785 241
rect 5800 97 5806 241
rect 5815 171 5828 241
rect 5880 237 5902 241
rect 5873 215 5902 229
rect 5955 215 5971 229
rect 6009 219 6015 227
rect 6022 225 6130 241
rect 5859 213 5971 215
rect 5857 185 5908 213
rect 5955 205 5989 213
rect 5962 203 5989 205
rect 5998 205 6015 219
rect 6060 205 6092 225
rect 6137 219 6143 227
rect 6151 219 6166 241
rect 6232 235 6251 238
rect 6137 213 6166 219
rect 6181 215 6197 229
rect 6232 216 6254 235
rect 6264 229 6280 230
rect 6263 227 6280 229
rect 6264 222 6280 227
rect 6254 215 6260 216
rect 6263 215 6292 222
rect 6181 214 6292 215
rect 6181 213 6298 214
rect 6137 205 6219 213
rect 6254 210 6260 213
rect 5998 203 6219 205
rect 5962 199 6034 203
rect 6062 201 6090 203
rect 5809 137 5828 171
rect 5873 184 5908 185
rect 5955 191 6087 199
rect 6090 191 6102 199
rect 5955 189 6034 191
rect 6115 189 6219 203
rect 5955 185 6052 189
rect 5873 177 5902 184
rect 5873 171 5890 177
rect 5873 168 5907 171
rect 5955 169 5971 185
rect 5972 181 6052 185
rect 6100 185 6219 189
rect 6100 181 6180 185
rect 5972 175 6180 181
rect 6181 175 6197 185
rect 6245 181 6260 196
rect 6263 184 6298 213
rect 5983 171 6093 175
rect 5874 165 5907 168
rect 5870 163 5907 165
rect 5870 162 5937 163
rect 5870 157 5901 162
rect 5907 157 5937 162
rect 5998 159 6013 171
rect 5870 153 5937 157
rect 5843 150 5937 153
rect 5843 143 5892 150
rect 5843 137 5873 143
rect 5892 138 5897 143
rect 5809 121 5889 137
rect 5901 129 5937 150
rect 6022 149 6052 158
rect 6075 153 6093 171
rect 6151 169 6197 175
rect 6232 171 6245 181
rect 6263 171 6280 184
rect 6113 163 6115 165
rect 6115 160 6118 163
rect 6118 158 6127 160
rect 6100 151 6130 158
rect 6100 149 6131 151
rect 6151 149 6187 169
rect 6232 168 6280 171
rect 6245 163 6279 168
rect 5998 145 6187 149
rect 6013 142 6187 145
rect 6006 139 6187 142
rect 6215 162 6279 163
rect 5809 119 5828 121
rect 5843 119 5877 121
rect 5809 103 5889 119
rect 5809 97 5828 103
rect 5479 71 5505 80
rect 5525 71 5628 81
rect 5479 69 5628 71
rect 5649 69 5684 81
rect 5318 67 5480 69
rect 5330 47 5349 67
rect 5364 65 5394 67
rect 5176 38 5211 39
rect 5219 38 5254 39
rect 5176 29 5205 38
rect 5219 29 5248 38
rect 5336 29 5349 47
rect 5401 51 5480 67
rect 5512 67 5684 69
rect 5512 51 5591 67
rect 5598 65 5628 67
rect 5401 43 5591 51
rect 5656 47 5662 67
rect 5401 39 5480 43
rect 5482 39 5510 43
rect 5512 39 5591 43
rect 5386 29 5394 39
rect 5413 31 5416 39
rect 5417 31 5435 39
rect 5480 31 5512 39
rect 5557 31 5575 39
rect 5413 29 5579 31
rect 5598 29 5609 39
rect 5671 29 5684 67
rect 5756 81 5785 97
rect 5799 81 5828 97
rect 5843 87 5873 103
rect 5901 81 5907 129
rect 5910 123 5929 129
rect 5944 123 5974 131
rect 5910 115 5974 123
rect 5910 99 5990 115
rect 6006 108 6068 139
rect 6084 108 6146 139
rect 6215 137 6264 162
rect 6279 137 6309 153
rect 6178 123 6208 131
rect 6215 129 6325 137
rect 6178 115 6223 123
rect 6017 104 6052 108
rect 5910 97 5929 99
rect 5944 97 5990 99
rect 5910 81 5990 97
rect 6022 92 6052 104
rect 6093 105 6130 108
rect 6093 103 6135 105
rect 6031 88 6038 92
rect 6038 87 6039 88
rect 5997 81 6007 87
rect 5756 69 5791 81
rect 5793 69 5834 81
rect 5756 39 5834 69
rect 5898 69 5929 81
rect 5944 69 6047 81
rect 6059 80 6076 97
rect 6100 92 6130 103
rect 6162 99 6224 115
rect 6162 97 6208 99
rect 6162 81 6224 97
rect 6236 81 6242 129
rect 6245 121 6325 129
rect 6245 119 6264 121
rect 6279 119 6313 121
rect 6245 103 6325 119
rect 6245 81 6264 103
rect 6279 87 6309 103
rect 6337 97 6343 171
rect 6346 97 6365 241
rect 6380 97 6386 241
rect 6395 171 6408 241
rect 6460 237 6482 241
rect 6453 215 6482 229
rect 6535 215 6551 229
rect 6589 219 6595 227
rect 6602 225 6710 241
rect 6439 213 6551 215
rect 6437 185 6488 213
rect 6535 205 6569 213
rect 6542 203 6569 205
rect 6578 205 6595 219
rect 6640 205 6672 225
rect 6717 219 6723 227
rect 6731 219 6746 241
rect 6812 235 6831 238
rect 6717 213 6746 219
rect 6761 215 6777 229
rect 6812 216 6834 235
rect 6844 229 6860 230
rect 6843 227 6860 229
rect 6844 222 6860 227
rect 6834 215 6840 216
rect 6843 215 6872 222
rect 6761 214 6872 215
rect 6761 213 6878 214
rect 6717 205 6799 213
rect 6834 210 6840 213
rect 6578 203 6799 205
rect 6542 199 6614 203
rect 6642 201 6670 203
rect 6389 137 6408 171
rect 6453 184 6488 185
rect 6535 191 6667 199
rect 6670 191 6682 199
rect 6535 189 6614 191
rect 6695 189 6799 203
rect 6535 185 6632 189
rect 6453 177 6482 184
rect 6453 171 6470 177
rect 6453 168 6487 171
rect 6535 169 6551 185
rect 6552 181 6632 185
rect 6680 185 6799 189
rect 6680 181 6760 185
rect 6552 175 6760 181
rect 6761 175 6777 185
rect 6825 181 6840 196
rect 6843 184 6878 213
rect 6563 171 6673 175
rect 6454 165 6487 168
rect 6450 163 6487 165
rect 6450 162 6517 163
rect 6450 157 6481 162
rect 6487 157 6517 162
rect 6578 159 6593 171
rect 6450 153 6517 157
rect 6423 150 6517 153
rect 6423 143 6472 150
rect 6423 137 6453 143
rect 6472 138 6477 143
rect 6389 121 6469 137
rect 6481 129 6517 150
rect 6602 149 6632 158
rect 6655 153 6673 171
rect 6731 169 6777 175
rect 6812 171 6825 181
rect 6843 171 6860 184
rect 6693 163 6695 165
rect 6695 160 6698 163
rect 6698 158 6707 160
rect 6680 151 6710 158
rect 6680 149 6711 151
rect 6731 149 6767 169
rect 6812 168 6860 171
rect 6825 163 6859 168
rect 6578 145 6767 149
rect 6593 142 6767 145
rect 6586 139 6767 142
rect 6795 162 6859 163
rect 6389 119 6408 121
rect 6423 119 6457 121
rect 6389 103 6469 119
rect 6389 97 6408 103
rect 6059 71 6085 80
rect 6105 71 6208 81
rect 6059 69 6208 71
rect 6229 69 6264 81
rect 5898 67 6060 69
rect 5910 47 5929 67
rect 5944 65 5974 67
rect 5756 38 5791 39
rect 5799 38 5834 39
rect 5756 29 5785 38
rect 5799 29 5828 38
rect 5916 29 5929 47
rect 5981 51 6060 67
rect 6092 67 6264 69
rect 6092 51 6171 67
rect 6178 65 6208 67
rect 5981 43 6171 51
rect 6236 47 6242 67
rect 5981 39 6060 43
rect 6062 39 6090 43
rect 6092 39 6171 43
rect 5966 29 5974 39
rect 5993 31 5996 39
rect 5997 31 6015 39
rect 6060 31 6092 39
rect 6137 31 6155 39
rect 5993 29 6159 31
rect 6178 29 6189 39
rect 6251 29 6264 67
rect 6336 81 6365 97
rect 6379 81 6408 97
rect 6423 87 6453 103
rect 6481 81 6487 129
rect 6490 123 6509 129
rect 6524 123 6554 131
rect 6490 115 6554 123
rect 6490 99 6570 115
rect 6586 108 6648 139
rect 6664 108 6726 139
rect 6795 137 6844 162
rect 6859 137 6889 153
rect 6758 123 6788 131
rect 6795 129 6905 137
rect 6758 115 6803 123
rect 6597 104 6632 108
rect 6490 97 6509 99
rect 6524 97 6570 99
rect 6490 81 6570 97
rect 6602 92 6632 104
rect 6673 105 6710 108
rect 6673 103 6715 105
rect 6611 88 6618 92
rect 6618 87 6619 88
rect 6577 81 6587 87
rect 6336 69 6371 81
rect 6373 69 6414 81
rect 6336 39 6414 69
rect 6478 69 6509 81
rect 6524 69 6627 81
rect 6639 80 6656 97
rect 6680 92 6710 103
rect 6742 99 6804 115
rect 6742 97 6788 99
rect 6742 81 6804 97
rect 6816 81 6822 129
rect 6825 121 6905 129
rect 6825 119 6844 121
rect 6859 119 6893 121
rect 6825 103 6905 119
rect 6825 81 6844 103
rect 6859 87 6889 103
rect 6917 97 6923 171
rect 6926 97 6945 241
rect 6960 97 6966 241
rect 6975 171 6988 241
rect 7040 237 7062 241
rect 7033 215 7062 229
rect 7115 215 7131 229
rect 7169 219 7175 227
rect 7182 225 7290 241
rect 7019 213 7131 215
rect 7017 185 7068 213
rect 7115 205 7149 213
rect 7122 203 7149 205
rect 7158 205 7175 219
rect 7220 205 7252 225
rect 7297 219 7303 227
rect 7311 219 7326 241
rect 7392 235 7411 238
rect 7297 213 7326 219
rect 7341 215 7357 229
rect 7392 216 7414 235
rect 7424 229 7440 230
rect 7423 227 7440 229
rect 7424 222 7440 227
rect 7414 215 7420 216
rect 7423 215 7452 222
rect 7341 214 7452 215
rect 7341 213 7458 214
rect 7297 205 7379 213
rect 7414 210 7420 213
rect 7158 203 7379 205
rect 7122 199 7194 203
rect 7222 201 7250 203
rect 6969 137 6988 171
rect 7033 184 7068 185
rect 7115 191 7247 199
rect 7250 191 7262 199
rect 7115 189 7194 191
rect 7275 189 7379 203
rect 7115 185 7212 189
rect 7033 177 7062 184
rect 7033 171 7050 177
rect 7033 168 7067 171
rect 7115 169 7131 185
rect 7132 181 7212 185
rect 7260 185 7379 189
rect 7260 181 7340 185
rect 7132 175 7340 181
rect 7341 175 7357 185
rect 7405 181 7420 196
rect 7423 184 7458 213
rect 7151 171 7253 175
rect 7034 165 7067 168
rect 7030 163 7067 165
rect 7030 162 7097 163
rect 7030 157 7061 162
rect 7067 157 7097 162
rect 7158 159 7173 171
rect 7030 153 7097 157
rect 7003 150 7097 153
rect 7003 143 7052 150
rect 7003 137 7033 143
rect 7052 138 7057 143
rect 6969 121 7049 137
rect 7061 129 7097 150
rect 7182 149 7212 158
rect 7235 153 7253 171
rect 7311 169 7357 175
rect 7392 171 7405 181
rect 7423 171 7440 184
rect 7273 163 7275 165
rect 7275 160 7278 163
rect 7278 158 7287 160
rect 7260 151 7290 158
rect 7260 149 7291 151
rect 7311 149 7347 169
rect 7392 168 7440 171
rect 7405 163 7439 168
rect 7158 145 7347 149
rect 7173 142 7347 145
rect 7166 139 7347 142
rect 7375 162 7439 163
rect 6969 119 6988 121
rect 7003 119 7037 121
rect 6969 103 7049 119
rect 6969 97 6988 103
rect 6639 71 6665 80
rect 6685 71 6788 81
rect 6639 69 6788 71
rect 6809 69 6844 81
rect 6478 67 6640 69
rect 6490 47 6509 67
rect 6524 65 6554 67
rect 6336 38 6371 39
rect 6379 38 6414 39
rect 6336 29 6365 38
rect 6379 29 6408 38
rect 6496 29 6509 47
rect 6561 51 6640 67
rect 6672 67 6844 69
rect 6672 51 6751 67
rect 6758 65 6788 67
rect 6561 43 6751 51
rect 6816 47 6822 67
rect 6561 39 6640 43
rect 6642 39 6670 43
rect 6672 39 6751 43
rect 6546 29 6554 39
rect 6573 31 6576 39
rect 6577 31 6595 39
rect 6640 31 6672 39
rect 6717 31 6735 39
rect 6573 29 6739 31
rect 6758 29 6769 39
rect 6831 29 6844 67
rect 6916 81 6945 97
rect 6959 81 6988 97
rect 7003 87 7033 103
rect 7061 81 7067 129
rect 7070 123 7089 129
rect 7104 123 7134 131
rect 7070 115 7134 123
rect 7070 99 7150 115
rect 7166 108 7228 139
rect 7244 108 7306 139
rect 7375 137 7424 162
rect 7439 137 7469 153
rect 7338 123 7368 131
rect 7375 129 7485 137
rect 7338 115 7383 123
rect 7177 105 7181 108
rect 7182 105 7212 108
rect 7181 104 7212 105
rect 7070 97 7089 99
rect 7104 97 7150 99
rect 7070 81 7150 97
rect 7182 92 7212 104
rect 7253 105 7259 108
rect 7260 105 7290 108
rect 7253 103 7295 105
rect 7191 88 7198 92
rect 7198 87 7199 88
rect 7157 81 7167 87
rect 7219 81 7235 97
rect 7260 92 7290 103
rect 7322 99 7384 115
rect 7322 97 7368 99
rect 7322 81 7384 97
rect 7396 81 7402 129
rect 7405 121 7485 129
rect 7405 119 7424 121
rect 7439 119 7473 121
rect 7405 103 7485 119
rect 7405 81 7424 103
rect 7439 87 7469 103
rect 7497 97 7503 171
rect 7506 97 7525 241
rect 7540 97 7546 241
rect 7555 171 7568 241
rect 7620 237 7642 241
rect 7613 215 7642 229
rect 7695 215 7711 229
rect 7749 219 7755 227
rect 7762 225 7870 241
rect 7599 213 7711 215
rect 7597 185 7648 213
rect 7695 205 7729 213
rect 7702 203 7729 205
rect 7738 205 7755 219
rect 7800 205 7832 225
rect 7877 219 7883 227
rect 7891 219 7906 241
rect 7972 235 7991 238
rect 7877 213 7906 219
rect 7921 215 7937 229
rect 7972 216 7994 235
rect 8004 229 8020 230
rect 8003 227 8020 229
rect 8004 222 8020 227
rect 7994 215 8000 216
rect 8003 215 8032 222
rect 7921 214 8032 215
rect 7921 213 8038 214
rect 7877 205 7959 213
rect 7994 210 8000 213
rect 7738 203 7959 205
rect 7702 199 7774 203
rect 7802 201 7830 203
rect 7549 137 7568 171
rect 7613 184 7648 185
rect 7695 191 7827 199
rect 7830 191 7842 199
rect 7695 189 7774 191
rect 7855 189 7959 203
rect 7695 185 7792 189
rect 7613 177 7642 184
rect 7613 171 7630 177
rect 7613 168 7647 171
rect 7695 169 7711 185
rect 7712 181 7792 185
rect 7840 185 7959 189
rect 7840 181 7920 185
rect 7712 175 7920 181
rect 7921 175 7937 185
rect 7985 181 8000 196
rect 8003 184 8038 213
rect 7723 171 7833 175
rect 7614 165 7647 168
rect 7610 163 7647 165
rect 7610 162 7677 163
rect 7610 157 7641 162
rect 7647 157 7677 162
rect 7738 159 7753 171
rect 7610 153 7677 157
rect 7583 150 7677 153
rect 7583 143 7632 150
rect 7583 137 7613 143
rect 7632 138 7637 143
rect 7549 121 7629 137
rect 7641 129 7677 150
rect 7762 149 7792 158
rect 7815 153 7833 171
rect 7891 169 7937 175
rect 7972 171 7985 181
rect 8003 171 8020 184
rect 7853 163 7855 165
rect 7855 160 7858 163
rect 7858 158 7867 160
rect 7840 151 7870 158
rect 7840 149 7871 151
rect 7891 149 7927 169
rect 7972 168 8020 171
rect 7985 163 8019 168
rect 7738 145 7927 149
rect 7753 142 7927 145
rect 7746 139 7927 142
rect 7955 162 8019 163
rect 7549 119 7568 121
rect 7583 119 7617 121
rect 7549 103 7629 119
rect 7549 97 7568 103
rect 6916 69 6951 81
rect 6953 69 6994 81
rect 6916 39 6994 69
rect 7058 69 7089 81
rect 7104 69 7207 81
rect 7219 80 7236 81
rect 7219 71 7245 80
rect 7265 71 7368 81
rect 7219 69 7368 71
rect 7389 69 7424 81
rect 7058 67 7220 69
rect 7070 47 7089 67
rect 7104 65 7134 67
rect 6916 38 6951 39
rect 6959 38 6994 39
rect 6916 29 6945 38
rect 6959 29 6988 38
rect 7076 29 7089 47
rect 7141 51 7220 67
rect 7252 67 7424 69
rect 7252 51 7331 67
rect 7338 65 7368 67
rect 7141 43 7331 51
rect 7396 47 7402 67
rect 7141 39 7220 43
rect 7222 39 7250 43
rect 7252 39 7331 43
rect 7126 29 7134 39
rect 7153 31 7156 39
rect 7157 31 7175 39
rect 7220 31 7252 39
rect 7297 31 7315 39
rect 7153 29 7319 31
rect 7338 29 7349 39
rect 7411 29 7424 67
rect 7496 81 7525 97
rect 7539 81 7568 97
rect 7583 87 7613 103
rect 7641 81 7647 129
rect 7650 123 7669 129
rect 7684 123 7714 131
rect 7650 115 7714 123
rect 7650 99 7730 115
rect 7746 108 7808 139
rect 7824 108 7886 139
rect 7955 137 8004 162
rect 8019 137 8049 153
rect 7918 123 7948 131
rect 7955 129 8065 137
rect 7918 115 7963 123
rect 7757 105 7761 108
rect 7762 105 7792 108
rect 7761 104 7792 105
rect 7650 97 7669 99
rect 7684 97 7730 99
rect 7650 81 7730 97
rect 7762 92 7792 104
rect 7833 105 7839 108
rect 7840 105 7870 108
rect 7833 103 7875 105
rect 7771 88 7778 92
rect 7778 87 7779 88
rect 7737 81 7747 87
rect 7799 81 7815 97
rect 7840 92 7870 103
rect 7902 99 7964 115
rect 7902 97 7948 99
rect 7902 81 7964 97
rect 7976 81 7982 129
rect 7985 121 8065 129
rect 7985 119 8004 121
rect 8019 119 8053 121
rect 7985 103 8065 119
rect 7985 81 8004 103
rect 8019 87 8049 103
rect 8077 97 8083 171
rect 8086 97 8105 241
rect 8120 97 8126 241
rect 8135 171 8148 241
rect 8200 237 8222 241
rect 8193 215 8222 229
rect 8275 215 8291 229
rect 8329 219 8335 227
rect 8342 225 8450 241
rect 8179 213 8291 215
rect 8177 185 8228 213
rect 8275 205 8309 213
rect 8282 203 8309 205
rect 8318 205 8335 219
rect 8380 205 8412 225
rect 8457 219 8463 227
rect 8471 219 8486 241
rect 8552 235 8571 238
rect 8457 213 8486 219
rect 8501 215 8517 229
rect 8552 216 8574 235
rect 8584 229 8600 230
rect 8583 227 8600 229
rect 8584 222 8600 227
rect 8574 215 8580 216
rect 8583 215 8612 222
rect 8501 214 8612 215
rect 8501 213 8618 214
rect 8457 205 8539 213
rect 8574 210 8580 213
rect 8318 203 8539 205
rect 8282 199 8354 203
rect 8382 201 8410 203
rect 8129 137 8148 171
rect 8193 184 8228 185
rect 8275 191 8407 199
rect 8410 191 8422 199
rect 8275 189 8354 191
rect 8435 189 8539 203
rect 8275 185 8372 189
rect 8193 177 8222 184
rect 8193 171 8210 177
rect 8193 168 8227 171
rect 8275 169 8291 185
rect 8292 181 8372 185
rect 8420 185 8539 189
rect 8420 181 8500 185
rect 8292 175 8500 181
rect 8501 175 8517 185
rect 8565 181 8580 196
rect 8583 184 8618 213
rect 8303 171 8413 175
rect 8194 165 8227 168
rect 8190 163 8227 165
rect 8190 162 8257 163
rect 8190 157 8221 162
rect 8227 157 8257 162
rect 8318 159 8333 171
rect 8190 153 8257 157
rect 8163 150 8257 153
rect 8163 143 8212 150
rect 8163 137 8193 143
rect 8212 138 8217 143
rect 8129 121 8209 137
rect 8221 129 8257 150
rect 8342 149 8372 158
rect 8395 153 8413 171
rect 8471 169 8517 175
rect 8552 171 8565 181
rect 8583 171 8600 184
rect 8433 163 8435 165
rect 8435 160 8438 163
rect 8438 158 8447 160
rect 8420 151 8450 158
rect 8420 149 8451 151
rect 8471 149 8507 169
rect 8552 168 8600 171
rect 8565 163 8599 168
rect 8318 145 8507 149
rect 8333 142 8507 145
rect 8326 139 8507 142
rect 8535 162 8599 163
rect 8129 119 8148 121
rect 8163 119 8197 121
rect 8129 103 8209 119
rect 8129 97 8148 103
rect 7496 69 7531 81
rect 7533 69 7574 81
rect 7496 39 7574 69
rect 7638 69 7669 81
rect 7684 69 7787 81
rect 7799 80 7816 81
rect 7799 71 7825 80
rect 7845 71 7948 81
rect 7799 69 7948 71
rect 7969 69 8004 81
rect 7638 67 7800 69
rect 7650 47 7669 67
rect 7684 65 7714 67
rect 7496 38 7531 39
rect 7539 38 7574 39
rect 7496 29 7525 38
rect 7539 29 7568 38
rect 7656 29 7669 47
rect 7721 51 7800 67
rect 7832 67 8004 69
rect 7832 51 7911 67
rect 7918 65 7948 67
rect 7721 43 7911 51
rect 7976 47 7982 67
rect 7721 39 7800 43
rect 7802 39 7830 43
rect 7832 39 7911 43
rect 7706 29 7714 39
rect 7733 31 7736 39
rect 7737 31 7755 39
rect 7800 31 7832 39
rect 7877 31 7895 39
rect 7733 29 7899 31
rect 7918 29 7929 39
rect 7991 29 8004 67
rect 8076 81 8105 97
rect 8119 81 8148 97
rect 8163 87 8193 103
rect 8221 81 8227 129
rect 8230 123 8249 129
rect 8264 123 8294 131
rect 8230 115 8294 123
rect 8230 99 8310 115
rect 8326 108 8388 139
rect 8404 108 8466 139
rect 8535 137 8584 162
rect 8599 137 8629 153
rect 8498 123 8528 131
rect 8535 129 8645 137
rect 8498 115 8543 123
rect 8337 104 8372 108
rect 8230 97 8249 99
rect 8264 97 8310 99
rect 8230 81 8310 97
rect 8342 92 8372 104
rect 8413 105 8450 108
rect 8413 103 8455 105
rect 8351 88 8358 92
rect 8358 87 8359 88
rect 8317 81 8327 87
rect 8076 69 8111 81
rect 8113 69 8154 81
rect 8076 39 8154 69
rect 8218 69 8249 81
rect 8264 69 8367 81
rect 8379 80 8396 97
rect 8420 92 8450 103
rect 8482 99 8544 115
rect 8482 97 8528 99
rect 8482 81 8544 97
rect 8556 81 8562 129
rect 8565 121 8645 129
rect 8565 119 8584 121
rect 8599 119 8633 121
rect 8565 103 8645 119
rect 8565 81 8584 103
rect 8599 87 8629 103
rect 8657 97 8663 171
rect 8666 97 8685 241
rect 8700 97 8706 241
rect 8715 171 8728 241
rect 8780 237 8802 241
rect 8773 215 8802 229
rect 8855 215 8871 229
rect 8909 219 8915 227
rect 8922 225 9030 241
rect 8759 213 8871 215
rect 8757 185 8808 213
rect 8855 205 8889 213
rect 8862 203 8889 205
rect 8898 205 8915 219
rect 8960 205 8992 225
rect 9037 219 9043 227
rect 9051 219 9066 241
rect 9132 235 9151 238
rect 9037 213 9066 219
rect 9081 215 9097 229
rect 9132 216 9154 235
rect 9164 229 9180 230
rect 9163 227 9180 229
rect 9164 222 9180 227
rect 9154 215 9160 216
rect 9163 215 9192 222
rect 9081 214 9192 215
rect 9081 213 9198 214
rect 9037 205 9119 213
rect 9154 210 9160 213
rect 8898 203 9119 205
rect 8862 199 8934 203
rect 8962 201 8990 203
rect 8709 137 8728 171
rect 8773 184 8808 185
rect 8855 191 8987 199
rect 8990 191 9002 199
rect 8855 189 8934 191
rect 9015 189 9119 203
rect 8855 185 8952 189
rect 8773 177 8802 184
rect 8773 171 8790 177
rect 8773 168 8807 171
rect 8855 169 8871 185
rect 8872 181 8952 185
rect 9000 185 9119 189
rect 9000 181 9080 185
rect 8872 175 9080 181
rect 9081 175 9097 185
rect 9145 181 9160 196
rect 9163 184 9198 213
rect 8883 171 8993 175
rect 8774 165 8807 168
rect 8770 163 8807 165
rect 8770 162 8837 163
rect 8770 157 8801 162
rect 8807 157 8837 162
rect 8898 159 8913 171
rect 8770 153 8837 157
rect 8743 150 8837 153
rect 8743 143 8792 150
rect 8743 137 8773 143
rect 8792 138 8797 143
rect 8709 121 8789 137
rect 8801 129 8837 150
rect 8922 149 8952 158
rect 8975 153 8993 171
rect 9051 169 9097 175
rect 9132 171 9145 181
rect 9163 171 9180 184
rect 9013 163 9015 165
rect 9015 160 9018 163
rect 9018 158 9027 160
rect 9000 151 9030 158
rect 9000 149 9031 151
rect 9051 149 9087 169
rect 9132 168 9180 171
rect 9145 163 9179 168
rect 8898 145 9087 149
rect 8913 142 9087 145
rect 8906 139 9087 142
rect 9115 162 9179 163
rect 8709 119 8728 121
rect 8743 119 8777 121
rect 8709 103 8789 119
rect 8709 97 8728 103
rect 8379 71 8405 80
rect 8425 71 8528 81
rect 8379 69 8528 71
rect 8549 69 8584 81
rect 8218 67 8380 69
rect 8230 47 8249 67
rect 8264 65 8294 67
rect 8076 38 8111 39
rect 8119 38 8154 39
rect 8076 29 8105 38
rect 8119 29 8148 38
rect 8236 29 8249 47
rect 8301 51 8380 67
rect 8412 67 8584 69
rect 8412 51 8491 67
rect 8498 65 8528 67
rect 8301 43 8491 51
rect 8556 47 8562 67
rect 8301 39 8380 43
rect 8382 39 8410 43
rect 8412 39 8491 43
rect 8286 29 8294 39
rect 8313 31 8316 39
rect 8317 31 8335 39
rect 8380 31 8412 39
rect 8457 31 8475 39
rect 8313 29 8479 31
rect 8498 29 8509 39
rect 8571 29 8584 67
rect 8656 81 8685 97
rect 8699 81 8728 97
rect 8743 87 8773 103
rect 8801 81 8807 129
rect 8810 123 8829 129
rect 8844 123 8874 131
rect 8810 115 8874 123
rect 8810 99 8890 115
rect 8906 108 8968 139
rect 8984 108 9046 139
rect 9115 137 9164 162
rect 9179 137 9209 153
rect 9078 123 9108 131
rect 9115 129 9225 137
rect 9078 115 9123 123
rect 8917 105 8921 108
rect 8922 105 8952 108
rect 8921 104 8952 105
rect 8810 97 8829 99
rect 8844 97 8890 99
rect 8810 81 8890 97
rect 8922 92 8952 104
rect 8993 105 8999 108
rect 9000 105 9030 108
rect 8993 103 9035 105
rect 8931 88 8938 92
rect 8938 87 8939 88
rect 8897 81 8907 87
rect 8959 81 8975 97
rect 9000 92 9030 103
rect 9062 99 9124 115
rect 9062 97 9108 99
rect 9062 81 9124 97
rect 9136 81 9142 129
rect 9145 121 9225 129
rect 9145 119 9164 121
rect 9179 119 9213 121
rect 9145 103 9225 119
rect 9145 81 9164 103
rect 9179 87 9209 103
rect 9237 97 9243 171
rect 9246 97 9265 241
rect 9280 97 9286 241
rect 9295 171 9308 241
rect 9360 237 9382 241
rect 9353 215 9382 229
rect 9435 215 9451 229
rect 9489 219 9495 227
rect 9502 225 9610 241
rect 9353 213 9451 215
rect 9337 205 9388 213
rect 9435 205 9469 213
rect 9337 193 9362 205
rect 9369 193 9388 205
rect 9442 203 9469 205
rect 9478 205 9495 219
rect 9540 205 9572 225
rect 9617 219 9623 227
rect 9631 219 9646 241
rect 9712 235 9731 238
rect 9617 213 9646 219
rect 9661 215 9677 229
rect 9712 216 9734 235
rect 9744 229 9760 230
rect 9743 227 9760 229
rect 9744 222 9760 227
rect 9734 215 9740 216
rect 9743 215 9772 222
rect 9661 214 9772 215
rect 9661 213 9778 214
rect 9617 205 9699 213
rect 9734 210 9740 213
rect 9478 203 9699 205
rect 9442 199 9514 203
rect 9542 201 9570 203
rect 9337 185 9388 193
rect 9435 191 9567 199
rect 9570 191 9581 199
rect 9435 189 9514 191
rect 9595 189 9699 203
rect 9743 205 9778 213
rect 9435 185 9532 189
rect 9289 137 9308 171
rect 9353 177 9382 185
rect 9353 171 9370 177
rect 9353 169 9387 171
rect 9435 169 9451 185
rect 9452 181 9532 185
rect 9580 185 9699 189
rect 9580 181 9660 185
rect 9452 175 9660 181
rect 9661 175 9677 185
rect 9725 181 9740 196
rect 9743 193 9744 205
rect 9751 193 9778 205
rect 9743 185 9778 193
rect 9743 184 9772 185
rect 9463 171 9573 175
rect 9354 165 9387 169
rect 9350 163 9387 165
rect 9350 162 9417 163
rect 9350 157 9381 162
rect 9387 157 9417 162
rect 9478 159 9493 171
rect 9350 153 9417 157
rect 9323 150 9417 153
rect 9323 143 9372 150
rect 9323 137 9353 143
rect 9372 138 9377 143
rect 9289 121 9369 137
rect 9381 129 9417 150
rect 9502 149 9532 158
rect 9555 153 9573 171
rect 9631 169 9677 175
rect 9712 171 9725 181
rect 9743 171 9760 184
rect 9712 169 9760 171
rect 9593 163 9595 165
rect 9595 161 9597 163
rect 9597 158 9607 161
rect 9580 151 9610 158
rect 9580 149 9611 151
rect 9631 149 9667 169
rect 9712 168 9759 169
rect 9725 163 9759 168
rect 9478 145 9667 149
rect 9493 142 9667 145
rect 9486 139 9667 142
rect 9695 162 9759 163
rect 9289 119 9308 121
rect 9323 119 9357 121
rect 9289 103 9369 119
rect 9289 97 9308 103
rect 8656 69 8691 81
rect 8693 69 8734 81
rect 8656 39 8734 69
rect 8798 69 8829 81
rect 8844 69 8947 81
rect 8959 80 8976 81
rect 8959 71 8985 80
rect 9005 71 9108 81
rect 8959 69 9108 71
rect 9129 69 9164 81
rect 8798 67 8960 69
rect 8810 47 8829 67
rect 8844 65 8874 67
rect 8656 38 8691 39
rect 8699 38 8734 39
rect 8656 29 8685 38
rect 8699 29 8728 38
rect 8816 29 8829 47
rect 8881 51 8960 67
rect 8992 67 9164 69
rect 8992 51 9071 67
rect 9078 65 9108 67
rect 8881 43 9071 51
rect 9136 47 9142 67
rect 8881 39 8960 43
rect 8962 39 8990 43
rect 8992 39 9071 43
rect 8866 29 8874 39
rect 8893 31 8896 39
rect 8897 31 8915 39
rect 8960 31 8992 39
rect 9037 31 9055 39
rect 8893 29 9059 31
rect 9078 29 9089 39
rect 9151 29 9164 67
rect 9236 81 9265 97
rect 9279 81 9308 97
rect 9323 87 9353 103
rect 9381 81 9387 129
rect 9390 123 9409 129
rect 9424 123 9454 131
rect 9390 115 9454 123
rect 9390 99 9470 115
rect 9486 108 9548 139
rect 9564 108 9626 139
rect 9695 137 9744 162
rect 9759 137 9789 153
rect 9658 123 9688 131
rect 9695 129 9805 137
rect 9658 115 9703 123
rect 9497 105 9501 108
rect 9502 105 9532 108
rect 9390 97 9409 99
rect 9424 97 9470 99
rect 9390 81 9470 97
rect 9501 95 9532 105
rect 9573 105 9579 108
rect 9580 105 9610 108
rect 9573 103 9615 105
rect 9502 92 9532 95
rect 9511 88 9518 92
rect 9518 87 9519 88
rect 9477 81 9487 87
rect 9539 81 9555 97
rect 9580 92 9610 103
rect 9642 99 9704 115
rect 9642 97 9688 99
rect 9642 81 9704 97
rect 9716 81 9722 129
rect 9725 121 9805 129
rect 9725 119 9744 121
rect 9759 119 9793 121
rect 9725 103 9805 119
rect 9725 81 9744 103
rect 9759 87 9789 103
rect 9817 97 9823 171
rect 9826 97 9845 241
rect 9860 97 9866 241
rect 9875 171 9888 241
rect 9940 237 9962 241
rect 9933 215 9962 229
rect 10015 215 10031 229
rect 10069 219 10075 227
rect 10082 225 10190 241
rect 9933 213 10031 215
rect 9917 205 9968 213
rect 10015 205 10049 213
rect 9917 193 9942 205
rect 9949 193 9968 205
rect 10022 203 10049 205
rect 10058 205 10075 219
rect 10120 205 10152 225
rect 10197 219 10203 227
rect 10211 219 10226 241
rect 10292 235 10311 238
rect 10197 213 10226 219
rect 10241 215 10257 229
rect 10292 216 10314 235
rect 10324 229 10340 230
rect 10323 227 10340 229
rect 10324 222 10340 227
rect 10314 215 10320 216
rect 10323 215 10352 222
rect 10241 214 10352 215
rect 10241 213 10358 214
rect 10197 205 10279 213
rect 10314 210 10320 213
rect 10058 203 10279 205
rect 10022 199 10094 203
rect 10122 201 10150 203
rect 9917 185 9968 193
rect 10015 191 10147 199
rect 10150 191 10161 199
rect 10015 189 10094 191
rect 10175 189 10279 203
rect 10323 205 10358 213
rect 10015 185 10112 189
rect 9869 137 9888 171
rect 9933 177 9962 185
rect 9933 171 9950 177
rect 9933 169 9967 171
rect 10015 169 10031 185
rect 10032 181 10112 185
rect 10160 185 10279 189
rect 10160 181 10240 185
rect 10032 175 10240 181
rect 10241 175 10257 185
rect 10305 181 10320 196
rect 10323 193 10324 205
rect 10331 193 10358 205
rect 10323 185 10358 193
rect 10323 184 10352 185
rect 10043 171 10153 175
rect 9934 165 9967 169
rect 9930 163 9967 165
rect 9930 162 9997 163
rect 9930 157 9961 162
rect 9967 157 9997 162
rect 10058 159 10073 171
rect 9930 153 9997 157
rect 9903 150 9997 153
rect 9903 143 9952 150
rect 9903 137 9933 143
rect 9952 138 9957 143
rect 9869 121 9949 137
rect 9961 129 9997 150
rect 10082 149 10112 158
rect 10135 153 10153 171
rect 10211 169 10257 175
rect 10292 171 10305 181
rect 10323 171 10340 184
rect 10292 169 10340 171
rect 10173 163 10175 165
rect 10175 161 10177 163
rect 10177 158 10187 161
rect 10160 151 10190 158
rect 10160 149 10191 151
rect 10211 149 10247 169
rect 10292 168 10339 169
rect 10305 163 10339 168
rect 10058 145 10247 149
rect 10073 142 10247 145
rect 10066 139 10247 142
rect 10275 162 10339 163
rect 9869 119 9888 121
rect 9903 119 9937 121
rect 9869 103 9949 119
rect 9869 97 9888 103
rect 9236 38 9271 81
rect 9273 73 9314 81
rect 9273 47 9288 73
rect 9295 47 9314 73
rect 9378 69 9409 81
rect 9424 69 9527 81
rect 9539 71 9565 81
rect 9585 71 9688 81
rect 9539 69 9688 71
rect 9709 69 9744 81
rect 9378 67 9540 69
rect 9390 47 9409 67
rect 9424 65 9454 67
rect 9273 39 9314 47
rect 9236 29 9265 38
rect 9279 29 9308 39
rect 9396 29 9409 47
rect 9461 51 9540 67
rect 9572 67 9744 69
rect 9572 51 9651 67
rect 9658 65 9688 67
rect 9461 43 9651 51
rect 9716 47 9722 67
rect 9461 39 9540 43
rect 9542 39 9570 43
rect 9572 39 9651 43
rect 9446 29 9454 39
rect 9473 31 9476 39
rect 9477 31 9495 39
rect 9540 31 9572 39
rect 9617 31 9635 39
rect 9473 29 9639 31
rect 9658 29 9669 39
rect 9731 29 9744 67
rect 9816 81 9845 97
rect 9859 81 9888 97
rect 9903 87 9933 103
rect 9961 81 9967 129
rect 9970 123 9989 129
rect 10004 123 10034 131
rect 9970 115 10034 123
rect 9970 99 10050 115
rect 10066 108 10128 139
rect 10144 108 10206 139
rect 10275 137 10324 162
rect 10339 137 10369 153
rect 10238 123 10268 131
rect 10275 129 10385 137
rect 10238 115 10283 123
rect 10077 105 10081 108
rect 10082 105 10112 108
rect 9970 97 9989 99
rect 10004 97 10050 99
rect 9970 81 10050 97
rect 10081 95 10112 105
rect 10153 105 10159 108
rect 10160 105 10190 108
rect 10153 103 10195 105
rect 10082 92 10112 95
rect 10091 88 10098 92
rect 10098 87 10099 88
rect 10057 81 10067 87
rect 10119 81 10135 97
rect 10160 92 10190 103
rect 10222 99 10284 115
rect 10222 97 10268 99
rect 10222 81 10284 97
rect 10296 81 10302 129
rect 10305 121 10385 129
rect 10305 119 10324 121
rect 10339 119 10373 121
rect 10305 103 10385 119
rect 10305 81 10324 103
rect 10339 87 10369 103
rect 10397 97 10403 171
rect 10406 97 10425 241
rect 10440 97 10446 241
rect 10455 171 10468 241
rect 10520 237 10542 241
rect 10513 215 10542 229
rect 10595 215 10611 229
rect 10649 219 10655 227
rect 10662 225 10770 241
rect 10513 213 10611 215
rect 10497 205 10548 213
rect 10595 205 10629 213
rect 10497 193 10522 205
rect 10529 193 10548 205
rect 10602 203 10629 205
rect 10638 205 10655 219
rect 10700 205 10732 225
rect 10777 219 10783 227
rect 10791 219 10806 241
rect 10872 235 10891 238
rect 10777 213 10806 219
rect 10821 215 10837 229
rect 10872 216 10894 235
rect 10904 229 10920 230
rect 10903 227 10920 229
rect 10904 222 10920 227
rect 10894 215 10900 216
rect 10903 215 10932 222
rect 10821 214 10932 215
rect 10821 213 10938 214
rect 10777 205 10859 213
rect 10894 210 10900 213
rect 10638 203 10859 205
rect 10602 199 10674 203
rect 10702 201 10730 203
rect 10497 185 10548 193
rect 10595 191 10727 199
rect 10730 191 10741 199
rect 10595 189 10674 191
rect 10755 189 10859 203
rect 10903 205 10938 213
rect 10595 185 10692 189
rect 10449 137 10468 171
rect 10513 177 10542 185
rect 10513 171 10530 177
rect 10513 169 10547 171
rect 10595 169 10611 185
rect 10612 181 10692 185
rect 10740 185 10859 189
rect 10740 181 10820 185
rect 10612 175 10820 181
rect 10821 175 10837 185
rect 10885 181 10900 196
rect 10903 193 10904 205
rect 10911 193 10938 205
rect 10903 185 10938 193
rect 10903 184 10932 185
rect 10623 171 10733 175
rect 10514 165 10547 169
rect 10510 163 10547 165
rect 10510 162 10577 163
rect 10510 157 10541 162
rect 10547 157 10577 162
rect 10638 159 10653 171
rect 10510 153 10577 157
rect 10483 150 10577 153
rect 10483 143 10532 150
rect 10483 137 10513 143
rect 10532 138 10537 143
rect 10449 121 10529 137
rect 10541 129 10577 150
rect 10662 149 10692 158
rect 10715 153 10733 171
rect 10791 169 10837 175
rect 10872 171 10885 181
rect 10903 171 10920 184
rect 10872 169 10920 171
rect 10753 163 10755 165
rect 10755 161 10757 163
rect 10757 158 10767 161
rect 10740 151 10770 158
rect 10740 149 10771 151
rect 10791 149 10827 169
rect 10872 168 10919 169
rect 10885 163 10919 168
rect 10638 145 10827 149
rect 10653 142 10827 145
rect 10646 139 10827 142
rect 10855 162 10919 163
rect 10449 119 10468 121
rect 10483 119 10517 121
rect 10449 103 10529 119
rect 10449 97 10468 103
rect 9816 73 9851 81
rect 9816 47 9817 73
rect 9824 47 9851 73
rect 9816 39 9851 47
rect 9853 73 9894 81
rect 9853 47 9868 73
rect 9875 47 9894 73
rect 9958 69 9989 81
rect 10004 69 10107 81
rect 10119 71 10145 81
rect 10165 71 10268 81
rect 10119 69 10268 71
rect 10289 69 10324 81
rect 9958 67 10120 69
rect 9970 47 9989 67
rect 10004 65 10034 67
rect 9853 39 9894 47
rect 9816 29 9845 39
rect 9859 29 9888 39
rect 9976 29 9989 47
rect 10041 51 10120 67
rect 10152 67 10324 69
rect 10152 51 10231 67
rect 10238 65 10268 67
rect 10041 43 10231 51
rect 10296 47 10302 67
rect 10041 39 10120 43
rect 10122 39 10150 43
rect 10152 39 10231 43
rect 10026 29 10034 39
rect 10053 31 10056 39
rect 10057 31 10075 39
rect 10120 31 10152 39
rect 10197 31 10215 39
rect 10053 29 10219 31
rect 10238 29 10249 39
rect 10311 29 10324 67
rect 10396 81 10425 97
rect 10439 81 10468 97
rect 10483 87 10513 103
rect 10541 81 10547 129
rect 10550 123 10569 129
rect 10584 123 10614 131
rect 10550 115 10614 123
rect 10550 99 10630 115
rect 10646 108 10708 139
rect 10724 108 10786 139
rect 10855 137 10904 162
rect 10919 137 10949 153
rect 10818 123 10848 131
rect 10855 129 10965 137
rect 10818 115 10863 123
rect 10657 105 10661 108
rect 10662 105 10692 108
rect 10550 97 10569 99
rect 10584 97 10630 99
rect 10550 81 10630 97
rect 10661 95 10692 105
rect 10733 105 10739 108
rect 10740 105 10770 108
rect 10733 103 10775 105
rect 10662 92 10692 95
rect 10671 88 10678 92
rect 10678 87 10679 88
rect 10637 81 10647 87
rect 10699 81 10715 97
rect 10740 92 10770 103
rect 10802 99 10864 115
rect 10802 97 10848 99
rect 10802 81 10864 97
rect 10876 81 10882 129
rect 10885 121 10965 129
rect 10885 119 10904 121
rect 10919 119 10953 121
rect 10885 103 10965 119
rect 10885 81 10904 103
rect 10919 87 10949 103
rect 10977 97 10983 171
rect 10986 97 11005 241
rect 11020 97 11026 241
rect 11035 171 11048 241
rect 11100 237 11122 241
rect 11093 215 11122 229
rect 11175 215 11191 229
rect 11229 219 11235 227
rect 11242 225 11350 241
rect 11093 213 11191 215
rect 11077 205 11128 213
rect 11175 205 11209 213
rect 11077 193 11102 205
rect 11109 193 11128 205
rect 11182 203 11209 205
rect 11218 205 11235 219
rect 11280 205 11312 225
rect 11357 219 11363 227
rect 11371 219 11386 241
rect 11452 235 11471 238
rect 11357 213 11386 219
rect 11401 215 11417 229
rect 11452 216 11474 235
rect 11484 229 11500 230
rect 11483 227 11500 229
rect 11484 222 11500 227
rect 11474 215 11480 216
rect 11483 215 11512 222
rect 11401 214 11512 215
rect 11401 213 11518 214
rect 11357 205 11439 213
rect 11474 210 11480 213
rect 11218 203 11439 205
rect 11182 199 11254 203
rect 11282 201 11310 203
rect 11077 185 11128 193
rect 11175 191 11307 199
rect 11310 191 11321 199
rect 11175 189 11254 191
rect 11335 189 11439 203
rect 11483 205 11518 213
rect 11175 185 11272 189
rect 11029 137 11048 171
rect 11093 177 11122 185
rect 11093 171 11110 177
rect 11093 169 11127 171
rect 11175 169 11191 185
rect 11192 181 11272 185
rect 11320 185 11439 189
rect 11320 181 11400 185
rect 11192 175 11400 181
rect 11401 175 11417 185
rect 11465 181 11480 196
rect 11483 193 11484 205
rect 11491 193 11518 205
rect 11483 185 11518 193
rect 11483 184 11512 185
rect 11203 171 11313 175
rect 11094 165 11127 169
rect 11090 163 11127 165
rect 11090 162 11157 163
rect 11090 157 11121 162
rect 11127 157 11157 162
rect 11218 159 11233 171
rect 11090 153 11157 157
rect 11063 150 11157 153
rect 11063 143 11112 150
rect 11063 137 11093 143
rect 11112 138 11117 143
rect 11029 121 11109 137
rect 11121 129 11157 150
rect 11242 149 11272 158
rect 11295 153 11313 171
rect 11371 169 11417 175
rect 11452 171 11465 181
rect 11483 171 11500 184
rect 11452 169 11500 171
rect 11333 163 11335 165
rect 11335 161 11337 163
rect 11337 158 11347 161
rect 11320 151 11350 158
rect 11320 149 11351 151
rect 11371 149 11407 169
rect 11452 168 11499 169
rect 11465 163 11499 168
rect 11218 145 11407 149
rect 11233 142 11407 145
rect 11226 139 11407 142
rect 11435 162 11499 163
rect 11029 119 11048 121
rect 11063 119 11097 121
rect 11029 103 11109 119
rect 11029 97 11048 103
rect 10396 73 10431 81
rect 10396 47 10397 73
rect 10404 47 10431 73
rect 10396 39 10431 47
rect 10433 73 10474 81
rect 10433 47 10448 73
rect 10455 47 10474 73
rect 10538 69 10569 81
rect 10584 69 10687 81
rect 10699 71 10725 81
rect 10745 71 10848 81
rect 10699 69 10848 71
rect 10869 69 10904 81
rect 10538 67 10700 69
rect 10550 47 10569 67
rect 10584 65 10614 67
rect 10433 39 10474 47
rect 10396 29 10425 39
rect 10439 29 10468 39
rect 10556 29 10569 47
rect 10621 51 10700 67
rect 10732 67 10904 69
rect 10732 51 10811 67
rect 10818 65 10848 67
rect 10621 43 10811 51
rect 10876 47 10882 67
rect 10621 39 10700 43
rect 10702 39 10730 43
rect 10732 39 10811 43
rect 10606 29 10614 39
rect 10633 31 10636 39
rect 10637 31 10655 39
rect 10700 31 10732 39
rect 10777 31 10795 39
rect 10633 29 10799 31
rect 10818 29 10829 39
rect 10891 29 10904 67
rect 10976 81 11005 97
rect 11019 81 11048 97
rect 11063 87 11093 103
rect 11121 81 11127 129
rect 11130 123 11149 129
rect 11164 123 11194 131
rect 11130 115 11194 123
rect 11130 99 11210 115
rect 11226 108 11288 139
rect 11304 108 11366 139
rect 11435 137 11484 162
rect 11499 137 11529 153
rect 11398 123 11428 131
rect 11435 129 11545 137
rect 11398 115 11443 123
rect 11237 105 11241 108
rect 11242 105 11272 108
rect 11130 97 11149 99
rect 11164 97 11210 99
rect 11130 81 11210 97
rect 11241 95 11272 105
rect 11313 105 11319 108
rect 11320 105 11350 108
rect 11313 103 11355 105
rect 11242 92 11272 95
rect 11251 88 11258 92
rect 11258 87 11259 88
rect 11217 81 11227 87
rect 11279 81 11295 97
rect 11320 92 11350 103
rect 11382 99 11444 115
rect 11382 97 11428 99
rect 11382 81 11444 97
rect 11456 81 11462 129
rect 11465 121 11545 129
rect 11465 119 11484 121
rect 11499 119 11533 121
rect 11465 103 11545 119
rect 11465 81 11484 103
rect 11499 87 11529 103
rect 11557 97 11563 171
rect 11566 97 11585 241
rect 11600 97 11606 241
rect 11615 171 11628 241
rect 11680 237 11702 241
rect 11673 215 11702 229
rect 11755 215 11771 229
rect 11809 219 11815 227
rect 11822 225 11930 241
rect 11673 213 11771 215
rect 11657 205 11708 213
rect 11755 205 11789 213
rect 11657 193 11682 205
rect 11689 193 11708 205
rect 11762 203 11789 205
rect 11798 205 11815 219
rect 11860 205 11892 225
rect 11937 219 11943 227
rect 11951 219 11966 241
rect 12032 235 12051 238
rect 11937 213 11966 219
rect 11981 215 11997 229
rect 12032 216 12054 235
rect 12064 229 12080 230
rect 12063 227 12080 229
rect 12064 222 12080 227
rect 12054 215 12060 216
rect 12063 215 12092 222
rect 11981 214 12092 215
rect 11981 213 12098 214
rect 11937 205 12019 213
rect 12054 210 12060 213
rect 11798 203 12019 205
rect 11762 199 11834 203
rect 11862 201 11890 203
rect 11657 185 11708 193
rect 11755 191 11887 199
rect 11890 191 11901 199
rect 11755 189 11834 191
rect 11915 189 12019 203
rect 12063 205 12098 213
rect 11755 185 11852 189
rect 11609 137 11628 171
rect 11673 177 11702 185
rect 11673 171 11690 177
rect 11673 169 11707 171
rect 11755 169 11771 185
rect 11772 181 11852 185
rect 11900 185 12019 189
rect 11900 181 11980 185
rect 11772 175 11980 181
rect 11981 175 11997 185
rect 12045 181 12060 196
rect 12063 193 12064 205
rect 12071 193 12098 205
rect 12063 185 12098 193
rect 12063 184 12092 185
rect 11783 171 11893 175
rect 11674 165 11707 169
rect 11670 163 11707 165
rect 11670 162 11737 163
rect 11670 157 11701 162
rect 11707 157 11737 162
rect 11798 159 11813 171
rect 11670 153 11737 157
rect 11643 150 11737 153
rect 11643 143 11692 150
rect 11643 137 11673 143
rect 11692 138 11697 143
rect 11609 121 11689 137
rect 11701 129 11737 150
rect 11822 149 11852 158
rect 11875 153 11893 171
rect 11951 169 11997 175
rect 12032 171 12045 181
rect 12063 171 12080 184
rect 12032 169 12080 171
rect 11913 163 11915 165
rect 11915 161 11917 163
rect 11917 158 11927 161
rect 11900 151 11930 158
rect 11900 149 11931 151
rect 11951 149 11987 169
rect 12032 168 12079 169
rect 12045 163 12079 168
rect 11798 145 11987 149
rect 11813 142 11987 145
rect 11806 139 11987 142
rect 12015 162 12079 163
rect 11609 119 11628 121
rect 11643 119 11677 121
rect 11609 103 11689 119
rect 11609 97 11628 103
rect 10976 73 11011 81
rect 10976 47 10977 73
rect 10984 47 11011 73
rect 10976 39 11011 47
rect 11013 73 11054 81
rect 11013 47 11028 73
rect 11035 47 11054 73
rect 11118 69 11149 81
rect 11164 69 11267 81
rect 11279 71 11305 81
rect 11325 71 11428 81
rect 11279 69 11428 71
rect 11449 69 11484 81
rect 11118 67 11280 69
rect 11130 47 11149 67
rect 11164 65 11194 67
rect 11013 39 11054 47
rect 10976 29 11005 39
rect 11019 29 11048 39
rect 11136 29 11149 47
rect 11201 51 11280 67
rect 11312 67 11484 69
rect 11312 51 11391 67
rect 11398 65 11428 67
rect 11201 43 11391 51
rect 11456 47 11462 67
rect 11201 39 11280 43
rect 11282 39 11310 43
rect 11312 39 11391 43
rect 11186 29 11194 39
rect 11213 31 11216 39
rect 11217 31 11235 39
rect 11280 31 11312 39
rect 11357 31 11375 39
rect 11213 29 11379 31
rect 11398 29 11409 39
rect 11471 29 11484 67
rect 11556 81 11585 97
rect 11599 81 11628 97
rect 11643 87 11673 103
rect 11701 81 11707 129
rect 11710 123 11729 129
rect 11744 123 11774 131
rect 11710 115 11774 123
rect 11710 99 11790 115
rect 11806 108 11868 139
rect 11884 108 11946 139
rect 12015 137 12064 162
rect 12079 137 12109 153
rect 11978 123 12008 131
rect 12015 129 12125 137
rect 11978 115 12023 123
rect 11817 105 11821 108
rect 11822 105 11852 108
rect 11710 97 11729 99
rect 11744 97 11790 99
rect 11710 81 11790 97
rect 11821 95 11852 105
rect 11893 105 11899 108
rect 11900 105 11930 108
rect 11893 103 11935 105
rect 11822 92 11852 95
rect 11831 88 11838 92
rect 11838 87 11839 88
rect 11797 81 11807 87
rect 11859 81 11875 97
rect 11900 92 11930 103
rect 11962 99 12024 115
rect 11962 97 12008 99
rect 11962 81 12024 97
rect 12036 81 12042 129
rect 12045 121 12125 129
rect 12045 119 12064 121
rect 12079 119 12113 121
rect 12045 103 12125 119
rect 12045 81 12064 103
rect 12079 87 12109 103
rect 12137 97 12143 171
rect 12146 97 12165 241
rect 12180 97 12186 241
rect 12195 171 12208 241
rect 12260 237 12282 241
rect 12253 215 12282 229
rect 12335 215 12351 229
rect 12389 219 12395 227
rect 12402 225 12510 241
rect 12253 213 12351 215
rect 12237 205 12288 213
rect 12335 205 12369 213
rect 12237 193 12262 205
rect 12269 193 12288 205
rect 12342 203 12369 205
rect 12378 205 12395 219
rect 12440 205 12472 225
rect 12517 219 12523 227
rect 12531 219 12546 241
rect 12612 235 12631 238
rect 12517 213 12546 219
rect 12561 215 12577 229
rect 12612 216 12634 235
rect 12644 229 12660 230
rect 12643 227 12660 229
rect 12644 222 12660 227
rect 12634 215 12640 216
rect 12643 215 12672 222
rect 12561 214 12672 215
rect 12561 213 12678 214
rect 12517 205 12599 213
rect 12634 210 12640 213
rect 12378 203 12599 205
rect 12342 199 12414 203
rect 12442 201 12470 203
rect 12237 185 12288 193
rect 12335 191 12467 199
rect 12470 191 12481 199
rect 12335 189 12414 191
rect 12495 189 12599 203
rect 12643 205 12678 213
rect 12335 185 12432 189
rect 12189 137 12208 171
rect 12253 177 12282 185
rect 12253 171 12270 177
rect 12253 169 12287 171
rect 12335 169 12351 185
rect 12352 181 12432 185
rect 12480 185 12599 189
rect 12480 181 12560 185
rect 12352 175 12560 181
rect 12561 175 12577 185
rect 12625 181 12640 196
rect 12643 193 12644 205
rect 12651 193 12678 205
rect 12643 185 12678 193
rect 12643 184 12672 185
rect 12363 171 12473 175
rect 12254 165 12287 169
rect 12250 163 12287 165
rect 12250 162 12317 163
rect 12250 157 12281 162
rect 12287 157 12317 162
rect 12378 159 12393 171
rect 12250 153 12317 157
rect 12223 150 12317 153
rect 12223 143 12272 150
rect 12223 137 12253 143
rect 12272 138 12277 143
rect 12189 121 12269 137
rect 12281 129 12317 150
rect 12402 149 12432 158
rect 12455 153 12473 171
rect 12531 169 12577 175
rect 12612 171 12625 181
rect 12643 171 12660 184
rect 12612 169 12660 171
rect 12493 163 12495 165
rect 12495 161 12497 163
rect 12497 158 12507 161
rect 12480 151 12510 158
rect 12480 149 12511 151
rect 12531 149 12567 169
rect 12612 168 12659 169
rect 12625 163 12659 168
rect 12378 145 12567 149
rect 12393 142 12567 145
rect 12386 139 12567 142
rect 12595 162 12659 163
rect 12189 119 12208 121
rect 12223 119 12257 121
rect 12189 103 12269 119
rect 12189 97 12208 103
rect 11556 73 11591 81
rect 11556 47 11557 73
rect 11564 47 11591 73
rect 11556 39 11591 47
rect 11593 73 11634 81
rect 11593 47 11608 73
rect 11615 47 11634 73
rect 11698 69 11729 81
rect 11744 69 11847 81
rect 11859 71 11885 81
rect 11905 71 12008 81
rect 11859 69 12008 71
rect 12029 69 12064 81
rect 11698 67 11860 69
rect 11710 47 11729 67
rect 11744 65 11774 67
rect 11593 39 11634 47
rect 11556 29 11585 39
rect 11599 29 11628 39
rect 11716 29 11729 47
rect 11781 51 11860 67
rect 11892 67 12064 69
rect 11892 51 11971 67
rect 11978 65 12008 67
rect 11781 43 11971 51
rect 12036 47 12042 67
rect 11781 39 11860 43
rect 11862 39 11890 43
rect 11892 39 11971 43
rect 11766 29 11774 39
rect 11793 31 11796 39
rect 11797 31 11815 39
rect 11860 31 11892 39
rect 11937 31 11955 39
rect 11793 29 11959 31
rect 11978 29 11989 39
rect 12051 29 12064 67
rect 12136 81 12165 97
rect 12179 81 12208 97
rect 12223 87 12253 103
rect 12281 81 12287 129
rect 12290 123 12309 129
rect 12324 123 12354 131
rect 12290 115 12354 123
rect 12290 99 12370 115
rect 12386 108 12448 139
rect 12464 108 12526 139
rect 12595 137 12644 162
rect 12659 137 12689 153
rect 12558 123 12588 131
rect 12595 129 12705 137
rect 12558 115 12603 123
rect 12397 105 12401 108
rect 12402 105 12432 108
rect 12290 97 12309 99
rect 12324 97 12370 99
rect 12290 81 12370 97
rect 12401 95 12432 105
rect 12473 105 12479 108
rect 12480 105 12510 108
rect 12473 103 12515 105
rect 12402 92 12432 95
rect 12411 88 12418 92
rect 12418 87 12419 88
rect 12377 81 12387 87
rect 12439 81 12455 97
rect 12480 92 12510 103
rect 12542 99 12604 115
rect 12542 97 12588 99
rect 12542 81 12604 97
rect 12616 81 12622 129
rect 12625 121 12705 129
rect 12625 119 12644 121
rect 12659 119 12693 121
rect 12625 103 12705 119
rect 12625 81 12644 103
rect 12659 87 12689 103
rect 12717 97 12723 171
rect 12726 97 12745 241
rect 12760 97 12766 241
rect 12775 171 12788 241
rect 12840 237 12862 241
rect 12833 215 12862 229
rect 12915 215 12931 229
rect 12969 219 12975 227
rect 12982 225 13090 241
rect 12833 213 12931 215
rect 12817 205 12868 213
rect 12915 205 12949 213
rect 12817 193 12842 205
rect 12849 193 12868 205
rect 12922 203 12949 205
rect 12958 205 12975 219
rect 13020 205 13052 225
rect 13097 219 13103 227
rect 13111 219 13126 241
rect 13192 235 13211 238
rect 13097 213 13126 219
rect 13141 215 13157 229
rect 13192 216 13214 235
rect 13224 229 13240 230
rect 13223 227 13240 229
rect 13224 222 13240 227
rect 13214 215 13220 216
rect 13223 215 13252 222
rect 13141 214 13252 215
rect 13141 213 13258 214
rect 13097 205 13179 213
rect 13214 210 13220 213
rect 12958 203 13179 205
rect 12922 199 12994 203
rect 13022 201 13050 203
rect 12817 185 12868 193
rect 12915 191 13047 199
rect 13050 191 13061 199
rect 12915 189 12994 191
rect 13075 189 13179 203
rect 13223 205 13258 213
rect 12915 185 13012 189
rect 12769 137 12788 171
rect 12833 177 12862 185
rect 12833 171 12850 177
rect 12833 169 12867 171
rect 12915 169 12931 185
rect 12932 181 13012 185
rect 13060 185 13179 189
rect 13060 181 13140 185
rect 12932 175 13140 181
rect 13141 175 13157 185
rect 13205 181 13220 196
rect 13223 193 13224 205
rect 13231 193 13258 205
rect 13223 185 13258 193
rect 13223 184 13252 185
rect 12943 171 13053 175
rect 12834 165 12867 169
rect 12830 163 12867 165
rect 12830 162 12897 163
rect 12830 157 12861 162
rect 12867 157 12897 162
rect 12958 159 12973 171
rect 12830 153 12897 157
rect 12803 150 12897 153
rect 12803 143 12852 150
rect 12803 137 12833 143
rect 12852 138 12857 143
rect 12769 121 12849 137
rect 12861 129 12897 150
rect 12982 149 13012 158
rect 13035 153 13053 171
rect 13111 169 13157 175
rect 13192 171 13205 181
rect 13223 171 13240 184
rect 13192 169 13240 171
rect 13073 163 13075 165
rect 13075 161 13077 163
rect 13077 158 13087 161
rect 13060 151 13090 158
rect 13060 149 13091 151
rect 13111 149 13147 169
rect 13192 168 13239 169
rect 13205 163 13239 168
rect 12958 145 13147 149
rect 12973 142 13147 145
rect 12966 139 13147 142
rect 13175 162 13239 163
rect 12769 119 12788 121
rect 12803 119 12837 121
rect 12769 103 12849 119
rect 12769 97 12788 103
rect 12136 73 12171 81
rect 12136 47 12137 73
rect 12144 47 12171 73
rect 12136 39 12171 47
rect 12173 73 12214 81
rect 12173 47 12188 73
rect 12195 47 12214 73
rect 12278 69 12309 81
rect 12324 69 12427 81
rect 12439 71 12465 81
rect 12485 71 12588 81
rect 12439 69 12588 71
rect 12609 69 12644 81
rect 12278 67 12440 69
rect 12290 47 12309 67
rect 12324 65 12354 67
rect 12173 39 12214 47
rect 12136 29 12165 39
rect 12179 29 12208 39
rect 12296 29 12309 47
rect 12361 51 12440 67
rect 12472 67 12644 69
rect 12472 51 12551 67
rect 12558 65 12588 67
rect 12361 43 12551 51
rect 12616 47 12622 67
rect 12361 39 12440 43
rect 12442 39 12470 43
rect 12472 39 12551 43
rect 12346 29 12354 39
rect 12373 31 12376 39
rect 12377 31 12395 39
rect 12440 31 12472 39
rect 12517 31 12535 39
rect 12373 29 12539 31
rect 12558 29 12569 39
rect 12631 29 12644 67
rect 12716 81 12745 97
rect 12759 81 12788 97
rect 12803 87 12833 103
rect 12861 81 12867 129
rect 12870 123 12889 129
rect 12904 123 12934 131
rect 12870 115 12934 123
rect 12870 99 12950 115
rect 12966 108 13028 139
rect 13044 108 13106 139
rect 13175 137 13224 162
rect 13239 137 13269 153
rect 13138 123 13168 131
rect 13175 129 13285 137
rect 13138 115 13183 123
rect 12977 105 12981 108
rect 12982 105 13012 108
rect 12870 97 12889 99
rect 12904 97 12950 99
rect 12870 81 12950 97
rect 12981 95 13012 105
rect 13053 105 13059 108
rect 13060 105 13090 108
rect 13053 103 13095 105
rect 12982 92 13012 95
rect 12991 88 12998 92
rect 12998 87 12999 88
rect 12957 81 12967 87
rect 13019 81 13035 97
rect 13060 92 13090 103
rect 13122 99 13184 115
rect 13122 97 13168 99
rect 13122 81 13184 97
rect 13196 81 13202 129
rect 13205 121 13285 129
rect 13205 119 13224 121
rect 13239 119 13273 121
rect 13205 103 13285 119
rect 13205 81 13224 103
rect 13239 87 13269 103
rect 13297 97 13303 171
rect 13306 97 13325 241
rect 13340 97 13346 241
rect 13355 171 13368 241
rect 13420 237 13442 241
rect 13413 215 13442 229
rect 13495 215 13511 229
rect 13549 219 13555 227
rect 13562 225 13670 241
rect 13413 213 13511 215
rect 13397 205 13448 213
rect 13495 205 13529 213
rect 13397 193 13422 205
rect 13429 193 13448 205
rect 13502 203 13529 205
rect 13538 205 13555 219
rect 13600 205 13632 225
rect 13677 219 13683 227
rect 13691 219 13706 241
rect 13772 235 13791 238
rect 13677 213 13706 219
rect 13721 215 13737 229
rect 13772 216 13794 235
rect 13804 229 13820 230
rect 13803 227 13820 229
rect 13804 222 13820 227
rect 13794 215 13800 216
rect 13803 215 13832 222
rect 13721 214 13832 215
rect 13721 213 13838 214
rect 13677 205 13759 213
rect 13794 210 13800 213
rect 13538 203 13759 205
rect 13502 199 13574 203
rect 13602 201 13630 203
rect 13397 185 13448 193
rect 13495 191 13627 199
rect 13630 191 13641 199
rect 13495 189 13574 191
rect 13655 189 13759 203
rect 13803 205 13838 213
rect 13495 185 13592 189
rect 13349 137 13368 171
rect 13413 177 13442 185
rect 13413 171 13430 177
rect 13413 169 13447 171
rect 13495 169 13511 185
rect 13512 181 13592 185
rect 13640 185 13759 189
rect 13640 181 13720 185
rect 13512 175 13720 181
rect 13721 175 13737 185
rect 13785 181 13800 196
rect 13803 193 13804 205
rect 13811 193 13838 205
rect 13803 185 13838 193
rect 13803 184 13832 185
rect 13523 171 13633 175
rect 13414 165 13447 169
rect 13410 163 13447 165
rect 13410 162 13477 163
rect 13410 157 13441 162
rect 13447 157 13477 162
rect 13538 159 13553 171
rect 13410 153 13477 157
rect 13383 150 13477 153
rect 13383 143 13432 150
rect 13383 137 13413 143
rect 13432 138 13437 143
rect 13349 121 13429 137
rect 13441 129 13477 150
rect 13562 149 13592 158
rect 13615 153 13633 171
rect 13691 169 13737 175
rect 13772 171 13785 181
rect 13803 171 13820 184
rect 13772 169 13820 171
rect 13653 163 13655 165
rect 13655 161 13657 163
rect 13657 158 13667 161
rect 13640 151 13670 158
rect 13640 149 13671 151
rect 13691 149 13727 169
rect 13772 168 13819 169
rect 13785 163 13819 168
rect 13538 145 13727 149
rect 13553 142 13727 145
rect 13546 139 13727 142
rect 13755 162 13819 163
rect 13349 119 13368 121
rect 13383 119 13417 121
rect 13349 103 13429 119
rect 13349 97 13368 103
rect 12716 73 12751 81
rect 12716 47 12717 73
rect 12724 47 12751 73
rect 12716 39 12751 47
rect 12753 73 12794 81
rect 12753 47 12768 73
rect 12775 47 12794 73
rect 12858 69 12889 81
rect 12904 69 13007 81
rect 13019 71 13045 81
rect 13065 71 13168 81
rect 13019 69 13168 71
rect 13189 69 13224 81
rect 12858 67 13020 69
rect 12870 47 12889 67
rect 12904 65 12934 67
rect 12753 39 12794 47
rect 12716 29 12745 39
rect 12759 29 12788 39
rect 12876 29 12889 47
rect 12941 51 13020 67
rect 13052 67 13224 69
rect 13052 51 13131 67
rect 13138 65 13168 67
rect 12941 43 13131 51
rect 13196 47 13202 67
rect 12941 39 13020 43
rect 13022 39 13050 43
rect 13052 39 13131 43
rect 12926 29 12934 39
rect 12953 31 12956 39
rect 12957 31 12975 39
rect 13020 31 13052 39
rect 13097 31 13115 39
rect 12953 29 13119 31
rect 13138 29 13149 39
rect 13211 29 13224 67
rect 13296 81 13325 97
rect 13339 81 13368 97
rect 13383 87 13413 103
rect 13441 81 13447 129
rect 13450 123 13469 129
rect 13484 123 13514 131
rect 13450 115 13514 123
rect 13450 99 13530 115
rect 13546 108 13608 139
rect 13624 108 13686 139
rect 13755 137 13804 162
rect 13819 137 13849 153
rect 13718 123 13748 131
rect 13755 129 13865 137
rect 13718 115 13763 123
rect 13557 105 13561 108
rect 13562 105 13592 108
rect 13450 97 13469 99
rect 13484 97 13530 99
rect 13450 81 13530 97
rect 13561 95 13592 105
rect 13633 105 13639 108
rect 13640 105 13670 108
rect 13633 103 13675 105
rect 13562 92 13592 95
rect 13571 88 13578 92
rect 13578 87 13579 88
rect 13537 81 13547 87
rect 13599 81 13615 97
rect 13640 92 13670 103
rect 13702 99 13764 115
rect 13702 97 13748 99
rect 13702 81 13764 97
rect 13776 81 13782 129
rect 13785 121 13865 129
rect 13785 119 13804 121
rect 13819 119 13853 121
rect 13785 103 13865 119
rect 13785 81 13804 103
rect 13819 87 13849 103
rect 13877 97 13883 171
rect 13886 97 13905 241
rect 13920 97 13926 241
rect 13935 171 13948 241
rect 14000 237 14022 241
rect 13993 215 14022 229
rect 14075 215 14091 229
rect 14129 219 14135 227
rect 14142 225 14250 241
rect 13993 213 14091 215
rect 13977 205 14028 213
rect 14075 205 14109 213
rect 13977 193 14002 205
rect 14009 193 14028 205
rect 14082 203 14109 205
rect 14118 205 14135 219
rect 14180 205 14212 225
rect 14257 219 14263 227
rect 14271 219 14286 241
rect 14352 235 14371 238
rect 14257 213 14286 219
rect 14301 215 14317 229
rect 14352 216 14374 235
rect 14384 229 14400 230
rect 14383 227 14400 229
rect 14384 222 14400 227
rect 14374 215 14380 216
rect 14383 215 14412 222
rect 14301 214 14412 215
rect 14301 213 14418 214
rect 14257 205 14339 213
rect 14374 210 14380 213
rect 14118 203 14339 205
rect 14082 199 14154 203
rect 14182 201 14210 203
rect 13977 185 14028 193
rect 14075 191 14207 199
rect 14210 191 14221 199
rect 14075 189 14154 191
rect 14235 189 14339 203
rect 14383 205 14418 213
rect 14075 185 14172 189
rect 13929 137 13948 171
rect 13993 177 14022 185
rect 13993 171 14010 177
rect 13993 169 14027 171
rect 14075 169 14091 185
rect 14092 181 14172 185
rect 14220 185 14339 189
rect 14220 181 14300 185
rect 14092 175 14300 181
rect 14301 175 14317 185
rect 14365 181 14380 196
rect 14383 193 14384 205
rect 14391 193 14418 205
rect 14383 185 14418 193
rect 14383 184 14412 185
rect 14103 171 14213 175
rect 13994 165 14027 169
rect 13990 163 14027 165
rect 13990 162 14057 163
rect 13990 157 14021 162
rect 14027 157 14057 162
rect 14118 159 14133 171
rect 13990 153 14057 157
rect 13963 150 14057 153
rect 13963 143 14012 150
rect 13963 137 13993 143
rect 14012 138 14017 143
rect 13929 121 14009 137
rect 14021 129 14057 150
rect 14142 149 14172 158
rect 14195 153 14213 171
rect 14271 169 14317 175
rect 14352 171 14365 181
rect 14383 171 14400 184
rect 14352 169 14400 171
rect 14233 163 14235 165
rect 14235 161 14237 163
rect 14237 158 14247 161
rect 14220 151 14250 158
rect 14220 149 14251 151
rect 14271 149 14307 169
rect 14352 168 14399 169
rect 14365 163 14399 168
rect 14118 145 14307 149
rect 14133 142 14307 145
rect 14126 139 14307 142
rect 14335 162 14399 163
rect 13929 119 13948 121
rect 13963 119 13997 121
rect 13929 103 14009 119
rect 13929 97 13948 103
rect 13296 73 13331 81
rect 13296 47 13297 73
rect 13304 47 13331 73
rect 13296 39 13331 47
rect 13333 73 13374 81
rect 13333 47 13348 73
rect 13355 47 13374 73
rect 13438 69 13469 81
rect 13484 69 13587 81
rect 13599 71 13625 81
rect 13645 71 13748 81
rect 13599 69 13748 71
rect 13769 69 13804 81
rect 13438 67 13600 69
rect 13450 47 13469 67
rect 13484 65 13514 67
rect 13333 39 13374 47
rect 13296 29 13325 39
rect 13339 29 13368 39
rect 13456 29 13469 47
rect 13521 51 13600 67
rect 13632 67 13804 69
rect 13632 51 13711 67
rect 13718 65 13748 67
rect 13521 43 13711 51
rect 13776 47 13782 67
rect 13521 39 13600 43
rect 13602 39 13630 43
rect 13632 39 13711 43
rect 13506 29 13514 39
rect 13533 31 13536 39
rect 13537 31 13555 39
rect 13600 31 13632 39
rect 13677 31 13695 39
rect 13533 29 13699 31
rect 13718 29 13729 39
rect 13791 29 13804 67
rect 13876 81 13905 97
rect 13919 81 13948 97
rect 13963 87 13993 103
rect 14021 81 14027 129
rect 14030 123 14049 129
rect 14064 123 14094 131
rect 14030 115 14094 123
rect 14030 99 14110 115
rect 14126 108 14188 139
rect 14204 108 14266 139
rect 14335 137 14384 162
rect 14399 137 14429 153
rect 14298 123 14328 131
rect 14335 129 14445 137
rect 14298 115 14343 123
rect 14137 104 14172 108
rect 14030 97 14049 99
rect 14064 97 14110 99
rect 14030 81 14110 97
rect 14142 92 14172 104
rect 14213 105 14250 108
rect 14213 103 14255 105
rect 14151 88 14158 92
rect 14158 87 14159 88
rect 14117 81 14127 87
rect 13876 73 13911 81
rect 13876 47 13877 73
rect 13884 47 13911 73
rect 13876 39 13911 47
rect 13913 73 13954 81
rect 13913 47 13928 73
rect 13935 47 13954 73
rect 14018 69 14049 81
rect 14064 69 14167 81
rect 14179 80 14196 97
rect 14220 92 14250 103
rect 14282 99 14344 115
rect 14282 97 14328 99
rect 14282 81 14344 97
rect 14356 81 14362 129
rect 14365 121 14445 129
rect 14365 119 14384 121
rect 14399 119 14433 121
rect 14365 103 14445 119
rect 14365 81 14384 103
rect 14399 87 14429 103
rect 14457 97 14463 171
rect 14466 97 14485 241
rect 14500 97 14506 241
rect 14515 171 14528 241
rect 14580 237 14602 241
rect 14573 215 14602 229
rect 14655 215 14671 229
rect 14709 219 14715 227
rect 14722 225 14830 241
rect 14573 213 14671 215
rect 14557 205 14608 213
rect 14655 205 14689 213
rect 14557 193 14582 205
rect 14589 193 14608 205
rect 14662 203 14689 205
rect 14698 205 14715 219
rect 14760 205 14792 225
rect 14837 219 14843 227
rect 14851 219 14866 241
rect 14932 235 14951 238
rect 14837 213 14866 219
rect 14881 215 14897 229
rect 14932 216 14954 235
rect 14964 229 14980 230
rect 14963 227 14980 229
rect 14964 222 14980 227
rect 14954 215 14960 216
rect 14963 215 14992 222
rect 14881 214 14992 215
rect 14881 213 14998 214
rect 14837 205 14919 213
rect 14954 210 14960 213
rect 14698 203 14919 205
rect 14662 199 14734 203
rect 14762 201 14790 203
rect 14557 185 14608 193
rect 14655 191 14787 199
rect 14790 191 14801 199
rect 14655 189 14734 191
rect 14815 189 14919 203
rect 14963 205 14998 213
rect 14655 185 14752 189
rect 14509 137 14528 171
rect 14573 177 14602 185
rect 14573 171 14590 177
rect 14573 169 14607 171
rect 14655 169 14671 185
rect 14672 181 14752 185
rect 14800 185 14919 189
rect 14800 181 14880 185
rect 14672 175 14880 181
rect 14881 175 14897 185
rect 14945 181 14960 196
rect 14963 193 14964 205
rect 14971 193 14998 205
rect 14963 185 14998 193
rect 14963 184 14992 185
rect 14683 171 14793 175
rect 14574 165 14607 169
rect 14570 163 14607 165
rect 14570 162 14637 163
rect 14570 157 14601 162
rect 14607 157 14637 162
rect 14698 159 14713 171
rect 14570 153 14637 157
rect 14543 150 14637 153
rect 14543 143 14592 150
rect 14543 137 14573 143
rect 14592 138 14597 143
rect 14509 121 14589 137
rect 14601 129 14637 150
rect 14722 149 14752 158
rect 14775 153 14793 171
rect 14851 169 14897 175
rect 14932 171 14945 181
rect 14963 171 14980 184
rect 14932 169 14980 171
rect 14813 163 14815 165
rect 14815 161 14817 163
rect 14817 158 14827 161
rect 14800 151 14830 158
rect 14800 149 14831 151
rect 14851 149 14887 169
rect 14932 168 14979 169
rect 14945 163 14979 168
rect 14698 145 14887 149
rect 14713 142 14887 145
rect 14706 139 14887 142
rect 14915 162 14979 163
rect 14509 119 14528 121
rect 14543 119 14577 121
rect 14509 103 14589 119
rect 14509 97 14528 103
rect 14179 71 14205 80
rect 14225 71 14328 81
rect 14179 69 14328 71
rect 14349 69 14384 81
rect 14018 67 14180 69
rect 14030 47 14049 67
rect 14064 65 14094 67
rect 13913 39 13954 47
rect 13876 29 13905 39
rect 13919 29 13948 39
rect 14036 29 14049 47
rect 14101 51 14180 67
rect 14212 67 14384 69
rect 14212 51 14291 67
rect 14298 65 14328 67
rect 14101 43 14291 51
rect 14356 47 14362 67
rect 14101 39 14180 43
rect 14182 39 14210 43
rect 14212 39 14291 43
rect 14086 29 14094 39
rect 14113 31 14116 39
rect 14117 31 14135 39
rect 14180 31 14212 39
rect 14257 31 14275 39
rect 14113 29 14279 31
rect 14298 29 14309 39
rect 14371 29 14384 67
rect 14456 81 14485 97
rect 14499 81 14528 97
rect 14543 87 14573 103
rect 14601 81 14607 129
rect 14610 123 14629 129
rect 14644 123 14674 131
rect 14610 115 14674 123
rect 14610 99 14690 115
rect 14706 108 14768 139
rect 14784 108 14846 139
rect 14915 137 14964 162
rect 14979 137 15009 153
rect 14878 123 14908 131
rect 14915 129 15025 137
rect 14878 115 14923 123
rect 14717 104 14752 108
rect 14610 97 14629 99
rect 14644 97 14690 99
rect 14610 81 14690 97
rect 14722 92 14752 104
rect 14793 105 14830 108
rect 14793 103 14835 105
rect 14731 88 14738 92
rect 14738 87 14739 88
rect 14697 81 14707 87
rect 14456 69 14491 81
rect 14493 69 14534 81
rect 14456 39 14534 69
rect 14598 69 14629 81
rect 14644 69 14747 81
rect 14759 80 14776 97
rect 14800 92 14830 103
rect 14862 99 14924 115
rect 14862 97 14908 99
rect 14862 81 14924 97
rect 14936 81 14942 129
rect 14945 121 15025 129
rect 14945 119 14964 121
rect 14979 119 15013 121
rect 14945 103 15025 119
rect 14945 81 14964 103
rect 14979 87 15009 103
rect 15037 97 15043 171
rect 15046 97 15065 241
rect 15080 97 15086 241
rect 15095 171 15108 241
rect 15160 237 15182 241
rect 15153 215 15182 229
rect 15235 215 15251 229
rect 15289 219 15295 227
rect 15302 225 15410 241
rect 15153 213 15251 215
rect 15137 205 15188 213
rect 15235 205 15269 213
rect 15137 193 15162 205
rect 15169 193 15188 205
rect 15242 203 15269 205
rect 15278 205 15295 219
rect 15340 205 15372 225
rect 15417 219 15423 227
rect 15431 219 15446 241
rect 15512 235 15531 238
rect 15417 213 15446 219
rect 15461 215 15477 229
rect 15512 216 15534 235
rect 15544 229 15560 230
rect 15543 227 15560 229
rect 15544 222 15560 227
rect 15534 215 15540 216
rect 15543 215 15572 222
rect 15461 214 15572 215
rect 15461 213 15578 214
rect 15417 205 15499 213
rect 15534 210 15540 213
rect 15278 203 15499 205
rect 15242 199 15314 203
rect 15342 201 15370 203
rect 15137 185 15188 193
rect 15235 191 15367 199
rect 15370 191 15381 199
rect 15235 189 15314 191
rect 15395 189 15499 203
rect 15543 205 15578 213
rect 15235 185 15332 189
rect 15089 137 15108 171
rect 15153 177 15182 185
rect 15153 171 15170 177
rect 15153 169 15187 171
rect 15235 169 15251 185
rect 15252 181 15332 185
rect 15380 185 15499 189
rect 15380 181 15460 185
rect 15252 175 15460 181
rect 15461 175 15477 185
rect 15525 181 15540 196
rect 15543 193 15544 205
rect 15551 193 15578 205
rect 15543 185 15578 193
rect 15543 184 15572 185
rect 15263 171 15373 175
rect 15154 165 15187 169
rect 15150 163 15187 165
rect 15150 162 15217 163
rect 15150 157 15181 162
rect 15187 157 15217 162
rect 15278 159 15293 171
rect 15150 153 15217 157
rect 15123 150 15217 153
rect 15123 143 15172 150
rect 15123 137 15153 143
rect 15172 138 15177 143
rect 15089 121 15169 137
rect 15181 129 15217 150
rect 15302 149 15332 158
rect 15355 153 15373 171
rect 15431 169 15477 175
rect 15512 171 15525 181
rect 15543 171 15560 184
rect 15512 169 15560 171
rect 15393 163 15395 165
rect 15395 161 15397 163
rect 15397 158 15407 161
rect 15380 151 15410 158
rect 15380 149 15411 151
rect 15431 149 15467 169
rect 15512 168 15559 169
rect 15525 163 15559 168
rect 15278 145 15467 149
rect 15293 142 15467 145
rect 15286 139 15467 142
rect 15495 162 15559 163
rect 15089 119 15108 121
rect 15123 119 15157 121
rect 15089 103 15169 119
rect 15089 97 15108 103
rect 14759 71 14785 80
rect 14805 71 14908 81
rect 14759 69 14908 71
rect 14929 69 14964 81
rect 14598 67 14760 69
rect 14610 47 14629 67
rect 14644 65 14674 67
rect 14456 38 14491 39
rect 14499 38 14534 39
rect 14456 29 14485 38
rect 14499 29 14528 38
rect 14616 29 14629 47
rect 14681 51 14760 67
rect 14792 67 14964 69
rect 14792 51 14871 67
rect 14878 65 14908 67
rect 14681 43 14871 51
rect 14936 47 14942 67
rect 14681 39 14760 43
rect 14762 39 14790 43
rect 14792 39 14871 43
rect 14666 29 14674 39
rect 14693 31 14696 39
rect 14697 31 14715 39
rect 14760 31 14792 39
rect 14837 31 14855 39
rect 14693 29 14859 31
rect 14878 29 14889 39
rect 14951 29 14964 67
rect 15036 81 15065 97
rect 15079 81 15108 97
rect 15123 87 15153 103
rect 15181 81 15187 129
rect 15190 123 15209 129
rect 15224 123 15254 131
rect 15190 115 15254 123
rect 15190 99 15270 115
rect 15286 108 15348 139
rect 15364 108 15426 139
rect 15495 137 15544 162
rect 15559 137 15589 153
rect 15458 123 15488 131
rect 15495 129 15605 137
rect 15458 115 15503 123
rect 15297 104 15332 108
rect 15190 97 15209 99
rect 15224 97 15270 99
rect 15190 81 15270 97
rect 15302 92 15332 104
rect 15373 105 15410 108
rect 15373 103 15415 105
rect 15311 88 15318 92
rect 15318 87 15319 88
rect 15277 81 15287 87
rect 15036 69 15071 81
rect 15073 69 15114 81
rect 15036 39 15114 69
rect 15178 69 15209 81
rect 15224 69 15327 81
rect 15339 80 15356 97
rect 15380 92 15410 103
rect 15442 99 15504 115
rect 15442 97 15488 99
rect 15442 81 15504 97
rect 15516 81 15522 129
rect 15525 121 15605 129
rect 15525 119 15544 121
rect 15559 119 15593 121
rect 15525 103 15605 119
rect 15525 81 15544 103
rect 15559 87 15589 103
rect 15617 97 15623 171
rect 15626 97 15645 241
rect 15660 97 15666 241
rect 15675 171 15688 241
rect 15740 237 15762 241
rect 15733 215 15762 229
rect 15815 215 15831 229
rect 15869 219 15875 227
rect 15882 225 15990 241
rect 15733 213 15831 215
rect 15717 205 15768 213
rect 15815 205 15849 213
rect 15717 193 15742 205
rect 15749 193 15768 205
rect 15822 203 15849 205
rect 15858 205 15875 219
rect 15920 205 15952 225
rect 15997 219 16003 227
rect 16011 219 16026 241
rect 16092 235 16111 238
rect 15997 213 16026 219
rect 16041 215 16057 229
rect 16092 216 16114 235
rect 16124 229 16140 230
rect 16123 227 16140 229
rect 16124 222 16140 227
rect 16114 215 16120 216
rect 16123 215 16152 222
rect 16041 214 16152 215
rect 16041 213 16158 214
rect 15997 205 16079 213
rect 16114 210 16120 213
rect 15858 203 16079 205
rect 15822 199 15894 203
rect 15922 201 15950 203
rect 15717 185 15768 193
rect 15815 191 15947 199
rect 15950 191 15961 199
rect 15815 189 15894 191
rect 15975 189 16079 203
rect 16123 205 16158 213
rect 15815 185 15912 189
rect 15669 137 15688 171
rect 15733 177 15762 185
rect 15733 171 15750 177
rect 15733 169 15767 171
rect 15815 169 15831 185
rect 15832 181 15912 185
rect 15960 185 16079 189
rect 15960 181 16040 185
rect 15832 175 16040 181
rect 16041 175 16057 185
rect 16105 181 16120 196
rect 16123 193 16124 205
rect 16131 193 16158 205
rect 16123 185 16158 193
rect 16123 184 16152 185
rect 15843 171 15953 175
rect 15734 165 15767 169
rect 15730 163 15767 165
rect 15730 162 15797 163
rect 15730 157 15761 162
rect 15767 157 15797 162
rect 15858 159 15873 171
rect 15730 153 15797 157
rect 15703 150 15797 153
rect 15703 143 15752 150
rect 15703 137 15733 143
rect 15752 138 15757 143
rect 15669 121 15749 137
rect 15761 129 15797 150
rect 15882 149 15912 158
rect 15935 153 15953 171
rect 16011 169 16057 175
rect 16092 171 16105 181
rect 16123 171 16140 184
rect 16092 169 16140 171
rect 15973 163 15975 165
rect 15975 161 15977 163
rect 15977 158 15987 161
rect 15960 151 15990 158
rect 15960 149 15991 151
rect 16011 149 16047 169
rect 16092 168 16139 169
rect 16105 163 16139 168
rect 15858 145 16047 149
rect 15873 142 16047 145
rect 15866 139 16047 142
rect 16075 162 16139 163
rect 15669 119 15688 121
rect 15703 119 15737 121
rect 15669 103 15749 119
rect 15669 97 15688 103
rect 15339 71 15365 80
rect 15385 71 15488 81
rect 15339 69 15488 71
rect 15509 69 15544 81
rect 15178 67 15340 69
rect 15190 47 15209 67
rect 15224 65 15254 67
rect 15036 38 15071 39
rect 15079 38 15114 39
rect 15036 29 15065 38
rect 15079 29 15108 38
rect 15196 29 15209 47
rect 15261 51 15340 67
rect 15372 67 15544 69
rect 15372 51 15451 67
rect 15458 65 15488 67
rect 15261 43 15451 51
rect 15516 47 15522 67
rect 15261 39 15340 43
rect 15342 39 15370 43
rect 15372 39 15451 43
rect 15246 29 15254 39
rect 15273 31 15276 39
rect 15277 31 15295 39
rect 15340 31 15372 39
rect 15417 31 15435 39
rect 15273 29 15439 31
rect 15458 29 15469 39
rect 15531 29 15544 67
rect 15616 81 15645 97
rect 15659 81 15688 97
rect 15703 87 15733 103
rect 15761 81 15767 129
rect 15770 123 15789 129
rect 15804 123 15834 131
rect 15770 115 15834 123
rect 15770 99 15850 115
rect 15866 108 15928 139
rect 15944 108 16006 139
rect 16075 137 16124 162
rect 16139 137 16169 153
rect 16038 123 16068 131
rect 16075 129 16185 137
rect 16038 115 16083 123
rect 15877 104 15912 108
rect 15770 97 15789 99
rect 15804 97 15850 99
rect 15770 81 15850 97
rect 15882 92 15912 104
rect 15953 105 15990 108
rect 15953 103 15995 105
rect 15891 88 15898 92
rect 15898 87 15899 88
rect 15857 81 15867 87
rect 15616 69 15651 81
rect 15653 69 15694 81
rect 15616 39 15694 69
rect 15758 69 15789 81
rect 15804 69 15907 81
rect 15919 80 15936 97
rect 15960 92 15990 103
rect 16022 99 16084 115
rect 16022 97 16068 99
rect 16022 81 16084 97
rect 16096 81 16102 129
rect 16105 121 16185 129
rect 16105 119 16124 121
rect 16139 119 16173 121
rect 16105 103 16185 119
rect 16105 81 16124 103
rect 16139 87 16169 103
rect 16197 97 16203 171
rect 16206 97 16225 241
rect 16240 97 16246 241
rect 16255 171 16268 241
rect 16320 237 16342 241
rect 16313 215 16342 229
rect 16395 215 16411 229
rect 16449 219 16455 227
rect 16462 225 16570 241
rect 16313 213 16411 215
rect 16297 205 16348 213
rect 16395 205 16429 213
rect 16297 193 16322 205
rect 16329 193 16348 205
rect 16402 203 16429 205
rect 16438 205 16455 219
rect 16500 205 16532 225
rect 16577 219 16583 227
rect 16591 219 16606 241
rect 16672 235 16691 238
rect 16577 213 16606 219
rect 16621 215 16637 229
rect 16672 216 16694 235
rect 16704 229 16720 230
rect 16703 227 16720 229
rect 16704 222 16720 227
rect 16694 215 16700 216
rect 16703 215 16732 222
rect 16621 214 16732 215
rect 16621 213 16738 214
rect 16577 205 16659 213
rect 16694 210 16700 213
rect 16438 203 16659 205
rect 16402 199 16474 203
rect 16502 201 16530 203
rect 16297 185 16348 193
rect 16395 191 16527 199
rect 16530 191 16541 199
rect 16395 189 16474 191
rect 16555 189 16659 203
rect 16703 205 16738 213
rect 16395 185 16492 189
rect 16249 137 16268 171
rect 16313 177 16342 185
rect 16313 171 16330 177
rect 16313 169 16347 171
rect 16395 169 16411 185
rect 16412 181 16492 185
rect 16540 185 16659 189
rect 16540 181 16620 185
rect 16412 175 16620 181
rect 16621 175 16637 185
rect 16685 181 16700 196
rect 16703 193 16704 205
rect 16711 193 16738 205
rect 16703 185 16738 193
rect 16703 184 16732 185
rect 16423 171 16533 175
rect 16314 165 16347 169
rect 16310 163 16347 165
rect 16310 162 16377 163
rect 16310 157 16341 162
rect 16347 157 16377 162
rect 16438 159 16453 171
rect 16310 153 16377 157
rect 16283 150 16377 153
rect 16283 143 16332 150
rect 16283 137 16313 143
rect 16332 138 16337 143
rect 16249 121 16329 137
rect 16341 129 16377 150
rect 16462 149 16492 158
rect 16515 153 16533 171
rect 16591 169 16637 175
rect 16672 171 16685 181
rect 16703 171 16720 184
rect 16672 169 16720 171
rect 16553 163 16555 165
rect 16555 161 16557 163
rect 16557 158 16567 161
rect 16540 151 16570 158
rect 16540 149 16571 151
rect 16591 149 16627 169
rect 16672 168 16719 169
rect 16685 163 16719 168
rect 16438 145 16627 149
rect 16453 142 16627 145
rect 16446 139 16627 142
rect 16655 162 16719 163
rect 16249 119 16268 121
rect 16283 119 16317 121
rect 16249 103 16329 119
rect 16249 97 16268 103
rect 15919 71 15945 80
rect 15965 71 16068 81
rect 15919 69 16068 71
rect 16089 69 16124 81
rect 15758 67 15920 69
rect 15770 47 15789 67
rect 15804 65 15834 67
rect 15616 38 15651 39
rect 15659 38 15694 39
rect 15616 29 15645 38
rect 15659 29 15688 38
rect 15776 29 15789 47
rect 15841 51 15920 67
rect 15952 67 16124 69
rect 15952 51 16031 67
rect 16038 65 16068 67
rect 15841 43 16031 51
rect 16096 47 16102 67
rect 15841 39 15920 43
rect 15922 39 15950 43
rect 15952 39 16031 43
rect 15826 29 15834 39
rect 15853 31 15856 39
rect 15857 31 15875 39
rect 15920 31 15952 39
rect 15997 31 16015 39
rect 15853 29 16019 31
rect 16038 29 16049 39
rect 16111 29 16124 67
rect 16196 81 16225 97
rect 16239 81 16268 97
rect 16283 87 16313 103
rect 16341 81 16347 129
rect 16350 123 16369 129
rect 16384 123 16414 131
rect 16350 115 16414 123
rect 16350 99 16430 115
rect 16446 108 16508 139
rect 16524 108 16586 139
rect 16655 137 16704 162
rect 16719 137 16749 153
rect 16618 123 16648 131
rect 16655 129 16765 137
rect 16618 115 16663 123
rect 16457 104 16492 108
rect 16350 97 16369 99
rect 16384 97 16430 99
rect 16350 81 16430 97
rect 16462 92 16492 104
rect 16533 105 16570 108
rect 16533 103 16575 105
rect 16471 88 16478 92
rect 16478 87 16479 88
rect 16437 81 16447 87
rect 16196 69 16231 81
rect 16233 69 16274 81
rect 16196 39 16274 69
rect 16338 69 16369 81
rect 16384 69 16487 81
rect 16499 80 16516 97
rect 16540 92 16570 103
rect 16602 99 16664 115
rect 16602 97 16648 99
rect 16602 81 16664 97
rect 16676 81 16682 129
rect 16685 121 16765 129
rect 16685 119 16704 121
rect 16719 119 16753 121
rect 16685 103 16765 119
rect 16685 81 16704 103
rect 16719 87 16749 103
rect 16777 97 16783 171
rect 16786 97 16805 241
rect 16820 97 16826 241
rect 16835 171 16848 241
rect 16900 237 16922 241
rect 16893 215 16922 229
rect 16975 215 16991 229
rect 17029 219 17035 227
rect 17042 225 17150 241
rect 16893 213 16991 215
rect 16877 205 16928 213
rect 16975 205 17009 213
rect 16877 193 16902 205
rect 16909 193 16928 205
rect 16982 203 17009 205
rect 17018 205 17035 219
rect 17080 205 17112 225
rect 17157 219 17163 227
rect 17171 219 17186 241
rect 17252 235 17271 238
rect 17157 213 17186 219
rect 17201 215 17217 229
rect 17252 216 17274 235
rect 17284 229 17300 230
rect 17283 227 17300 229
rect 17284 222 17300 227
rect 17274 215 17280 216
rect 17283 215 17312 222
rect 17201 214 17312 215
rect 17201 213 17318 214
rect 17157 205 17239 213
rect 17274 210 17280 213
rect 17018 203 17239 205
rect 16982 199 17054 203
rect 17082 201 17110 203
rect 16877 185 16928 193
rect 16975 191 17107 199
rect 17110 191 17121 199
rect 16975 189 17054 191
rect 17135 189 17239 203
rect 17283 205 17318 213
rect 16975 185 17072 189
rect 16829 137 16848 171
rect 16893 177 16922 185
rect 16893 171 16910 177
rect 16893 169 16927 171
rect 16975 169 16991 185
rect 16992 181 17072 185
rect 17120 185 17239 189
rect 17120 181 17200 185
rect 16992 175 17200 181
rect 17201 175 17217 185
rect 17265 181 17280 196
rect 17283 193 17284 205
rect 17291 193 17318 205
rect 17283 185 17318 193
rect 17283 184 17312 185
rect 17003 171 17113 175
rect 16894 165 16927 169
rect 16890 163 16927 165
rect 16890 162 16957 163
rect 16890 157 16921 162
rect 16927 157 16957 162
rect 17018 159 17033 171
rect 16890 153 16957 157
rect 16863 150 16957 153
rect 16863 143 16912 150
rect 16863 137 16893 143
rect 16912 138 16917 143
rect 16829 121 16909 137
rect 16921 129 16957 150
rect 17042 149 17072 158
rect 17095 153 17113 171
rect 17171 169 17217 175
rect 17252 171 17265 181
rect 17283 171 17300 184
rect 17252 169 17300 171
rect 17133 163 17135 165
rect 17135 161 17137 163
rect 17137 158 17147 161
rect 17120 151 17150 158
rect 17120 149 17151 151
rect 17171 149 17207 169
rect 17252 168 17299 169
rect 17265 163 17299 168
rect 17018 145 17207 149
rect 17033 142 17207 145
rect 17026 139 17207 142
rect 17235 162 17299 163
rect 16829 119 16848 121
rect 16863 119 16897 121
rect 16829 103 16909 119
rect 16829 97 16848 103
rect 16499 71 16525 80
rect 16545 71 16648 81
rect 16499 69 16648 71
rect 16669 69 16704 81
rect 16338 67 16500 69
rect 16350 47 16369 67
rect 16384 65 16414 67
rect 16196 38 16231 39
rect 16239 38 16274 39
rect 16196 29 16225 38
rect 16239 29 16268 38
rect 16356 29 16369 47
rect 16421 51 16500 67
rect 16532 67 16704 69
rect 16532 51 16611 67
rect 16618 65 16648 67
rect 16421 43 16611 51
rect 16676 47 16682 67
rect 16421 39 16500 43
rect 16502 39 16530 43
rect 16532 39 16611 43
rect 16406 29 16414 39
rect 16433 31 16436 39
rect 16437 31 16455 39
rect 16500 31 16532 39
rect 16577 31 16595 39
rect 16433 29 16599 31
rect 16618 29 16629 39
rect 16691 29 16704 67
rect 16776 81 16805 97
rect 16819 81 16848 97
rect 16863 87 16893 103
rect 16921 81 16927 129
rect 16930 123 16949 129
rect 16964 123 16994 131
rect 16930 115 16994 123
rect 16930 99 17010 115
rect 17026 108 17088 139
rect 17104 108 17166 139
rect 17235 137 17284 162
rect 17299 137 17329 153
rect 17198 123 17228 131
rect 17235 129 17345 137
rect 17198 115 17243 123
rect 17037 104 17072 108
rect 16930 97 16949 99
rect 16964 97 17010 99
rect 16930 81 17010 97
rect 17042 92 17072 104
rect 17113 105 17150 108
rect 17113 103 17155 105
rect 17051 88 17058 92
rect 17058 87 17059 88
rect 17017 81 17027 87
rect 16776 69 16811 81
rect 16813 69 16854 81
rect 16776 39 16854 69
rect 16918 69 16949 81
rect 16964 69 17067 81
rect 17079 80 17096 97
rect 17120 92 17150 103
rect 17182 99 17244 115
rect 17182 97 17228 99
rect 17182 81 17244 97
rect 17256 81 17262 129
rect 17265 121 17345 129
rect 17265 119 17284 121
rect 17299 119 17333 121
rect 17265 103 17345 119
rect 17265 81 17284 103
rect 17299 87 17329 103
rect 17357 97 17363 171
rect 17366 97 17385 241
rect 17400 97 17406 241
rect 17415 171 17428 241
rect 17480 237 17502 241
rect 17473 215 17502 229
rect 17555 215 17571 229
rect 17609 219 17615 227
rect 17622 225 17730 241
rect 17473 213 17571 215
rect 17457 205 17508 213
rect 17555 205 17589 213
rect 17457 193 17482 205
rect 17489 193 17508 205
rect 17562 203 17589 205
rect 17598 205 17615 219
rect 17660 205 17692 225
rect 17737 219 17743 227
rect 17751 219 17766 241
rect 17832 235 17851 238
rect 17737 213 17766 219
rect 17781 215 17797 229
rect 17832 216 17854 235
rect 17864 229 17880 230
rect 17863 227 17880 229
rect 17864 222 17880 227
rect 17854 215 17860 216
rect 17863 215 17892 222
rect 17781 214 17892 215
rect 17781 213 17898 214
rect 17737 205 17819 213
rect 17854 210 17860 213
rect 17598 203 17819 205
rect 17562 199 17634 203
rect 17662 201 17690 203
rect 17457 185 17508 193
rect 17555 191 17687 199
rect 17690 191 17701 199
rect 17555 189 17634 191
rect 17715 189 17819 203
rect 17863 205 17898 213
rect 17555 185 17652 189
rect 17409 137 17428 171
rect 17473 177 17502 185
rect 17473 171 17490 177
rect 17473 169 17507 171
rect 17555 169 17571 185
rect 17572 181 17652 185
rect 17700 185 17819 189
rect 17700 181 17780 185
rect 17572 175 17780 181
rect 17781 175 17797 185
rect 17845 181 17860 196
rect 17863 193 17864 205
rect 17871 193 17898 205
rect 17863 185 17898 193
rect 17863 184 17892 185
rect 17583 171 17693 175
rect 17474 165 17507 169
rect 17470 163 17507 165
rect 17470 162 17537 163
rect 17470 157 17501 162
rect 17507 157 17537 162
rect 17598 159 17613 171
rect 17470 153 17537 157
rect 17443 150 17537 153
rect 17443 143 17492 150
rect 17443 137 17473 143
rect 17492 138 17497 143
rect 17409 121 17489 137
rect 17501 129 17537 150
rect 17622 149 17652 158
rect 17675 153 17693 171
rect 17751 169 17797 175
rect 17832 171 17845 181
rect 17863 171 17880 184
rect 17832 169 17880 171
rect 17713 163 17715 165
rect 17715 161 17717 163
rect 17717 158 17727 161
rect 17700 151 17730 158
rect 17700 149 17731 151
rect 17751 149 17787 169
rect 17832 168 17879 169
rect 17845 163 17879 168
rect 17598 145 17787 149
rect 17613 142 17787 145
rect 17606 139 17787 142
rect 17815 162 17879 163
rect 17409 119 17428 121
rect 17443 119 17477 121
rect 17409 103 17489 119
rect 17409 97 17428 103
rect 17079 71 17105 80
rect 17125 71 17228 81
rect 17079 69 17228 71
rect 17249 69 17284 81
rect 16918 67 17080 69
rect 16930 47 16949 67
rect 16964 65 16994 67
rect 16776 38 16811 39
rect 16819 38 16854 39
rect 16776 29 16805 38
rect 16819 29 16848 38
rect 16936 29 16949 47
rect 17001 51 17080 67
rect 17112 67 17284 69
rect 17112 51 17191 67
rect 17198 65 17228 67
rect 17001 43 17191 51
rect 17256 47 17262 67
rect 17001 39 17080 43
rect 17082 39 17110 43
rect 17112 39 17191 43
rect 16986 29 16994 39
rect 17013 31 17016 39
rect 17017 31 17035 39
rect 17080 31 17112 39
rect 17157 31 17175 39
rect 17013 29 17179 31
rect 17198 29 17209 39
rect 17271 29 17284 67
rect 17356 81 17385 97
rect 17399 81 17428 97
rect 17443 87 17473 103
rect 17501 81 17507 129
rect 17510 123 17529 129
rect 17544 123 17574 131
rect 17510 115 17574 123
rect 17510 99 17590 115
rect 17606 108 17668 139
rect 17684 108 17746 139
rect 17815 137 17864 162
rect 17879 137 17909 153
rect 17778 123 17808 131
rect 17815 129 17925 137
rect 17778 115 17823 123
rect 17617 104 17652 108
rect 17510 97 17529 99
rect 17544 97 17590 99
rect 17510 81 17590 97
rect 17622 92 17652 104
rect 17693 105 17730 108
rect 17693 103 17735 105
rect 17631 88 17638 92
rect 17638 87 17639 88
rect 17597 81 17607 87
rect 17356 69 17391 81
rect 17393 69 17434 81
rect 17356 39 17434 69
rect 17498 69 17529 81
rect 17544 69 17647 81
rect 17659 80 17676 97
rect 17700 92 17730 103
rect 17762 99 17824 115
rect 17762 97 17808 99
rect 17762 81 17824 97
rect 17836 81 17842 129
rect 17845 121 17925 129
rect 17845 119 17864 121
rect 17879 119 17913 121
rect 17845 103 17925 119
rect 17845 81 17864 103
rect 17879 87 17909 103
rect 17937 97 17943 171
rect 17946 97 17965 241
rect 17980 97 17986 241
rect 17995 171 18008 241
rect 18060 237 18082 241
rect 18053 215 18082 229
rect 18135 215 18151 229
rect 18189 219 18195 227
rect 18202 225 18310 241
rect 18053 213 18151 215
rect 18037 205 18088 213
rect 18135 205 18169 213
rect 18037 193 18062 205
rect 18069 193 18088 205
rect 18142 203 18169 205
rect 18178 205 18195 219
rect 18240 205 18272 225
rect 18317 219 18323 227
rect 18331 219 18346 241
rect 18412 235 18431 238
rect 18317 213 18346 219
rect 18361 215 18377 229
rect 18412 216 18434 235
rect 18444 229 18460 230
rect 18443 227 18460 229
rect 18444 222 18460 227
rect 18434 215 18440 216
rect 18443 215 18472 222
rect 18361 214 18472 215
rect 18361 213 18478 214
rect 18317 205 18399 213
rect 18434 210 18440 213
rect 18178 203 18399 205
rect 18142 199 18214 203
rect 18242 201 18270 203
rect 18037 185 18088 193
rect 18135 191 18267 199
rect 18270 191 18281 199
rect 18135 189 18214 191
rect 18295 189 18399 203
rect 18443 205 18478 213
rect 18135 185 18232 189
rect 17989 137 18008 171
rect 18053 177 18082 185
rect 18053 171 18070 177
rect 18053 169 18087 171
rect 18135 169 18151 185
rect 18152 181 18232 185
rect 18280 185 18399 189
rect 18280 181 18360 185
rect 18152 175 18360 181
rect 18361 175 18377 185
rect 18425 181 18440 196
rect 18443 193 18444 205
rect 18451 193 18478 205
rect 18443 185 18478 193
rect 18443 184 18472 185
rect 18163 171 18273 175
rect 18054 165 18087 169
rect 18050 163 18087 165
rect 18050 162 18117 163
rect 18050 157 18081 162
rect 18087 157 18117 162
rect 18178 159 18193 171
rect 18050 153 18117 157
rect 18023 150 18117 153
rect 18023 143 18072 150
rect 18023 137 18053 143
rect 18072 138 18077 143
rect 17989 121 18069 137
rect 18081 129 18117 150
rect 18202 149 18232 158
rect 18255 153 18273 171
rect 18331 169 18377 175
rect 18412 171 18425 181
rect 18443 171 18460 184
rect 18412 169 18460 171
rect 18293 163 18295 165
rect 18295 161 18297 163
rect 18297 158 18307 161
rect 18280 151 18310 158
rect 18280 149 18311 151
rect 18331 149 18367 169
rect 18412 168 18459 169
rect 18425 163 18459 168
rect 18178 145 18367 149
rect 18193 142 18367 145
rect 18186 139 18367 142
rect 18395 162 18459 163
rect 17989 119 18008 121
rect 18023 119 18057 121
rect 17989 103 18069 119
rect 17989 97 18008 103
rect 17659 71 17685 80
rect 17705 71 17808 81
rect 17659 69 17808 71
rect 17829 69 17864 81
rect 17498 67 17660 69
rect 17510 47 17529 67
rect 17544 65 17574 67
rect 17356 38 17391 39
rect 17399 38 17434 39
rect 17356 29 17385 38
rect 17399 29 17428 38
rect 17516 29 17529 47
rect 17581 51 17660 67
rect 17692 67 17864 69
rect 17692 51 17771 67
rect 17778 65 17808 67
rect 17581 43 17771 51
rect 17836 47 17842 67
rect 17581 39 17660 43
rect 17662 39 17690 43
rect 17692 39 17771 43
rect 17566 29 17574 39
rect 17593 31 17596 39
rect 17597 31 17615 39
rect 17660 31 17692 39
rect 17737 31 17755 39
rect 17593 29 17759 31
rect 17778 29 17789 39
rect 17851 29 17864 67
rect 17936 81 17965 97
rect 17979 81 18008 97
rect 18023 87 18053 103
rect 18081 81 18087 129
rect 18090 123 18109 129
rect 18124 123 18154 131
rect 18090 115 18154 123
rect 18090 99 18170 115
rect 18186 108 18248 139
rect 18264 108 18326 139
rect 18395 137 18444 162
rect 18459 137 18489 153
rect 18358 123 18388 131
rect 18395 129 18505 137
rect 18358 115 18403 123
rect 18197 104 18232 108
rect 18090 97 18109 99
rect 18124 97 18170 99
rect 18090 81 18170 97
rect 18202 92 18232 104
rect 18273 105 18310 108
rect 18273 103 18315 105
rect 18211 88 18218 92
rect 18218 87 18219 88
rect 18177 81 18187 87
rect 17936 69 17971 81
rect 17973 69 18014 81
rect 17936 39 18014 69
rect 18078 69 18109 81
rect 18124 69 18227 81
rect 18239 80 18256 97
rect 18280 92 18310 103
rect 18342 99 18404 115
rect 18342 97 18388 99
rect 18342 81 18404 97
rect 18416 81 18422 129
rect 18425 121 18505 129
rect 18425 119 18444 121
rect 18459 119 18493 121
rect 18425 103 18505 119
rect 18425 81 18444 103
rect 18459 87 18489 103
rect 18517 97 18523 171
rect 18532 97 18545 241
rect 18239 71 18265 80
rect 18285 71 18388 81
rect 18239 69 18388 71
rect 18409 69 18444 81
rect 18078 67 18240 69
rect 18090 47 18109 67
rect 18124 65 18154 67
rect 17936 38 17971 39
rect 17979 38 18014 39
rect 17936 29 17965 38
rect 17979 29 18008 38
rect 18096 29 18109 47
rect 18161 51 18240 67
rect 18272 67 18444 69
rect 18272 51 18351 67
rect 18358 65 18388 67
rect 18161 43 18351 51
rect 18416 47 18422 67
rect 18161 39 18240 43
rect 18242 39 18270 43
rect 18272 39 18351 43
rect 18146 29 18154 39
rect 18173 31 18176 39
rect 18177 31 18195 39
rect 18240 31 18272 39
rect 18317 31 18335 39
rect 18173 29 18339 31
rect 18358 29 18369 39
rect 18431 29 18444 67
rect 18516 81 18545 97
rect 18516 38 18551 81
rect 18516 29 18545 38
rect 4596 28 18545 29
rect -1 22 18545 28
rect 0 15 18545 22
rect 0 14 4631 15
rect 15 0 28 14
rect 43 -4 73 14
rect 116 0 159 14
rect 166 1 174 14
rect 207 1 345 14
rect 378 1 386 14
rect 129 -18 159 0
rect 222 -2 330 1
rect 222 -4 252 -2
rect 300 -4 330 -2
rect 393 -18 423 14
rect 451 0 464 14
rect 479 -4 509 14
rect 546 0 565 14
rect 580 0 586 14
rect 595 0 608 14
rect 623 -4 653 14
rect 696 0 739 14
rect 746 1 754 14
rect 787 1 925 14
rect 958 1 966 14
rect 709 -18 739 0
rect 802 -2 910 1
rect 802 -4 832 -2
rect 880 -4 910 -2
rect 973 -18 1003 14
rect 1031 0 1044 14
rect 1059 -4 1089 14
rect 1126 0 1145 14
rect 1160 0 1166 14
rect 1175 0 1188 14
rect 1203 -4 1233 14
rect 1276 0 1319 14
rect 1326 1 1334 14
rect 1367 1 1505 14
rect 1538 1 1546 14
rect 1289 -18 1319 0
rect 1382 -2 1490 1
rect 1382 -4 1412 -2
rect 1460 -4 1490 -2
rect 1553 -18 1583 14
rect 1611 0 1624 14
rect 1639 -4 1669 14
rect 1706 0 1725 14
rect 1740 0 1746 14
rect 1755 0 1768 14
rect 1783 -4 1813 14
rect 1856 0 1899 14
rect 1906 1 1914 14
rect 1947 1 2085 14
rect 2118 1 2126 14
rect 1869 -18 1899 0
rect 1962 -2 2070 1
rect 1962 -4 1992 -2
rect 2040 -4 2070 -2
rect 2133 -18 2163 14
rect 2191 0 2204 14
rect 2219 -4 2249 14
rect 2286 0 2305 14
rect 2320 0 2326 14
rect 2335 0 2348 14
rect 2363 -4 2393 14
rect 2436 0 2479 14
rect 2486 1 2494 14
rect 2527 1 2665 14
rect 2698 1 2706 14
rect 2449 -18 2479 0
rect 2542 -2 2650 1
rect 2542 -4 2572 -2
rect 2620 -4 2650 -2
rect 2713 -18 2743 14
rect 2771 0 2784 14
rect 2799 -4 2829 14
rect 2866 0 2885 14
rect 2900 0 2906 14
rect 2915 0 2928 14
rect 2943 -4 2973 14
rect 3016 0 3059 14
rect 3066 1 3074 14
rect 3107 1 3245 14
rect 3278 1 3286 14
rect 3029 -18 3059 0
rect 3122 -2 3230 1
rect 3122 -4 3152 -2
rect 3200 -4 3230 -2
rect 3293 -18 3323 14
rect 3351 0 3364 14
rect 3379 -4 3409 14
rect 3446 0 3465 14
rect 3480 0 3486 14
rect 3495 0 3508 14
rect 3523 -4 3553 14
rect 3596 0 3639 14
rect 3646 1 3654 14
rect 3687 1 3825 14
rect 3858 1 3866 14
rect 3609 -18 3639 0
rect 3702 -2 3810 1
rect 3702 -4 3732 -2
rect 3780 -4 3810 -2
rect 3873 -18 3903 14
rect 3931 0 3944 14
rect 3959 -4 3989 14
rect 4026 0 4045 14
rect 4060 0 4066 14
rect 4075 0 4088 14
rect 4103 -4 4133 14
rect 4176 0 4219 14
rect 4226 1 4234 14
rect 4267 1 4405 14
rect 4438 1 4446 14
rect 4189 -18 4219 0
rect 4282 -2 4390 1
rect 4282 -4 4312 -2
rect 4360 -4 4390 -2
rect 4453 -18 4483 14
rect 4511 0 4524 14
rect 4539 -4 4569 14
rect 4606 0 4625 14
rect 4640 1 4646 15
rect 4655 1 4668 15
rect 4683 -3 4713 15
rect 4756 1 4799 15
rect 4806 2 4814 15
rect 4847 2 4985 15
rect 5018 2 5026 15
rect 4769 -17 4799 1
rect 4862 -1 4970 2
rect 4862 -3 4892 -1
rect 4940 -3 4970 -1
rect 5033 -17 5063 15
rect 5091 1 5104 15
rect 5119 -3 5149 15
rect 5186 1 5205 15
rect 5220 1 5226 15
rect 5235 1 5248 15
rect 5263 -3 5293 15
rect 5336 1 5379 15
rect 5386 2 5394 15
rect 5427 2 5565 15
rect 5598 2 5606 15
rect 5349 -17 5379 1
rect 5442 -1 5550 2
rect 5442 -3 5472 -1
rect 5520 -3 5550 -1
rect 5613 -17 5643 15
rect 5671 1 5684 15
rect 5699 -3 5729 15
rect 5766 1 5785 15
rect 5800 1 5806 15
rect 5815 1 5828 15
rect 5843 -3 5873 15
rect 5916 1 5959 15
rect 5966 2 5974 15
rect 6007 2 6145 15
rect 6178 2 6186 15
rect 5929 -17 5959 1
rect 6022 -1 6130 2
rect 6022 -3 6052 -1
rect 6100 -3 6130 -1
rect 6193 -17 6223 15
rect 6251 1 6264 15
rect 6279 -3 6309 15
rect 6346 1 6365 15
rect 6380 1 6386 15
rect 6395 1 6408 15
rect 6423 -3 6453 15
rect 6496 1 6539 15
rect 6546 2 6554 15
rect 6587 2 6725 15
rect 6758 2 6766 15
rect 6509 -17 6539 1
rect 6602 -1 6710 2
rect 6602 -3 6632 -1
rect 6680 -3 6710 -1
rect 6773 -17 6803 15
rect 6831 1 6844 15
rect 6859 -3 6889 15
rect 6926 1 6945 15
rect 6960 1 6966 15
rect 6975 1 6988 15
rect 7003 -3 7033 15
rect 7076 1 7119 15
rect 7126 2 7134 15
rect 7167 2 7305 15
rect 7338 2 7346 15
rect 7089 -17 7119 1
rect 7182 -1 7290 2
rect 7182 -3 7212 -1
rect 7260 -3 7290 -1
rect 7353 -17 7383 15
rect 7411 1 7424 15
rect 7439 -3 7469 15
rect 7506 1 7525 15
rect 7540 1 7546 15
rect 7555 1 7568 15
rect 7583 -3 7613 15
rect 7656 1 7699 15
rect 7706 2 7714 15
rect 7747 2 7885 15
rect 7918 2 7926 15
rect 7669 -17 7699 1
rect 7762 -1 7870 2
rect 7762 -3 7792 -1
rect 7840 -3 7870 -1
rect 7933 -17 7963 15
rect 7991 1 8004 15
rect 8019 -3 8049 15
rect 8086 1 8105 15
rect 8120 1 8126 15
rect 8135 1 8148 15
rect 8163 -3 8193 15
rect 8236 1 8279 15
rect 8286 2 8294 15
rect 8327 2 8465 15
rect 8498 2 8506 15
rect 8249 -17 8279 1
rect 8342 -1 8450 2
rect 8342 -3 8372 -1
rect 8420 -3 8450 -1
rect 8513 -17 8543 15
rect 8571 1 8584 15
rect 8599 -3 8629 15
rect 8666 1 8685 15
rect 8700 1 8706 15
rect 8715 1 8728 15
rect 8743 -3 8773 15
rect 8816 1 8859 15
rect 8866 2 8874 15
rect 8907 2 9045 15
rect 9078 2 9086 15
rect 8829 -17 8859 1
rect 8922 -1 9030 2
rect 8922 -3 8952 -1
rect 9000 -3 9030 -1
rect 9093 -17 9123 15
rect 9151 1 9164 15
rect 9179 -3 9209 15
rect 9246 1 9265 15
rect 9280 1 9286 15
rect 9295 1 9308 15
rect 9323 -3 9353 15
rect 9396 1 9439 15
rect 9446 2 9454 15
rect 9487 2 9625 15
rect 9658 2 9666 15
rect 9409 -17 9439 1
rect 9502 -1 9610 2
rect 9502 -3 9532 -1
rect 9580 -3 9610 -1
rect 9673 -17 9703 15
rect 9731 1 9744 15
rect 9759 -3 9789 15
rect 9826 1 9845 15
rect 9860 1 9866 15
rect 9875 1 9888 15
rect 9903 -3 9933 15
rect 9976 1 10019 15
rect 10026 2 10034 15
rect 10067 2 10205 15
rect 10238 2 10246 15
rect 9989 -17 10019 1
rect 10082 -1 10190 2
rect 10082 -3 10112 -1
rect 10160 -3 10190 -1
rect 10253 -17 10283 15
rect 10311 1 10324 15
rect 10339 -3 10369 15
rect 10406 1 10425 15
rect 10440 1 10446 15
rect 10455 1 10468 15
rect 10483 -3 10513 15
rect 10556 1 10599 15
rect 10606 2 10614 15
rect 10647 2 10785 15
rect 10818 2 10826 15
rect 10569 -17 10599 1
rect 10662 -1 10770 2
rect 10662 -3 10692 -1
rect 10740 -3 10770 -1
rect 10833 -17 10863 15
rect 10891 1 10904 15
rect 10919 -3 10949 15
rect 10986 1 11005 15
rect 11020 1 11026 15
rect 11035 1 11048 15
rect 11063 -3 11093 15
rect 11136 1 11179 15
rect 11186 2 11194 15
rect 11227 2 11365 15
rect 11398 2 11406 15
rect 11149 -17 11179 1
rect 11242 -1 11350 2
rect 11242 -3 11272 -1
rect 11320 -3 11350 -1
rect 11413 -17 11443 15
rect 11471 1 11484 15
rect 11499 -3 11529 15
rect 11566 1 11585 15
rect 11600 1 11606 15
rect 11615 1 11628 15
rect 11643 -3 11673 15
rect 11716 1 11759 15
rect 11766 2 11774 15
rect 11807 2 11945 15
rect 11978 2 11986 15
rect 11729 -17 11759 1
rect 11822 -1 11930 2
rect 11822 -3 11852 -1
rect 11900 -3 11930 -1
rect 11993 -17 12023 15
rect 12051 1 12064 15
rect 12079 -3 12109 15
rect 12146 1 12165 15
rect 12180 1 12186 15
rect 12195 1 12208 15
rect 12223 -3 12253 15
rect 12296 1 12339 15
rect 12346 2 12354 15
rect 12387 2 12525 15
rect 12558 2 12566 15
rect 12309 -17 12339 1
rect 12402 -1 12510 2
rect 12402 -3 12432 -1
rect 12480 -3 12510 -1
rect 12573 -17 12603 15
rect 12631 1 12644 15
rect 12659 -3 12689 15
rect 12726 1 12745 15
rect 12760 1 12766 15
rect 12775 1 12788 15
rect 12803 -3 12833 15
rect 12876 1 12919 15
rect 12926 2 12934 15
rect 12967 2 13105 15
rect 13138 2 13146 15
rect 12889 -17 12919 1
rect 12982 -1 13090 2
rect 12982 -3 13012 -1
rect 13060 -3 13090 -1
rect 13153 -17 13183 15
rect 13211 1 13224 15
rect 13239 -3 13269 15
rect 13306 1 13325 15
rect 13340 1 13346 15
rect 13355 1 13368 15
rect 13383 -3 13413 15
rect 13456 1 13499 15
rect 13506 2 13514 15
rect 13547 2 13685 15
rect 13718 2 13726 15
rect 13469 -17 13499 1
rect 13562 -1 13670 2
rect 13562 -3 13592 -1
rect 13640 -3 13670 -1
rect 13733 -17 13763 15
rect 13791 1 13804 15
rect 13819 -3 13849 15
rect 13886 1 13905 15
rect 13920 1 13926 15
rect 13935 1 13948 15
rect 13963 -3 13993 15
rect 14036 1 14079 15
rect 14086 2 14094 15
rect 14127 2 14265 15
rect 14298 2 14306 15
rect 14049 -17 14079 1
rect 14142 -1 14250 2
rect 14142 -3 14172 -1
rect 14220 -3 14250 -1
rect 14313 -17 14343 15
rect 14371 1 14384 15
rect 14399 -3 14429 15
rect 14466 1 14485 15
rect 14500 1 14506 15
rect 14515 1 14528 15
rect 14543 -3 14573 15
rect 14616 1 14659 15
rect 14666 2 14674 15
rect 14707 2 14845 15
rect 14878 2 14886 15
rect 14629 -17 14659 1
rect 14722 -1 14830 2
rect 14722 -3 14752 -1
rect 14800 -3 14830 -1
rect 14893 -17 14923 15
rect 14951 1 14964 15
rect 14979 -3 15009 15
rect 15046 1 15065 15
rect 15080 1 15086 15
rect 15095 1 15108 15
rect 15123 -3 15153 15
rect 15196 1 15239 15
rect 15246 2 15254 15
rect 15287 2 15425 15
rect 15458 2 15466 15
rect 15209 -17 15239 1
rect 15302 -1 15410 2
rect 15302 -3 15332 -1
rect 15380 -3 15410 -1
rect 15473 -17 15503 15
rect 15531 1 15544 15
rect 15559 -3 15589 15
rect 15626 1 15645 15
rect 15660 1 15666 15
rect 15675 1 15688 15
rect 15703 -3 15733 15
rect 15776 1 15819 15
rect 15826 2 15834 15
rect 15867 2 16005 15
rect 16038 2 16046 15
rect 15789 -17 15819 1
rect 15882 -1 15990 2
rect 15882 -3 15912 -1
rect 15960 -3 15990 -1
rect 16053 -17 16083 15
rect 16111 1 16124 15
rect 16139 -3 16169 15
rect 16206 1 16225 15
rect 16240 1 16246 15
rect 16255 1 16268 15
rect 16283 -3 16313 15
rect 16356 1 16399 15
rect 16406 2 16414 15
rect 16447 2 16585 15
rect 16618 2 16626 15
rect 16369 -17 16399 1
rect 16462 -1 16570 2
rect 16462 -3 16492 -1
rect 16540 -3 16570 -1
rect 16633 -17 16663 15
rect 16691 1 16704 15
rect 16719 -3 16749 15
rect 16786 1 16805 15
rect 16820 1 16826 15
rect 16835 1 16848 15
rect 16863 -3 16893 15
rect 16936 1 16979 15
rect 16986 2 16994 15
rect 17027 2 17165 15
rect 17198 2 17206 15
rect 16949 -17 16979 1
rect 17042 -1 17150 2
rect 17042 -3 17072 -1
rect 17120 -3 17150 -1
rect 17213 -17 17243 15
rect 17271 1 17284 15
rect 17299 -3 17329 15
rect 17366 1 17385 15
rect 17400 1 17406 15
rect 17415 1 17428 15
rect 17443 -3 17473 15
rect 17516 1 17559 15
rect 17566 2 17574 15
rect 17607 2 17745 15
rect 17778 2 17786 15
rect 17529 -17 17559 1
rect 17622 -1 17730 2
rect 17622 -3 17652 -1
rect 17700 -3 17730 -1
rect 17793 -17 17823 15
rect 17851 1 17864 15
rect 17879 -3 17909 15
rect 17946 1 17965 15
rect 17980 1 17986 15
rect 17995 1 18008 15
rect 18023 -3 18053 15
rect 18096 1 18139 15
rect 18146 2 18154 15
rect 18187 2 18325 15
rect 18358 2 18366 15
rect 18109 -17 18139 1
rect 18202 -1 18310 2
rect 18202 -3 18232 -1
rect 18280 -3 18310 -1
rect 18373 -17 18403 15
rect 18431 1 18444 15
rect 18459 -3 18489 15
rect 18532 1 18545 15
<< pwell >>
rect 4612 7560 4640 7574
rect 4612 7516 4640 7530
rect 4612 7290 4640 7304
rect 4612 7246 4640 7260
rect 4612 7020 4640 7034
rect 4612 6976 4640 6990
rect 4612 6750 4640 6764
rect 4612 6706 4640 6720
rect 4612 6480 4640 6494
rect 4612 6436 4640 6450
rect 4612 6210 4640 6224
rect 4612 6166 4640 6180
rect 4612 5940 4640 5954
rect 4612 5896 4640 5910
rect 4612 5670 4640 5684
rect 4612 5626 4640 5640
rect 4612 5400 4640 5414
rect 4612 5356 4640 5370
rect 4612 5130 4640 5144
rect 4612 5086 4640 5100
rect 4612 4860 4640 4874
rect 4612 4816 4640 4830
rect 4612 4590 4640 4604
rect 4612 4546 4640 4560
rect 4612 4320 4640 4334
rect 4612 4276 4640 4290
rect 4612 4050 4640 4064
rect 4612 4006 4640 4020
rect 4612 3780 4640 3794
rect 4612 3736 4640 3750
rect 4612 3510 4640 3524
rect 4612 3466 4640 3480
rect 4612 3240 4640 3254
rect 4612 3196 4640 3210
rect 4612 2970 4640 2984
rect 4612 2926 4640 2940
rect 4612 2700 4640 2714
rect 4612 2656 4640 2670
rect 4612 2430 4640 2444
rect 4612 2386 4640 2400
rect 4612 2160 4640 2174
rect 4612 2116 4640 2130
rect 4612 1890 4640 1904
rect 4612 1846 4640 1860
rect 4612 1620 4640 1634
rect 4612 1576 4640 1590
rect 4612 1350 4640 1364
rect 4612 1306 4640 1320
rect 4612 1080 4640 1094
rect 4612 1036 4640 1050
rect 4612 810 4640 824
rect 4612 766 4640 780
rect 4612 540 4640 554
rect 4612 496 4640 510
rect 4612 270 4640 284
rect 4612 226 4640 240
rect 74 184 89 212
rect 464 184 479 213
rect 4714 184 4729 212
rect 5104 184 5119 213
rect 0 38 15 80
rect 537 38 552 80
rect 580 38 595 80
rect 4640 38 4655 80
rect 5177 38 5192 80
rect 5220 38 5235 80
rect 4612 0 4640 14
<< ndiffc >>
rect 74 184 89 212
rect 464 184 479 213
rect 654 184 669 212
rect 1044 184 1059 213
rect 1234 184 1249 212
rect 1624 184 1639 213
rect 1814 184 1829 212
rect 2204 184 2219 213
rect 2394 184 2409 212
rect 2784 184 2799 213
rect 2974 184 2989 212
rect 3364 184 3379 213
rect 3554 184 3569 212
rect 3944 184 3959 213
rect 4134 184 4149 212
rect 4524 184 4539 213
rect 4714 185 4729 213
rect 5104 184 5119 213
rect 5294 184 5309 212
rect 5684 184 5699 213
rect 5874 184 5889 212
rect 6264 184 6279 213
rect 6454 184 6469 212
rect 6844 184 6859 213
rect 7034 184 7049 212
rect 7424 184 7439 213
rect 7614 184 7629 212
rect 8004 184 8019 213
rect 8194 184 8209 212
rect 8584 184 8599 213
rect 8774 184 8789 212
rect 9164 184 9179 213
rect 9354 185 9369 213
rect 9744 185 9759 214
rect 9934 185 9949 213
rect 10324 185 10339 214
rect 10514 185 10529 213
rect 10904 185 10919 214
rect 11094 185 11109 213
rect 11484 185 11499 214
rect 11674 185 11689 213
rect 12064 185 12079 214
rect 12254 185 12269 213
rect 12644 185 12659 214
rect 12834 185 12849 213
rect 13224 185 13239 214
rect 13414 185 13429 213
rect 13804 185 13819 214
rect 13994 185 14009 213
rect 14384 185 14399 214
rect 14574 185 14589 213
rect 14964 185 14979 214
rect 15154 185 15169 213
rect 15544 185 15559 214
rect 15734 185 15749 213
rect 16124 185 16139 214
rect 16314 185 16329 213
rect 16704 185 16719 214
rect 16894 185 16909 213
rect 17284 185 17299 214
rect 17474 185 17489 213
rect 17864 185 17879 214
rect 18054 185 18069 213
rect 18444 185 18459 214
rect 0 38 15 80
rect 537 38 552 80
rect 580 38 595 80
rect 1117 38 1132 80
rect 1160 38 1175 80
rect 1697 38 1712 80
rect 1740 38 1755 80
rect 2277 38 2292 80
rect 2320 38 2335 80
rect 2857 38 2872 80
rect 2900 38 2915 80
rect 3437 38 3452 80
rect 3480 38 3495 80
rect 4017 38 4032 80
rect 4060 38 4075 80
rect 4597 38 4612 80
rect 4640 39 4655 81
rect 5177 38 5192 80
rect 5220 38 5235 80
rect 5757 38 5772 80
rect 5800 38 5815 80
rect 6337 38 6352 80
rect 6380 38 6395 80
rect 6917 38 6932 80
rect 6960 38 6975 80
rect 7497 38 7512 80
rect 7540 38 7555 80
rect 8077 38 8092 80
rect 8120 38 8135 80
rect 8657 38 8672 80
rect 8700 38 8715 80
rect 9237 38 9252 80
rect 9280 39 9295 81
rect 9817 39 9832 81
rect 9860 39 9875 81
rect 10397 39 10412 81
rect 10440 39 10455 81
rect 10977 39 10992 81
rect 11020 39 11035 81
rect 11557 39 11572 81
rect 11600 39 11615 81
rect 12137 39 12152 81
rect 12180 39 12195 81
rect 12717 39 12732 81
rect 12760 39 12775 81
rect 13297 39 13312 81
rect 13340 39 13355 81
rect 13877 39 13892 81
rect 13920 39 13935 81
rect 14457 38 14472 80
rect 14500 38 14515 80
rect 15037 38 15052 80
rect 15080 38 15095 80
rect 15617 38 15632 80
rect 15660 38 15675 80
rect 16197 38 16212 80
rect 16240 38 16255 80
rect 16777 38 16792 80
rect 16820 38 16835 80
rect 17357 38 17372 80
rect 17400 38 17415 80
rect 17937 38 17952 80
rect 17980 38 17995 80
rect 18517 38 18532 80
<< poly >>
rect 0 8610 30 8640
rect 4561 8610 4708 8640
rect 9222 8610 9315 8640
rect 13841 8610 13988 8640
rect 0 8340 30 8370
rect 4567 8340 4701 8370
rect 9222 8340 9310 8370
rect 13847 8340 13981 8370
rect 0 8070 30 8100
rect 4571 8070 4694 8100
rect 9198 8070 9318 8100
rect 13851 8070 13974 8100
rect 0 7800 30 7830
rect 4574 7800 4724 7830
rect 9215 7800 9310 7830
rect 13854 7800 14004 7830
rect 0 7530 30 7560
rect 4558 7530 4711 7560
rect 9209 7530 9318 7560
rect 13838 7530 13991 7560
rect 0 7260 30 7290
rect 4556 7260 4739 7290
rect 9212 7260 9318 7290
rect 13836 7260 14019 7290
rect 0 6990 30 7020
rect 4554 6990 4707 7020
rect 9222 6990 9332 7020
rect 13834 6990 13987 7020
rect 0 6720 30 6750
rect 4563 6720 4759 6750
rect 9212 6720 9318 6750
rect 13843 6720 14039 6750
rect 0 6450 30 6480
rect 4572 6450 4700 6480
rect 9212 6450 9312 6480
rect 13852 6450 13980 6480
rect 0 6180 30 6210
rect 4575 6180 4747 6210
rect 9212 6180 9349 6210
rect 13855 6180 14027 6210
rect 0 5910 30 5940
rect 4563 5910 4729 5940
rect 9215 5910 9344 5940
rect 13843 5910 14009 5940
rect 0 5640 30 5670
rect 4560 5640 4732 5670
rect 9212 5640 9329 5670
rect 13840 5640 14012 5670
rect 0 5370 30 5400
rect 4563 5370 4700 5400
rect 9212 5370 9323 5400
rect 13843 5370 13980 5400
rect 0 5100 30 5130
rect 4572 5100 4706 5130
rect 9209 5100 9310 5130
rect 13852 5100 13986 5130
rect 0 4830 30 4860
rect 4544 4830 4694 4860
rect 9212 4830 9335 4860
rect 13824 4830 13974 4860
rect 0 4560 30 4590
rect 4561 4560 4714 4590
rect 9221 4560 9335 4590
rect 13841 4560 13994 4590
rect 0 4290 30 4320
rect 4568 4290 4703 4320
rect 9209 4290 9318 4320
rect 13848 4290 13983 4320
rect 0 4020 30 4050
rect 4566 4020 4736 4050
rect 9215 4020 9318 4050
rect 13846 4020 14016 4050
rect 0 3750 30 3780
rect 4563 3750 4719 3780
rect 9203 3750 9323 3780
rect 13843 3750 13999 3780
rect 0 3480 30 3510
rect 4561 3480 4713 3510
rect 9212 3480 9310 3510
rect 13841 3480 13993 3510
rect 0 3210 30 3240
rect 4563 3210 4714 3240
rect 9212 3210 9315 3240
rect 13843 3210 13994 3240
rect 0 2940 30 2970
rect 4565 2940 4704 2970
rect 9206 2940 9318 2970
rect 13845 2940 13984 2970
rect 0 2670 30 2700
rect 4553 2670 4697 2700
rect 9209 2670 9312 2700
rect 13833 2670 13977 2700
rect 0 2400 30 2430
rect 4553 2400 4701 2430
rect 9212 2400 9315 2430
rect 13833 2400 13981 2430
rect 0 2130 30 2160
rect 4562 2130 4697 2160
rect 9209 2130 9310 2160
rect 13842 2130 13977 2160
rect 0 1860 30 1890
rect 4564 1860 4695 1890
rect 9212 1860 9315 1890
rect 13844 1860 13975 1890
rect 0 1590 30 1620
rect 4566 1590 4721 1620
rect 9209 1590 9318 1620
rect 13846 1590 14001 1620
rect 0 1320 30 1350
rect 4569 1320 4706 1350
rect 9201 1320 9324 1350
rect 13849 1320 13986 1350
rect 0 1050 30 1080
rect 4549 1050 4695 1080
rect 9211 1050 9313 1080
rect 13829 1050 13975 1080
rect 0 780 30 810
rect 4564 780 4713 810
rect 9207 780 9326 810
rect 13844 780 13993 810
rect 0 509 30 539
rect 4577 510 4701 540
rect 9203 511 9328 541
rect 13857 510 13981 540
rect 4631 270 4698 271
rect 0 240 30 270
rect 4570 241 4698 270
rect 9209 241 9337 271
rect 13850 241 13978 271
rect 4570 240 4631 241
<< metal1 >>
rect 0 8596 15 8610
rect 4576 8596 4671 8610
rect 9217 8596 9321 8610
rect 13856 8596 13951 8610
rect 0 8472 15 8506
rect 4505 8472 4691 8506
rect 9137 8472 9314 8506
rect 13785 8472 13971 8506
rect 0 8370 15 8384
rect 4573 8370 4670 8384
rect 9238 8370 9295 8384
rect 13853 8370 13950 8384
rect 0 8326 15 8340
rect 4578 8326 4678 8340
rect 9232 8326 9304 8340
rect 13858 8326 13958 8340
rect 0 8202 15 8236
rect 4502 8202 4701 8236
rect 9145 8202 9308 8236
rect 13782 8202 13981 8236
rect 0 8100 15 8114
rect 4578 8100 4688 8114
rect 9232 8100 9298 8114
rect 13858 8100 13968 8114
rect 0 8056 15 8070
rect 4581 8056 4663 8070
rect 9235 8056 9336 8070
rect 13861 8056 13943 8070
rect 0 7932 15 7966
rect 4505 7932 4727 7966
rect 9143 7932 9305 7966
rect 13785 7932 14007 7966
rect 0 7830 15 7844
rect 4582 7830 4666 7844
rect 9237 7830 9301 7844
rect 13862 7830 13946 7844
rect 0 7786 15 7800
rect 4575 7786 4685 7800
rect 9229 7786 9315 7800
rect 13855 7786 13965 7800
rect 0 7662 15 7696
rect 4640 7662 4655 7696
rect 9143 7662 9308 7696
rect 13920 7662 13935 7696
rect 0 7560 15 7574
rect 4612 7560 4655 7574
rect 9229 7560 9298 7574
rect 13892 7560 13935 7574
rect 0 7516 15 7530
rect 4612 7516 4655 7530
rect 9223 7516 9324 7530
rect 13892 7516 13935 7530
rect 0 7392 15 7426
rect 4504 7392 4727 7426
rect 9143 7392 9314 7426
rect 13784 7392 14007 7426
rect 0 7290 15 7304
rect 4612 7290 4655 7304
rect 9223 7290 9307 7304
rect 13892 7290 13935 7304
rect 0 7246 15 7260
rect 4612 7246 4655 7260
rect 9235 7246 9324 7260
rect 13892 7246 13935 7260
rect 0 7122 15 7156
rect 4496 7122 4683 7156
rect 9140 7122 9314 7156
rect 13776 7122 13963 7156
rect 0 7020 15 7034
rect 4612 7020 4655 7034
rect 9232 7020 9301 7034
rect 13892 7020 13935 7034
rect 0 6976 15 6990
rect 4612 6976 4655 6990
rect 9232 6976 9321 6990
rect 13892 6976 13935 6990
rect 0 6852 15 6886
rect 4505 6852 4734 6886
rect 9132 6852 9308 6886
rect 13785 6852 14014 6886
rect 0 6750 15 6764
rect 4612 6750 4655 6764
rect 9229 6750 9295 6764
rect 13892 6750 13935 6764
rect 0 6706 15 6720
rect 4612 6706 4655 6720
rect 9229 6706 9315 6720
rect 13892 6706 13935 6720
rect 0 6582 15 6616
rect 4502 6582 4705 6616
rect 9126 6582 9305 6616
rect 13782 6582 13985 6616
rect 0 6480 15 6494
rect 4612 6480 4655 6494
rect 9217 6480 9295 6494
rect 13892 6480 13935 6494
rect 0 6436 15 6450
rect 4612 6436 4655 6450
rect 9232 6436 9298 6450
rect 13892 6436 13935 6450
rect 0 6312 15 6346
rect 4505 6312 4722 6346
rect 9145 6312 9325 6346
rect 13785 6312 14002 6346
rect 0 6210 15 6224
rect 4612 6210 4655 6224
rect 9220 6210 9315 6224
rect 13892 6210 13935 6224
rect 0 6166 15 6180
rect 4612 6166 4655 6180
rect 9235 6166 9315 6180
rect 13892 6166 13935 6180
rect 0 6042 15 6076
rect 4499 6042 4731 6076
rect 9143 6042 9305 6076
rect 13779 6042 14011 6076
rect 0 5940 15 5954
rect 4612 5940 4655 5954
rect 9217 5940 9312 5954
rect 13892 5940 13935 5954
rect 0 5896 15 5910
rect 4612 5896 4655 5910
rect 9229 5896 9312 5910
rect 13892 5896 13935 5910
rect 0 5772 15 5806
rect 4505 5772 4740 5806
rect 9140 5772 9295 5806
rect 13785 5772 14020 5806
rect 0 5670 15 5684
rect 4612 5670 4655 5684
rect 9223 5670 9307 5684
rect 13892 5670 13935 5684
rect 0 5626 15 5640
rect 4612 5626 4655 5640
rect 9232 5626 9324 5640
rect 13892 5626 13935 5640
rect 0 5502 15 5536
rect 4505 5502 4728 5536
rect 9137 5502 9317 5536
rect 13785 5502 14008 5536
rect 0 5400 15 5414
rect 4612 5400 4655 5414
rect 9220 5400 9301 5414
rect 13892 5400 13935 5414
rect 0 5356 15 5370
rect 4612 5356 4655 5370
rect 9232 5356 9336 5370
rect 13892 5356 13935 5370
rect 0 5232 15 5266
rect 4496 5232 4728 5266
rect 9123 5232 9311 5266
rect 13776 5232 14008 5266
rect 0 5130 15 5144
rect 4612 5130 4655 5144
rect 9232 5130 9298 5144
rect 13892 5130 13935 5144
rect 0 5086 15 5100
rect 4612 5086 4655 5100
rect 9237 5086 9295 5100
rect 13892 5086 13935 5100
rect 0 4962 15 4996
rect 4502 4962 4746 4996
rect 9140 4962 9308 4996
rect 13782 4962 14026 4996
rect 0 4860 15 4874
rect 4612 4860 4655 4874
rect 9237 4860 9298 4874
rect 13892 4860 13935 4874
rect 0 4816 15 4830
rect 4612 4816 4655 4830
rect 9223 4816 9312 4830
rect 13892 4816 13935 4830
rect 0 4692 15 4726
rect 4505 4692 4716 4726
rect 9132 4692 9299 4726
rect 13785 4692 13996 4726
rect 0 4590 15 4604
rect 4612 4590 4655 4604
rect 9229 4590 9310 4604
rect 13892 4590 13935 4604
rect 0 4546 15 4560
rect 4612 4546 4655 4560
rect 9220 4546 9324 4560
rect 13892 4546 13935 4560
rect 0 4422 15 4456
rect 4503 4422 4753 4456
rect 9132 4422 9302 4456
rect 13783 4422 14033 4456
rect 0 4320 15 4334
rect 4612 4320 4655 4334
rect 9229 4320 9307 4334
rect 13892 4320 13935 4334
rect 0 4276 15 4290
rect 4612 4276 4655 4290
rect 9232 4276 9315 4290
rect 13892 4276 13935 4290
rect 0 4152 15 4186
rect 4505 4152 4724 4186
rect 9143 4152 9302 4186
rect 13785 4152 14004 4186
rect 0 4050 15 4064
rect 4612 4050 4655 4064
rect 9232 4050 9307 4064
rect 13892 4050 13935 4064
rect 0 4006 15 4020
rect 4612 4006 4655 4020
rect 9229 4006 9312 4020
rect 13892 4006 13935 4020
rect 0 3882 15 3916
rect 4503 3882 4731 3916
rect 9137 3882 9302 3916
rect 13783 3882 14011 3916
rect 0 3780 15 3794
rect 4612 3780 4655 3794
rect 9220 3780 9298 3794
rect 13892 3780 13935 3794
rect 0 3736 15 3750
rect 4612 3736 4655 3750
rect 9232 3736 9310 3750
rect 13892 3736 13935 3750
rect 0 3612 15 3646
rect 4505 3612 4736 3646
rect 9137 3612 9305 3646
rect 13785 3612 14016 3646
rect 0 3510 15 3524
rect 4612 3510 4655 3524
rect 9220 3510 9295 3524
rect 13892 3510 13935 3524
rect 0 3466 15 3480
rect 4612 3466 4655 3480
rect 9235 3466 9321 3480
rect 13892 3466 13935 3480
rect 0 3342 15 3376
rect 4496 3342 4727 3376
rect 9137 3342 9302 3376
rect 13776 3342 14007 3376
rect 0 3240 15 3254
rect 4612 3240 4655 3254
rect 9232 3240 9321 3254
rect 13892 3240 13935 3254
rect 0 3196 15 3210
rect 4612 3196 4655 3210
rect 9232 3196 9330 3210
rect 13892 3196 13935 3210
rect 0 3072 15 3106
rect 4502 3072 4741 3106
rect 9143 3072 9322 3106
rect 13782 3072 14021 3106
rect 0 2970 15 2984
rect 4612 2970 4655 2984
rect 9223 2970 9298 2984
rect 13892 2970 13935 2984
rect 0 2926 15 2940
rect 4612 2926 4655 2940
rect 9223 2926 9315 2940
rect 13892 2926 13935 2940
rect 0 2802 15 2836
rect 4502 2802 4734 2836
rect 9140 2802 9308 2836
rect 13782 2802 14014 2836
rect 0 2700 15 2714
rect 4612 2700 4655 2714
rect 9223 2700 9301 2714
rect 13892 2700 13935 2714
rect 0 2656 15 2670
rect 4612 2656 4655 2670
rect 9232 2656 9321 2670
rect 13892 2656 13935 2670
rect 0 2532 15 2566
rect 4505 2532 4736 2566
rect 9140 2532 9305 2566
rect 13785 2532 14016 2566
rect 0 2430 15 2444
rect 4612 2430 4655 2444
rect 9220 2430 9295 2444
rect 13892 2430 13935 2444
rect 0 2386 15 2400
rect 4612 2386 4655 2400
rect 9232 2386 9310 2400
rect 13892 2386 13935 2400
rect 0 2262 15 2296
rect 4497 2262 4740 2296
rect 9140 2262 9314 2296
rect 13777 2262 14020 2296
rect 0 2160 15 2174
rect 4612 2160 4655 2174
rect 9235 2160 9310 2174
rect 13892 2160 13935 2174
rect 0 2116 15 2130
rect 4612 2116 4655 2130
rect 9229 2116 9295 2130
rect 13892 2116 13935 2130
rect 0 1992 15 2026
rect 4505 1992 4710 2026
rect 9143 1992 9317 2026
rect 13785 1992 13990 2026
rect 0 1890 15 1904
rect 4612 1890 4655 1904
rect 9223 1890 9321 1904
rect 13892 1890 13935 1904
rect 0 1846 15 1860
rect 4612 1846 4655 1860
rect 9217 1846 9321 1860
rect 13892 1846 13935 1860
rect 0 1722 15 1756
rect 4505 1722 4688 1756
rect 9126 1722 9311 1756
rect 13785 1722 13968 1756
rect 0 1620 15 1634
rect 4612 1620 4655 1634
rect 9223 1620 9295 1634
rect 13892 1620 13935 1634
rect 0 1576 15 1590
rect 4612 1576 4655 1590
rect 9223 1576 9307 1590
rect 13892 1576 13935 1590
rect 0 1452 15 1486
rect 4501 1452 4708 1486
rect 9141 1452 9319 1486
rect 13781 1452 13988 1486
rect 0 1350 15 1364
rect 4612 1350 4655 1364
rect 9227 1350 9309 1364
rect 13892 1350 13935 1364
rect 0 1306 15 1320
rect 4612 1306 4655 1320
rect 9227 1306 9306 1320
rect 13892 1306 13935 1320
rect 0 1182 15 1216
rect 4505 1182 4701 1216
rect 9135 1182 9317 1216
rect 13785 1182 13981 1216
rect 0 1080 15 1094
rect 4612 1080 4655 1094
rect 9226 1080 9307 1094
rect 13892 1080 13935 1094
rect 0 1036 15 1050
rect 4612 1036 4655 1050
rect 9212 1036 9304 1050
rect 13892 1036 13935 1050
rect 0 912 15 946
rect 4505 912 4725 946
rect 9138 912 9320 946
rect 13785 912 14005 946
rect 0 810 15 824
rect 4612 810 4655 824
rect 9214 810 9327 824
rect 13892 810 13935 824
rect 0 766 15 780
rect 4612 766 4655 780
rect 9211 766 9311 780
rect 13892 766 13935 780
rect 0 642 15 676
rect 4505 642 4741 676
rect 9145 642 9372 676
rect 13785 642 14021 676
rect 0 540 15 554
rect 4612 540 4655 554
rect 9211 541 9330 555
rect 13892 540 13935 554
rect 0 495 15 509
rect 4612 496 4655 510
rect 9234 497 9303 511
rect 13892 496 13935 510
rect 0 371 15 405
rect 4505 372 4683 406
rect 9145 373 9330 407
rect 13785 372 13963 406
rect 4631 284 4640 285
rect 0 270 15 283
rect 4612 271 4655 284
rect 9233 271 9295 285
rect 13892 271 13935 284
rect 4612 270 4631 271
rect 4631 240 4655 241
rect 0 226 15 240
rect 4612 227 4655 240
rect 9237 227 9297 241
rect 13892 227 13935 241
rect 4612 226 4631 227
rect 4631 136 4705 137
rect 0 102 15 136
rect 4505 103 4705 136
rect 9140 103 9313 137
rect 13785 103 13985 137
rect 4505 102 4631 103
rect 4631 14 4655 15
rect 0 0 15 14
rect 4612 1 4655 14
rect 9238 1 9307 15
rect 13892 1 13935 15
rect 4612 0 4631 1
use 10T_1x8_magic  10T_1x8_magic_0
timestamp 1658881652
transform 1 0 0 0 1 7830
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_1
timestamp 1658881652
transform 1 0 0 0 1 7560
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_2
timestamp 1658881652
transform 1 0 0 0 1 8370
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_3
timestamp 1658881652
transform 1 0 0 0 1 8100
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_4
timestamp 1658881652
transform 1 0 0 0 1 6480
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_5
timestamp 1658881652
transform 1 0 0 0 1 6750
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_6
timestamp 1658881652
transform 1 0 0 0 1 7290
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_7
timestamp 1658881652
transform 1 0 0 0 1 7020
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_8
timestamp 1658881652
transform 1 0 0 0 1 4590
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_9
timestamp 1658881652
transform 1 0 0 0 1 4320
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_10
timestamp 1658881652
transform 1 0 0 0 1 4860
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_11
timestamp 1658881652
transform 1 0 0 0 1 5130
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_12
timestamp 1658881652
transform 1 0 0 0 1 5400
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_13
timestamp 1658881652
transform 1 0 0 0 1 5670
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_14
timestamp 1658881652
transform 1 0 0 0 1 6210
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_15
timestamp 1658881652
transform 1 0 0 0 1 5940
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_16
timestamp 1658881652
transform 1 0 0 0 1 0
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_17
timestamp 1658881652
transform 1 0 0 0 1 540
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_18
timestamp 1658881652
transform 1 0 0 0 1 270
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_19
timestamp 1658881652
transform 1 0 0 0 1 1080
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_20
timestamp 1658881652
transform 1 0 0 0 1 810
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_21
timestamp 1658881652
transform 1 0 0 0 1 1620
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_22
timestamp 1658881652
transform 1 0 0 0 1 1350
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_23
timestamp 1658881652
transform 1 0 0 0 1 2160
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_24
timestamp 1658881652
transform 1 0 0 0 1 1890
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_25
timestamp 1658881652
transform 1 0 0 0 1 2700
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_26
timestamp 1658881652
transform 1 0 0 0 1 2430
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_27
timestamp 1658881652
transform 1 0 0 0 1 3240
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_28
timestamp 1658881652
transform 1 0 0 0 1 2970
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_29
timestamp 1658881652
transform 1 0 0 0 1 3780
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_30
timestamp 1658881652
transform 1 0 0 0 1 3510
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_31
timestamp 1658881652
transform 1 0 0 0 1 4050
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_32
timestamp 1658881652
transform 1 0 4640 0 1 271
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_33
timestamp 1658881652
transform 1 0 4640 0 1 1
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_34
timestamp 1658881652
transform 1 0 4640 0 1 810
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_35
timestamp 1658881652
transform 1 0 4640 0 1 540
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_36
timestamp 1658881652
transform 1 0 4640 0 1 1350
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_37
timestamp 1658881652
transform 1 0 4640 0 1 1080
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_38
timestamp 1658881652
transform 1 0 4640 0 1 1890
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_39
timestamp 1658881652
transform 1 0 4640 0 1 2160
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_40
timestamp 1658881652
transform 1 0 4640 0 1 1620
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_41
timestamp 1658881652
transform 1 0 4640 0 1 2430
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_42
timestamp 1658881652
transform 1 0 4640 0 1 2700
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_43
timestamp 1658881652
transform 1 0 4640 0 1 2970
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_44
timestamp 1658881652
transform 1 0 4640 0 1 3240
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_45
timestamp 1658881652
transform 1 0 4640 0 1 3780
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_46
timestamp 1658881652
transform 1 0 4640 0 1 3510
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_47
timestamp 1658881652
transform 1 0 4640 0 1 4050
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_48
timestamp 1658881652
transform 1 0 4640 0 1 4320
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_49
timestamp 1658881652
transform 1 0 4640 0 1 4590
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_50
timestamp 1658881652
transform 1 0 4640 0 1 4860
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_51
timestamp 1658881652
transform 1 0 4640 0 1 5130
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_52
timestamp 1658881652
transform 1 0 4640 0 1 5400
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_53
timestamp 1658881652
transform 1 0 4640 0 1 5670
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_54
timestamp 1658881652
transform 1 0 4640 0 1 5940
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_55
timestamp 1658881652
transform 1 0 4640 0 1 6210
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_56
timestamp 1658881652
transform 1 0 4640 0 1 6480
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_57
timestamp 1658881652
transform 1 0 4640 0 1 6750
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_58
timestamp 1658881652
transform 1 0 4640 0 1 7020
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_59
timestamp 1658881652
transform 1 0 4640 0 1 7290
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_60
timestamp 1658881652
transform 1 0 4640 0 1 7560
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_61
timestamp 1658881652
transform 1 0 4640 0 1 7830
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_62
timestamp 1658881652
transform 1 0 4640 0 1 8100
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_63
timestamp 1658881652
transform 1 0 4640 0 1 8370
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_64
timestamp 1658881652
transform 1 0 9280 0 1 1
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_65
timestamp 1658881652
transform 1 0 9280 0 1 271
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_66
timestamp 1658881652
transform 1 0 13920 0 1 271
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_67
timestamp 1658881652
transform 1 0 13920 0 1 1
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_68
timestamp 1658881652
transform 1 0 9280 0 1 540
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_69
timestamp 1658881652
transform 1 0 13920 0 1 540
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_70
timestamp 1658881652
transform 1 0 9280 0 1 810
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_71
timestamp 1658881652
transform 1 0 13920 0 1 810
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_72
timestamp 1658881652
transform 1 0 9280 0 1 1080
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_73
timestamp 1658881652
transform 1 0 13920 0 1 1080
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_74
timestamp 1658881652
transform 1 0 9280 0 1 1350
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_75
timestamp 1658881652
transform 1 0 13920 0 1 1350
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_76
timestamp 1658881652
transform 1 0 9280 0 1 1620
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_77
timestamp 1658881652
transform 1 0 9280 0 1 1890
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_78
timestamp 1658881652
transform 1 0 13920 0 1 1890
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_79
timestamp 1658881652
transform 1 0 13920 0 1 1620
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_80
timestamp 1658881652
transform 1 0 9280 0 1 2160
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_81
timestamp 1658881652
transform 1 0 13920 0 1 2160
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_82
timestamp 1658881652
transform 1 0 9280 0 1 2430
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_83
timestamp 1658881652
transform 1 0 13920 0 1 2430
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_84
timestamp 1658881652
transform 1 0 9280 0 1 2700
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_85
timestamp 1658881652
transform 1 0 13920 0 1 2700
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_86
timestamp 1658881652
transform 1 0 9280 0 1 2970
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_87
timestamp 1658881652
transform 1 0 13920 0 1 2970
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_88
timestamp 1658881652
transform 1 0 9280 0 1 3240
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_89
timestamp 1658881652
transform 1 0 13920 0 1 3240
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_90
timestamp 1658881652
transform 1 0 9280 0 1 3780
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_91
timestamp 1658881652
transform 1 0 9280 0 1 3510
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_92
timestamp 1658881652
transform 1 0 13920 0 1 3780
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_93
timestamp 1658881652
transform 1 0 13920 0 1 3510
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_94
timestamp 1658881652
transform 1 0 9280 0 1 4050
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_95
timestamp 1658881652
transform 1 0 13920 0 1 4050
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_96
timestamp 1658881652
transform 1 0 9280 0 1 4320
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_97
timestamp 1658881652
transform 1 0 13920 0 1 4320
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_98
timestamp 1658881652
transform 1 0 9280 0 1 4590
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_99
timestamp 1658881652
transform 1 0 13920 0 1 4590
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_100
timestamp 1658881652
transform 1 0 9280 0 1 4860
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_101
timestamp 1658881652
transform 1 0 13920 0 1 4860
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_102
timestamp 1658881652
transform 1 0 9280 0 1 5130
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_103
timestamp 1658881652
transform 1 0 13920 0 1 5130
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_104
timestamp 1658881652
transform 1 0 9280 0 1 5400
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_105
timestamp 1658881652
transform 1 0 9280 0 1 5670
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_106
timestamp 1658881652
transform 1 0 13920 0 1 5400
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_107
timestamp 1658881652
transform 1 0 13920 0 1 5670
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_108
timestamp 1658881652
transform 1 0 9280 0 1 5940
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_109
timestamp 1658881652
transform 1 0 13920 0 1 5940
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_110
timestamp 1658881652
transform 1 0 9280 0 1 6210
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_111
timestamp 1658881652
transform 1 0 13920 0 1 6210
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_112
timestamp 1658881652
transform 1 0 9280 0 1 6480
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_113
timestamp 1658881652
transform 1 0 13920 0 1 6480
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_114
timestamp 1658881652
transform 1 0 9280 0 1 6750
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_115
timestamp 1658881652
transform 1 0 13920 0 1 6750
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_116
timestamp 1658881652
transform 1 0 9280 0 1 7290
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_117
timestamp 1658881652
transform 1 0 9280 0 1 7020
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_118
timestamp 1658881652
transform 1 0 13920 0 1 7020
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_119
timestamp 1658881652
transform 1 0 13920 0 1 7290
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_120
timestamp 1658881652
transform 1 0 9280 0 1 7560
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_121
timestamp 1658881652
transform 1 0 13920 0 1 7560
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_122
timestamp 1658881652
transform 1 0 9280 0 1 7830
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_123
timestamp 1658881652
transform 1 0 13920 0 1 7830
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_124
timestamp 1658881652
transform 1 0 9280 0 1 8100
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_125
timestamp 1658881652
transform 1 0 13920 0 1 8100
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_126
timestamp 1658881652
transform 1 0 9280 0 1 8370
box -7 -18 4631 312
use 10T_1x8_magic  10T_1x8_magic_127
timestamp 1658881652
transform 1 0 13920 0 1 8370
box -7 -18 4631 312
<< labels >>
rlabel locali 4640 39 4655 81 1 RBL1_8
port 17 ns signal output
rlabel locali 5177 38 5192 80 1 RBL0_8
port 18 ns signal output
rlabel locali 5220 38 5235 80 1 RBL1_9
port 19 ns signal output
rlabel locali 5757 38 5772 80 1 RBL0_9
port 20 ns signal output
rlabel locali 5800 38 5815 80 1 RBL1_10
port 21 ns signal output
rlabel locali 6337 38 6352 80 1 RBL0_10
port 22 ns signal output
rlabel locali 6380 38 6395 80 1 RBL1_11
port 23 ns signal output
rlabel locali 6917 38 6932 80 1 RBL0_11
port 24 ns signal output
rlabel locali 6960 38 6975 80 1 RBL1_12
port 25 ns signal output
rlabel locali 7497 38 7512 80 1 RBL0_12
port 26 ns signal output
rlabel locali 7540 38 7555 80 1 RBL1_13
port 27 ns signal output
rlabel locali 8077 38 8092 80 1 RBL0_13
port 28 ns signal output
rlabel locali 8120 38 8135 80 1 RBL1_14
port 29 ns signal output
rlabel locali 8657 38 8672 80 1 RBL0_14
port 30 ns signal output
rlabel locali 8700 38 8715 80 1 RBL1_15
port 31 ns signal output
rlabel locali 9237 38 9252 80 1 RBL0_15
port 32 ns signal output
rlabel poly 0 8610 30 8640 1 WWL_0
port 33 ew signal input
rlabel metal1 0 8472 15 8506 1 RWL_0
port 34 ew signal input
rlabel poly 0 8340 30 8370 1 WWL_1
port 35 ew signal input
rlabel metal1 0 8202 15 8236 1 RWL_1
port 36 ew signal input
rlabel poly 0 8070 30 8100 1 WWL_2
port 37 ew signal input
rlabel metal1 0 7932 15 7966 1 RWL_2
port 38 ew signal input
rlabel poly 0 7800 30 7830 1 WWL_3
port 39 ew signal input
rlabel metal1 0 7662 15 7696 1 RWL_3
port 40 ew signal input
rlabel poly 0 7530 30 7560 1 WWL_4
port 41 ew signal input
rlabel metal1 0 7392 15 7426 1 RWL_4
port 42 ew signal input
rlabel poly 0 7260 30 7290 1 WWL_5
port 43 ew signal input
rlabel metal1 0 7122 15 7156 1 RWL_5
port 44 ew signal input
rlabel poly 0 6990 30 7020 1 WWL_6
port 45 ew signal input
rlabel metal1 0 6852 15 6886 1 RWL_6
port 46 ew signal input
rlabel poly 0 6720 30 6750 1 WWL_7
port 47 ew signal input
rlabel metal1 0 6582 15 6616 1 RWL_7
port 48 ew signal input
rlabel poly 0 6450 30 6480 1 WWL_8
port 49 ew signal input
rlabel metal1 0 6312 15 6346 1 RWL_8
port 50 ew signal input
rlabel poly 0 6180 30 6210 1 WWL_9
port 51 ew signal input
rlabel metal1 0 6042 15 6076 1 RWL_9
port 52 ew signal input
rlabel poly 0 5910 30 5940 1 WWL_10
port 53 ew signal input
rlabel metal1 0 5772 15 5806 1 RWL_10
port 54 ew signal input
rlabel poly 0 5640 30 5670 1 WWL_11
port 55 ew signal input
rlabel metal1 0 5502 15 5536 1 RWL_11
port 56 ew signal input
rlabel poly 0 5370 30 5400 1 WWL_12
port 57 ew signal input
rlabel metal1 0 5232 15 5266 1 RWL_12
port 58 ew signal input
rlabel poly 0 5100 30 5130 1 WWL_13
port 59 ew signal input
rlabel metal1 0 4962 15 4996 1 RWL_13
port 60 ew signal input
rlabel poly 0 4830 30 4860 1 WWL_14
port 61 ew signal input
rlabel metal1 0 4692 15 4726 1 RWL_14
port 62 ew signal input
rlabel poly 0 4560 30 4590 1 WWL_15
port 63 ew signal input
rlabel metal1 0 4422 15 4456 1 RWL_15
port 64 ew signal input
rlabel poly 0 4290 30 4320 1 WWL_16
port 65 ew signal input
rlabel metal1 0 4152 15 4186 1 RWL_16
port 66 ew signal input
rlabel poly 0 4020 30 4050 1 WWL_17
port 67 ew signal input
rlabel metal1 0 3882 15 3916 1 RWL_17
port 68 ew signal input
rlabel poly 0 3750 30 3780 1 WWL_18
port 69 ew signal input
rlabel metal1 0 3612 15 3646 1 RWL_18
port 70 ew signal input
rlabel poly 0 3480 30 3510 1 WWL_19
port 71 ew signal input
rlabel metal1 0 3342 15 3376 1 RWL_19
port 72 ew signal input
rlabel poly 0 3210 30 3240 1 WWL_20
port 73 ew signal input
rlabel metal1 0 3072 15 3106 1 RWL_20
port 74 ew signal input
rlabel poly 0 2940 30 2970 1 WWL_21
port 75 ew signal input
rlabel metal1 0 2802 15 2836 1 RWL_21
port 76 ew signal input
rlabel poly 0 2670 30 2700 1 WWL_22
port 77 ew signal input
rlabel metal1 0 2532 15 2566 1 RWL_22
port 78 ew signal input
rlabel poly 0 2400 30 2430 1 WWL_23
port 79 ew signal input
rlabel metal1 0 2262 15 2296 1 RWL_23
port 80 ew signal input
rlabel poly 0 2130 30 2160 1 WWL_24
port 81 ew signal input
rlabel metal1 0 1992 15 2026 1 RWL_24
port 82 ew signal input
rlabel poly 0 1860 30 1890 1 WWL_25
port 83 ew signal input
rlabel metal1 0 1722 15 1756 1 RWL_25
port 84 ew signal input
rlabel poly 0 1590 30 1620 1 WWL_26
port 85 ew signal input
rlabel metal1 0 1452 15 1486 1 RWL_26
port 86 ew signal input
rlabel poly 0 1320 30 1350 1 WWL_27
port 87 ew signal input
rlabel metal1 0 1182 15 1216 1 RWL_27
port 88 ew signal input
rlabel poly 0 1050 30 1080 1 WWL_28
port 89 ew signal input
rlabel metal1 0 912 15 946 1 RWL_28
port 90 ew signal input
rlabel poly 0 780 30 810 1 WWL_29
port 91 ew signal input
rlabel metal1 0 642 15 676 1 RWL_29
port 92 ew signal input
rlabel locali 9280 39 9295 81 1 RBL1_16
port 97 ns signal output
rlabel locali 9817 39 9832 81 1 RBL0_16
port 98 ns signal output
rlabel locali 9860 39 9875 81 1 RBL1_17
port 99 ns signal output
rlabel locali 10397 39 10412 81 1 RBL0_17
port 101 ns signal output
rlabel locali 10440 39 10455 81 1 RBL1_18
port 102 ns signal output
rlabel locali 10977 39 10992 81 1 RBL0_18
port 103 ns signal output
rlabel locali 11020 39 11035 81 1 RBL1_19
port 104 ns signal output
rlabel locali 11557 39 11572 81 1 RBL0_19
port 105 ns signal output
rlabel locali 11600 39 11615 81 1 RBL1_20
port 106 ns signal output
rlabel locali 12137 39 12152 81 1 RBL0_20
port 107 ns signal output
rlabel locali 12180 39 12195 81 1 RBL1_21
port 108 ns signal output
rlabel locali 12717 39 12732 81 1 RBL0_21
port 109 ns signal output
rlabel locali 12760 39 12775 81 1 RBL1_22
port 110 ns signal output
rlabel locali 13297 39 13312 81 1 RBL0_22
port 111 ns signal output
rlabel locali 13340 39 13355 81 1 RBL1_23
port 112 ns signal output
rlabel locali 13877 39 13892 81 1 RBL0_23
port 113 ns signal output
rlabel locali 13920 39 13935 81 1 RBL1_24
port 114 ns signal output
rlabel locali 14457 38 14472 80 1 RBL0_24
port 115 ns signal output
rlabel locali 14500 38 14515 80 1 RBL1_25
port 116 ns signal output
rlabel locali 15037 38 15052 80 1 RBL0_25
port 117 ns signal output
rlabel locali 15080 38 15095 80 1 RBL1_26
port 118 ns signal output
rlabel locali 15617 38 15632 80 1 RBL0_26
port 119 ns signal output
rlabel locali 15660 38 15675 80 1 RBL1_27
port 120 ns signal output
rlabel locali 16197 38 16212 80 1 RBL0_27
port 121 ns signal output
rlabel locali 16240 38 16255 80 1 RBL1_28
port 122 ns signal output
rlabel locali 16777 38 16792 80 1 RBL0_28
port 123 ns signal output
rlabel locali 16820 38 16835 80 1 RBL1_29
port 124 ns signal output
rlabel locali 17357 38 17372 80 1 RBL0_29
port 125 ns signal output
rlabel locali 17400 38 17415 80 1 RBL1_30
port 126 ns signal output
rlabel locali 17937 38 17952 80 1 RBL0_30
port 127 ns signal output
rlabel locali 17980 38 17995 80 1 RBL1_31
port 128 ns signal output
rlabel locali 18517 38 18532 80 1 RBL0_31
port 129 ns signal output
rlabel locali 5104 184 5119 213 1 WBL_8
port 146 ns signal input
rlabel locali 4714 185 4729 213 1 WBLb_8
port 147 ns signal input
rlabel locali 5684 184 5699 213 1 WBL_9
port 148 ns signal input
rlabel locali 5294 184 5309 212 1 WBLb_9
port 149 ns signal input
rlabel locali 6264 184 6279 213 1 WBL_10
port 150 ns signal input
rlabel locali 5874 184 5889 212 1 WBLb_10
port 151 ns signal input
rlabel locali 6844 184 6859 213 1 WBL_11
port 152 ns signal input
rlabel locali 6454 184 6469 212 1 WBLb_11
port 153 ns signal input
rlabel locali 7424 184 7439 213 1 WBL_12
port 154 ns signal input
rlabel locali 7034 184 7049 212 1 WBLb_12
port 155 ns signal input
rlabel locali 8004 184 8019 213 1 WBL_13
port 156 ns signal input
rlabel locali 7614 184 7629 212 1 WBLb_13
port 157 ns signal input
rlabel locali 8584 184 8599 213 1 WBL_14
port 158 ns signal input
rlabel locali 8194 184 8209 212 1 WBLb_14
port 159 ns signal input
rlabel locali 9164 184 9179 213 1 WBL_15
port 160 ns signal input
rlabel locali 8774 184 8789 212 1 WBLb_15
port 161 ns signal input
rlabel locali 9744 185 9759 214 1 WBL_16
port 130 ns signal input
rlabel locali 9354 185 9369 213 1 WBLb_16
port 131 ns signal input
rlabel locali 10324 185 10339 214 1 WBL_17
port 132 ns signal input
rlabel locali 9934 185 9949 213 1 WBLb_17
port 133 ns signal input
rlabel locali 10904 185 10919 214 1 WBL_18
port 134 ns signal input
rlabel locali 10514 185 10529 213 1 WBLb_18
port 135 ns signal input
rlabel locali 11484 185 11499 214 1 WBL_19
port 136 ns signal input
rlabel locali 11094 185 11109 213 1 WBLb_19
port 137 ns signal input
rlabel locali 12064 185 12079 214 1 WBL_20
port 138 ns signal input
rlabel locali 11674 185 11689 213 1 WBLb_20
port 139 ns signal input
rlabel locali 12644 185 12659 214 1 WBL_21
port 140 ns signal input
rlabel locali 12254 185 12269 213 1 WBLb_21
port 141 ns signal input
rlabel locali 13224 185 13239 214 1 WBL_22
port 142 ns signal input
rlabel locali 12834 185 12849 213 1 WBLb_22
port 143 ns signal input
rlabel locali 13804 185 13819 214 1 WBL_23
port 144 ns signal input
rlabel locali 13414 185 13429 213 1 WBLb_23
port 145 ns signal input
rlabel locali 13994 185 14009 213 1 WBLb_24
port 147 ns signal input
rlabel locali 14384 185 14399 214 1 WBL_24
port 146 ns signal input
rlabel locali 14964 185 14979 214 1 WBL_25
port 148 ns signal input
rlabel locali 14574 185 14589 213 1 WBLb_25
port 149 ns signal input
rlabel locali 15544 185 15559 214 1 WBL_26
port 150 ns signal input
rlabel locali 15154 185 15169 213 1 WBLb_26
port 151 ns signal input
rlabel locali 16124 185 16139 214 1 WBL_27
port 152 ns signal input
rlabel locali 15734 185 15749 213 1 WBLb_27
port 153 ns signal input
rlabel locali 16704 185 16719 214 1 WBL_28
port 154 ns signal input
rlabel locali 16314 185 16329 213 1 WBLb_28
port 155 ns signal input
rlabel locali 17284 185 17299 214 1 WBL_29
port 156 ns signal input
rlabel locali 16894 185 16909 213 1 WBLb_29
port 157 ns signal input
rlabel locali 17864 185 17879 214 1 WBL_30
port 158 ns signal input
rlabel locali 17474 185 17489 213 1 WBLb_30
port 159 ns signal input
rlabel locali 18444 185 18459 214 1 WBL_31
port 160 ns signal input
rlabel locali 18054 185 18069 213 1 WBLb_31
port 161 ns signal input
rlabel metal1 0 8596 15 8610 1 VDD
port 162 ew power bidirectional abutment
rlabel metal1 0 8370 15 8384 1 GND
port 163 ew ground bidirectional abutment
rlabel metal1 0 8326 15 8340 1 VDD
port 162 ew power bidirectional abutment
rlabel metal1 0 8100 15 8114 1 GND
port 163 ew ground bidirectional abutment
rlabel metal1 0 8056 15 8070 1 VDD
port 162 ew power bidirectional abutment
rlabel metal1 0 7830 15 7844 1 GND
port 163 ew ground bidirectional abutment
rlabel metal1 0 7786 15 7800 1 VDD
port 162 ew power bidirectional abutment
rlabel metal1 0 7560 15 7574 1 GND
port 163 ew ground bidirectional abutment
rlabel metal1 0 7516 15 7530 1 VDD
port 162 ew power bidirectional abutment
rlabel metal1 0 7290 15 7304 1 GND
port 163 ew ground bidirectional abutment
rlabel metal1 0 7246 15 7260 1 VDD
port 162 ew power bidirectional abutment
rlabel metal1 0 7020 15 7034 1 GND
port 163 ew ground bidirectional abutment
rlabel metal1 0 6976 15 6990 1 VDD
port 162 ew power bidirectional abutment
rlabel metal1 0 6750 15 6764 1 GND
port 163 ew ground bidirectional abutment
rlabel metal1 0 6706 15 6720 1 VDD
port 162 ew power bidirectional abutment
rlabel metal1 0 6480 15 6494 1 GND
port 163 ew ground bidirectional abutment
rlabel metal1 0 6436 15 6450 1 VDD
port 162 ew power bidirectional abutment
rlabel metal1 0 6210 15 6224 1 GND
port 163 ew ground bidirectional abutment
rlabel metal1 0 6166 15 6180 1 VDD
port 162 ew power bidirectional abutment
rlabel metal1 0 5940 15 5954 1 GND
port 163 ew ground bidirectional abutment
rlabel metal1 0 5896 15 5910 1 VDD
port 162 ew power bidirectional abutment
rlabel metal1 0 5670 15 5684 1 GND
port 163 ew ground bidirectional abutment
rlabel metal1 0 5626 15 5640 1 VDD
port 162 ew power bidirectional abutment
rlabel metal1 0 5400 15 5414 1 GND
port 163 ew ground bidirectional abutment
rlabel metal1 0 5356 15 5370 1 VDD
port 162 ew power bidirectional abutment
rlabel metal1 0 5130 15 5144 1 GND
port 163 ew ground bidirectional abutment
rlabel metal1 0 5086 15 5100 1 VDD
port 162 ew power bidirectional abutment
rlabel metal1 0 4860 15 4874 1 GND
port 163 ew ground bidirectional abutment
rlabel metal1 0 4816 15 4830 1 VDD
port 162 ew power bidirectional abutment
rlabel metal1 0 4590 15 4604 1 GND
port 163 ew ground bidirectional abutment
rlabel metal1 0 4546 15 4560 1 VDD
port 162 ew power bidirectional abutment
rlabel metal1 0 4320 15 4334 1 GND
port 163 ew ground bidirectional abutment
rlabel metal1 0 4276 15 4290 1 VDD
port 162 ew power bidirectional abutment
rlabel metal1 0 4050 15 4064 1 GND
port 163 ew ground bidirectional abutment
rlabel metal1 0 4006 15 4020 1 VDD
port 162 ew power bidirectional abutment
rlabel metal1 0 3780 15 3794 1 GND
port 163 ew ground bidirectional abutment
rlabel metal1 0 3736 15 3750 1 VDD
port 162 ew power bidirectional abutment
rlabel metal1 0 3510 15 3524 1 GND
port 163 ew ground bidirectional abutment
rlabel metal1 0 3466 15 3480 1 VDD
port 162 ew power bidirectional abutment
rlabel metal1 0 3240 15 3254 1 GND
port 163 ew ground bidirectional abutment
rlabel metal1 0 3196 15 3210 1 VDD
port 162 ew power bidirectional abutment
rlabel metal1 0 2926 15 2940 1 VDD
port 162 ew power bidirectional abutment
rlabel metal1 0 2970 15 2984 1 GND
port 163 ew ground bidirectional abutment
rlabel metal1 0 2700 15 2714 1 GND
port 163 ew ground bidirectional abutment
rlabel metal1 0 2656 15 2670 1 VDD
port 162 ew power bidirectional abutment
rlabel metal1 0 2430 15 2444 1 GND
port 163 ew ground bidirectional abutment
rlabel metal1 0 2386 15 2400 1 VDD
port 162 ew power bidirectional abutment
rlabel metal1 0 2160 15 2174 1 GND
port 163 ew ground bidirectional abutment
rlabel metal1 0 2116 15 2130 1 VDD
port 162 ew power bidirectional abutment
rlabel metal1 0 1890 15 1904 1 GND
port 163 ew ground bidirectional abutment
rlabel metal1 0 1846 15 1860 1 VDD
port 162 ew power bidirectional abutment
rlabel metal1 0 1620 15 1634 1 GND
port 163 ew ground bidirectional abutment
rlabel metal1 0 1576 15 1590 1 VDD
port 162 ew power bidirectional abutment
rlabel metal1 0 1350 15 1364 1 GND
port 163 ew ground bidirectional abutment
rlabel metal1 0 1306 15 1320 1 VDD
port 162 ew power bidirectional abutment
rlabel metal1 0 1080 15 1094 1 GND
port 163 ew ground bidirectional abutment
rlabel metal1 0 1036 15 1050 1 VDD
port 162 ew power bidirectional abutment
rlabel metal1 0 810 15 824 1 GND
port 163 ew ground bidirectional abutment
rlabel metal1 0 766 15 780 1 VDD
port 162 ew power bidirectional abutment
rlabel metal1 0 540 15 554 1 GND
port 163 ew ground bidirectional abutment
rlabel locali 0 38 15 80 1 RBL1_0
port 1 ns signal output
rlabel locali 537 38 552 80 1 RBL0_0
port 2 ns signal output
rlabel locali 580 38 595 80 1 RBL1_1
port 3 ns signal output
rlabel locali 1117 38 1132 80 1 RBL0_1
port 4 ns signal output
rlabel locali 1160 38 1175 80 1 RBL1_2
port 5 ns signal output
rlabel locali 1697 38 1712 80 1 RBL0_2
port 6 ns signal output
rlabel locali 1740 38 1755 80 1 RBL1_3
port 7 ns signal output
rlabel locali 2277 38 2292 80 1 RBL0_3
port 8 ns signal output
rlabel locali 2320 38 2335 80 1 RBL1_4
port 9 ns signal output
rlabel locali 2857 38 2872 80 1 RBL0_4
port 10 ns signal output
rlabel locali 2900 38 2915 80 1 RBL1_5
port 11 ns signal output
rlabel locali 3437 38 3452 80 1 RBL0_5
port 12 ns signal output
rlabel locali 3480 38 3495 80 1 RBL1_6
port 13 ns signal output
rlabel locali 4017 38 4032 80 1 RBL0_6
port 14 ns signal output
rlabel locali 4060 38 4075 80 1 RBL1_7
port 15 ns signal output
rlabel locali 4597 38 4612 80 1 RBL0_7
port 16 ns signal output
rlabel poly 0 240 30 270 1 WWL_31
port 95 ew signal input
rlabel metal1 0 102 15 136 1 RWL_31
port 96 ew signal input
rlabel locali 464 184 479 213 1 WBL_0
port 130 ns signal input
rlabel locali 74 184 89 212 1 WBLb_0
port 131 ns signal input
rlabel locali 1044 184 1059 213 1 WBL_1
port 132 ns signal input
rlabel locali 654 184 669 212 1 WBLb_1
port 133 ns signal input
rlabel locali 1624 184 1639 213 1 WBL_2
port 134 ns signal input
rlabel locali 1234 184 1249 212 1 WBLb_2
port 135 ns signal input
rlabel locali 2204 184 2219 213 1 WBL_3
port 136 ns signal input
rlabel locali 1814 184 1829 212 1 WBLb_3
port 137 ns signal input
rlabel locali 2784 184 2799 213 1 WBL_4
port 138 ns signal input
rlabel locali 2394 184 2409 212 1 WBLb_4
port 139 ns signal input
rlabel locali 3364 184 3379 213 1 WBL_5
port 140 ns signal input
rlabel locali 2974 184 2989 212 1 WBLb_5
port 141 ns signal input
rlabel locali 3944 184 3959 213 1 WBL_6
port 142 ns signal input
rlabel locali 3554 184 3569 212 1 WBLb_6
port 143 ns signal input
rlabel locali 4524 184 4539 213 1 WBL_7
port 144 ns signal input
rlabel locali 4134 184 4149 212 1 WBLb_7
port 145 ns signal input
rlabel metal1 0 226 15 240 1 VDD
port 162 ew power bidirectional abutment
rlabel metal1 0 0 15 14 1 GND
port 163 ew ground bidirectional abutment
rlabel space 0 269 15 283 1 GND
port 163 ew ground bidirectional abutment
rlabel metal1 0 371 15 405 1 RWL_30
port 94 ew signal input
rlabel metal1 0 495 15 509 1 VDD
port 162 ew power bidirectional abutment
rlabel poly 0 509 30 539 1 WWL_30
port 93 ew signal input
<< end >>
