magic
tech sky130A
magscale 1 2
timestamp 1658883737
<< nwell >>
rect 198 144 351 240
rect 778 144 931 240
rect 1358 144 1511 240
rect 1938 144 2091 240
rect 2518 144 2671 240
rect 3098 144 3251 240
rect 3678 144 3831 240
rect 4258 144 4411 240
<< pwell >>
rect 0 98 170 270
rect 382 98 750 270
rect 962 98 1330 270
rect 1542 98 1910 270
rect 2122 98 2490 270
rect 2702 98 3070 270
rect 3282 98 3650 270
rect 3862 98 4230 270
rect 4442 98 4612 270
rect 0 0 4612 98
<< nmos >>
rect 107 184 137 212
rect 415 184 445 212
rect 687 184 717 212
rect 995 184 1025 212
rect 1267 184 1297 212
rect 1575 184 1605 212
rect 1847 184 1877 212
rect 2155 184 2185 212
rect 2427 184 2457 212
rect 2735 184 2765 212
rect 3007 184 3037 212
rect 3315 184 3345 212
rect 3587 184 3617 212
rect 3895 184 3925 212
rect 4167 184 4197 212
rect 4475 184 4505 212
rect 43 38 73 80
rect 479 38 509 80
rect 623 38 653 80
rect 1059 38 1089 80
rect 1203 38 1233 80
rect 1639 38 1669 80
rect 1783 38 1813 80
rect 2219 38 2249 80
rect 2363 38 2393 80
rect 2799 38 2829 80
rect 2943 38 2973 80
rect 3379 38 3409 80
rect 3523 38 3553 80
rect 3959 38 3989 80
rect 4103 38 4133 80
rect 4539 38 4569 80
<< npd >>
rect 222 38 252 80
rect 300 38 330 80
rect 802 38 832 80
rect 880 38 910 80
rect 1382 38 1412 80
rect 1460 38 1490 80
rect 1962 38 1992 80
rect 2040 38 2070 80
rect 2542 38 2572 80
rect 2620 38 2650 80
rect 3122 38 3152 80
rect 3200 38 3230 80
rect 3702 38 3732 80
rect 3780 38 3810 80
rect 4282 38 4312 80
rect 4360 38 4390 80
<< npass >>
rect 129 38 159 66
rect 393 38 423 66
rect 709 38 739 66
rect 973 38 1003 66
rect 1289 38 1319 66
rect 1553 38 1583 66
rect 1869 38 1899 66
rect 2133 38 2163 66
rect 2449 38 2479 66
rect 2713 38 2743 66
rect 3029 38 3059 66
rect 3293 38 3323 66
rect 3609 38 3639 66
rect 3873 38 3903 66
rect 4189 38 4219 66
rect 4453 38 4483 66
<< ppu >>
rect 222 174 252 202
rect 300 174 330 202
rect 802 174 832 202
rect 880 174 910 202
rect 1382 174 1412 202
rect 1460 174 1490 202
rect 1962 174 1992 202
rect 2040 174 2070 202
rect 2542 174 2572 202
rect 2620 174 2650 202
rect 3122 174 3152 202
rect 3200 174 3230 202
rect 3702 174 3732 202
rect 3780 174 3810 202
rect 4282 174 4312 202
rect 4360 174 4390 202
<< ndiff >>
rect 89 184 107 212
rect 137 184 155 212
rect 397 184 415 212
rect 445 184 464 212
rect 669 184 687 212
rect 717 184 735 212
rect 977 184 995 212
rect 1025 184 1044 212
rect 1249 184 1267 212
rect 1297 184 1315 212
rect 1557 184 1575 212
rect 1605 184 1624 212
rect 1829 184 1847 212
rect 1877 184 1895 212
rect 2137 184 2155 212
rect 2185 184 2204 212
rect 2409 184 2427 212
rect 2457 184 2475 212
rect 2717 184 2735 212
rect 2765 184 2784 212
rect 2989 184 3007 212
rect 3037 184 3055 212
rect 3297 184 3315 212
rect 3345 184 3364 212
rect 3569 184 3587 212
rect 3617 184 3635 212
rect 3877 184 3895 212
rect 3925 184 3944 212
rect 4149 184 4167 212
rect 4197 184 4215 212
rect 4457 184 4475 212
rect 4505 184 4524 212
rect 15 38 43 80
rect 73 66 98 80
rect 197 70 222 80
rect 73 38 129 66
rect 159 38 193 66
tri 207 63 214 70 ne
rect 214 38 222 70
rect 252 38 300 80
rect 330 70 355 80
rect 330 38 338 70
rect 454 66 479 80
rect 359 38 393 66
rect 423 38 479 66
rect 509 38 537 80
rect 595 38 623 80
rect 653 66 678 80
rect 777 70 802 80
rect 653 38 709 66
rect 739 38 773 66
tri 787 63 794 70 ne
rect 794 38 802 70
rect 832 38 880 80
rect 910 70 935 80
rect 910 38 918 70
rect 1034 66 1059 80
rect 939 38 973 66
rect 1003 38 1059 66
rect 1089 38 1117 80
rect 1175 38 1203 80
rect 1233 66 1258 80
rect 1357 70 1382 80
rect 1233 38 1289 66
rect 1319 38 1353 66
tri 1367 63 1374 70 ne
rect 1374 38 1382 70
rect 1412 38 1460 80
rect 1490 70 1515 80
rect 1490 38 1498 70
rect 1614 66 1639 80
rect 1519 38 1553 66
rect 1583 38 1639 66
rect 1669 38 1697 80
rect 1755 38 1783 80
rect 1813 66 1838 80
rect 1937 70 1962 80
rect 1813 38 1869 66
rect 1899 38 1933 66
tri 1947 63 1954 70 ne
rect 1954 38 1962 70
rect 1992 38 2040 80
rect 2070 70 2095 80
rect 2070 38 2078 70
rect 2194 66 2219 80
rect 2099 38 2133 66
rect 2163 38 2219 66
rect 2249 38 2277 80
rect 2335 38 2363 80
rect 2393 66 2418 80
rect 2517 70 2542 80
rect 2393 38 2449 66
rect 2479 38 2513 66
tri 2527 63 2534 70 ne
rect 2534 38 2542 70
rect 2572 38 2620 80
rect 2650 70 2675 80
rect 2650 38 2658 70
rect 2774 66 2799 80
rect 2679 38 2713 66
rect 2743 38 2799 66
rect 2829 38 2857 80
rect 2915 38 2943 80
rect 2973 66 2998 80
rect 3097 70 3122 80
rect 2973 38 3029 66
rect 3059 38 3093 66
tri 3107 63 3114 70 ne
rect 3114 38 3122 70
rect 3152 38 3200 80
rect 3230 70 3255 80
rect 3230 38 3238 70
rect 3354 66 3379 80
rect 3259 38 3293 66
rect 3323 38 3379 66
rect 3409 38 3437 80
rect 3495 38 3523 80
rect 3553 66 3578 80
rect 3677 70 3702 80
rect 3553 38 3609 66
rect 3639 38 3673 66
tri 3687 63 3694 70 ne
rect 3694 38 3702 70
rect 3732 38 3780 80
rect 3810 70 3835 80
rect 3810 38 3818 70
rect 3934 66 3959 80
rect 3839 38 3873 66
rect 3903 38 3959 66
rect 3989 38 4017 80
rect 4075 38 4103 80
rect 4133 66 4158 80
rect 4257 70 4282 80
rect 4133 38 4189 66
rect 4219 38 4253 66
tri 4267 63 4274 70 ne
rect 4274 38 4282 70
rect 4312 38 4360 80
rect 4390 70 4415 80
rect 4390 38 4398 70
rect 4514 66 4539 80
rect 4419 38 4453 66
rect 4483 38 4539 66
rect 4569 38 4597 80
rect 166 14 193 38
rect 260 16 292 38
rect 260 14 262 16
rect 290 14 292 16
rect 359 14 386 38
rect 166 0 260 14
rect 292 0 386 14
rect 746 14 773 38
rect 840 16 872 38
rect 840 14 842 16
rect 870 14 872 16
rect 939 14 966 38
rect 746 0 840 14
rect 872 0 966 14
rect 1326 14 1353 38
rect 1420 16 1452 38
rect 1420 14 1422 16
rect 1450 14 1452 16
rect 1519 14 1546 38
rect 1326 0 1420 14
rect 1452 0 1546 14
rect 1906 14 1933 38
rect 2000 16 2032 38
rect 2000 14 2002 16
rect 2030 14 2032 16
rect 2099 14 2126 38
rect 1906 0 2000 14
rect 2032 0 2126 14
rect 2486 14 2513 38
rect 2580 16 2612 38
rect 2580 14 2582 16
rect 2610 14 2612 16
rect 2679 14 2706 38
rect 2486 0 2580 14
rect 2612 0 2706 14
rect 3066 14 3093 38
rect 3160 16 3192 38
rect 3160 14 3162 16
rect 3190 14 3192 16
rect 3259 14 3286 38
rect 3066 0 3160 14
rect 3192 0 3286 14
rect 3646 14 3673 38
rect 3740 16 3772 38
rect 3740 14 3742 16
rect 3770 14 3772 16
rect 3839 14 3866 38
rect 3646 0 3740 14
rect 3772 0 3866 14
rect 4226 14 4253 38
rect 4320 16 4352 38
rect 4320 14 4322 16
rect 4350 14 4352 16
rect 4419 14 4446 38
rect 4226 0 4320 14
rect 4352 0 4446 14
<< pdiff >>
rect 260 224 262 226
rect 290 224 292 226
rect 260 202 292 224
rect 213 174 222 202
rect 252 174 300 202
rect 330 174 339 202
tri 339 174 351 186 sw
rect 840 224 842 226
rect 870 224 872 226
rect 840 202 872 224
rect 793 174 802 202
rect 832 174 880 202
rect 910 174 919 202
tri 919 174 931 186 sw
rect 1420 224 1422 226
rect 1450 224 1452 226
rect 1420 202 1452 224
rect 1373 174 1382 202
rect 1412 174 1460 202
rect 1490 174 1499 202
tri 1499 174 1511 186 sw
rect 2000 224 2002 226
rect 2030 224 2032 226
rect 2000 202 2032 224
rect 1953 174 1962 202
rect 1992 174 2040 202
rect 2070 174 2079 202
tri 2079 174 2091 186 sw
rect 2580 224 2582 226
rect 2610 224 2612 226
rect 2580 202 2612 224
rect 2533 174 2542 202
rect 2572 174 2620 202
rect 2650 174 2659 202
tri 2659 174 2671 186 sw
rect 3160 224 3162 226
rect 3190 224 3192 226
rect 3160 202 3192 224
rect 3113 174 3122 202
rect 3152 174 3200 202
rect 3230 174 3239 202
tri 3239 174 3251 186 sw
rect 3740 224 3742 226
rect 3770 224 3772 226
rect 3740 202 3772 224
rect 3693 174 3702 202
rect 3732 174 3780 202
rect 3810 174 3819 202
tri 3819 174 3831 186 sw
rect 4320 224 4322 226
rect 4350 224 4352 226
rect 4320 202 4352 224
rect 4273 174 4282 202
rect 4312 174 4360 202
rect 4390 174 4399 202
tri 4399 174 4411 186 sw
<< ndiffc >>
rect 74 184 89 212
rect 155 184 170 212
rect 382 184 397 212
rect 464 184 479 213
rect 654 184 669 212
rect 735 184 750 212
rect 962 184 977 212
rect 1044 184 1059 213
rect 1234 184 1249 212
rect 1315 184 1330 212
rect 1542 184 1557 212
rect 1624 184 1639 213
rect 1814 184 1829 212
rect 1895 184 1910 212
rect 2122 184 2137 212
rect 2204 184 2219 213
rect 2394 184 2409 212
rect 2475 184 2490 212
rect 2702 184 2717 212
rect 2784 184 2799 213
rect 2974 184 2989 212
rect 3055 184 3070 212
rect 3282 184 3297 212
rect 3364 184 3379 213
rect 3554 184 3569 212
rect 3635 184 3650 212
rect 3862 184 3877 212
rect 3944 184 3959 213
rect 4134 184 4149 212
rect 4215 184 4230 212
rect 4442 184 4457 212
rect 4524 184 4539 213
rect 0 38 15 80
rect 197 63 207 70
tri 207 63 214 70 sw
rect 197 38 214 63
rect 338 38 355 70
rect 537 38 552 80
rect 580 38 595 80
rect 777 63 787 70
tri 787 63 794 70 sw
rect 777 38 794 63
rect 918 38 935 70
rect 1117 38 1132 80
rect 1160 38 1175 80
rect 1357 63 1367 70
tri 1367 63 1374 70 sw
rect 1357 38 1374 63
rect 1498 38 1515 70
rect 1697 38 1712 80
rect 1740 38 1755 80
rect 1937 63 1947 70
tri 1947 63 1954 70 sw
rect 1937 38 1954 63
rect 2078 38 2095 70
rect 2277 38 2292 80
rect 2320 38 2335 80
rect 2517 63 2527 70
tri 2527 63 2534 70 sw
rect 2517 38 2534 63
rect 2658 38 2675 70
rect 2857 38 2872 80
rect 2900 38 2915 80
rect 3097 63 3107 70
tri 3107 63 3114 70 sw
rect 3097 38 3114 63
rect 3238 38 3255 70
rect 3437 38 3452 80
rect 3480 38 3495 80
rect 3677 63 3687 70
tri 3687 63 3694 70 sw
rect 3677 38 3694 63
rect 3818 38 3835 70
rect 4017 38 4032 80
rect 4060 38 4075 80
rect 4257 63 4267 70
tri 4267 63 4274 70 sw
rect 4257 38 4274 63
rect 4398 38 4415 70
rect 4597 38 4612 80
rect 260 0 292 14
rect 840 0 872 14
rect 1420 0 1452 14
rect 2000 0 2032 14
rect 2580 0 2612 14
rect 3160 0 3192 14
rect 3740 0 3772 14
rect 4320 0 4352 14
<< pdiffc >>
rect 260 226 292 240
rect 198 174 213 202
rect 339 186 351 202
tri 339 174 351 186 ne
rect 840 226 872 240
rect 778 174 793 202
rect 919 186 931 202
tri 919 174 931 186 ne
rect 1420 226 1452 240
rect 1358 174 1373 202
rect 1499 186 1511 202
tri 1499 174 1511 186 ne
rect 2000 226 2032 240
rect 1938 174 1953 202
rect 2079 186 2091 202
tri 2079 174 2091 186 ne
rect 2580 226 2612 240
rect 2518 174 2533 202
rect 2659 186 2671 202
tri 2659 174 2671 186 ne
rect 3160 226 3192 240
rect 3098 174 3113 202
rect 3239 186 3251 202
tri 3239 174 3251 186 ne
rect 3740 226 3772 240
rect 3678 174 3693 202
rect 3819 186 3831 202
tri 3819 174 3831 186 ne
rect 4320 226 4352 240
rect 4258 174 4273 202
rect 4399 186 4411 202
tri 4399 174 4411 186 ne
<< psubdiffcont >>
rect 262 14 290 16
rect 842 14 870 16
rect 1422 14 1450 16
rect 2002 14 2030 16
rect 2582 14 2610 16
rect 3162 14 3190 16
rect 3742 14 3770 16
rect 4322 14 4350 16
<< nsubdiffcont >>
rect 262 224 290 226
rect 842 224 870 226
rect 1422 224 1450 226
rect 2002 224 2030 226
rect 2582 224 2610 226
rect 3162 224 3190 226
rect 3742 224 3770 226
rect 4322 224 4350 226
<< poly >>
rect 0 240 4612 270
rect 107 212 137 240
rect 222 202 252 224
rect 300 202 330 224
rect 415 212 445 240
rect 107 162 137 184
rect 687 212 717 240
rect 802 202 832 224
rect 880 202 910 224
rect 995 212 1025 240
rect 222 141 252 174
rect 43 80 73 102
rect 129 80 144 114
rect 222 80 252 107
rect 300 141 330 174
rect 415 162 445 184
rect 687 162 717 184
rect 1267 212 1297 240
rect 1382 202 1412 224
rect 1460 202 1490 224
rect 1575 212 1605 240
rect 802 141 832 174
rect 300 80 330 107
rect 408 80 423 114
rect 479 80 509 102
rect 623 80 653 102
rect 709 80 724 114
rect 802 80 832 107
rect 880 141 910 174
rect 995 162 1025 184
rect 1267 162 1297 184
rect 1847 212 1877 240
rect 1962 202 1992 224
rect 2040 202 2070 224
rect 2155 212 2185 240
rect 1382 141 1412 174
rect 880 80 910 107
rect 988 80 1003 114
rect 1059 80 1089 102
rect 1203 80 1233 102
rect 1289 80 1304 114
rect 1382 80 1412 107
rect 1460 141 1490 174
rect 1575 162 1605 184
rect 1847 162 1877 184
rect 2427 212 2457 240
rect 2542 202 2572 224
rect 2620 202 2650 224
rect 2735 212 2765 240
rect 1962 141 1992 174
rect 1460 80 1490 107
rect 1568 80 1583 114
rect 1639 80 1669 102
rect 1783 80 1813 102
rect 1869 80 1884 114
rect 1962 80 1992 107
rect 2040 141 2070 174
rect 2155 162 2185 184
rect 2427 162 2457 184
rect 3007 212 3037 240
rect 3122 202 3152 224
rect 3200 202 3230 224
rect 3315 212 3345 240
rect 2542 141 2572 174
rect 2040 80 2070 107
rect 2148 80 2163 114
rect 2219 80 2249 102
rect 2363 80 2393 102
rect 2449 80 2464 114
rect 2542 80 2572 107
rect 2620 141 2650 174
rect 2735 162 2765 184
rect 3007 162 3037 184
rect 3587 212 3617 240
rect 3702 202 3732 224
rect 3780 202 3810 224
rect 3895 212 3925 240
rect 3122 141 3152 174
rect 2620 80 2650 107
rect 2728 80 2743 114
rect 2799 80 2829 102
rect 2943 80 2973 102
rect 3029 80 3044 114
rect 3122 80 3152 107
rect 3200 141 3230 174
rect 3315 162 3345 184
rect 3587 162 3617 184
rect 4167 212 4197 240
rect 4282 202 4312 224
rect 4360 202 4390 224
rect 4475 212 4505 240
rect 3702 141 3732 174
rect 3200 80 3230 107
rect 3308 80 3323 114
rect 3379 80 3409 102
rect 3523 80 3553 102
rect 3609 80 3624 114
rect 3702 80 3732 107
rect 3780 141 3810 174
rect 3895 162 3925 184
rect 4167 162 4197 184
rect 4282 141 4312 174
rect 3780 80 3810 107
rect 3888 80 3903 114
rect 3959 80 3989 102
rect 4103 80 4133 102
rect 4189 80 4204 114
rect 4282 80 4312 107
rect 4360 141 4390 174
rect 4475 162 4505 184
rect 4360 80 4390 107
rect 4468 80 4483 114
rect 4539 80 4569 102
rect 129 66 159 80
rect 393 66 423 80
rect 709 66 739 80
rect 973 66 1003 80
rect 1289 66 1319 80
rect 1553 66 1583 80
rect 1869 66 1899 80
rect 2133 66 2163 80
rect 2449 66 2479 80
rect 2713 66 2743 80
rect 3029 66 3059 80
rect 3293 66 3323 80
rect 3609 66 3639 80
rect 3873 66 3903 80
rect 4189 66 4219 80
rect 4453 66 4483 80
rect 43 16 73 38
rect 129 16 159 38
rect 222 16 252 38
rect 300 16 330 38
rect 393 16 423 38
rect 479 16 509 38
rect 623 16 653 38
rect 709 16 739 38
rect 802 16 832 38
rect 880 16 910 38
rect 973 16 1003 38
rect 1059 16 1089 38
rect 1203 16 1233 38
rect 1289 16 1319 38
rect 1382 16 1412 38
rect 1460 16 1490 38
rect 1553 16 1583 38
rect 1639 16 1669 38
rect 1783 16 1813 38
rect 1869 16 1899 38
rect 1962 16 1992 38
rect 2040 16 2070 38
rect 2133 16 2163 38
rect 2219 16 2249 38
rect 2363 16 2393 38
rect 2449 16 2479 38
rect 2542 16 2572 38
rect 2620 16 2650 38
rect 2713 16 2743 38
rect 2799 16 2829 38
rect 2943 16 2973 38
rect 3029 16 3059 38
rect 3122 16 3152 38
rect 3200 16 3230 38
rect 3293 16 3323 38
rect 3379 16 3409 38
rect 3523 16 3553 38
rect 3609 16 3639 38
rect 3702 16 3732 38
rect 3780 16 3810 38
rect 3873 16 3903 38
rect 3959 16 3989 38
rect 4103 16 4133 38
rect 4189 16 4219 38
rect 4282 16 4312 38
rect 4360 16 4390 38
rect 4453 16 4483 38
rect 4539 16 4569 38
<< polycont >>
rect 43 102 73 136
rect 144 80 174 114
rect 222 107 252 141
rect 300 107 330 141
rect 378 80 408 114
rect 479 102 509 136
rect 623 102 653 136
rect 724 80 754 114
rect 802 107 832 141
rect 880 107 910 141
rect 958 80 988 114
rect 1059 102 1089 136
rect 1203 102 1233 136
rect 1304 80 1334 114
rect 1382 107 1412 141
rect 1460 107 1490 141
rect 1538 80 1568 114
rect 1639 102 1669 136
rect 1783 102 1813 136
rect 1884 80 1914 114
rect 1962 107 1992 141
rect 2040 107 2070 141
rect 2118 80 2148 114
rect 2219 102 2249 136
rect 2363 102 2393 136
rect 2464 80 2494 114
rect 2542 107 2572 141
rect 2620 107 2650 141
rect 2698 80 2728 114
rect 2799 102 2829 136
rect 2943 102 2973 136
rect 3044 80 3074 114
rect 3122 107 3152 141
rect 3200 107 3230 141
rect 3278 80 3308 114
rect 3379 102 3409 136
rect 3523 102 3553 136
rect 3624 80 3654 114
rect 3702 107 3732 141
rect 3780 107 3810 141
rect 3858 80 3888 114
rect 3959 102 3989 136
rect 4103 102 4133 136
rect 4204 80 4234 114
rect 4282 107 4312 141
rect 4360 107 4390 141
rect 4438 80 4468 114
rect 4539 102 4569 136
<< corelocali >>
rect 0 80 15 270
tri 80 234 102 256 se
rect 102 249 117 270
tri 102 234 117 249 nw
rect 436 249 451 270
tri 74 228 80 234 se
rect 80 228 89 234
rect 74 212 89 228
tri 89 221 102 234 nw
rect 243 226 260 240
rect 292 226 309 240
tri 436 234 451 249 ne
tri 451 234 473 256 sw
rect 74 176 89 184
rect 155 212 215 226
rect 170 202 215 212
rect 170 184 198 202
tri 74 161 89 176 ne
tri 89 161 111 183 sw
rect 155 174 198 184
rect 213 198 215 202
rect 337 212 397 226
tri 451 221 464 234 ne
rect 464 228 473 234
tri 473 228 479 234 sw
rect 337 202 382 212
rect 213 174 287 198
rect 155 170 287 174
tri 287 170 315 198 sw
rect 337 188 339 202
tri 337 186 339 188 ne
rect 351 184 382 202
rect 351 174 397 184
rect 464 213 479 228
tri 89 149 101 161 ne
rect 101 156 111 161
tri 111 156 116 161 sw
rect 0 0 15 38
rect 101 0 116 156
rect 155 114 183 170
tri 275 152 293 170 ne
rect 293 150 315 170
tri 315 150 335 170 sw
tri 351 156 369 174 ne
rect 174 80 183 114
rect 217 141 259 142
rect 217 107 222 141
rect 252 107 259 141
rect 217 98 259 107
rect 293 141 335 150
rect 293 107 300 141
rect 330 107 335 141
rect 293 102 335 107
rect 369 114 397 174
tri 442 161 464 183 se
rect 464 176 479 184
tri 464 161 479 176 nw
tri 436 155 442 161 se
rect 442 155 451 161
rect 155 70 183 80
tri 183 70 207 94 sw
rect 155 38 197 70
tri 214 62 215 63 sw
rect 214 38 215 62
tri 217 61 254 98 ne
rect 254 70 259 98
tri 259 70 285 96 sw
rect 369 80 378 114
rect 369 70 397 80
rect 254 61 338 70
tri 254 42 273 61 ne
rect 273 42 338 61
rect 155 16 215 38
rect 337 38 338 42
rect 355 38 397 70
rect 337 16 397 38
rect 243 0 260 14
rect 292 0 309 14
rect 436 0 451 155
tri 451 148 464 161 nw
rect 537 80 552 270
rect 537 0 552 38
rect 580 80 595 270
tri 660 234 682 256 se
rect 682 249 697 270
tri 682 234 697 249 nw
rect 1016 249 1031 270
tri 654 228 660 234 se
rect 660 228 669 234
rect 654 212 669 228
tri 669 221 682 234 nw
rect 823 226 840 240
rect 872 226 889 240
tri 1016 234 1031 249 ne
tri 1031 234 1053 256 sw
rect 654 176 669 184
rect 735 212 795 226
rect 750 202 795 212
rect 750 184 778 202
tri 654 161 669 176 ne
tri 669 161 691 183 sw
rect 735 174 778 184
rect 793 198 795 202
rect 917 212 977 226
tri 1031 221 1044 234 ne
rect 1044 228 1053 234
tri 1053 228 1059 234 sw
rect 917 202 962 212
rect 793 174 867 198
rect 735 170 867 174
tri 867 170 895 198 sw
rect 917 188 919 202
tri 917 186 919 188 ne
rect 931 184 962 202
rect 931 174 977 184
rect 1044 213 1059 228
tri 669 149 681 161 ne
rect 681 156 691 161
tri 691 156 696 161 sw
rect 580 0 595 38
rect 681 0 696 156
rect 735 114 763 170
tri 855 152 873 170 ne
rect 873 150 895 170
tri 895 150 915 170 sw
tri 931 156 949 174 ne
rect 754 80 763 114
rect 797 141 839 142
rect 797 107 802 141
rect 832 107 839 141
rect 797 98 839 107
rect 873 141 915 150
rect 873 107 880 141
rect 910 107 915 141
rect 873 102 915 107
rect 949 114 977 174
tri 1022 161 1044 183 se
rect 1044 176 1059 184
tri 1044 161 1059 176 nw
tri 1016 155 1022 161 se
rect 1022 155 1031 161
rect 735 70 763 80
tri 763 70 787 94 sw
rect 735 38 777 70
tri 794 62 795 63 sw
rect 794 38 795 62
tri 797 61 834 98 ne
rect 834 70 839 98
tri 839 70 865 96 sw
rect 949 80 958 114
rect 949 70 977 80
rect 834 61 918 70
tri 834 42 853 61 ne
rect 853 42 918 61
rect 735 16 795 38
rect 917 38 918 42
rect 935 38 977 70
rect 917 16 977 38
rect 823 0 840 14
rect 872 0 889 14
rect 1016 0 1031 155
tri 1031 148 1044 161 nw
rect 1117 80 1132 270
rect 1117 0 1132 38
rect 1160 80 1175 270
tri 1240 234 1262 256 se
rect 1262 249 1277 270
tri 1262 234 1277 249 nw
rect 1596 249 1611 270
tri 1234 228 1240 234 se
rect 1240 228 1249 234
rect 1234 212 1249 228
tri 1249 221 1262 234 nw
rect 1403 226 1420 240
rect 1452 226 1469 240
tri 1596 234 1611 249 ne
tri 1611 234 1633 256 sw
rect 1234 176 1249 184
rect 1315 212 1375 226
rect 1330 202 1375 212
rect 1330 184 1358 202
tri 1234 161 1249 176 ne
tri 1249 161 1271 183 sw
rect 1315 174 1358 184
rect 1373 198 1375 202
rect 1497 212 1557 226
tri 1611 221 1624 234 ne
rect 1624 228 1633 234
tri 1633 228 1639 234 sw
rect 1497 202 1542 212
rect 1373 174 1447 198
rect 1315 170 1447 174
tri 1447 170 1475 198 sw
rect 1497 188 1499 202
tri 1497 186 1499 188 ne
rect 1511 184 1542 202
rect 1511 174 1557 184
rect 1624 213 1639 228
tri 1249 149 1261 161 ne
rect 1261 156 1271 161
tri 1271 156 1276 161 sw
rect 1160 0 1175 38
rect 1261 0 1276 156
rect 1315 114 1343 170
tri 1435 152 1453 170 ne
rect 1453 150 1475 170
tri 1475 150 1495 170 sw
tri 1511 156 1529 174 ne
rect 1334 80 1343 114
rect 1377 141 1419 142
rect 1377 107 1382 141
rect 1412 107 1419 141
rect 1377 98 1419 107
rect 1453 141 1495 150
rect 1453 107 1460 141
rect 1490 107 1495 141
rect 1453 102 1495 107
rect 1529 114 1557 174
tri 1602 161 1624 183 se
rect 1624 176 1639 184
tri 1624 161 1639 176 nw
tri 1596 155 1602 161 se
rect 1602 155 1611 161
rect 1315 70 1343 80
tri 1343 70 1367 94 sw
rect 1315 38 1357 70
tri 1374 62 1375 63 sw
rect 1374 38 1375 62
tri 1377 61 1414 98 ne
rect 1414 70 1419 98
tri 1419 70 1445 96 sw
rect 1529 80 1538 114
rect 1529 70 1557 80
rect 1414 61 1498 70
tri 1414 42 1433 61 ne
rect 1433 42 1498 61
rect 1315 16 1375 38
rect 1497 38 1498 42
rect 1515 38 1557 70
rect 1497 16 1557 38
rect 1403 0 1420 14
rect 1452 0 1469 14
rect 1596 0 1611 155
tri 1611 148 1624 161 nw
rect 1697 80 1712 270
rect 1697 0 1712 38
rect 1740 80 1755 270
tri 1820 234 1842 256 se
rect 1842 249 1857 270
tri 1842 234 1857 249 nw
rect 2176 249 2191 270
tri 1814 228 1820 234 se
rect 1820 228 1829 234
rect 1814 212 1829 228
tri 1829 221 1842 234 nw
rect 1983 226 2000 240
rect 2032 226 2049 240
tri 2176 234 2191 249 ne
tri 2191 234 2213 256 sw
rect 1814 176 1829 184
rect 1895 212 1955 226
rect 1910 202 1955 212
rect 1910 184 1938 202
tri 1814 161 1829 176 ne
tri 1829 161 1851 183 sw
rect 1895 174 1938 184
rect 1953 198 1955 202
rect 2077 212 2137 226
tri 2191 221 2204 234 ne
rect 2204 228 2213 234
tri 2213 228 2219 234 sw
rect 2077 202 2122 212
rect 1953 174 2027 198
rect 1895 170 2027 174
tri 2027 170 2055 198 sw
rect 2077 188 2079 202
tri 2077 186 2079 188 ne
rect 2091 184 2122 202
rect 2091 174 2137 184
rect 2204 213 2219 228
tri 1829 149 1841 161 ne
rect 1841 156 1851 161
tri 1851 156 1856 161 sw
rect 1740 0 1755 38
rect 1841 0 1856 156
rect 1895 114 1923 170
tri 2015 152 2033 170 ne
rect 2033 150 2055 170
tri 2055 150 2075 170 sw
tri 2091 156 2109 174 ne
rect 1914 80 1923 114
rect 1957 141 1999 142
rect 1957 107 1962 141
rect 1992 107 1999 141
rect 1957 98 1999 107
rect 2033 141 2075 150
rect 2033 107 2040 141
rect 2070 107 2075 141
rect 2033 102 2075 107
rect 2109 114 2137 174
tri 2182 161 2204 183 se
rect 2204 176 2219 184
tri 2204 161 2219 176 nw
tri 2176 155 2182 161 se
rect 2182 155 2191 161
rect 1895 70 1923 80
tri 1923 70 1947 94 sw
rect 1895 38 1937 70
tri 1954 62 1955 63 sw
rect 1954 38 1955 62
tri 1957 61 1994 98 ne
rect 1994 70 1999 98
tri 1999 70 2025 96 sw
rect 2109 80 2118 114
rect 2109 70 2137 80
rect 1994 61 2078 70
tri 1994 42 2013 61 ne
rect 2013 42 2078 61
rect 1895 16 1955 38
rect 2077 38 2078 42
rect 2095 38 2137 70
rect 2077 16 2137 38
rect 1983 0 2000 14
rect 2032 0 2049 14
rect 2176 0 2191 155
tri 2191 148 2204 161 nw
rect 2277 80 2292 270
rect 2277 0 2292 38
rect 2320 80 2335 270
tri 2400 234 2422 256 se
rect 2422 249 2437 270
tri 2422 234 2437 249 nw
rect 2756 249 2771 270
tri 2394 228 2400 234 se
rect 2400 228 2409 234
rect 2394 212 2409 228
tri 2409 221 2422 234 nw
rect 2563 226 2580 240
rect 2612 226 2629 240
tri 2756 234 2771 249 ne
tri 2771 234 2793 256 sw
rect 2394 176 2409 184
rect 2475 212 2535 226
rect 2490 202 2535 212
rect 2490 184 2518 202
tri 2394 161 2409 176 ne
tri 2409 161 2431 183 sw
rect 2475 174 2518 184
rect 2533 198 2535 202
rect 2657 212 2717 226
tri 2771 221 2784 234 ne
rect 2784 228 2793 234
tri 2793 228 2799 234 sw
rect 2657 202 2702 212
rect 2533 174 2607 198
rect 2475 170 2607 174
tri 2607 170 2635 198 sw
rect 2657 188 2659 202
tri 2657 186 2659 188 ne
rect 2671 184 2702 202
rect 2671 174 2717 184
rect 2784 213 2799 228
tri 2409 149 2421 161 ne
rect 2421 156 2431 161
tri 2431 156 2436 161 sw
rect 2320 0 2335 38
rect 2421 0 2436 156
rect 2475 114 2503 170
tri 2595 152 2613 170 ne
rect 2613 150 2635 170
tri 2635 150 2655 170 sw
tri 2671 156 2689 174 ne
rect 2494 80 2503 114
rect 2537 141 2579 142
rect 2537 107 2542 141
rect 2572 107 2579 141
rect 2537 98 2579 107
rect 2613 141 2655 150
rect 2613 107 2620 141
rect 2650 107 2655 141
rect 2613 102 2655 107
rect 2689 114 2717 174
tri 2762 161 2784 183 se
rect 2784 176 2799 184
tri 2784 161 2799 176 nw
tri 2756 155 2762 161 se
rect 2762 155 2771 161
rect 2475 70 2503 80
tri 2503 70 2527 94 sw
rect 2475 38 2517 70
tri 2534 62 2535 63 sw
rect 2534 38 2535 62
tri 2537 61 2574 98 ne
rect 2574 70 2579 98
tri 2579 70 2605 96 sw
rect 2689 80 2698 114
rect 2689 70 2717 80
rect 2574 61 2658 70
tri 2574 42 2593 61 ne
rect 2593 42 2658 61
rect 2475 16 2535 38
rect 2657 38 2658 42
rect 2675 38 2717 70
rect 2657 16 2717 38
rect 2563 0 2580 14
rect 2612 0 2629 14
rect 2756 0 2771 155
tri 2771 148 2784 161 nw
rect 2857 80 2872 270
rect 2857 0 2872 38
rect 2900 80 2915 270
tri 2980 234 3002 256 se
rect 3002 249 3017 270
tri 3002 234 3017 249 nw
rect 3336 249 3351 270
tri 2974 228 2980 234 se
rect 2980 228 2989 234
rect 2974 212 2989 228
tri 2989 221 3002 234 nw
rect 3143 226 3160 240
rect 3192 226 3209 240
tri 3336 234 3351 249 ne
tri 3351 234 3373 256 sw
rect 2974 176 2989 184
rect 3055 212 3115 226
rect 3070 202 3115 212
rect 3070 184 3098 202
tri 2974 161 2989 176 ne
tri 2989 161 3011 183 sw
rect 3055 174 3098 184
rect 3113 198 3115 202
rect 3237 212 3297 226
tri 3351 221 3364 234 ne
rect 3364 228 3373 234
tri 3373 228 3379 234 sw
rect 3237 202 3282 212
rect 3113 174 3187 198
rect 3055 170 3187 174
tri 3187 170 3215 198 sw
rect 3237 188 3239 202
tri 3237 186 3239 188 ne
rect 3251 184 3282 202
rect 3251 174 3297 184
rect 3364 213 3379 228
tri 2989 149 3001 161 ne
rect 3001 156 3011 161
tri 3011 156 3016 161 sw
rect 2900 0 2915 38
rect 3001 0 3016 156
rect 3055 114 3083 170
tri 3175 152 3193 170 ne
rect 3193 150 3215 170
tri 3215 150 3235 170 sw
tri 3251 156 3269 174 ne
rect 3074 80 3083 114
rect 3117 141 3159 142
rect 3117 107 3122 141
rect 3152 107 3159 141
rect 3117 98 3159 107
rect 3193 141 3235 150
rect 3193 107 3200 141
rect 3230 107 3235 141
rect 3193 102 3235 107
rect 3269 114 3297 174
tri 3342 161 3364 183 se
rect 3364 176 3379 184
tri 3364 161 3379 176 nw
tri 3336 155 3342 161 se
rect 3342 155 3351 161
rect 3055 70 3083 80
tri 3083 70 3107 94 sw
rect 3055 38 3097 70
tri 3114 62 3115 63 sw
rect 3114 38 3115 62
tri 3117 61 3154 98 ne
rect 3154 70 3159 98
tri 3159 70 3185 96 sw
rect 3269 80 3278 114
rect 3269 70 3297 80
rect 3154 61 3238 70
tri 3154 42 3173 61 ne
rect 3173 42 3238 61
rect 3055 16 3115 38
rect 3237 38 3238 42
rect 3255 38 3297 70
rect 3237 16 3297 38
rect 3143 0 3160 14
rect 3192 0 3209 14
rect 3336 0 3351 155
tri 3351 148 3364 161 nw
rect 3437 80 3452 270
rect 3437 0 3452 38
rect 3480 80 3495 270
tri 3560 234 3582 256 se
rect 3582 249 3597 270
tri 3582 234 3597 249 nw
rect 3916 249 3931 270
tri 3554 228 3560 234 se
rect 3560 228 3569 234
rect 3554 212 3569 228
tri 3569 221 3582 234 nw
rect 3723 226 3740 240
rect 3772 226 3789 240
tri 3916 234 3931 249 ne
tri 3931 234 3953 256 sw
rect 3554 176 3569 184
rect 3635 212 3695 226
rect 3650 202 3695 212
rect 3650 184 3678 202
tri 3554 161 3569 176 ne
tri 3569 161 3591 183 sw
rect 3635 174 3678 184
rect 3693 198 3695 202
rect 3817 212 3877 226
tri 3931 221 3944 234 ne
rect 3944 228 3953 234
tri 3953 228 3959 234 sw
rect 3817 202 3862 212
rect 3693 174 3767 198
rect 3635 170 3767 174
tri 3767 170 3795 198 sw
rect 3817 188 3819 202
tri 3817 186 3819 188 ne
rect 3831 184 3862 202
rect 3831 174 3877 184
rect 3944 213 3959 228
tri 3569 149 3581 161 ne
rect 3581 156 3591 161
tri 3591 156 3596 161 sw
rect 3480 0 3495 38
rect 3581 0 3596 156
rect 3635 114 3663 170
tri 3755 152 3773 170 ne
rect 3773 150 3795 170
tri 3795 150 3815 170 sw
tri 3831 156 3849 174 ne
rect 3654 80 3663 114
rect 3697 141 3739 142
rect 3697 107 3702 141
rect 3732 107 3739 141
rect 3697 98 3739 107
rect 3773 141 3815 150
rect 3773 107 3780 141
rect 3810 107 3815 141
rect 3773 102 3815 107
rect 3849 114 3877 174
tri 3922 161 3944 183 se
rect 3944 176 3959 184
tri 3944 161 3959 176 nw
tri 3916 155 3922 161 se
rect 3922 155 3931 161
rect 3635 70 3663 80
tri 3663 70 3687 94 sw
rect 3635 38 3677 70
tri 3694 62 3695 63 sw
rect 3694 38 3695 62
tri 3697 61 3734 98 ne
rect 3734 70 3739 98
tri 3739 70 3765 96 sw
rect 3849 80 3858 114
rect 3849 70 3877 80
rect 3734 61 3818 70
tri 3734 42 3753 61 ne
rect 3753 42 3818 61
rect 3635 16 3695 38
rect 3817 38 3818 42
rect 3835 38 3877 70
rect 3817 16 3877 38
rect 3723 0 3740 14
rect 3772 0 3789 14
rect 3916 0 3931 155
tri 3931 148 3944 161 nw
rect 4017 80 4032 270
rect 4017 0 4032 38
rect 4060 80 4075 270
tri 4140 234 4162 256 se
rect 4162 249 4177 270
tri 4162 234 4177 249 nw
rect 4496 249 4511 270
tri 4134 228 4140 234 se
rect 4140 228 4149 234
rect 4134 212 4149 228
tri 4149 221 4162 234 nw
rect 4303 226 4320 240
rect 4352 226 4369 240
tri 4496 234 4511 249 ne
tri 4511 234 4533 256 sw
rect 4134 176 4149 184
rect 4215 212 4275 226
rect 4230 202 4275 212
rect 4230 184 4258 202
tri 4134 161 4149 176 ne
tri 4149 161 4171 183 sw
rect 4215 174 4258 184
rect 4273 198 4275 202
rect 4397 212 4457 226
tri 4511 221 4524 234 ne
rect 4524 228 4533 234
tri 4533 228 4539 234 sw
rect 4397 202 4442 212
rect 4273 174 4347 198
rect 4215 170 4347 174
tri 4347 170 4375 198 sw
rect 4397 188 4399 202
tri 4397 186 4399 188 ne
rect 4411 184 4442 202
rect 4411 174 4457 184
rect 4524 213 4539 228
tri 4149 149 4161 161 ne
rect 4161 156 4171 161
tri 4171 156 4176 161 sw
rect 4060 0 4075 38
rect 4161 0 4176 156
rect 4215 114 4243 170
tri 4335 152 4353 170 ne
rect 4353 150 4375 170
tri 4375 150 4395 170 sw
tri 4411 156 4429 174 ne
rect 4234 80 4243 114
rect 4277 141 4319 142
rect 4277 107 4282 141
rect 4312 107 4319 141
rect 4277 98 4319 107
rect 4353 141 4395 150
rect 4353 107 4360 141
rect 4390 107 4395 141
rect 4353 102 4395 107
rect 4429 114 4457 174
tri 4502 161 4524 183 se
rect 4524 176 4539 184
tri 4524 161 4539 176 nw
tri 4496 155 4502 161 se
rect 4502 155 4511 161
rect 4215 70 4243 80
tri 4243 70 4267 94 sw
rect 4215 38 4257 70
tri 4274 62 4275 63 sw
rect 4274 38 4275 62
tri 4277 61 4314 98 ne
rect 4314 70 4319 98
tri 4319 70 4345 96 sw
rect 4429 80 4438 114
rect 4429 70 4457 80
rect 4314 61 4398 70
tri 4314 42 4333 61 ne
rect 4333 42 4398 61
rect 4215 16 4275 38
rect 4397 38 4398 42
rect 4415 38 4457 70
rect 4397 16 4457 38
rect 4303 0 4320 14
rect 4352 0 4369 14
rect 4496 0 4511 155
tri 4511 148 4524 161 nw
rect 4597 80 4612 270
rect 4597 0 4612 38
<< viali >>
rect 260 226 292 240
rect 43 102 73 136
rect 260 0 292 14
rect 479 102 509 136
rect 840 226 872 240
rect 623 102 653 136
rect 840 0 872 14
rect 1059 102 1089 136
rect 1420 226 1452 240
rect 1203 102 1233 136
rect 1420 0 1452 14
rect 1639 102 1669 136
rect 2000 226 2032 240
rect 1783 102 1813 136
rect 2000 0 2032 14
rect 2219 102 2249 136
rect 2580 226 2612 240
rect 2363 102 2393 136
rect 2580 0 2612 14
rect 2799 102 2829 136
rect 3160 226 3192 240
rect 2943 102 2973 136
rect 3160 0 3192 14
rect 3379 102 3409 136
rect 3740 226 3772 240
rect 3523 102 3553 136
rect 3740 0 3772 14
rect 3959 102 3989 136
rect 4320 226 4352 240
rect 4103 102 4133 136
rect 4320 0 4352 14
rect 4539 102 4569 136
<< metal1 >>
rect 0 226 260 240
rect 292 226 840 240
rect 872 226 1420 240
rect 1452 226 2000 240
rect 2032 226 2580 240
rect 2612 226 3160 240
rect 3192 226 3740 240
rect 3772 226 4320 240
rect 4352 226 4612 240
rect 0 102 43 136
rect 73 102 479 136
rect 509 102 623 136
rect 653 102 1059 136
rect 1089 102 1203 136
rect 1233 102 1639 136
rect 1669 102 1783 136
rect 1813 102 2219 136
rect 2249 102 2363 136
rect 2393 102 2799 136
rect 2829 102 2943 136
rect 2973 102 3379 136
rect 3409 102 3523 136
rect 3553 102 3959 136
rect 3989 102 4103 136
rect 4133 102 4539 136
rect 0 0 260 14
rect 292 0 840 14
rect 872 0 1420 14
rect 1452 0 2000 14
rect 2032 0 2580 14
rect 2612 0 3160 14
rect 3192 0 3740 14
rect 3772 0 4320 14
rect 4352 0 4612 14
<< labels >>
rlabel poly 0 240 30 270 1 WWL
port 17 ew signal input
rlabel metal1 0 102 15 136 1 RWL
port 18 ew signal input
rlabel corelocali 74 184 89 212 1 WBLb_0
port 19 ns signal input
rlabel corelocali 464 184 479 213 1 WBL_0
port 20 ns signal input
rlabel corelocali 0 38 15 80 1 RBL1_0
port 1 ns signal output
rlabel corelocali 537 38 552 80 1 RBL0_0
port 2 ns signal output
rlabel corelocali 654 184 669 212 1 WBLb_1
port 21 ns signal input
rlabel corelocali 1044 184 1059 213 1 WBL_1
port 22 ns signal input
rlabel corelocali 580 38 595 80 1 RBL1_1
port 3 ns signal output
rlabel corelocali 1117 38 1132 80 1 RBL0_1
port 4 ns signal output
rlabel corelocali 1234 184 1249 212 1 WBLb_2
port 23 ns signal input
rlabel corelocali 1624 184 1639 213 1 WBL_2
port 24 ns signal input
rlabel corelocali 1160 38 1175 80 1 RBL1_2
port 5 ns signal output
rlabel corelocali 1697 38 1712 80 1 RBL0_2
port 6 ns signal output
rlabel corelocali 1814 184 1829 212 1 WBLb_3
port 25 ns signal input
rlabel corelocali 2204 184 2219 213 1 WBL_3
port 26 ns signal input
rlabel corelocali 1740 38 1755 80 1 RBL1_3
port 7 ns signal output
rlabel corelocali 2277 38 2292 80 1 RBL0_3
port 8 ns signal output
rlabel corelocali 2394 184 2409 212 1 WBLb_4
port 27 ns signal input
rlabel corelocali 2784 184 2799 213 1 WBL_4
port 28 ns signal input
rlabel corelocali 2320 38 2335 80 1 RBL1_4
port 8 ns signal output
rlabel corelocali 2857 38 2872 80 1 RBL0_4
port 10 ns signal output
rlabel corelocali 2974 184 2989 212 1 WBLb_5
port 29 ns signal input
rlabel corelocali 3364 184 3379 213 1 WBL_5
port 30 ns signal input
rlabel corelocali 2900 38 2915 80 1 RBL1_5
port 11 ns signal output
rlabel corelocali 3437 38 3452 80 1 RBL0_5
port 12 ns signal output
rlabel corelocali 3554 184 3569 212 1 WBLb_6
port 31 ns signal input
rlabel corelocali 3944 184 3959 213 1 WBL_6
port 32 ns signal input
rlabel corelocali 3480 38 3495 80 1 RBL1_6
port 13 ns signal output
rlabel corelocali 4017 38 4032 80 1 RBL0_6
port 14 ns signal output
rlabel corelocali 4134 184 4149 212 1 WBLb_7
port 33 ns signal input
rlabel corelocali 4524 184 4539 213 1 WBL_7
port 34 ns signal input
rlabel corelocali 4060 38 4075 80 1 RBL1_7
port 15 ns signal output
rlabel corelocali 4597 38 4612 80 1 RBL0_7
port 16 ns signal output
rlabel metal1 0 226 15 240 1 VDD
port 35 ns power bidirectional abutment
rlabel metal1 0 0 15 14 1 GND
port 36 ns ground bidirectional abutment
rlabel poly 0 240 552 270 1 10T_toy_magic_7/WWL
rlabel locali 479 102 509 136 1 10T_toy_magic_7/RWL
rlabel locali 43 102 73 136 1 10T_toy_magic_7/RWL
rlabel locali 464 184 479 213 1 10T_toy_magic_7/WBL
rlabel locali 74 184 89 212 1 10T_toy_magic_7/WBLb
rlabel locali 537 38 552 80 1 10T_toy_magic_7/RBL0
rlabel locali 0 38 15 80 1 10T_toy_magic_7/RBL1
rlabel metal1 260 226 292 240 1 10T_toy_magic_7/VDD
rlabel metal1 260 0 292 14 7 10T_toy_magic_7/GND
rlabel polycont 222 107 252 141 1 10T_toy_magic_7/junc0
rlabel polycont 300 107 330 141 1 10T_toy_magic_7/junc1
rlabel ndiff 73 38 129 66 1 10T_toy_magic_7/RWL1_junc
rlabel ndiff 423 38 479 66 1 10T_toy_magic_7/RWL0_junc
rlabel poly 580 240 1132 270 1 10T_toy_magic_6/WWL
rlabel locali 1059 102 1089 136 1 10T_toy_magic_6/RWL
rlabel locali 623 102 653 136 1 10T_toy_magic_6/RWL
rlabel locali 1044 184 1059 213 1 10T_toy_magic_6/WBL
rlabel locali 654 184 669 212 1 10T_toy_magic_6/WBLb
rlabel locali 1117 38 1132 80 1 10T_toy_magic_6/RBL0
rlabel locali 580 38 595 80 1 10T_toy_magic_6/RBL1
rlabel metal1 840 226 872 240 1 10T_toy_magic_6/VDD
rlabel metal1 840 0 872 14 7 10T_toy_magic_6/GND
rlabel polycont 802 107 832 141 1 10T_toy_magic_6/junc0
rlabel polycont 880 107 910 141 1 10T_toy_magic_6/junc1
rlabel ndiff 653 38 709 66 1 10T_toy_magic_6/RWL1_junc
rlabel ndiff 1003 38 1059 66 1 10T_toy_magic_6/RWL0_junc
rlabel poly 1160 240 1712 270 1 10T_toy_magic_5/WWL
rlabel locali 1639 102 1669 136 1 10T_toy_magic_5/RWL
rlabel locali 1203 102 1233 136 1 10T_toy_magic_5/RWL
rlabel locali 1624 184 1639 213 1 10T_toy_magic_5/WBL
rlabel locali 1234 184 1249 212 1 10T_toy_magic_5/WBLb
rlabel locali 1697 38 1712 80 1 10T_toy_magic_5/RBL0
rlabel locali 1160 38 1175 80 1 10T_toy_magic_5/RBL1
rlabel metal1 1420 226 1452 240 1 10T_toy_magic_5/VDD
rlabel metal1 1420 0 1452 14 7 10T_toy_magic_5/GND
rlabel polycont 1382 107 1412 141 1 10T_toy_magic_5/junc0
rlabel polycont 1460 107 1490 141 1 10T_toy_magic_5/junc1
rlabel ndiff 1233 38 1289 66 1 10T_toy_magic_5/RWL1_junc
rlabel ndiff 1583 38 1639 66 1 10T_toy_magic_5/RWL0_junc
rlabel poly 1740 240 2292 270 1 10T_toy_magic_4/WWL
rlabel locali 2219 102 2249 136 1 10T_toy_magic_4/RWL
rlabel locali 1783 102 1813 136 1 10T_toy_magic_4/RWL
rlabel locali 2204 184 2219 213 1 10T_toy_magic_4/WBL
rlabel locali 1814 184 1829 212 1 10T_toy_magic_4/WBLb
rlabel locali 2277 38 2292 80 1 10T_toy_magic_4/RBL0
rlabel locali 1740 38 1755 80 1 10T_toy_magic_4/RBL1
rlabel metal1 2000 226 2032 240 1 10T_toy_magic_4/VDD
rlabel metal1 2000 0 2032 14 7 10T_toy_magic_4/GND
rlabel polycont 1962 107 1992 141 1 10T_toy_magic_4/junc0
rlabel polycont 2040 107 2070 141 1 10T_toy_magic_4/junc1
rlabel ndiff 1813 38 1869 66 1 10T_toy_magic_4/RWL1_junc
rlabel ndiff 2163 38 2219 66 1 10T_toy_magic_4/RWL0_junc
rlabel poly 2320 240 2872 270 1 10T_toy_magic_3/WWL
rlabel locali 2799 102 2829 136 1 10T_toy_magic_3/RWL
rlabel locali 2363 102 2393 136 1 10T_toy_magic_3/RWL
rlabel locali 2784 184 2799 213 1 10T_toy_magic_3/WBL
rlabel locali 2394 184 2409 212 1 10T_toy_magic_3/WBLb
rlabel locali 2857 38 2872 80 1 10T_toy_magic_3/RBL0
rlabel locali 2320 38 2335 80 1 10T_toy_magic_3/RBL1
rlabel metal1 2580 226 2612 240 1 10T_toy_magic_3/VDD
rlabel metal1 2580 0 2612 14 7 10T_toy_magic_3/GND
rlabel polycont 2542 107 2572 141 1 10T_toy_magic_3/junc0
rlabel polycont 2620 107 2650 141 1 10T_toy_magic_3/junc1
rlabel ndiff 2393 38 2449 66 1 10T_toy_magic_3/RWL1_junc
rlabel ndiff 2743 38 2799 66 1 10T_toy_magic_3/RWL0_junc
rlabel poly 2900 240 3452 270 1 10T_toy_magic_2/WWL
rlabel locali 3379 102 3409 136 1 10T_toy_magic_2/RWL
rlabel locali 2943 102 2973 136 1 10T_toy_magic_2/RWL
rlabel locali 3364 184 3379 213 1 10T_toy_magic_2/WBL
rlabel locali 2974 184 2989 212 1 10T_toy_magic_2/WBLb
rlabel locali 3437 38 3452 80 1 10T_toy_magic_2/RBL0
rlabel locali 2900 38 2915 80 1 10T_toy_magic_2/RBL1
rlabel metal1 3160 226 3192 240 1 10T_toy_magic_2/VDD
rlabel metal1 3160 0 3192 14 7 10T_toy_magic_2/GND
rlabel polycont 3122 107 3152 141 1 10T_toy_magic_2/junc0
rlabel polycont 3200 107 3230 141 1 10T_toy_magic_2/junc1
rlabel ndiff 2973 38 3029 66 1 10T_toy_magic_2/RWL1_junc
rlabel ndiff 3323 38 3379 66 1 10T_toy_magic_2/RWL0_junc
rlabel poly 4060 240 4612 270 1 10T_toy_magic_1/WWL
rlabel locali 4539 102 4569 136 1 10T_toy_magic_1/RWL
rlabel locali 4103 102 4133 136 1 10T_toy_magic_1/RWL
rlabel locali 4524 184 4539 213 1 10T_toy_magic_1/WBL
rlabel locali 4134 184 4149 212 1 10T_toy_magic_1/WBLb
rlabel locali 4597 38 4612 80 1 10T_toy_magic_1/RBL0
rlabel locali 4060 38 4075 80 1 10T_toy_magic_1/RBL1
rlabel metal1 4320 226 4352 240 1 10T_toy_magic_1/VDD
rlabel metal1 4320 0 4352 14 7 10T_toy_magic_1/GND
rlabel polycont 4282 107 4312 141 1 10T_toy_magic_1/junc0
rlabel polycont 4360 107 4390 141 1 10T_toy_magic_1/junc1
rlabel ndiff 4133 38 4189 66 1 10T_toy_magic_1/RWL1_junc
rlabel ndiff 4483 38 4539 66 1 10T_toy_magic_1/RWL0_junc
rlabel poly 3480 240 4032 270 1 10T_toy_magic_0/WWL
rlabel locali 3959 102 3989 136 1 10T_toy_magic_0/RWL
rlabel locali 3523 102 3553 136 1 10T_toy_magic_0/RWL
rlabel locali 3944 184 3959 213 1 10T_toy_magic_0/WBL
rlabel locali 3554 184 3569 212 1 10T_toy_magic_0/WBLb
rlabel locali 4017 38 4032 80 1 10T_toy_magic_0/RBL0
rlabel locali 3480 38 3495 80 1 10T_toy_magic_0/RBL1
rlabel metal1 3740 226 3772 240 1 10T_toy_magic_0/VDD
rlabel metal1 3740 0 3772 14 7 10T_toy_magic_0/GND
rlabel polycont 3702 107 3732 141 1 10T_toy_magic_0/junc0
rlabel polycont 3780 107 3810 141 1 10T_toy_magic_0/junc1
rlabel ndiff 3553 38 3609 66 1 10T_toy_magic_0/RWL1_junc
rlabel ndiff 3903 38 3959 66 1 10T_toy_magic_0/RWL0_junc
<< end >>
