* HSPICE file created from 10T_32x32_magic.ext - technology: sky130A

.subckt x10T_toy_magic WWL RWL0 RWL1 WBL WBLb RBL0 RBL1 VDD GND
M1000 VDD junc0 junc1 VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15
M1001 WBL WWL junc0 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15
M1002 junc1 WWL WBLb GND sky130_fd_pr__nfet_01v8 w=1 l=0.15
M1003 GND junc0 junc1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15
M1004 RWL0_junc junc0 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15
M1005 RBL0 RWL0 RWL0_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15
M1006 GND junc1 RWL1_junc GND sky130_fd_pr__nfet_01v8 w=1 l=0.15
M1007 RWL1_junc RWL1 RBL1 GND sky130_fd_pr__nfet_01v8 w=1 l=0.15
M1008 junc0 junc1 GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.15
M1009 junc0 junc1 VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.15
.ends

.subckt x10T_1x8_magic RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4
+ RBL1_5 RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL RWL WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x0/RBL0
+ x5/WBLb x5/RBL1 x4/WBLb x7/WBL x5/RBL0 x4/RBL1 x1/WBLb x4/RBL0 x6/WBL x1/RBL1 x1/RBL0
+ x7/WBLb x3/WBL x5/WWL x7/RBL1 x6/WBLb x7/RBL0 x2/WBL x6/RBL1 x6/RBL0 x0/WBL x5/VDD
+ x3/WBLb x5/WBL x3/RBL1 x2/WBLb x4/WBL x3/RBL0 x2/RBL1 x0/WBLb x2/RBL0 x1/WBL x0/RBL1
+ VSUBS
X10T_toy_magic_0 x5/WWL RWL RWL x0/WBL x0/WBLb x0/RBL0 x0/RBL1 x5/VDD VSUBS x10T_toy_magic
X10T_toy_magic_1 x5/WWL RWL RWL x1/WBL x1/WBLb x1/RBL0 x1/RBL1 x5/VDD VSUBS x10T_toy_magic
X10T_toy_magic_3 x5/WWL RWL RWL x2/WBL x2/WBLb x2/RBL0 x2/RBL1 x5/VDD VSUBS x10T_toy_magic
X10T_toy_magic_2 x5/WWL RWL RWL x6/WBL x6/WBLb x6/RBL0 x6/RBL1 x5/VDD VSUBS x10T_toy_magic
X10T_toy_magic_4 x5/WWL RWL RWL x4/WBL x4/WBLb x4/RBL0 x4/RBL1 x5/VDD VSUBS x10T_toy_magic
X10T_toy_magic_5 x5/WWL RWL RWL x7/WBL x7/WBLb x7/RBL0 x7/RBL1 x5/VDD VSUBS x10T_toy_magic
X10T_toy_magic_6 x5/WWL RWL RWL x3/WBL x3/WBLb x3/RBL0 x3/RBL1 x5/VDD VSUBS x10T_toy_magic
X10T_toy_magic_7 x5/WWL RWL RWL x5/WBL x5/WBLb x5/RBL0 x5/RBL1 x5/VDD VSUBS x10T_toy_magic
.ends

.subckt x10T_32x32_magic RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL0_3 RBL1_4
+ RBL0_4 RBL1_5 RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10
+ RBL0_10 RBL1_11 RBL0_11 RBL1_12 RBL0_12 RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15
+ RBL0_15 WWL_0 RWL_0 WWL_1 RWL_1 WWL_2 RWL_2 WWL_3 RWL_3 WWL_4 RWL_4 WWL_5 RWL_5
+ WWL_6 RWL_6 WWL_7 RWL_7 WWL_8 RWL_8 WWL_9 RWL_9 WWL_10 RWL_10 WWL_11 RWL_11 WWL_12
+ RWL_12 WWL_13 RWL_13 WWL_14 RWL_14 WWL_15 RWL_15 WWL_16 RWL_16 WWL_17 RWL_17 WWL_18
+ RWL_18 WWL_19 RWL_19 WWL_20 RWL_20 WWL_21 RWL_21 WWL_22 RWL_22 WWL_23 RWL_23 WWL_24
+ RWL_24 WWL_25 RWL_25 WWL_26 RWL_26 WWL_27 RWL_27 WWL_28 RWL_28 WWL_29 RWL_29 WWL_30
+ RWL_30 WWL_31 RWL_31 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL0_19
+ RBL1_20 RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 RBL1_24 RBL0_24
+ RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL0_27 RBL1_28 RBL0_28 RBL1_29 RBL0_29
+ RBL1_30 RBL0_30 RBL1_31 RBL0_31 WBL_0 WBLb_0 WBL_1 WBLb_1 WBL_2 WBLb_2 WBL_3 WBLb_19
+ WBL_4 WBLb_4 WBL_5 WBLb_5 WBL_22 WBLb_6 WBL_23 WBLb_7 WBL_24 WBLb_8 WBL_25 WBLb_9
+ WBL_26 WBLb_10 WBL_11 WBLb_11 WBL_12 WBLb_12 WBL_13 WBLb_13 WBL_14 WBLb_30 WBL_15
+ WBLb_31 VDD GND
X10T_1x8_magic_0 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_2 RWL_2 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND RBL0_6
+ x0/WBLb RBL1_0 x1/WBLb x2/WBL RBL0_0 RBL1_3 x3/WBLb RBL0_3 x4/WBL RBL1_7 RBL0_7
+ x2/WBLb x5/WBL x6/WWL RBL1_2 x4/WBLb RBL0_2 x7/WBL RBL1_5 RBL0_5 x8/WBL x6/VDD x5/WBLb
+ x0/WBL RBL1_1 x7/WBLb x1/WBL RBL0_1 RBL1_4 x8/WBLb RBL0_4 x3/WBL RBL1_6 VSUBS x10T_1x8_magic
X10T_1x8_magic_1 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_3 RWL_3 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x9/RBL0
+ x10/WBLb x10/RBL1 x11/WBLb x12/WBL x10/RBL0 x11/RBL1 x13/WBLb x11/RBL0 x14/WBL x13/RBL1
+ x13/RBL0 x12/WBLb x15/WBL x16/WWL x12/RBL1 x14/WBLb x12/RBL0 x17/WBL x14/RBL1 x14/RBL0
+ x9/WBL x16/VDD x15/WBLb x10/WBL x15/RBL1 x17/WBLb x11/WBL x15/RBL0 x17/RBL1 x9/WBLb
+ x17/RBL0 x13/WBL x9/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_2 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_0 RWL_0 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x18/RBL0
+ x19/WBLb x19/RBL1 x20/WBLb x21/WBL x19/RBL0 x20/RBL1 x22/WBLb x20/RBL0 x23/WBL x22/RBL1
+ x22/RBL0 x21/WBLb x24/WBL x25/WWL x21/RBL1 x23/WBLb x21/RBL0 x26/WBL x23/RBL1 x23/RBL0
+ x18/WBL x25/VDD x24/WBLb x19/WBL x24/RBL1 x26/WBLb x20/WBL x24/RBL0 x26/RBL1 x18/WBLb
+ x26/RBL0 x22/WBL x18/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_3 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_1 RWL_1 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x27/RBL0
+ x28/WBLb x28/RBL1 x29/WBLb x30/WBL x28/RBL0 x29/RBL1 x31/WBLb x29/RBL0 x32/WBL x31/RBL1
+ x31/RBL0 x30/WBLb x33/WBL x34/WWL x30/RBL1 x32/WBLb x30/RBL0 x35/WBL x32/RBL1 x32/RBL0
+ x27/WBL x34/VDD x33/WBLb x28/WBL x33/RBL1 x35/WBLb x29/WBL x33/RBL0 x35/RBL1 x27/WBLb
+ x35/RBL0 x31/WBL x27/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_4 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_7 RWL_7 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND RBL0_6
+ x36/WBLb RBL1_0 x37/WBLb x38/WBL RBL0_0 RBL1_3 x39/WBLb RBL0_3 x40/WBL RBL1_7 RBL0_7
+ x38/WBLb x41/WBL x42/WWL RBL1_2 x40/WBLb RBL0_2 x43/WBL RBL1_5 RBL0_5 x44/WBL x42/VDD
+ x41/WBLb x36/WBL RBL1_1 x43/WBLb x37/WBL RBL0_1 RBL1_4 x44/WBLb RBL0_4 x39/WBL RBL1_6
+ VSUBS x10T_1x8_magic
X10T_1x8_magic_5 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_6 RWL_6 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x45/RBL0
+ x46/WBLb x46/RBL1 x47/WBLb x48/WBL x46/RBL0 x47/RBL1 x49/WBLb x47/RBL0 x50/WBL x49/RBL1
+ x49/RBL0 x48/WBLb x51/WBL x52/WWL x48/RBL1 x50/WBLb x48/RBL0 x53/WBL x50/RBL1 x50/RBL0
+ x45/WBL x52/VDD x51/WBLb x46/WBL x51/RBL1 x53/WBLb x47/WBL x51/RBL0 x53/RBL1 x45/WBLb
+ x53/RBL0 x49/WBL x45/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_6 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_4 RWL_4 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x54/RBL0
+ WBLb_0 x55/RBL1 WBLb_3 WBL_2 x55/RBL0 x56/RBL1 WBLb_7 x56/RBL0 WBL_5 x57/RBL1 x57/RBL0
+ WBLb_2 WBL_1 x58/WWL x59/RBL1 WBLb_5 x59/RBL0 WBL_4 x60/RBL1 x60/RBL0 WBL_6 x58/VDD
+ WBLb_1 WBL_0 x61/RBL1 WBLb_4 WBL_3 x61/RBL0 x62/RBL1 WBLb_6 x62/RBL0 WBL_7 x54/RBL1
+ VSUBS x10T_1x8_magic
X10T_1x8_magic_7 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_5 RWL_5 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x63/RBL0
+ x64/WBLb x64/RBL1 x65/WBLb x66/WBL x64/RBL0 x65/RBL1 x67/WBLb x65/RBL0 x68/WBL x67/RBL1
+ x67/RBL0 x66/WBLb x69/WBL x70/WWL x66/RBL1 x68/WBLb x66/RBL0 x71/WBL x68/RBL1 x68/RBL0
+ x63/WBL x70/VDD x69/WBLb x64/WBL x69/RBL1 x71/WBLb x65/WBL x69/RBL0 x71/RBL1 x63/WBLb
+ x71/RBL0 x67/WBL x63/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_90 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x72/WWL RWL_17 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x72/VDD VSUBS x73/RBL0 WBLb_16 x74/RBL1 x75/WBLb x76/WBL x74/RBL0
+ x75/RBL1 x77/WBLb x75/RBL0 x78/WBL x77/RBL1 x77/RBL0 x76/WBLb x79/WBL x80/WWL x76/RBL1
+ x78/WBLb x76/RBL0 x81/WBL RBL1_21 x78/RBL0 x73/WBL x80/VDD x79/WBLb x74/WBL x79/RBL1
+ x81/WBLb x75/WBL x79/RBL0 x81/RBL1 x73/WBLb x81/RBL0 x77/WBL x73/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_8 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_14 RWL_14 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND RBL0_6
+ WBLb_0 RBL1_0 WBLb_3 WBL_2 RBL0_0 RBL1_3 WBLb_7 RBL0_3 WBL_5 RBL1_7 RBL0_7 WBLb_2
+ WBL_1 x82/WWL RBL1_2 WBLb_5 RBL0_2 WBL_4 RBL1_5 RBL0_5 WBL_6 x82/VDD WBLb_1 WBL_0
+ RBL1_1 WBLb_4 WBL_3 RBL0_1 RBL1_4 WBLb_6 RBL0_4 WBL_7 RBL1_6 VSUBS x10T_1x8_magic
X10T_1x8_magic_80 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x83/WWL RWL_23 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 VDD VSUBS RBL0_22 WBLb_16 RBL1_16 WBLb_19 WBL_18 RBL0_16 RBL1_19
+ WBLb_23 RBL0_19 WBL_21 RBL1_23 RBL0_23 WBLb_18 WBL_17 x84/WWL RBL1_18 WBLb_21 RBL0_18
+ WBL_20 RBL1_21 RBL0_21 WBL_22 VDD WBLb_17 WBL_16 RBL1_17 WBLb_20 WBL_19 RBL0_17
+ RBL1_20 WBLb_22 RBL0_20 WBL_23 RBL1_22 VSUBS x10T_1x8_magic
X10T_1x8_magic_91 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x85/WWL RWL_18 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x85/VDD VSUBS x86/RBL0 WBLb_16 x87/RBL1 x88/WBLb x89/WBL x87/RBL0
+ x88/RBL1 x90/WBLb x88/RBL0 x91/WBL x90/RBL1 x90/RBL0 x89/WBLb x92/WBL x93/WWL x89/RBL1
+ x91/WBLb x89/RBL0 x94/WBL RBL1_21 x91/RBL0 x86/WBL x93/VDD x92/WBLb x87/WBL x92/RBL1
+ x94/WBLb x88/WBL x92/RBL0 x94/RBL1 x86/WBLb x94/RBL0 x90/WBL x86/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_70 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x95/WWL RWL_28 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x95/VDD VSUBS RBL0_22 WBLb_16 RBL1_16 x96/WBLb x97/WBL RBL0_16
+ RBL1_19 x98/WBLb RBL0_19 x99/WBL RBL1_23 RBL0_23 x97/WBLb x100/WBL x101/WWL RBL1_18
+ x99/WBLb RBL0_18 x102/WBL RBL1_21 RBL0_21 x103/WBL x101/VDD x100/WBLb x104/WBL RBL1_17
+ x102/WBLb x96/WBL RBL0_17 RBL1_20 x103/WBLb RBL0_20 x98/WBL RBL1_22 VSUBS x10T_1x8_magic
X10T_1x8_magic_81 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x84/WWL RWL_23 WBLb_24 WBL_24
+ WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29 WBLb_30
+ WBL_30 WBLb_31 WBL_31 VDD VSUBS RBL0_30 WBLb_24 RBL1_24 WBLb_27 WBL_26 RBL0_24 RBL1_27
+ WBLb_31 RBL0_27 WBL_29 RBL1_31 RBL0_31 WBLb_26 WBL_25 x105/WWL RBL1_26 WBLb_29 RBL0_26
+ WBL_28 RBL1_29 RBL0_29 WBL_30 VDD WBLb_25 WBL_24 RBL1_25 WBLb_28 WBL_27 RBL0_25
+ RBL1_28 WBLb_30 RBL0_28 WBL_31 RBL1_30 VSUBS x10T_1x8_magic
X10T_1x8_magic_92 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x80/WWL RWL_17 WBLb_24 WBL_24
+ WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29 WBLb_30
+ WBL_30 WBLb_31 WBL_31 x80/VDD VSUBS x106/RBL0 x107/WBLb x107/RBL1 x108/WBLb x109/WBL
+ x107/RBL0 x108/RBL1 x110/WBLb x108/RBL0 x111/WBL x110/RBL1 x110/RBL0 x109/WBLb x112/WBL
+ x107/WWL x109/RBL1 x111/WBLb x109/RBL0 x113/WBL x111/RBL1 x111/RBL0 x106/WBL x107/VDD
+ x112/WBLb x107/WBL x112/RBL1 x113/WBLb x108/WBL x112/RBL0 x113/RBL1 x106/WBLb x113/RBL0
+ x110/WBL x106/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_9 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_15 RWL_15 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x114/RBL0
+ x115/WBLb x115/RBL1 x116/WBLb x117/WBL x115/RBL0 x116/RBL1 x118/WBLb x116/RBL0 x119/WBL
+ x118/RBL1 x118/RBL0 x117/WBLb x120/WBL x121/WWL x117/RBL1 x119/WBLb x117/RBL0 x122/WBL
+ x119/RBL1 x119/RBL0 x114/WBL x121/VDD x120/WBLb x115/WBL x120/RBL1 x122/WBLb x116/WBL
+ x120/RBL0 x122/RBL1 x114/WBLb x122/RBL0 x118/WBL x114/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_60 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x16/WWL x16/RWL WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x16/VDD VSUBS x123/RBL0 x124/WBLb x124/RBL1 x125/WBLb x126/WBL x124/RBL0
+ x125/RBL1 x127/WBLb x125/RBL0 x128/WBL x127/RBL1 x127/RBL0 x126/WBLb x129/WBL x130/WWL
+ x126/RBL1 x128/WBLb x126/RBL0 x131/WBL x128/RBL1 x128/RBL0 x123/WBL x130/VDD x129/WBLb
+ x124/WBL x129/RBL1 x131/WBLb x125/WBL x129/RBL0 x131/RBL1 x123/WBLb x131/RBL0 x127/WBL
+ x123/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_71 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x101/WWL RWL_28 WBLb_24
+ WBL_24 WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29
+ WBLb_30 WBL_30 WBLb_31 WBL_31 x101/VDD VSUBS RBL0_30 x132/WBLb RBL1_24 x133/WBLb
+ x134/WBL RBL0_24 RBL1_27 x135/WBLb RBL0_27 x136/WBL RBL1_31 RBL0_31 x134/WBLb x137/WBL
+ x132/WWL RBL1_26 x136/WBLb RBL0_26 x138/WBL RBL1_29 RBL0_29 x139/WBL x132/VDD x137/WBLb
+ x132/WBL RBL1_25 x138/WBLb x133/WBL RBL0_25 RBL1_28 x139/WBLb RBL0_28 x135/WBL RBL1_30
+ VSUBS x10T_1x8_magic
X10T_1x8_magic_82 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x140/WWL RWL_22 WBLb_16
+ WBL_16 WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21
+ WBLb_22 WBL_22 WBLb_23 WBL_23 x140/VDD VSUBS x141/RBL0 WBLb_16 x142/RBL1 x143/WBLb
+ x144/WBL x142/RBL0 x143/RBL1 x145/WBLb x143/RBL0 x146/WBL x145/RBL1 x145/RBL0 x144/WBLb
+ x147/WBL x148/WWL x144/RBL1 x146/WBLb x144/RBL0 x149/WBL RBL1_21 x146/RBL0 x141/WBL
+ x148/VDD x147/WBLb x142/WBL x147/RBL1 x149/WBLb x143/WBL x147/RBL0 x149/RBL1 x141/WBLb
+ x149/RBL0 x145/WBL x141/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_93 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x93/WWL RWL_18 WBLb_24 WBL_24
+ WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29 WBLb_30
+ WBL_30 WBLb_31 WBL_31 x93/VDD VSUBS x150/RBL0 x151/WBLb x151/RBL1 x152/WBLb x153/WBL
+ x151/RBL0 x152/RBL1 x154/WBLb x152/RBL0 x155/WBL x154/RBL1 x154/RBL0 x153/WBLb x156/WBL
+ x151/WWL x153/RBL1 x155/WBLb x153/RBL0 x157/WBL x155/RBL1 x155/RBL0 x150/WBL x151/VDD
+ x156/WBLb x151/WBL x156/RBL1 x157/WBLb x152/WBL x156/RBL0 x157/RBL1 x150/WBLb x157/RBL0
+ x154/WBL x150/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_61 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x6/WWL RWL_2 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x6/VDD VSUBS RBL0_14 x158/WBLb RBL1_8 x159/WBLb x160/WBL RBL0_8 RBL1_11
+ x161/WBLb RBL0_11 x162/WBL RBL1_15 RBL0_15 x160/WBLb x163/WBL x164/WWL RBL1_10 x162/WBLb
+ RBL0_10 x165/WBL RBL1_13 RBL0_13 x166/WBL x164/VDD x163/WBLb x158/WBL RBL1_9 x165/WBLb
+ x159/WBL RBL0_9 RBL1_12 x166/WBLb RBL0_12 x161/WBL RBL1_14 VSUBS x10T_1x8_magic
X10T_1x8_magic_72 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x167/WWL RWL_27 WBLb_16
+ WBL_16 WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21
+ WBLb_22 WBL_22 WBLb_23 WBL_23 x167/VDD VSUBS x168/RBL0 WBLb_16 x169/RBL1 x170/WBLb
+ x171/WBL x169/RBL0 x170/RBL1 x172/WBLb x170/RBL0 x173/WBL x172/RBL1 x172/RBL0 x171/WBLb
+ x174/WBL x175/WWL x171/RBL1 x173/WBLb x171/RBL0 x176/WBL RBL1_21 x173/RBL0 x168/WBL
+ x175/VDD x174/WBLb x169/WBL x174/RBL1 x176/WBLb x170/WBL x174/RBL0 x176/RBL1 x168/WBLb
+ x176/RBL0 x172/WBL x168/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_83 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x148/WWL RWL_22 WBLb_24
+ WBL_24 WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29
+ WBLb_30 WBL_30 WBLb_31 WBL_31 x148/VDD VSUBS x177/RBL0 x178/WBLb x178/RBL1 x179/WBLb
+ x180/WBL x178/RBL0 x179/RBL1 x181/WBLb x179/RBL0 x182/WBL x181/RBL1 x181/RBL0 x180/WBLb
+ x183/WBL x178/WWL x180/RBL1 x182/WBLb x180/RBL0 x184/WBL x182/RBL1 x182/RBL0 x177/WBL
+ x178/VDD x183/WBLb x178/WBL x183/RBL1 x184/WBLb x179/WBL x183/RBL0 x184/RBL1 x177/WBLb
+ x184/RBL0 x181/WBL x177/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_94 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x185/WWL RWL_16 WBLb_16
+ WBL_16 WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21
+ WBLb_22 WBL_22 WBLb_23 WBL_23 x185/VDD VSUBS x186/RBL0 WBLb_16 x187/RBL1 x188/WBLb
+ x189/WBL x187/RBL0 x188/RBL1 x190/WBLb x188/RBL0 x191/WBL x190/RBL1 x190/RBL0 x189/WBLb
+ x192/WBL x193/WWL x189/RBL1 x191/WBLb x189/RBL0 x194/WBL RBL1_21 x191/RBL0 x186/WBL
+ x193/VDD x192/WBLb x187/WBL x192/RBL1 x194/WBLb x188/WBL x192/RBL0 x194/RBL1 x186/WBLb
+ x194/RBL0 x190/WBL x186/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_50 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x195/WWL RWL_13 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x195/VDD VSUBS x196/RBL0 x197/WBLb x197/RBL1 x198/WBLb x199/WBL x197/RBL0
+ x198/RBL1 x200/WBLb x198/RBL0 x201/WBL x200/RBL1 x200/RBL0 x199/WBLb x202/WBL x203/WWL
+ x199/RBL1 x201/WBLb x199/RBL0 x204/WBL x201/RBL1 x201/RBL0 x196/WBL x203/VDD x202/WBLb
+ x197/WBL x202/RBL1 x204/WBLb x198/WBL x202/RBL0 x204/RBL1 x196/WBLb x204/RBL0 x200/WBL
+ x196/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_62 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x34/WWL RWL_1 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x34/VDD VSUBS x205/RBL0 x206/WBLb x206/RBL1 x207/WBLb x208/WBL x206/RBL0
+ x207/RBL1 x209/WBLb x207/RBL0 x210/WBL x209/RBL1 x209/RBL0 x208/WBLb x211/WBL x212/WWL
+ x208/RBL1 x210/WBLb x208/RBL0 x213/WBL x210/RBL1 x210/RBL0 x205/WBL x212/VDD x211/WBLb
+ x206/WBL x211/RBL1 x213/WBLb x207/WBL x211/RBL0 x213/RBL1 x205/WBLb x213/RBL0 x209/WBL
+ x205/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_120 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x130/WWL x16/RWL WBLb_16
+ WBL_16 WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21
+ WBLb_22 WBL_22 WBLb_23 WBL_23 x130/VDD VSUBS x214/RBL0 WBLb_16 x215/RBL1 x216/WBLb
+ x217/WBL x215/RBL0 x216/RBL1 x218/WBLb x216/RBL0 x219/WBL x218/RBL1 x218/RBL0 x217/WBLb
+ x220/WBL x221/WWL x217/RBL1 x219/WBLb x217/RBL0 x222/WBL RBL1_21 x219/RBL0 x214/WBL
+ x221/VDD x220/WBLb x215/WBL x220/RBL1 x222/WBLb x216/WBL x220/RBL0 x222/RBL1 x214/WBLb
+ x222/RBL0 x218/WBL x214/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_73 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x175/WWL RWL_27 WBLb_24
+ WBL_24 WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29
+ WBLb_30 WBL_30 WBLb_31 WBL_31 x175/VDD VSUBS x223/RBL0 x224/WBLb x224/RBL1 x225/WBLb
+ x226/WBL x224/RBL0 x225/RBL1 x227/WBLb x225/RBL0 x228/WBL x227/RBL1 x227/RBL0 x226/WBLb
+ x229/WBL x224/WWL x226/RBL1 x228/WBLb x226/RBL0 x230/WBL x228/RBL1 x228/RBL0 x223/WBL
+ x224/VDD x229/WBLb x224/WBL x229/RBL1 x230/WBLb x225/WBL x229/RBL0 x230/RBL1 x223/WBLb
+ x230/RBL0 x227/WBL x223/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_40 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x231/WWL RWL_25 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x231/VDD VSUBS x232/RBL0 WBLb_8 x233/RBL1 WBLb_11 WBL_10 x233/RBL0
+ x234/RBL1 WBLb_15 x234/RBL0 WBL_13 x235/RBL1 x235/RBL0 WBLb_10 WBL_9 x236/WWL x237/RBL1
+ WBLb_13 x237/RBL0 WBL_12 x238/RBL1 x238/RBL0 WBL_14 x236/VDD WBLb_9 WBL_8 x239/RBL1
+ WBLb_12 WBL_11 x239/RBL0 x240/RBL1 WBLb_14 x240/RBL0 WBL_15 x232/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_84 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x241/WWL RWL_21 WBLb_16
+ WBL_16 WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21
+ WBLb_22 WBL_22 WBLb_23 WBL_23 x241/VDD VSUBS x242/RBL0 WBLb_16 x243/RBL1 x244/WBLb
+ x245/WBL x243/RBL0 x244/RBL1 x246/WBLb x244/RBL0 x247/WBL x246/RBL1 x246/RBL0 x245/WBLb
+ x248/WBL x249/WWL x245/RBL1 x247/WBLb x245/RBL0 x250/WBL RBL1_21 x247/RBL0 x242/WBL
+ x249/VDD x248/WBLb x243/WBL x248/RBL1 x250/WBLb x244/WBL x248/RBL0 x250/RBL1 x242/WBLb
+ x250/RBL0 x246/WBL x242/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_95 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x193/WWL RWL_16 WBLb_24
+ WBL_24 WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29
+ WBLb_30 WBL_30 WBLb_31 WBL_31 x193/VDD VSUBS x251/RBL0 x252/WBLb x252/RBL1 x253/WBLb
+ x254/WBL x252/RBL0 x253/RBL1 x255/WBLb x253/RBL0 x256/WBL x255/RBL1 x255/RBL0 x254/WBLb
+ x257/WBL x252/WWL x254/RBL1 x256/WBLb x254/RBL0 x258/WBL x256/RBL1 x256/RBL0 x251/WBL
+ x252/VDD x257/WBLb x252/WBL x257/RBL1 x258/WBLb x253/WBL x257/RBL0 x258/RBL1 x251/WBLb
+ x258/RBL0 x255/WBL x251/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_51 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x259/WWL RWL_12 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x259/VDD VSUBS RBL0_14 x260/WBLb RBL1_8 x261/WBLb x262/WBL RBL0_8
+ RBL1_11 x263/WBLb RBL0_11 x264/WBL RBL1_15 RBL0_15 x262/WBLb x265/WBL x266/WWL RBL1_10
+ x264/WBLb RBL0_10 x267/WBL RBL1_13 RBL0_13 x268/WBL x266/VDD x265/WBLb x260/WBL
+ RBL1_9 x267/WBLb x261/WBL RBL0_9 RBL1_12 x268/WBLb RBL0_12 x263/WBL RBL1_14 VSUBS
+ x10T_1x8_magic
X10T_1x8_magic_63 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x25/WWL RWL_0 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x25/VDD VSUBS x269/RBL0 x270/WBLb x270/RBL1 x271/WBLb x272/WBL x270/RBL0
+ x271/RBL1 x273/WBLb x271/RBL0 x274/WBL x273/RBL1 x273/RBL0 x272/WBLb x275/WBL x276/WWL
+ x272/RBL1 x274/WBLb x272/RBL0 x277/WBL x274/RBL1 x274/RBL0 x269/WBL x276/VDD x275/WBLb
+ x270/WBL x275/RBL1 x277/WBLb x271/WBL x275/RBL0 x277/RBL1 x269/WBLb x277/RBL0 x273/WBL
+ x269/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_121 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x221/WWL x221/RWL WBLb_24
+ WBL_24 WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29
+ WBLb_30 WBL_30 WBLb_31 WBL_31 x221/VDD VSUBS x278/RBL0 x279/WBLb x279/RBL1 x280/WBLb
+ x281/WBL x279/RBL0 x280/RBL1 x282/WBLb x280/RBL0 x283/WBL x282/RBL1 x282/RBL0 x281/WBLb
+ x284/WBL x279/WWL x281/RBL1 x283/WBLb x281/RBL0 x285/WBL x283/RBL1 x283/RBL0 x278/WBL
+ x279/VDD x284/WBLb x279/WBL x284/RBL1 x285/WBLb x280/WBL x284/RBL0 x285/RBL1 x278/WBLb
+ x285/RBL0 x282/WBL x278/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_74 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x286/WWL RWL_26 WBLb_16
+ WBL_16 WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21
+ WBLb_22 WBL_22 WBLb_23 WBL_23 x286/VDD VSUBS x287/RBL0 WBLb_16 x288/RBL1 x289/WBLb
+ x290/WBL x288/RBL0 x289/RBL1 x291/WBLb x289/RBL0 x292/WBL x291/RBL1 x291/RBL0 x290/WBLb
+ x293/WBL x294/WWL x290/RBL1 x292/WBLb x290/RBL0 x295/WBL RBL1_21 x292/RBL0 x287/WBL
+ x294/VDD x293/WBLb x288/WBL x293/RBL1 x295/WBLb x289/WBL x293/RBL0 x295/RBL1 x287/WBLb
+ x295/RBL0 x291/WBL x287/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_41 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x296/WWL RWL_22 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x296/VDD VSUBS x297/RBL0 x298/WBLb x298/RBL1 x299/WBLb x300/WBL x298/RBL0
+ x299/RBL1 x301/WBLb x299/RBL0 x302/WBL x301/RBL1 x301/RBL0 x300/WBLb x303/WBL x140/WWL
+ x300/RBL1 x302/WBLb x300/RBL0 x304/WBL x302/RBL1 x302/RBL0 x297/WBL x140/VDD x303/WBLb
+ x298/WBL x303/RBL1 x304/WBLb x299/WBL x303/RBL0 x304/RBL1 x297/WBLb x304/RBL0 x301/WBL
+ x297/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_85 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x249/WWL RWL_21 WBLb_24
+ WBL_24 WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29
+ WBLb_30 WBL_30 WBLb_31 WBL_31 x249/VDD VSUBS x305/RBL0 x306/WBLb x306/RBL1 x307/WBLb
+ x308/WBL x306/RBL0 x307/RBL1 x309/WBLb x307/RBL0 x310/WBL x309/RBL1 x309/RBL0 x308/WBLb
+ x311/WBL x306/WWL x308/RBL1 x310/WBLb x308/RBL0 x312/WBL x310/RBL1 x310/RBL0 x305/WBL
+ x306/VDD x311/WBLb x306/WBL x311/RBL1 x312/WBLb x307/WBL x311/RBL0 x312/RBL1 x305/WBLb
+ x312/RBL0 x309/WBL x305/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_30 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_18 RWL_18 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x313/RBL0
+ x314/WBLb x314/RBL1 x315/WBLb x316/WBL x314/RBL0 x315/RBL1 x317/WBLb x315/RBL0 x318/WBL
+ x317/RBL1 x317/RBL0 x316/WBLb x319/WBL x320/WWL x316/RBL1 x318/WBLb x316/RBL0 x321/WBL
+ x318/RBL1 x318/RBL0 x313/WBL x320/VDD x319/WBLb x314/WBL x319/RBL1 x321/WBLb x315/WBL
+ x319/RBL0 x321/RBL1 x313/WBLb x321/RBL0 x317/WBL x313/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_96 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x322/WWL RWL_15 WBLb_16
+ WBL_16 WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21
+ WBLb_22 WBL_22 WBLb_23 WBL_23 x322/VDD VSUBS x323/RBL0 WBLb_16 x324/RBL1 x325/WBLb
+ x326/WBL x324/RBL0 x325/RBL1 x327/WBLb x325/RBL0 x328/WBL x327/RBL1 x327/RBL0 x326/WBLb
+ x329/WBL x330/WWL x326/RBL1 x328/WBLb x326/RBL0 x331/WBL RBL1_21 x328/RBL0 x323/WBL
+ x330/VDD x329/WBLb x324/WBL x329/RBL1 x331/WBLb x325/WBL x329/RBL0 x331/RBL1 x323/WBLb
+ x331/RBL0 x327/WBL x323/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_52 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x332/WWL RWL_11 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x332/VDD VSUBS x333/RBL0 x334/WBLb x334/RBL1 x335/WBLb x336/WBL x334/RBL0
+ x335/RBL1 x337/WBLb x335/RBL0 x338/WBL x337/RBL1 x337/RBL0 x336/WBLb x339/WBL x340/WWL
+ x336/RBL1 x338/WBLb x336/RBL0 x341/WBL x338/RBL1 x338/RBL0 x333/WBL x340/VDD x339/WBLb
+ x334/WBL x339/RBL1 x341/WBLb x335/WBL x339/RBL0 x341/RBL1 x333/WBLb x341/RBL0 x337/WBL
+ x333/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_110 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x342/WWL RWL_8 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x342/VDD VSUBS x343/RBL0 WBLb_16 x344/RBL1 x345/WBLb x346/WBL
+ x344/RBL0 x345/RBL1 x347/WBLb x345/RBL0 x348/WBL x347/RBL1 x347/RBL0 x346/WBLb x349/WBL
+ x350/WWL x346/RBL1 x348/WBLb x346/RBL0 x351/WBL RBL1_21 x348/RBL0 x343/WBL x350/VDD
+ x349/WBLb x344/WBL x349/RBL1 x351/WBLb x345/WBL x349/RBL0 x351/RBL1 x343/WBLb x351/RBL0
+ x347/WBL x343/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_122 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x164/WWL RWL_2 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x164/VDD VSUBS RBL0_22 WBLb_16 RBL1_16 x352/WBLb x353/WBL
+ RBL0_16 RBL1_19 x354/WBLb RBL0_19 x355/WBL RBL1_23 RBL0_23 x353/WBLb x356/WBL x357/WWL
+ RBL1_18 x355/WBLb RBL0_18 x358/WBL RBL1_21 RBL0_21 x359/WBL x357/VDD x356/WBLb x360/WBL
+ RBL1_17 x358/WBLb x352/WBL RBL0_17 RBL1_20 x359/WBLb RBL0_20 x354/WBL RBL1_22 VSUBS
+ x10T_1x8_magic
X10T_1x8_magic_64 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x361/WWL RWL_31 WBLb_16
+ WBL_16 WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21
+ WBLb_22 WBL_22 WBLb_23 WBL_23 x361/VDD VSUBS x362/RBL0 WBLb_16 x363/RBL1 x364/WBLb
+ x365/WBL x363/RBL0 x364/RBL1 x366/WBLb x364/RBL0 x367/WBL x366/RBL1 x366/RBL0 x365/WBLb
+ x368/WBL x369/WWL x365/RBL1 x367/WBLb x365/RBL0 x370/WBL RBL1_21 x367/RBL0 x362/WBL
+ x369/VDD x368/WBLb x363/WBL x368/RBL1 x370/WBLb x364/WBL x368/RBL0 x370/RBL1 x362/WBLb
+ x370/RBL0 x366/WBL x362/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_20 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_28 RWL_28 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND RBL0_6
+ x371/WBLb RBL1_0 x372/WBLb x373/WBL RBL0_0 RBL1_3 x374/WBLb RBL0_3 x375/WBL RBL1_7
+ RBL0_7 x373/WBLb x376/WBL x377/WWL RBL1_2 x375/WBLb RBL0_2 x378/WBL RBL1_5 RBL0_5
+ x379/WBL x377/VDD x376/WBLb x371/WBL RBL1_1 x378/WBLb x372/WBL RBL0_1 RBL1_4 x379/WBLb
+ RBL0_4 x374/WBL RBL1_6 VSUBS x10T_1x8_magic
X10T_1x8_magic_75 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x294/WWL RWL_26 WBLb_24
+ WBL_24 WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29
+ WBLb_30 WBL_30 WBLb_31 WBL_31 x294/VDD VSUBS x380/RBL0 x381/WBLb x381/RBL1 x382/WBLb
+ x383/WBL x381/RBL0 x382/RBL1 x384/WBLb x382/RBL0 x385/WBL x384/RBL1 x384/RBL0 x383/WBLb
+ x386/WBL x381/WWL x383/RBL1 x385/WBLb x383/RBL0 x387/WBL x385/RBL1 x385/RBL0 x380/WBL
+ x381/VDD x386/WBLb x381/WBL x386/RBL1 x387/WBLb x382/WBL x386/RBL0 x387/RBL1 x380/WBLb
+ x387/RBL0 x384/WBL x380/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_42 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x388/WWL RWL_21 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x388/VDD VSUBS x389/RBL0 x390/WBLb x390/RBL1 x391/WBLb x392/WBL x390/RBL0
+ x391/RBL1 x393/WBLb x391/RBL0 x394/WBL x393/RBL1 x393/RBL0 x392/WBLb x395/WBL x241/WWL
+ x392/RBL1 x394/WBLb x392/RBL0 x396/WBL x394/RBL1 x394/RBL0 x389/WBL x241/VDD x395/WBLb
+ x390/WBL x395/RBL1 x396/WBLb x391/WBL x395/RBL0 x396/RBL1 x389/WBLb x396/RBL0 x393/WBL
+ x389/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_86 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x397/WWL RWL_20 WBLb_16
+ WBL_16 WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21
+ WBLb_22 WBL_22 WBLb_23 WBL_23 VDD VSUBS x398/RBL0 WBLb_16 x399/RBL1 x400/WBLb x401/WBL
+ x399/RBL0 x400/RBL1 x402/WBLb x400/RBL0 x403/WBL x402/RBL1 x402/RBL0 x401/WBLb x404/WBL
+ x405/WWL x401/RBL1 x403/WBLb x401/RBL0 x406/WBL RBL1_21 x403/RBL0 x398/WBL VDD x404/WBLb
+ x399/WBL x404/RBL1 x406/WBLb x400/WBL x404/RBL0 x406/RBL1 x398/WBLb x406/RBL0 x402/WBL
+ x398/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_31 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_16 RWL_16 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x407/RBL0
+ x408/WBLb x408/RBL1 x409/WBLb x410/WBL x408/RBL0 x409/RBL1 x411/WBLb x409/RBL0 x412/WBL
+ x411/RBL1 x411/RBL0 x410/WBLb x413/WBL x414/WWL x410/RBL1 x412/WBLb x410/RBL0 x415/WBL
+ x412/RBL1 x412/RBL0 x407/WBL x414/VDD x413/WBLb x408/WBL x413/RBL1 x415/WBLb x409/WBL
+ x413/RBL0 x415/RBL1 x407/WBLb x415/RBL0 x411/WBL x407/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_97 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x330/WWL RWL_15 WBLb_24
+ WBL_24 WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29
+ WBLb_30 WBL_30 WBLb_31 WBL_31 x330/VDD VSUBS x416/RBL0 x417/WBLb x417/RBL1 x418/WBLb
+ x419/WBL x417/RBL0 x418/RBL1 x420/WBLb x418/RBL0 x421/WBL x420/RBL1 x420/RBL0 x419/WBLb
+ x422/WBL x417/WWL x419/RBL1 x421/WBLb x419/RBL0 x423/WBL x421/RBL1 x421/RBL0 x416/WBL
+ x417/VDD x422/WBLb x417/WBL x422/RBL1 x423/WBLb x418/WBL x422/RBL0 x423/RBL1 x416/WBLb
+ x423/RBL0 x420/WBL x416/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_100 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x203/WWL RWL_13 WBLb_16
+ WBL_16 WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21
+ WBLb_22 WBL_22 WBLb_23 WBL_23 x203/VDD VSUBS x424/RBL0 WBLb_16 x425/RBL1 x426/WBLb
+ x427/WBL x425/RBL0 x426/RBL1 x428/WBLb x426/RBL0 x429/WBL x428/RBL1 x428/RBL0 x427/WBLb
+ x430/WBL x431/WWL x427/RBL1 x429/WBLb x427/RBL0 x432/WBL RBL1_21 x429/RBL0 x424/WBL
+ x431/VDD x430/WBLb x425/WBL x430/RBL1 x432/WBLb x426/WBL x430/RBL0 x432/RBL1 x424/WBLb
+ x432/RBL0 x428/WBL x424/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_53 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x433/WWL RWL_10 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x433/VDD VSUBS x434/RBL0 x435/WBLb x435/RBL1 x436/WBLb x437/WBL x435/RBL0
+ x436/RBL1 x438/WBLb x436/RBL0 x439/WBL x438/RBL1 x438/RBL0 x437/WBLb x440/WBL x441/WWL
+ x437/RBL1 x439/WBLb x437/RBL0 x442/WBL x439/RBL1 x439/RBL0 x434/WBL x441/VDD x440/WBLb
+ x435/WBL x440/RBL1 x442/WBLb x436/WBL x440/RBL0 x442/RBL1 x434/WBLb x442/RBL0 x438/WBL
+ x434/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_111 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x350/WWL RWL_8 WBLb_24 WBL_24
+ WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29 WBLb_30
+ WBL_30 WBLb_31 WBL_31 x350/VDD VSUBS x443/RBL0 x444/WBLb x444/RBL1 x445/WBLb x446/WBL
+ x444/RBL0 x445/RBL1 x447/WBLb x445/RBL0 x448/WBL x447/RBL1 x447/RBL0 x446/WBLb x449/WBL
+ x444/WWL x446/RBL1 x448/WBLb x446/RBL0 x450/WBL x448/RBL1 x448/RBL0 x443/WBL x444/VDD
+ x449/WBLb x444/WBL x449/RBL1 x450/WBLb x445/WBL x449/RBL0 x450/RBL1 x443/WBLb x450/RBL0
+ x447/WBL x443/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_123 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x357/WWL RWL_2 WBLb_24 WBL_24
+ WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29 WBLb_30
+ WBL_30 WBLb_31 WBL_31 x357/VDD VSUBS RBL0_30 x451/WBLb RBL1_24 x452/WBLb x453/WBL
+ RBL0_24 RBL1_27 x454/WBLb RBL0_27 x455/WBL RBL1_31 RBL0_31 x453/WBLb x456/WBL x451/WWL
+ RBL1_26 x455/WBLb RBL0_26 x457/WBL RBL1_29 RBL0_29 x458/WBL x451/VDD x456/WBLb x451/WBL
+ RBL1_25 x457/WBLb x452/WBL RBL0_25 RBL1_28 x458/WBLb RBL0_28 x454/WBL RBL1_30 VSUBS
+ x10T_1x8_magic
X10T_1x8_magic_112 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x459/WWL RWL_7 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x459/VDD VSUBS RBL0_22 WBLb_16 RBL1_16 x460/WBLb x461/WBL
+ RBL0_16 RBL1_19 x462/WBLb RBL0_19 x463/WBL RBL1_23 RBL0_23 x461/WBLb x464/WBL x465/WWL
+ RBL1_18 x463/WBLb RBL0_18 x466/WBL RBL1_21 RBL0_21 x467/WBL x465/VDD x464/WBLb x468/WBL
+ RBL1_17 x466/WBLb x460/WBL RBL0_17 RBL1_20 x467/WBLb RBL0_20 x462/WBL RBL1_22 VSUBS
+ x10T_1x8_magic
X10T_1x8_magic_32 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x469/WWL RWL_30 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x469/VDD VSUBS x470/RBL0 x471/WBLb x471/RBL1 x472/WBLb x473/WBL x471/RBL0
+ x472/RBL1 x474/WBLb x472/RBL0 x475/WBL x474/RBL1 x474/RBL0 x473/WBLb x476/WBL x477/WWL
+ x473/RBL1 x475/WBLb x473/RBL0 x478/WBL x475/RBL1 x475/RBL0 x470/WBL x477/VDD x476/WBLb
+ x471/WBL x476/RBL1 x478/WBLb x472/WBL x476/RBL0 x478/RBL1 x470/WBLb x478/RBL0 x474/WBL
+ x470/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_65 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x477/WWL RWL_30 WBLb_16
+ WBL_16 WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21
+ WBLb_22 WBL_22 WBLb_23 WBL_23 x477/VDD VSUBS x479/RBL0 WBLb_16 x480/RBL1 x481/WBLb
+ x482/WBL x480/RBL0 x481/RBL1 x483/WBLb x481/RBL0 x484/WBL x483/RBL1 x483/RBL0 x482/WBLb
+ x485/WBL x486/WWL x482/RBL1 x484/WBLb x482/RBL0 x487/WBL RBL1_21 x484/RBL0 x479/WBL
+ x486/VDD x485/WBLb x480/WBL x485/RBL1 x487/WBLb x481/WBL x485/RBL0 x487/RBL1 x479/WBLb
+ x487/RBL0 x483/WBL x479/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_21 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_25 RWL_25 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x488/RBL0
+ WBLb_0 x489/RBL1 WBLb_3 WBL_2 x489/RBL0 x490/RBL1 WBLb_7 x490/RBL0 WBL_5 x491/RBL1
+ x491/RBL0 WBLb_2 WBL_1 x231/WWL x492/RBL1 WBLb_5 x492/RBL0 WBL_4 x493/RBL1 x493/RBL0
+ WBL_6 x231/VDD WBLb_1 WBL_0 x494/RBL1 WBLb_4 WBL_3 x494/RBL0 x495/RBL1 WBLb_6 x495/RBL0
+ WBL_7 x488/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_76 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x236/WWL RWL_25 WBLb_16
+ WBL_16 WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21
+ WBLb_22 WBL_22 WBLb_23 WBL_23 x236/VDD VSUBS x496/RBL0 WBLb_16 x497/RBL1 WBLb_19
+ WBL_18 x497/RBL0 x498/RBL1 WBLb_23 x498/RBL0 WBL_21 x499/RBL1 x499/RBL0 WBLb_18
+ WBL_17 x500/WWL x501/RBL1 WBLb_21 x501/RBL0 WBL_20 RBL1_21 x502/RBL0 WBL_22 x500/VDD
+ WBLb_17 WBL_16 x503/RBL1 WBLb_20 WBL_19 x503/RBL0 x504/RBL1 WBLb_22 x504/RBL0 WBL_23
+ x496/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_43 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x505/WWL RWL_20 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 VDD VSUBS x506/RBL0 x507/WBLb x507/RBL1 x508/WBLb x509/WBL x507/RBL0
+ x508/RBL1 x510/WBLb x508/RBL0 x511/WBL x510/RBL1 x510/RBL0 x509/WBLb x512/WBL x397/WWL
+ x509/RBL1 x511/WBLb x509/RBL0 x513/WBL x511/RBL1 x511/RBL0 x506/WBL VDD x512/WBLb
+ x507/WBL x512/RBL1 x513/WBLb x508/WBL x512/RBL0 x513/RBL1 x506/WBLb x513/RBL0 x510/WBL
+ x506/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_87 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x405/WWL RWL_20 WBLb_24
+ WBL_24 WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29
+ WBLb_30 WBL_30 WBLb_31 WBL_31 VDD VSUBS x514/RBL0 x515/WBLb x515/RBL1 x516/WBLb
+ x517/WBL x515/RBL0 x516/RBL1 x518/WBLb x516/RBL0 x519/WBL x518/RBL1 x518/RBL0 x517/WBLb
+ x520/WBL x515/WWL x517/RBL1 x519/WBLb x517/RBL0 x521/WBL x519/RBL1 x519/RBL0 x514/WBL
+ VDD x520/WBLb x515/WBL x520/RBL1 x521/WBLb x516/WBL x520/RBL0 x521/RBL1 x514/WBLb
+ x521/RBL0 x518/WBL x514/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_98 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x522/WWL RWL_14 WBLb_16
+ WBL_16 WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21
+ WBLb_22 WBL_22 WBLb_23 WBL_23 x522/VDD VSUBS RBL0_22 WBLb_16 RBL1_16 WBLb_19 WBL_18
+ RBL0_16 RBL1_19 WBLb_23 RBL0_19 WBL_21 RBL1_23 RBL0_23 WBLb_18 WBL_17 x523/WWL RBL1_18
+ WBLb_21 RBL0_18 WBL_20 RBL1_21 RBL0_21 WBL_22 x523/VDD WBLb_17 WBL_16 RBL1_17 WBLb_20
+ WBL_19 RBL0_17 RBL1_20 WBLb_22 RBL0_20 WBL_23 RBL1_22 VSUBS x10T_1x8_magic
X10T_1x8_magic_10 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_13 RWL_13 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x524/RBL0
+ x525/WBLb x525/RBL1 x526/WBLb x527/WBL x525/RBL0 x526/RBL1 x528/WBLb x526/RBL0 x529/WBL
+ x528/RBL1 x528/RBL0 x527/WBLb x530/WBL x195/WWL x527/RBL1 x529/WBLb x527/RBL0 x531/WBL
+ x529/RBL1 x529/RBL0 x524/WBL x195/VDD x530/WBLb x525/WBL x530/RBL1 x531/WBLb x526/WBL
+ x530/RBL0 x531/RBL1 x524/WBLb x531/RBL0 x528/WBL x524/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_101 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x431/WWL RWL_13 WBLb_24
+ WBL_24 WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29
+ WBLb_30 WBL_30 WBLb_31 WBL_31 x431/VDD VSUBS x532/RBL0 x533/WBLb x533/RBL1 x534/WBLb
+ x535/WBL x533/RBL0 x534/RBL1 x536/WBLb x534/RBL0 x537/WBL x536/RBL1 x536/RBL0 x535/WBLb
+ x538/WBL x533/WWL x535/RBL1 x537/WBLb x535/RBL0 x539/WBL x537/RBL1 x537/RBL0 x532/WBL
+ x533/VDD x538/WBLb x533/WBL x538/RBL1 x539/WBLb x534/WBL x538/RBL0 x539/RBL1 x532/WBLb
+ x539/RBL0 x536/WBL x532/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_54 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x540/WWL RWL_9 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x540/VDD VSUBS RBL0_14 WBLb_8 RBL1_8 WBLb_11 WBL_10 RBL0_8 RBL1_11
+ WBLb_15 RBL0_11 WBL_13 RBL1_15 RBL0_15 WBLb_10 WBL_9 x541/WWL RBL1_10 WBLb_13 RBL0_10
+ WBL_12 RBL1_13 RBL0_13 WBL_14 x541/VDD WBLb_9 WBL_8 RBL1_9 WBLb_12 WBL_11 RBL0_9
+ RBL1_12 WBLb_14 RBL0_12 WBL_15 RBL1_14 VSUBS x10T_1x8_magic
X10T_1x8_magic_124 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x212/WWL RWL_1 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x212/VDD VSUBS x542/RBL0 WBLb_16 x543/RBL1 x544/WBLb x545/WBL
+ x543/RBL0 x544/RBL1 x546/WBLb x544/RBL0 x547/WBL x546/RBL1 x546/RBL0 x545/WBLb x548/WBL
+ x549/WWL x545/RBL1 x547/WBLb x545/RBL0 x550/WBL RBL1_21 x547/RBL0 x542/WBL x549/VDD
+ x548/WBLb x543/WBL x548/RBL1 x550/WBLb x544/WBL x548/RBL0 x550/RBL1 x542/WBLb x550/RBL0
+ x546/WBL x542/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_113 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x465/WWL RWL_7 WBLb_24 WBL_24
+ WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29 WBLb_30
+ WBL_30 WBLb_31 WBL_31 x465/VDD VSUBS RBL0_30 x551/WBLb RBL1_24 x552/WBLb x553/WBL
+ RBL0_24 RBL1_27 x554/WBLb RBL0_27 x555/WBL RBL1_31 RBL0_31 x553/WBLb x556/WBL x551/WWL
+ RBL1_26 x555/WBLb RBL0_26 x557/WBL RBL1_29 RBL0_29 x558/WBL x551/VDD x556/WBLb x551/WBL
+ RBL1_25 x557/WBLb x552/WBL RBL0_25 RBL1_28 x558/WBLb RBL0_28 x554/WBL RBL1_30 VSUBS
+ x10T_1x8_magic
X10T_1x8_magic_33 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x559/WWL RWL_31 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x559/VDD VSUBS x560/RBL0 x561/WBLb x561/RBL1 x562/WBLb x563/WBL x561/RBL0
+ x562/RBL1 x564/WBLb x562/RBL0 x565/WBL x564/RBL1 x564/RBL0 x563/WBLb x566/WBL x361/WWL
+ x563/RBL1 x565/WBLb x563/RBL0 x567/WBL x565/RBL1 x565/RBL0 x560/WBL x361/VDD x566/WBLb
+ x561/WBL x566/RBL1 x567/WBLb x562/WBL x566/RBL0 x567/RBL1 x560/WBLb x567/RBL0 x564/WBL
+ x560/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_66 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x486/WWL RWL_30 WBLb_24
+ WBL_24 WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29
+ WBLb_30 WBL_30 WBLb_31 WBL_31 x486/VDD VSUBS x568/RBL0 x569/WBLb x569/RBL1 x570/WBLb
+ x571/WBL x569/RBL0 x570/RBL1 x572/WBLb x570/RBL0 x573/WBL x572/RBL1 x572/RBL0 x571/WBLb
+ x574/WBL x569/WWL x571/RBL1 x573/WBLb x571/RBL0 x575/WBL x573/RBL1 x573/RBL0 x568/WBL
+ x569/VDD x574/WBLb x569/WBL x574/RBL1 x575/WBLb x570/WBL x574/RBL0 x575/RBL1 x568/WBLb
+ x575/RBL0 x572/WBL x568/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_22 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_26 RWL_26 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x576/RBL0
+ x577/WBLb x577/RBL1 x578/WBLb x579/WBL x577/RBL0 x578/RBL1 x580/WBLb x578/RBL0 x581/WBL
+ x580/RBL1 x580/RBL0 x579/WBLb x582/WBL x583/WWL x579/RBL1 x581/WBLb x579/RBL0 x584/WBL
+ x581/RBL1 x581/RBL0 x576/WBL x583/VDD x582/WBLb x577/WBL x582/RBL1 x584/WBLb x578/WBL
+ x582/RBL0 x584/RBL1 x576/WBLb x584/RBL0 x580/WBL x576/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_77 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x585/WWL RWL_24 WBLb_16
+ WBL_16 WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21
+ WBLb_22 WBL_22 WBLb_23 WBL_23 x585/VDD VSUBS x586/RBL0 WBLb_16 x587/RBL1 x588/WBLb
+ x589/WBL x587/RBL0 x588/RBL1 x590/WBLb x588/RBL0 x591/WBL x590/RBL1 x590/RBL0 x589/WBLb
+ x592/WBL x593/WWL x589/RBL1 x591/WBLb x589/RBL0 x594/WBL RBL1_21 x591/RBL0 x586/WBL
+ x593/VDD x592/WBLb x587/WBL x592/RBL1 x594/WBLb x588/WBL x592/RBL0 x594/RBL1 x586/WBLb
+ x594/RBL0 x590/WBL x586/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_44 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x595/WWL RWL_19 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x595/VDD VSUBS x596/RBL0 x597/WBLb x597/RBL1 x598/WBLb x599/WBL x597/RBL0
+ x598/RBL1 x600/WBLb x598/RBL0 x601/WBL x600/RBL1 x600/RBL0 x599/WBLb x602/WBL x603/WWL
+ x599/RBL1 x601/WBLb x599/RBL0 x604/WBL x601/RBL1 x601/RBL0 x596/WBL x603/VDD x602/WBLb
+ x597/WBL x602/RBL1 x604/WBLb x598/WBL x602/RBL0 x604/RBL1 x596/WBLb x604/RBL0 x600/WBL
+ x596/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_88 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x603/WWL RWL_19 WBLb_16
+ WBL_16 WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21
+ WBLb_22 WBL_22 WBLb_23 WBL_23 x603/VDD VSUBS x605/RBL0 WBLb_16 x606/RBL1 x607/WBLb
+ x608/WBL x606/RBL0 x607/RBL1 x609/WBLb x607/RBL0 x610/WBL x609/RBL1 x609/RBL0 x608/WBLb
+ x611/WBL x612/WWL x608/RBL1 x610/WBLb x608/RBL0 x613/WBL RBL1_21 x610/RBL0 x605/WBL
+ x612/VDD x611/WBLb x606/WBL x611/RBL1 x613/WBLb x607/WBL x611/RBL0 x613/RBL1 x605/WBLb
+ x613/RBL0 x609/WBL x605/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_99 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x523/WWL RWL_14 WBLb_24
+ WBL_24 WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29
+ WBLb_30 WBL_30 WBLb_31 WBL_31 x523/VDD VSUBS RBL0_30 WBLb_24 RBL1_24 WBLb_27 WBL_26
+ RBL0_24 RBL1_27 WBLb_31 RBL0_27 WBL_29 RBL1_31 RBL0_31 WBLb_26 WBL_25 x614/WWL RBL1_26
+ WBLb_29 RBL0_26 WBL_28 RBL1_29 RBL0_29 WBL_30 x614/VDD WBLb_25 WBL_24 RBL1_25 WBLb_28
+ WBL_27 RBL0_25 RBL1_28 WBLb_30 RBL0_28 WBL_31 RBL1_30 VSUBS x10T_1x8_magic
X10T_1x8_magic_11 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_12 RWL_12 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND RBL0_6
+ x615/WBLb RBL1_0 x616/WBLb x617/WBL RBL0_0 RBL1_3 x618/WBLb RBL0_3 x619/WBL RBL1_7
+ RBL0_7 x617/WBLb x620/WBL x259/WWL RBL1_2 x619/WBLb RBL0_2 x621/WBL RBL1_5 RBL0_5
+ x622/WBL x259/VDD x620/WBLb x615/WBL RBL1_1 x621/WBLb x616/WBL RBL0_1 RBL1_4 x622/WBLb
+ RBL0_4 x618/WBL RBL1_6 VSUBS x10T_1x8_magic
X10T_1x8_magic_102 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x266/WWL RWL_12 WBLb_16
+ WBL_16 WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21
+ WBLb_22 WBL_22 WBLb_23 WBL_23 x266/VDD VSUBS RBL0_22 WBLb_16 RBL1_16 x623/WBLb x624/WBL
+ RBL0_16 RBL1_19 x625/WBLb RBL0_19 x626/WBL RBL1_23 RBL0_23 x624/WBLb x627/WBL x628/WWL
+ RBL1_18 x626/WBLb RBL0_18 x629/WBL RBL1_21 RBL0_21 x630/WBL x628/VDD x627/WBLb x631/WBL
+ RBL1_17 x629/WBLb x623/WBL RBL0_17 RBL1_20 x630/WBLb RBL0_20 x625/WBL RBL1_22 VSUBS
+ x10T_1x8_magic
X10T_1x8_magic_55 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x632/WWL RWL_8 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x632/VDD VSUBS x633/RBL0 x634/WBLb x634/RBL1 x635/WBLb x636/WBL x634/RBL0
+ x635/RBL1 x637/WBLb x635/RBL0 x638/WBL x637/RBL1 x637/RBL0 x636/WBLb x639/WBL x342/WWL
+ x636/RBL1 x638/WBLb x636/RBL0 x640/WBL x638/RBL1 x638/RBL0 x633/WBL x342/VDD x639/WBLb
+ x634/WBL x639/RBL1 x640/WBLb x635/WBL x639/RBL0 x640/RBL1 x633/WBLb x640/RBL0 x637/WBL
+ x633/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_12 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_11 RWL_11 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x641/RBL0
+ x642/WBLb x642/RBL1 x643/WBLb x644/WBL x642/RBL0 x643/RBL1 x645/WBLb x643/RBL0 x646/WBL
+ x645/RBL1 x645/RBL0 x644/WBLb x647/WBL x332/WWL x644/RBL1 x646/WBLb x644/RBL0 x648/WBL
+ x646/RBL1 x646/RBL0 x641/WBL x332/VDD x647/WBLb x642/WBL x647/RBL1 x648/WBLb x643/WBL
+ x647/RBL0 x648/RBL1 x641/WBLb x648/RBL0 x645/WBL x641/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_125 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x549/WWL RWL_1 WBLb_24 WBL_24
+ WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29 WBLb_30
+ WBL_30 WBLb_31 WBL_31 x549/VDD VSUBS x649/RBL0 x650/WBLb x650/RBL1 x651/WBLb x652/WBL
+ x650/RBL0 x651/RBL1 x653/WBLb x651/RBL0 x654/WBL x653/RBL1 x653/RBL0 x652/WBLb x655/WBL
+ x650/WWL x652/RBL1 x654/WBLb x652/RBL0 x656/WBL x654/RBL1 x654/RBL0 x649/WBL x650/VDD
+ x655/WBLb x650/WBL x655/RBL1 x656/WBLb x651/WBL x655/RBL0 x656/RBL1 x649/WBLb x656/RBL0
+ x653/WBL x649/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_114 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x657/WWL RWL_6 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x657/VDD VSUBS x658/RBL0 WBLb_16 x659/RBL1 x660/WBLb x661/WBL
+ x659/RBL0 x660/RBL1 x662/WBLb x660/RBL0 x663/WBL x662/RBL1 x662/RBL0 x661/WBLb x664/WBL
+ x665/WWL x661/RBL1 x663/WBLb x661/RBL0 x666/WBL RBL1_21 x663/RBL0 x658/WBL x665/VDD
+ x664/WBLb x659/WBL x664/RBL1 x666/WBLb x660/WBL x664/RBL0 x666/RBL1 x658/WBLb x666/RBL0
+ x662/WBL x658/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_56 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x42/WWL RWL_7 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x42/VDD VSUBS RBL0_14 x667/WBLb RBL1_8 x668/WBLb x669/WBL RBL0_8
+ RBL1_11 x670/WBLb RBL0_11 x671/WBL RBL1_15 RBL0_15 x669/WBLb x672/WBL x459/WWL RBL1_10
+ x671/WBLb RBL0_10 x673/WBL RBL1_13 RBL0_13 x674/WBL x459/VDD x672/WBLb x667/WBL
+ RBL1_9 x673/WBLb x668/WBL RBL0_9 RBL1_12 x674/WBLb RBL0_12 x670/WBL RBL1_14 VSUBS
+ x10T_1x8_magic
X10T_1x8_magic_67 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x369/WWL RWL_31 WBLb_24
+ WBL_24 WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29
+ WBLb_30 WBL_30 WBLb_31 WBL_31 x369/VDD VSUBS x675/RBL0 x676/WBLb x676/RBL1 x677/WBLb
+ x678/WBL x676/RBL0 x677/RBL1 x679/WBLb x677/RBL0 x680/WBL x679/RBL1 x679/RBL0 x678/WBLb
+ x681/WBL x676/WWL x678/RBL1 x680/WBLb x678/RBL0 x682/WBL x680/RBL1 x680/RBL0 x675/WBL
+ x676/VDD x681/WBLb x676/WBL x681/RBL1 x682/WBLb x677/WBL x681/RBL0 x682/RBL1 x675/WBLb
+ x682/RBL0 x679/WBL x675/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_34 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x377/WWL RWL_28 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x377/VDD VSUBS RBL0_14 x683/WBLb RBL1_8 x684/WBLb x685/WBL RBL0_8
+ RBL1_11 x686/WBLb RBL0_11 x687/WBL RBL1_15 RBL0_15 x685/WBLb x688/WBL x95/WWL RBL1_10
+ x687/WBLb RBL0_10 x689/WBL RBL1_13 RBL0_13 x690/WBL x95/VDD x688/WBLb x683/WBL RBL1_9
+ x689/WBLb x684/WBL RBL0_9 RBL1_12 x690/WBLb RBL0_12 x686/WBL RBL1_14 VSUBS x10T_1x8_magic
X10T_1x8_magic_78 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x593/WWL RWL_24 WBLb_24
+ WBL_24 WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29
+ WBLb_30 WBL_30 WBLb_31 WBL_31 x593/VDD VSUBS x691/RBL0 x692/WBLb x692/RBL1 x693/WBLb
+ x694/WBL x692/RBL0 x693/RBL1 x695/WBLb x693/RBL0 x696/WBL x695/RBL1 x695/RBL0 x694/WBLb
+ x697/WBL x692/WWL x694/RBL1 x696/WBLb x694/RBL0 x698/WBL x696/RBL1 x696/RBL0 x691/WBL
+ x692/VDD x697/WBLb x692/WBL x697/RBL1 x698/WBLb x693/WBL x697/RBL0 x698/RBL1 x691/WBLb
+ x698/RBL0 x695/WBL x691/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_23 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_23 RWL_23 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND RBL0_6
+ WBLb_0 RBL1_0 WBLb_3 WBL_2 RBL0_0 RBL1_3 WBLb_7 RBL0_3 WBL_5 RBL1_7 RBL0_7 WBLb_2
+ WBL_1 x699/WWL RBL1_2 WBLb_5 RBL0_2 WBL_4 RBL1_5 RBL0_5 WBL_6 VDD WBLb_1 WBL_0 RBL1_1
+ WBLb_4 WBL_3 RBL0_1 RBL1_4 WBLb_6 RBL0_4 WBL_7 RBL1_6 VSUBS x10T_1x8_magic
X10T_1x8_magic_89 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x612/WWL RWL_19 WBLb_24
+ WBL_24 WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29
+ WBLb_30 WBL_30 WBLb_31 WBL_31 x612/VDD VSUBS x700/RBL0 x701/WBLb x701/RBL1 x702/WBLb
+ x703/WBL x701/RBL0 x702/RBL1 x704/WBLb x702/RBL0 x705/WBL x704/RBL1 x704/RBL0 x703/WBLb
+ x706/WBL x701/WWL x703/RBL1 x705/WBLb x703/RBL0 x707/WBL x705/RBL1 x705/RBL0 x700/WBL
+ x701/VDD x706/WBLb x701/WBL x706/RBL1 x707/WBLb x702/WBL x706/RBL0 x707/RBL1 x700/WBLb
+ x707/RBL0 x704/WBL x700/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_45 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x708/WWL RWL_17 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x708/VDD VSUBS x709/RBL0 x710/WBLb x710/RBL1 x711/WBLb x712/WBL x710/RBL0
+ x711/RBL1 x713/WBLb x711/RBL0 x714/WBL x713/RBL1 x713/RBL0 x712/WBLb x715/WBL x72/WWL
+ x712/RBL1 x714/WBLb x712/RBL0 x716/WBL x714/RBL1 x714/RBL0 x709/WBL x72/VDD x715/WBLb
+ x710/WBL x715/RBL1 x716/WBLb x711/WBL x715/RBL0 x716/RBL1 x709/WBLb x716/RBL0 x713/WBL
+ x709/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_103 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x628/WWL RWL_12 WBLb_24
+ WBL_24 WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29
+ WBLb_30 WBL_30 WBLb_31 WBL_31 x628/VDD VSUBS RBL0_30 x717/WBLb RBL1_24 x718/WBLb
+ x719/WBL RBL0_24 RBL1_27 x720/WBLb RBL0_27 x721/WBL RBL1_31 RBL0_31 x719/WBLb x722/WBL
+ x717/WWL RBL1_26 x721/WBLb RBL0_26 x723/WBL RBL1_29 RBL0_29 x724/WBL x717/VDD x722/WBLb
+ x717/WBL RBL1_25 x723/WBLb x718/WBL RBL0_25 RBL1_28 x724/WBLb RBL0_28 x720/WBL RBL1_30
+ VSUBS x10T_1x8_magic
X10T_1x8_magic_126 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x276/WWL RWL_0 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x276/VDD VSUBS x725/RBL0 WBLb_16 x726/RBL1 x727/WBLb x728/WBL
+ x726/RBL0 x727/RBL1 x729/WBLb x727/RBL0 x730/WBL x729/RBL1 x729/RBL0 x728/WBLb x731/WBL
+ x732/WWL x728/RBL1 x730/WBLb x728/RBL0 x733/WBL RBL1_21 x730/RBL0 x725/WBL x732/VDD
+ x731/WBLb x726/WBL x731/RBL1 x733/WBLb x727/WBL x731/RBL0 x733/RBL1 x725/WBLb x733/RBL0
+ x729/WBL x725/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_115 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x665/WWL RWL_6 WBLb_24 WBL_24
+ WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29 WBLb_30
+ WBL_30 WBLb_31 WBL_31 x665/VDD VSUBS x734/RBL0 x735/WBLb x735/RBL1 x736/WBLb x737/WBL
+ x735/RBL0 x736/RBL1 x738/WBLb x736/RBL0 x739/WBL x738/RBL1 x738/RBL0 x737/WBLb x740/WBL
+ x735/WWL x737/RBL1 x739/WBLb x737/RBL0 x741/WBL x739/RBL1 x739/RBL0 x734/WBL x735/VDD
+ x740/WBLb x735/WBL x740/RBL1 x741/WBLb x736/WBL x740/RBL0 x741/RBL1 x734/WBLb x741/RBL0
+ x738/WBL x734/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_57 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x52/WWL RWL_6 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x52/VDD VSUBS x742/RBL0 x743/WBLb x743/RBL1 x744/WBLb x745/WBL x743/RBL0
+ x744/RBL1 x746/WBLb x744/RBL0 x747/WBL x746/RBL1 x746/RBL0 x745/WBLb x748/WBL x657/WWL
+ x745/RBL1 x747/WBLb x745/RBL0 x749/WBL x747/RBL1 x747/RBL0 x742/WBL x657/VDD x748/WBLb
+ x743/WBL x748/RBL1 x749/WBLb x744/WBL x748/RBL0 x749/RBL1 x742/WBLb x749/RBL0 x746/WBL
+ x742/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_35 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x750/WWL RWL_29 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x750/VDD VSUBS x751/RBL0 x752/WBLb x752/RBL1 x753/WBLb x754/WBL x752/RBL0
+ x753/RBL1 x755/WBLb x753/RBL0 x756/WBL x755/RBL1 x755/RBL0 x754/WBLb x757/WBL x758/WWL
+ x754/RBL1 x756/WBLb x754/RBL0 x759/WBL x756/RBL1 x756/RBL0 x751/WBL x758/VDD x757/WBLb
+ x752/WBL x757/RBL1 x759/WBLb x753/WBL x757/RBL0 x759/RBL1 x751/WBLb x759/RBL0 x755/WBL
+ x751/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_68 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x758/WWL RWL_29 WBLb_16
+ WBL_16 WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21
+ WBLb_22 WBL_22 WBLb_23 WBL_23 x758/VDD VSUBS x760/RBL0 WBLb_16 x761/RBL1 x762/WBLb
+ x763/WBL x761/RBL0 x762/RBL1 x764/WBLb x762/RBL0 x765/WBL x764/RBL1 x764/RBL0 x763/WBLb
+ x766/WBL x767/WWL x763/RBL1 x765/WBLb x763/RBL0 x768/WBL RBL1_21 x765/RBL0 x760/WBL
+ x767/VDD x766/WBLb x761/WBL x766/RBL1 x768/WBLb x762/WBL x766/RBL0 x768/RBL1 x760/WBLb
+ x768/RBL0 x764/WBL x760/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_79 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x500/WWL RWL_25 WBLb_24
+ WBL_24 WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29
+ WBLb_30 WBL_30 WBLb_31 WBL_31 x500/VDD VSUBS x769/RBL0 WBLb_24 x770/RBL1 WBLb_27
+ WBL_26 x770/RBL0 x771/RBL1 WBLb_31 x771/RBL0 WBL_29 x772/RBL1 x772/RBL0 WBLb_26
+ WBL_25 x770/WWL x773/RBL1 WBLb_29 x773/RBL0 WBL_28 x774/RBL1 x774/RBL0 WBL_30 x770/VDD
+ WBLb_25 WBL_24 x775/RBL1 WBLb_28 WBL_27 x775/RBL0 x776/RBL1 WBLb_30 x776/RBL0 WBL_31
+ x769/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_24 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_24 RWL_24 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x777/RBL0
+ x778/WBLb x778/RBL1 x779/WBLb x780/WBL x778/RBL0 x779/RBL1 x781/WBLb x779/RBL0 x782/WBL
+ x781/RBL1 x781/RBL0 x780/WBLb x783/WBL x784/WWL x780/RBL1 x782/WBLb x780/RBL0 x785/WBL
+ x782/RBL1 x782/RBL0 x777/WBL x784/VDD x783/WBLb x778/WBL x783/RBL1 x785/WBLb x779/WBL
+ x783/RBL0 x785/RBL1 x777/WBLb x785/RBL0 x781/WBL x777/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_46 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x320/WWL RWL_18 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x320/VDD VSUBS x786/RBL0 x787/WBLb x787/RBL1 x788/WBLb x789/WBL x787/RBL0
+ x788/RBL1 x790/WBLb x788/RBL0 x791/WBL x790/RBL1 x790/RBL0 x789/WBLb x792/WBL x85/WWL
+ x789/RBL1 x791/WBLb x789/RBL0 x793/WBL x791/RBL1 x791/RBL0 x786/WBL x85/VDD x792/WBLb
+ x787/WBL x792/RBL1 x793/WBLb x788/WBL x792/RBL0 x793/RBL1 x786/WBLb x793/RBL0 x790/WBL
+ x786/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_104 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x340/WWL RWL_11 WBLb_16
+ WBL_16 WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21
+ WBLb_22 WBL_22 WBLb_23 WBL_23 x340/VDD VSUBS x794/RBL0 WBLb_16 x795/RBL1 x796/WBLb
+ x797/WBL x795/RBL0 x796/RBL1 x798/WBLb x796/RBL0 x799/WBL x798/RBL1 x798/RBL0 x797/WBLb
+ x800/WBL x801/WWL x797/RBL1 x799/WBLb x797/RBL0 x802/WBL RBL1_21 x799/RBL0 x794/WBL
+ x801/VDD x800/WBLb x795/WBL x800/RBL1 x802/WBLb x796/WBL x800/RBL0 x802/RBL1 x794/WBLb
+ x802/RBL0 x798/WBL x794/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_13 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_10 RWL_10 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x803/RBL0
+ x804/WBLb x804/RBL1 x805/WBLb x806/WBL x804/RBL0 x805/RBL1 x807/WBLb x805/RBL0 x808/WBL
+ x807/RBL1 x807/RBL0 x806/WBLb x809/WBL x433/WWL x806/RBL1 x808/WBLb x806/RBL0 x810/WBL
+ x808/RBL1 x808/RBL0 x803/WBL x433/VDD x809/WBLb x804/WBL x809/RBL1 x810/WBLb x805/WBL
+ x809/RBL0 x810/RBL1 x803/WBLb x810/RBL0 x807/WBL x803/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_127 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x732/WWL RWL_0 WBLb_24 WBL_24
+ WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29 WBLb_30
+ WBL_30 WBLb_31 WBL_31 x732/VDD VSUBS x811/RBL0 x812/WBLb x812/RBL1 x813/WBLb x814/WBL
+ x812/RBL0 x813/RBL1 x815/WBLb x813/RBL0 x816/WBL x815/RBL1 x815/RBL0 x814/WBLb x817/WBL
+ x812/WWL x814/RBL1 x816/WBLb x814/RBL0 x818/WBL x816/RBL1 x816/RBL0 x811/WBL x812/VDD
+ x817/WBLb x812/WBL x817/RBL1 x818/WBLb x813/WBL x817/RBL0 x818/RBL1 x811/WBLb x818/RBL0
+ x815/WBL x811/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_116 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x819/WWL RWL_4 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x819/VDD VSUBS x820/RBL0 WBLb_16 x821/RBL1 WBLb_19 WBL_18
+ x821/RBL0 x822/RBL1 WBLb_23 x822/RBL0 WBL_21 x823/RBL1 x823/RBL0 WBLb_18 WBL_17
+ x824/WWL x825/RBL1 WBLb_21 x825/RBL0 WBL_20 RBL1_21 x826/RBL0 WBL_22 x824/VDD WBLb_17
+ WBL_16 x827/RBL1 WBLb_20 WBL_19 x827/RBL0 x828/RBL1 WBLb_22 x828/RBL0 WBL_23 x820/RBL1
+ VSUBS x10T_1x8_magic
X10T_1x8_magic_58 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x70/WWL RWL_5 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x70/VDD VSUBS x829/RBL0 x830/WBLb x830/RBL1 x831/WBLb x832/WBL x830/RBL0
+ x831/RBL1 x833/WBLb x831/RBL0 x834/WBL x833/RBL1 x833/RBL0 x832/WBLb x835/WBL x836/WWL
+ x832/RBL1 x834/WBLb x832/RBL0 x837/WBL x834/RBL1 x834/RBL0 x829/WBL x836/VDD x835/WBLb
+ x830/WBL x835/RBL1 x837/WBLb x831/WBL x835/RBL0 x837/RBL1 x829/WBLb x837/RBL0 x833/WBL
+ x829/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_69 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x767/WWL RWL_29 WBLb_24
+ WBL_24 WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29
+ WBLb_30 WBL_30 WBLb_31 WBL_31 x767/VDD VSUBS x838/RBL0 x839/WBLb x839/RBL1 x840/WBLb
+ x841/WBL x839/RBL0 x840/RBL1 x842/WBLb x840/RBL0 x843/WBL x842/RBL1 x842/RBL0 x841/WBLb
+ x844/WBL x839/WWL x841/RBL1 x843/WBLb x841/RBL0 x845/WBL x843/RBL1 x843/RBL0 x838/WBL
+ x839/VDD x844/WBLb x839/WBL x844/RBL1 x845/WBLb x840/WBL x844/RBL0 x845/RBL1 x838/WBLb
+ x845/RBL0 x842/WBL x838/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_36 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x583/WWL RWL_26 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x583/VDD VSUBS x846/RBL0 x847/WBLb x847/RBL1 x848/WBLb x849/WBL x847/RBL0
+ x848/RBL1 x850/WBLb x848/RBL0 x851/WBL x850/RBL1 x850/RBL0 x849/WBLb x852/WBL x286/WWL
+ x849/RBL1 x851/WBLb x849/RBL0 x853/WBL x851/RBL1 x851/RBL0 x846/WBL x286/VDD x852/WBLb
+ x847/WBL x852/RBL1 x853/WBLb x848/WBL x852/RBL0 x853/RBL1 x846/WBLb x853/RBL0 x850/WBL
+ x846/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_25 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_21 RWL_21 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x854/RBL0
+ x855/WBLb x855/RBL1 x856/WBLb x857/WBL x855/RBL0 x856/RBL1 x858/WBLb x856/RBL0 x859/WBL
+ x858/RBL1 x858/RBL0 x857/WBLb x860/WBL x388/WWL x857/RBL1 x859/WBLb x857/RBL0 x861/WBL
+ x859/RBL1 x859/RBL0 x854/WBL x388/VDD x860/WBLb x855/WBL x860/RBL1 x861/WBLb x856/WBL
+ x860/RBL0 x861/RBL1 x854/WBLb x861/RBL0 x858/WBL x854/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_47 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x414/WWL RWL_16 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x414/VDD VSUBS x862/RBL0 x863/WBLb x863/RBL1 x864/WBLb x865/WBL x863/RBL0
+ x864/RBL1 x866/WBLb x864/RBL0 x867/WBL x866/RBL1 x866/RBL0 x865/WBLb x868/WBL x185/WWL
+ x865/RBL1 x867/WBLb x865/RBL0 x869/WBL x867/RBL1 x867/RBL0 x862/WBL x185/VDD x868/WBLb
+ x863/WBL x868/RBL1 x869/WBLb x864/WBL x868/RBL0 x869/RBL1 x862/WBLb x869/RBL0 x866/WBL
+ x862/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_105 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x441/WWL RWL_10 WBLb_16
+ WBL_16 WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21
+ WBLb_22 WBL_22 WBLb_23 WBL_23 x441/VDD VSUBS x870/RBL0 WBLb_16 x871/RBL1 x872/WBLb
+ x873/WBL x871/RBL0 x872/RBL1 x874/WBLb x872/RBL0 x875/WBL x874/RBL1 x874/RBL0 x873/WBLb
+ x876/WBL x877/WWL x873/RBL1 x875/WBLb x873/RBL0 x878/WBL RBL1_21 x875/RBL0 x870/WBL
+ x877/VDD x876/WBLb x871/WBL x876/RBL1 x878/WBLb x872/WBL x876/RBL0 x878/RBL1 x870/WBLb
+ x878/RBL0 x874/WBL x870/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_14 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_8 RWL_8 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x879/RBL0
+ x880/WBLb x880/RBL1 x881/WBLb x882/WBL x880/RBL0 x881/RBL1 x883/WBLb x881/RBL0 x884/WBL
+ x883/RBL1 x883/RBL0 x882/WBLb x885/WBL x632/WWL x882/RBL1 x884/WBLb x882/RBL0 x886/WBL
+ x884/RBL1 x884/RBL0 x879/WBL x632/VDD x885/WBLb x880/WBL x885/RBL1 x886/WBLb x881/WBL
+ x885/RBL0 x886/RBL1 x879/WBLb x886/RBL0 x883/WBL x879/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_59 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x58/WWL RWL_4 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x58/VDD VSUBS x887/RBL0 WBLb_8 x888/RBL1 WBLb_11 WBL_10 x888/RBL0
+ x889/RBL1 WBLb_15 x889/RBL0 WBL_13 x890/RBL1 x890/RBL0 WBLb_10 WBL_9 x819/WWL x891/RBL1
+ WBLb_13 x891/RBL0 WBL_12 x892/RBL1 x892/RBL0 WBL_14 x819/VDD WBLb_9 WBL_8 x893/RBL1
+ WBLb_12 WBL_11 x893/RBL0 x894/RBL1 WBLb_14 x894/RBL0 WBL_15 x887/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_117 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x836/WWL RWL_5 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x836/VDD VSUBS x895/RBL0 WBLb_16 x896/RBL1 x897/WBLb x898/WBL
+ x896/RBL0 x897/RBL1 x899/WBLb x897/RBL0 x900/WBL x899/RBL1 x899/RBL0 x898/WBLb x901/WBL
+ x902/WWL x898/RBL1 x900/WBLb x898/RBL0 x903/WBL RBL1_21 x900/RBL0 x895/WBL x902/VDD
+ x901/WBLb x896/WBL x901/RBL1 x903/WBLb x897/WBL x901/RBL0 x903/RBL1 x895/WBLb x903/RBL0
+ x899/WBL x895/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_37 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x904/WWL RWL_27 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x904/VDD VSUBS x905/RBL0 x906/WBLb x906/RBL1 x907/WBLb x908/WBL x906/RBL0
+ x907/RBL1 x909/WBLb x907/RBL0 x910/WBL x909/RBL1 x909/RBL0 x908/WBLb x911/WBL x167/WWL
+ x908/RBL1 x910/WBLb x908/RBL0 x912/WBL x910/RBL1 x910/RBL0 x905/WBL x167/VDD x911/WBLb
+ x906/WBL x911/RBL1 x912/WBLb x907/WBL x911/RBL0 x912/RBL1 x905/WBLb x912/RBL0 x909/WBL
+ x905/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_26 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_22 RWL_22 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x913/RBL0
+ x914/WBLb x914/RBL1 x915/WBLb x916/WBL x914/RBL0 x915/RBL1 x917/WBLb x915/RBL0 x918/WBL
+ x917/RBL1 x917/RBL0 x916/WBLb x919/WBL x296/WWL x916/RBL1 x918/WBLb x916/RBL0 x920/WBL
+ x918/RBL1 x918/RBL0 x913/WBL x296/VDD x919/WBLb x914/WBL x919/RBL1 x920/WBLb x915/WBL
+ x919/RBL0 x920/RBL1 x913/WBLb x920/RBL0 x917/WBL x913/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_48 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x121/WWL RWL_15 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x121/VDD VSUBS x921/RBL0 x922/WBLb x922/RBL1 x923/WBLb x924/WBL x922/RBL0
+ x923/RBL1 x925/WBLb x923/RBL0 x926/WBL x925/RBL1 x925/RBL0 x924/WBLb x927/WBL x322/WWL
+ x924/RBL1 x926/WBLb x924/RBL0 x928/WBL x926/RBL1 x926/RBL0 x921/WBL x322/VDD x927/WBLb
+ x922/WBL x927/RBL1 x928/WBLb x923/WBL x927/RBL0 x928/RBL1 x921/WBLb x928/RBL0 x925/WBL
+ x921/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_106 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x801/WWL RWL_11 WBLb_24
+ WBL_24 WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29
+ WBLb_30 WBL_30 WBLb_31 WBL_31 x801/VDD VSUBS x929/RBL0 x930/WBLb x930/RBL1 x931/WBLb
+ x932/WBL x930/RBL0 x931/RBL1 x933/WBLb x931/RBL0 x934/WBL x933/RBL1 x933/RBL0 x932/WBLb
+ x935/WBL x930/WWL x932/RBL1 x934/WBLb x932/RBL0 x936/WBL x934/RBL1 x934/RBL0 x929/WBL
+ x930/VDD x935/WBLb x930/WBL x935/RBL1 x936/WBLb x931/WBL x935/RBL0 x936/RBL1 x929/WBLb
+ x936/RBL0 x933/WBL x929/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_15 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_9 RWL_9 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND RBL0_6
+ WBLb_0 RBL1_0 WBLb_3 WBL_2 RBL0_0 RBL1_3 WBLb_7 RBL0_3 WBL_5 RBL1_7 RBL0_7 WBLb_2
+ WBL_1 x540/WWL RBL1_2 WBLb_5 RBL0_2 WBL_4 RBL1_5 RBL0_5 WBL_6 x540/VDD WBLb_1 WBL_0
+ RBL1_1 WBLb_4 WBL_3 RBL0_1 RBL1_4 WBLb_6 RBL0_4 WBL_7 RBL1_6 VSUBS x10T_1x8_magic
X10T_1x8_magic_118 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x902/WWL RWL_5 WBLb_24 WBL_24
+ WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29 WBLb_30
+ WBL_30 WBLb_31 WBL_31 x902/VDD VSUBS x937/RBL0 x938/WBLb x938/RBL1 x939/WBLb x940/WBL
+ x938/RBL0 x939/RBL1 x941/WBLb x939/RBL0 x942/WBL x941/RBL1 x941/RBL0 x940/WBLb x943/WBL
+ x938/WWL x940/RBL1 x942/WBLb x940/RBL0 x944/WBL x942/RBL1 x942/RBL0 x937/WBL x938/VDD
+ x943/WBLb x938/WBL x943/RBL1 x944/WBLb x939/WBL x943/RBL0 x944/RBL1 x937/WBLb x944/RBL0
+ x941/WBL x937/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_16 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_31 RWL_31 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x945/RBL0
+ x946/WBLb x946/RBL1 x947/WBLb x948/WBL x946/RBL0 x947/RBL1 x949/WBLb x947/RBL0 x950/WBL
+ x949/RBL1 x949/RBL0 x948/WBLb x951/WBL x559/WWL x948/RBL1 x950/WBLb x948/RBL0 x952/WBL
+ x950/RBL1 x950/RBL0 x945/WBL x559/VDD x951/WBLb x946/WBL x951/RBL1 x952/WBLb x947/WBL
+ x951/RBL0 x952/RBL1 x945/WBLb x952/RBL0 x949/WBL x945/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_38 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x784/WWL RWL_24 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x784/VDD VSUBS x953/RBL0 x954/WBLb x954/RBL1 x955/WBLb x956/WBL x954/RBL0
+ x955/RBL1 x957/WBLb x955/RBL0 x958/WBL x957/RBL1 x957/RBL0 x956/WBLb x959/WBL x585/WWL
+ x956/RBL1 x958/WBLb x956/RBL0 x960/WBL x958/RBL1 x958/RBL0 x953/WBL x585/VDD x959/WBLb
+ x954/WBL x959/RBL1 x960/WBLb x955/WBL x959/RBL0 x960/RBL1 x953/WBLb x960/RBL0 x957/WBL
+ x953/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_27 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_19 RWL_19 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x961/RBL0
+ x962/WBLb x962/RBL1 x963/WBLb x964/WBL x962/RBL0 x963/RBL1 x965/WBLb x963/RBL0 x966/WBL
+ x965/RBL1 x965/RBL0 x964/WBLb x967/WBL x595/WWL x964/RBL1 x966/WBLb x964/RBL0 x968/WBL
+ x966/RBL1 x966/RBL0 x961/WBL x595/VDD x967/WBLb x962/WBL x967/RBL1 x968/WBLb x963/WBL
+ x967/RBL0 x968/RBL1 x961/WBLb x968/RBL0 x965/WBL x961/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_49 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x82/WWL RWL_14 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 x82/VDD VSUBS RBL0_14 WBLb_8 RBL1_8 WBLb_11 WBL_10 RBL0_8 RBL1_11
+ WBLb_15 RBL0_11 WBL_13 RBL1_15 RBL0_15 WBLb_10 WBL_9 x522/WWL RBL1_10 WBLb_13 RBL0_10
+ WBL_12 RBL1_13 RBL0_13 WBL_14 x522/VDD WBLb_9 WBL_8 RBL1_9 WBLb_12 WBL_11 RBL0_9
+ RBL1_12 WBLb_14 RBL0_12 WBL_15 RBL1_14 VSUBS x10T_1x8_magic
X10T_1x8_magic_107 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x877/WWL RWL_10 WBLb_24
+ WBL_24 WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29
+ WBLb_30 WBL_30 WBLb_31 WBL_31 x877/VDD VSUBS x969/RBL0 x970/WBLb x970/RBL1 x971/WBLb
+ x972/WBL x970/RBL0 x971/RBL1 x973/WBLb x971/RBL0 x974/WBL x973/RBL1 x973/RBL0 x972/WBLb
+ x975/WBL x970/WWL x972/RBL1 x974/WBLb x972/RBL0 x976/WBL x974/RBL1 x974/RBL0 x969/WBL
+ x970/VDD x975/WBLb x970/WBL x975/RBL1 x976/WBLb x971/WBL x975/RBL0 x976/RBL1 x969/WBLb
+ x976/RBL0 x973/WBL x969/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_119 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x824/WWL RWL_4 WBLb_24 WBL_24
+ WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29 WBLb_30
+ WBL_30 WBLb_31 WBL_31 x824/VDD VSUBS x977/RBL0 WBLb_24 x978/RBL1 WBLb_27 WBL_26
+ x978/RBL0 x979/RBL1 WBLb_31 x979/RBL0 WBL_29 x980/RBL1 x980/RBL0 WBLb_26 WBL_25
+ x978/WWL x981/RBL1 WBLb_29 x981/RBL0 WBL_28 x982/RBL1 x982/RBL0 WBL_30 x978/VDD
+ WBLb_25 WBL_24 x983/RBL1 WBLb_28 WBL_27 x983/RBL0 x984/RBL1 WBLb_30 x984/RBL0 WBL_31
+ x977/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_17 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_29 RWL_29 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x985/RBL0
+ x986/WBLb x986/RBL1 x987/WBLb x988/WBL x986/RBL0 x987/RBL1 x989/WBLb x987/RBL0 x990/WBL
+ x989/RBL1 x989/RBL0 x988/WBLb x991/WBL x750/WWL x988/RBL1 x990/WBLb x988/RBL0 x992/WBL
+ x990/RBL1 x990/RBL0 x985/WBL x750/VDD x991/WBLb x986/WBL x991/RBL1 x992/WBLb x987/WBL
+ x991/RBL0 x992/RBL1 x985/WBLb x992/RBL0 x989/WBL x985/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_39 RBL1_8 RBL0_8 RBL1_9 RBL0_9 RBL1_10 RBL0_10 RBL1_11 RBL1_12 RBL0_12
+ RBL1_13 RBL0_13 RBL1_14 RBL0_14 RBL1_15 RBL0_15 x699/WWL RWL_23 WBLb_8 WBL_8 WBLb_9
+ WBL_9 WBLb_10 WBL_10 WBLb_11 WBL_11 WBLb_12 WBL_12 WBLb_13 WBL_13 WBLb_14 WBL_14
+ WBLb_15 WBL_15 VDD VSUBS RBL0_14 WBLb_8 RBL1_8 WBLb_11 WBL_10 RBL0_8 RBL1_11 WBLb_15
+ RBL0_11 WBL_13 RBL1_15 RBL0_15 WBLb_10 WBL_9 x83/WWL RBL1_10 WBLb_13 RBL0_10 WBL_12
+ RBL1_13 RBL0_13 WBL_14 VDD WBLb_9 WBL_8 RBL1_9 WBLb_12 WBL_11 RBL0_9 RBL1_12 WBLb_14
+ RBL0_12 WBL_15 RBL1_14 VSUBS x10T_1x8_magic
X10T_1x8_magic_28 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_20 RWL_20 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x993/RBL0
+ x994/WBLb x994/RBL1 x995/WBLb x996/WBL x994/RBL0 x995/RBL1 x997/WBLb x995/RBL0 x998/WBL
+ x997/RBL1 x997/RBL0 x996/WBLb x999/WBL x505/WWL x996/RBL1 x998/WBLb x996/RBL0 x1000/WBL
+ x998/RBL1 x998/RBL0 x993/WBL VDD x999/WBLb x994/WBL x999/RBL1 x1000/WBLb x995/WBL
+ x999/RBL0 x1000/RBL1 x993/WBLb x1000/RBL0 x997/WBL x993/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_108 RBL1_16 RBL0_16 RBL1_17 RBL0_17 RBL1_18 RBL0_18 RBL1_19 RBL1_20
+ RBL0_20 RBL1_21 RBL0_21 RBL1_22 RBL0_22 RBL1_23 RBL0_23 x541/WWL RWL_9 WBLb_16 WBL_16
+ WBLb_17 WBL_17 WBLb_18 WBL_18 WBLb_19 WBL_19 WBLb_20 WBL_20 WBLb_21 WBL_21 WBLb_22
+ WBL_22 WBLb_23 WBL_23 x541/VDD VSUBS RBL0_22 WBLb_16 RBL1_16 WBLb_19 WBL_18 RBL0_16
+ RBL1_19 WBLb_23 RBL0_19 WBL_21 RBL1_23 RBL0_23 WBLb_18 WBL_17 x1001/WWL RBL1_18
+ WBLb_21 RBL0_18 WBL_20 RBL1_21 RBL0_21 WBL_22 x1001/VDD WBLb_17 WBL_16 RBL1_17 WBLb_20
+ WBL_19 RBL0_17 RBL1_20 WBLb_22 RBL0_20 WBL_23 RBL1_22 VSUBS x10T_1x8_magic
X10T_1x8_magic_18 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_30 RWL_30 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x1002/RBL0
+ x1003/WBLb x1003/RBL1 x1004/WBLb x1005/WBL x1003/RBL0 x1004/RBL1 x1006/WBLb x1004/RBL0
+ x1007/WBL x1006/RBL1 x1006/RBL0 x1005/WBLb x1008/WBL x469/WWL x1005/RBL1 x1007/WBLb
+ x1005/RBL0 x1009/WBL x1007/RBL1 x1007/RBL0 x1002/WBL x469/VDD x1008/WBLb x1003/WBL
+ x1008/RBL1 x1009/WBLb x1004/WBL x1008/RBL0 x1009/RBL1 x1002/WBLb x1009/RBL0 x1006/WBL
+ x1002/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_29 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_17 RWL_17 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x1010/RBL0
+ x1011/WBLb x1011/RBL1 x1012/WBLb x1013/WBL x1011/RBL0 x1012/RBL1 x1014/WBLb x1012/RBL0
+ x1015/WBL x1014/RBL1 x1014/RBL0 x1013/WBLb x1016/WBL x708/WWL x1013/RBL1 x1015/WBLb
+ x1013/RBL0 x1017/WBL x1015/RBL1 x1015/RBL0 x1010/WBL x708/VDD x1016/WBLb x1011/WBL
+ x1016/RBL1 x1017/WBLb x1012/WBL x1016/RBL0 x1017/RBL1 x1010/WBLb x1017/RBL0 x1014/WBL
+ x1010/RBL1 VSUBS x10T_1x8_magic
X10T_1x8_magic_109 RBL1_24 RBL0_24 RBL1_25 RBL0_25 RBL1_26 RBL0_26 RBL1_27 RBL1_28
+ RBL0_28 RBL1_29 RBL0_29 RBL1_30 RBL0_30 RBL1_31 RBL0_31 x1001/WWL RWL_9 WBLb_24
+ WBL_24 WBLb_25 WBL_25 WBLb_26 WBL_26 WBLb_27 WBL_27 WBLb_28 WBL_28 WBLb_29 WBL_29
+ WBLb_30 WBL_30 WBLb_31 WBL_31 x1001/VDD VSUBS RBL0_30 WBLb_24 RBL1_24 WBLb_27 WBL_26
+ RBL0_24 RBL1_27 WBLb_31 RBL0_27 WBL_29 RBL1_31 RBL0_31 WBLb_26 WBL_25 x1018/WWL
+ RBL1_26 WBLb_29 RBL0_26 WBL_28 RBL1_29 RBL0_29 WBL_30 x1018/VDD WBLb_25 WBL_24 RBL1_25
+ WBLb_28 WBL_27 RBL0_25 RBL1_28 WBLb_30 RBL0_28 WBL_31 RBL1_30 VSUBS x10T_1x8_magic
X10T_1x8_magic_19 RBL1_0 RBL0_0 RBL1_1 RBL0_1 RBL1_2 RBL0_2 RBL1_3 RBL1_4 RBL0_4 RBL1_5
+ RBL0_5 RBL1_6 RBL0_6 RBL1_7 RBL0_7 WWL_27 RWL_27 WBLb_0 WBL_0 WBLb_1 WBL_1 WBLb_2
+ WBL_2 WBLb_3 WBL_3 WBLb_4 WBL_4 WBLb_5 WBL_5 WBLb_6 WBL_6 WBLb_7 WBL_7 VDD GND x1019/RBL0
+ x1020/WBLb x1020/RBL1 x1021/WBLb x1022/WBL x1020/RBL0 x1021/RBL1 x1023/WBLb x1021/RBL0
+ x1024/WBL x1023/RBL1 x1023/RBL0 x1022/WBLb x1025/WBL x904/WWL x1022/RBL1 x1024/WBLb
+ x1022/RBL0 x1026/WBL x1024/RBL1 x1024/RBL0 x1019/WBL x904/VDD x1025/WBLb x1020/WBL
+ x1025/RBL1 x1026/WBLb x1021/WBL x1025/RBL0 x1026/RBL1 x1019/WBLb x1026/RBL0 x1023/WBL
+ x1019/RBL1 VSUBS x10T_1x8_magic
.ends

